magic
tech scmos
magscale 1 30
timestamp 1719895877
<< checkpaint >>
rect 47800 171700 61200 180850
rect 18300 145440 61200 171700
rect 18300 145200 44800 145440
rect 47800 145200 61200 145440
rect 61300 145200 74700 180850
rect 74800 145200 88200 180850
rect 88300 146970 101700 180850
rect 101900 146970 115100 180850
rect 88300 145200 115100 146970
rect 115300 145200 128700 180850
rect 128800 171700 142200 180850
rect 128800 145440 171700 171700
rect 128800 145200 142200 145440
rect 145200 145200 171700 145440
rect 18300 142200 44650 145200
rect 9150 128800 44800 142200
rect 101100 140200 103040 145200
rect 145440 142200 171700 145200
rect 145200 128800 180850 142200
rect 9150 115300 44800 128700
rect 145200 115300 180850 128700
rect 9150 101800 44800 115200
rect 145200 101800 180850 115200
rect 9150 88300 44800 101700
rect 145200 88300 180850 101700
rect 9150 74900 44800 88100
rect 45930 85530 47165 85855
rect 45055 77480 47165 85530
rect 145200 74800 180850 88200
rect 9150 61300 44800 74700
rect 145200 61300 180850 74700
rect 9150 47800 44800 61200
rect 145200 47800 180850 61200
rect 18300 44800 44560 47800
rect 97740 45875 100710 47165
rect 99000 45640 100610 45875
rect 145440 44800 171700 47800
rect 18300 44560 44800 44800
rect 47800 44560 61200 44800
rect 18300 18300 61200 44560
rect 47800 9150 61200 18300
rect 61300 9150 74700 44800
rect 74800 9150 88200 44800
rect 88300 9150 101700 44800
rect 101800 9150 115200 44800
rect 115300 9150 128700 44800
rect 128800 44560 142200 44800
rect 145200 44560 171700 44800
rect 128800 18300 171700 44560
rect 128800 9150 142200 18300
<< error_p >>
rect 46660 140300 77250 140440
rect 90420 140300 101100 140440
rect 46660 140260 101100 140300
rect 105100 140260 132000 140440
rect 46660 136360 143140 136540
rect 46660 132460 143140 132640
rect 46660 128560 143140 128740
rect 46660 124660 143140 124840
rect 46660 120760 143140 120940
rect 46660 116860 142840 117040
rect 46660 112960 142840 113140
rect 46660 109060 142840 109240
rect 48000 105160 143140 105340
rect 48570 101260 143140 101440
rect 48000 97360 143140 97540
rect 47160 93460 143140 93640
rect 47160 89560 143140 89740
rect 47160 85660 143140 85840
rect 47160 81760 143140 81940
rect 47160 77860 143140 78040
rect 47160 73960 143140 74140
rect 46660 70060 143090 70240
rect 46660 66160 143090 66340
rect 46660 62260 143090 62440
rect 46660 58360 143090 58540
rect 46660 54460 143140 54640
rect 46660 50560 143140 50740
rect 48000 46660 60000 46840
rect 72000 46660 84000 46840
rect 120000 46800 143140 46840
rect 142200 46660 143140 46800
<< error_s >>
rect 44065 171030 44145 171040
rect 44385 171030 44465 171040
rect 44705 171030 44785 171040
rect 45025 171030 45105 171040
rect 45345 171030 45425 171040
rect 45665 171030 45745 171040
rect 45985 171030 46065 171040
rect 46305 171030 46385 171040
rect 46625 171030 46705 171040
rect 46945 171030 47025 171040
rect 47265 171030 47345 171040
rect 47585 171030 47665 171040
rect 47905 171030 47985 171040
rect 48225 171030 48305 171040
rect 48500 171030 48605 171100
rect 44145 170950 44155 171030
rect 44465 170950 44475 171030
rect 44785 170950 44795 171030
rect 45105 170950 45115 171030
rect 45425 170950 45435 171030
rect 45745 170950 45755 171030
rect 46065 170950 46075 171030
rect 46385 170950 46395 171030
rect 46705 170950 46715 171030
rect 47025 170950 47035 171030
rect 47345 170950 47355 171030
rect 47665 170950 47675 171030
rect 47985 170950 47995 171030
rect 48305 170950 48315 171030
rect 48500 171020 48640 171030
rect 48710 171020 48790 171030
rect 60060 171020 60140 171030
rect 60210 171020 60290 171030
rect 60360 171020 60440 171030
rect 60610 171029 60690 171039
rect 60930 171029 61010 171039
rect 61350 171029 61430 171039
rect 61670 171029 61750 171039
rect 43060 170940 43140 170950
rect 43380 170940 43460 170950
rect 43140 170860 43150 170940
rect 43460 170860 43470 170940
rect 43905 170870 43985 170880
rect 44225 170870 44305 170880
rect 44545 170870 44625 170880
rect 44865 170870 44945 170880
rect 45185 170870 45265 170880
rect 45505 170870 45585 170880
rect 45825 170870 45905 170880
rect 46145 170870 46225 170880
rect 46465 170870 46545 170880
rect 46785 170870 46865 170880
rect 47105 170870 47185 170880
rect 47425 170870 47505 170880
rect 47745 170870 47825 170880
rect 48065 170870 48145 170880
rect 43985 170790 43995 170870
rect 44305 170790 44315 170870
rect 44625 170790 44635 170870
rect 44945 170790 44955 170870
rect 45265 170790 45275 170870
rect 45585 170790 45595 170870
rect 45905 170790 45915 170870
rect 46225 170790 46235 170870
rect 46545 170790 46555 170870
rect 46865 170790 46875 170870
rect 47185 170790 47195 170870
rect 47505 170790 47515 170870
rect 47825 170790 47835 170870
rect 48145 170790 48155 170870
rect 48500 170850 48605 171020
rect 48640 170940 48650 171020
rect 48790 170940 48800 171020
rect 49180 170960 49210 170990
rect 49300 170960 49330 170990
rect 49420 170960 49450 170990
rect 49540 170960 49570 170990
rect 49660 170960 49690 170990
rect 49780 170960 49810 170990
rect 49900 170960 49930 170990
rect 50020 170960 50050 170990
rect 50140 170960 50170 170990
rect 50260 170960 50290 170990
rect 50380 170960 50410 170990
rect 50500 170960 50530 170990
rect 50620 170960 50650 170990
rect 50740 170960 50770 170990
rect 50860 170960 50890 170990
rect 50980 170960 51010 170990
rect 51100 170960 51130 170990
rect 51220 170960 51250 170990
rect 51340 170960 51370 170990
rect 51460 170960 51490 170990
rect 51580 170960 51610 170990
rect 51700 170960 51730 170990
rect 51820 170960 51850 170990
rect 51940 170960 51970 170990
rect 52060 170960 52090 170990
rect 52180 170960 52210 170990
rect 52300 170960 52330 170990
rect 52420 170960 52450 170990
rect 52540 170960 52570 170990
rect 52660 170960 52690 170990
rect 52780 170960 52810 170990
rect 52900 170960 52930 170990
rect 53020 170960 53050 170990
rect 53140 170960 53170 170990
rect 53260 170960 53290 170990
rect 53380 170960 53410 170990
rect 53500 170960 53530 170990
rect 53620 170960 53650 170990
rect 53740 170960 53770 170990
rect 53860 170960 53890 170990
rect 53980 170960 54010 170990
rect 54100 170960 54130 170990
rect 54220 170960 54250 170990
rect 54340 170960 54370 170990
rect 54460 170960 54490 170990
rect 54580 170960 54610 170990
rect 54700 170960 54730 170990
rect 54820 170960 54850 170990
rect 54940 170960 54970 170990
rect 55060 170960 55090 170990
rect 55180 170960 55210 170990
rect 55300 170960 55330 170990
rect 55420 170960 55450 170990
rect 55540 170960 55570 170990
rect 55660 170960 55690 170990
rect 55780 170960 55810 170990
rect 55900 170960 55930 170990
rect 56020 170960 56050 170990
rect 56140 170960 56170 170990
rect 56260 170960 56290 170990
rect 56380 170960 56410 170990
rect 56500 170960 56530 170990
rect 56620 170960 56650 170990
rect 56740 170960 56770 170990
rect 56860 170960 56890 170990
rect 56980 170960 57010 170990
rect 57100 170960 57130 170990
rect 57220 170960 57250 170990
rect 57340 170960 57370 170990
rect 57460 170960 57490 170990
rect 57580 170960 57610 170990
rect 57700 170960 57730 170990
rect 57820 170960 57850 170990
rect 57940 170960 57970 170990
rect 58060 170960 58090 170990
rect 58180 170960 58210 170990
rect 58300 170960 58330 170990
rect 58420 170960 58450 170990
rect 58540 170960 58570 170990
rect 58660 170960 58690 170990
rect 58780 170960 58810 170990
rect 58900 170960 58930 170990
rect 59020 170960 59050 170990
rect 59140 170960 59170 170990
rect 59260 170960 59290 170990
rect 59380 170960 59410 170990
rect 59500 170960 59530 170990
rect 59620 170960 59650 170990
rect 59740 170960 59770 170990
rect 49060 170930 49120 170960
rect 49180 170930 49240 170960
rect 49300 170930 49360 170960
rect 49420 170930 49480 170960
rect 49540 170930 49600 170960
rect 49660 170930 49720 170960
rect 49780 170930 49840 170960
rect 49900 170930 49960 170960
rect 50020 170930 50080 170960
rect 50140 170930 50200 170960
rect 50260 170930 50320 170960
rect 50380 170930 50440 170960
rect 50500 170930 50560 170960
rect 50620 170930 50680 170960
rect 50740 170930 50800 170960
rect 50860 170930 50920 170960
rect 50980 170930 51040 170960
rect 51100 170930 51160 170960
rect 51220 170930 51280 170960
rect 51340 170930 51400 170960
rect 51460 170930 51520 170960
rect 51580 170930 51640 170960
rect 51700 170930 51760 170960
rect 51820 170930 51880 170960
rect 51940 170930 52000 170960
rect 52060 170930 52120 170960
rect 52180 170930 52240 170960
rect 52300 170930 52360 170960
rect 52420 170930 52480 170960
rect 52540 170930 52600 170960
rect 52660 170930 52720 170960
rect 52780 170930 52840 170960
rect 52900 170930 52960 170960
rect 53020 170930 53080 170960
rect 53140 170930 53200 170960
rect 53260 170930 53320 170960
rect 53380 170930 53440 170960
rect 53500 170930 53560 170960
rect 53620 170930 53680 170960
rect 53740 170930 53800 170960
rect 53860 170930 53920 170960
rect 53980 170930 54040 170960
rect 54100 170930 54160 170960
rect 54220 170930 54280 170960
rect 54340 170930 54400 170960
rect 54460 170930 54520 170960
rect 54580 170930 54640 170960
rect 54700 170930 54760 170960
rect 54820 170930 54880 170960
rect 54940 170930 55000 170960
rect 55060 170930 55120 170960
rect 55180 170930 55240 170960
rect 55300 170930 55360 170960
rect 55420 170930 55480 170960
rect 55540 170930 55600 170960
rect 55660 170930 55720 170960
rect 55780 170930 55840 170960
rect 55900 170930 55960 170960
rect 56020 170930 56080 170960
rect 56140 170930 56200 170960
rect 56260 170930 56320 170960
rect 56380 170930 56440 170960
rect 56500 170930 56560 170960
rect 56620 170930 56680 170960
rect 56740 170930 56800 170960
rect 56860 170930 56920 170960
rect 56980 170930 57040 170960
rect 57100 170930 57160 170960
rect 57220 170930 57280 170960
rect 57340 170930 57400 170960
rect 57460 170930 57520 170960
rect 57580 170930 57640 170960
rect 57700 170930 57760 170960
rect 57820 170930 57880 170960
rect 57940 170930 58000 170960
rect 58060 170930 58120 170960
rect 58180 170930 58240 170960
rect 58300 170930 58360 170960
rect 58420 170930 58480 170960
rect 58540 170930 58600 170960
rect 58660 170930 58720 170960
rect 58780 170930 58840 170960
rect 58900 170930 58960 170960
rect 59020 170930 59080 170960
rect 59140 170930 59200 170960
rect 59260 170930 59320 170960
rect 59380 170930 59440 170960
rect 59500 170930 59560 170960
rect 59620 170930 59680 170960
rect 59740 170930 59800 170960
rect 60140 170940 60150 171020
rect 60290 170940 60300 171020
rect 60440 170940 60450 171020
rect 60690 170949 60700 171029
rect 61010 170949 61020 171029
rect 61430 170949 61440 171029
rect 61750 170949 61760 171029
rect 62060 171020 62140 171030
rect 62210 171020 62290 171030
rect 73560 171020 73640 171030
rect 73710 171020 73790 171030
rect 73860 171020 73940 171030
rect 74110 171029 74190 171039
rect 74430 171029 74510 171039
rect 74850 171029 74930 171039
rect 75170 171029 75250 171039
rect 62140 170940 62150 171020
rect 62290 170940 62300 171020
rect 62680 170960 62710 170990
rect 73245 170960 73270 170990
rect 62560 170930 62620 170960
rect 62680 170930 62740 170960
rect 73245 170930 73300 170960
rect 73640 170940 73650 171020
rect 73790 170940 73800 171020
rect 73940 170940 73950 171020
rect 74190 170949 74200 171029
rect 74510 170949 74520 171029
rect 74930 170949 74940 171029
rect 75250 170949 75260 171029
rect 75560 171020 75640 171030
rect 75710 171020 75790 171030
rect 87060 171020 87140 171030
rect 87210 171020 87290 171030
rect 87360 171020 87440 171030
rect 87610 171029 87690 171039
rect 87930 171029 88010 171039
rect 88350 171029 88430 171039
rect 88670 171029 88750 171039
rect 75640 170940 75650 171020
rect 75790 170940 75800 171020
rect 76180 170960 76210 170990
rect 86745 170960 86770 170990
rect 76060 170930 76120 170960
rect 76180 170930 76240 170960
rect 86745 170930 86800 170960
rect 87140 170940 87150 171020
rect 87290 170940 87300 171020
rect 87440 170940 87450 171020
rect 87690 170949 87700 171029
rect 88010 170949 88020 171029
rect 88430 170949 88440 171029
rect 88750 170949 88760 171029
rect 89060 171020 89140 171030
rect 89210 171020 89290 171030
rect 100560 171020 100640 171030
rect 100710 171020 100790 171030
rect 100860 171020 100940 171030
rect 101110 171029 101190 171039
rect 101430 171029 101510 171039
rect 101850 171029 101930 171039
rect 102170 171029 102250 171039
rect 114610 171029 114690 171039
rect 114930 171029 115010 171039
rect 115350 171029 115430 171039
rect 115670 171029 115750 171039
rect 89140 170940 89150 171020
rect 89290 170940 89300 171020
rect 89680 170960 89710 170990
rect 100245 170960 100270 170990
rect 89560 170930 89620 170960
rect 89680 170930 89740 170960
rect 100245 170930 100300 170960
rect 100640 170940 100650 171020
rect 100790 170940 100800 171020
rect 100940 170940 100950 171020
rect 101190 170949 101200 171029
rect 101510 170949 101520 171029
rect 101930 170949 101940 171029
rect 102250 170949 102260 171029
rect 114690 170949 114700 171029
rect 115010 170949 115020 171029
rect 115430 170949 115440 171029
rect 115750 170949 115760 171029
rect 116060 171020 116140 171030
rect 116210 171020 116290 171030
rect 127560 171020 127640 171030
rect 127710 171020 127790 171030
rect 127860 171020 127940 171030
rect 128110 171029 128190 171039
rect 128430 171029 128510 171039
rect 128850 171029 128930 171039
rect 129170 171029 129250 171039
rect 141825 171030 141905 171040
rect 142145 171030 142200 171040
rect 145345 171030 145425 171040
rect 145665 171030 145745 171040
rect 145985 171030 146065 171040
rect 116140 170940 116150 171020
rect 116290 170940 116300 171020
rect 116680 170960 116710 170990
rect 127245 170960 127270 170990
rect 116560 170930 116620 170960
rect 116680 170930 116740 170960
rect 127245 170930 127300 170960
rect 127640 170940 127650 171020
rect 127790 170940 127800 171020
rect 127940 170940 127950 171020
rect 128190 170949 128200 171029
rect 128510 170949 128520 171029
rect 128930 170949 128940 171029
rect 129250 170949 129260 171029
rect 129560 171020 129640 171030
rect 129710 171020 129790 171030
rect 141060 171020 141140 171030
rect 141210 171020 141290 171030
rect 141360 171020 141440 171030
rect 129640 170940 129650 171020
rect 129790 170940 129800 171020
rect 130180 170960 130210 170990
rect 140740 170960 140770 170990
rect 130060 170930 130120 170960
rect 130180 170930 130240 170960
rect 140740 170930 140800 170960
rect 141140 170940 141150 171020
rect 141290 170940 141300 171020
rect 141440 170940 141450 171020
rect 141905 170950 141915 171030
rect 145425 170950 145435 171030
rect 145745 170950 145755 171030
rect 146065 170950 146075 171030
rect 146540 170940 146620 170950
rect 146860 170940 146940 170950
rect 48500 170840 48640 170850
rect 48710 170840 48790 170850
rect 49180 170840 49210 170870
rect 49300 170840 49330 170870
rect 49420 170840 49450 170870
rect 49540 170840 49570 170870
rect 49660 170840 49690 170870
rect 49780 170840 49810 170870
rect 49900 170840 49930 170870
rect 50020 170840 50050 170870
rect 50140 170840 50170 170870
rect 50260 170840 50290 170870
rect 50380 170840 50410 170870
rect 50500 170840 50530 170870
rect 50620 170840 50650 170870
rect 50740 170840 50770 170870
rect 50860 170840 50890 170870
rect 50980 170840 51010 170870
rect 51100 170840 51130 170870
rect 51220 170840 51250 170870
rect 51340 170840 51370 170870
rect 51460 170840 51490 170870
rect 51580 170840 51610 170870
rect 51700 170840 51730 170870
rect 51820 170840 51850 170870
rect 51940 170840 51970 170870
rect 52060 170840 52090 170870
rect 52180 170840 52210 170870
rect 52300 170840 52330 170870
rect 52420 170840 52450 170870
rect 52540 170840 52570 170870
rect 52660 170840 52690 170870
rect 52780 170840 52810 170870
rect 52900 170840 52930 170870
rect 53020 170840 53050 170870
rect 53140 170840 53170 170870
rect 53260 170840 53290 170870
rect 53380 170840 53410 170870
rect 53500 170840 53530 170870
rect 53620 170840 53650 170870
rect 53740 170840 53770 170870
rect 53860 170840 53890 170870
rect 53980 170840 54010 170870
rect 54100 170840 54130 170870
rect 54220 170840 54250 170870
rect 54340 170840 54370 170870
rect 54460 170840 54490 170870
rect 54580 170840 54610 170870
rect 54700 170840 54730 170870
rect 54820 170840 54850 170870
rect 54940 170840 54970 170870
rect 55060 170840 55090 170870
rect 55180 170840 55210 170870
rect 55300 170840 55330 170870
rect 55420 170840 55450 170870
rect 55540 170840 55570 170870
rect 55660 170840 55690 170870
rect 55780 170840 55810 170870
rect 55900 170840 55930 170870
rect 56020 170840 56050 170870
rect 56140 170840 56170 170870
rect 56260 170840 56290 170870
rect 56380 170840 56410 170870
rect 56500 170840 56530 170870
rect 56620 170840 56650 170870
rect 56740 170840 56770 170870
rect 56860 170840 56890 170870
rect 56980 170840 57010 170870
rect 57100 170840 57130 170870
rect 57220 170840 57250 170870
rect 57340 170840 57370 170870
rect 57460 170840 57490 170870
rect 57580 170840 57610 170870
rect 57700 170840 57730 170870
rect 57820 170840 57850 170870
rect 57940 170840 57970 170870
rect 58060 170840 58090 170870
rect 58180 170840 58210 170870
rect 58300 170840 58330 170870
rect 58420 170840 58450 170870
rect 58540 170840 58570 170870
rect 58660 170840 58690 170870
rect 58780 170840 58810 170870
rect 58900 170840 58930 170870
rect 59020 170840 59050 170870
rect 59140 170840 59170 170870
rect 59260 170840 59290 170870
rect 59380 170840 59410 170870
rect 59500 170840 59530 170870
rect 59620 170840 59650 170870
rect 59740 170840 59770 170870
rect 60770 170869 60850 170879
rect 61090 170869 61170 170879
rect 61510 170869 61590 170879
rect 61830 170869 61910 170879
rect 60060 170840 60140 170850
rect 60210 170840 60290 170850
rect 60360 170840 60440 170850
rect 42950 170780 42980 170790
rect 43220 170780 43300 170790
rect 42980 170700 42990 170780
rect 43300 170700 43310 170780
rect 44065 170710 44145 170720
rect 44385 170710 44465 170720
rect 44705 170710 44785 170720
rect 45025 170710 45105 170720
rect 45345 170710 45425 170720
rect 45665 170710 45745 170720
rect 45985 170710 46065 170720
rect 46305 170710 46385 170720
rect 46625 170710 46705 170720
rect 46945 170710 47025 170720
rect 47265 170710 47345 170720
rect 47585 170710 47665 170720
rect 47905 170710 47985 170720
rect 48225 170710 48305 170720
rect 44145 170630 44155 170710
rect 44465 170630 44475 170710
rect 44785 170630 44795 170710
rect 45105 170630 45115 170710
rect 45425 170630 45435 170710
rect 45745 170630 45755 170710
rect 46065 170630 46075 170710
rect 46385 170630 46395 170710
rect 46705 170630 46715 170710
rect 47025 170630 47035 170710
rect 47345 170630 47355 170710
rect 47665 170630 47675 170710
rect 47985 170630 47995 170710
rect 48305 170630 48315 170710
rect 48500 170670 48605 170840
rect 48640 170760 48650 170840
rect 48790 170760 48800 170840
rect 49060 170810 49120 170840
rect 49180 170810 49240 170840
rect 49300 170810 49360 170840
rect 49420 170810 49480 170840
rect 49540 170810 49600 170840
rect 49660 170810 49720 170840
rect 49780 170810 49840 170840
rect 49900 170810 49960 170840
rect 50020 170810 50080 170840
rect 50140 170810 50200 170840
rect 50260 170810 50320 170840
rect 50380 170810 50440 170840
rect 50500 170810 50560 170840
rect 50620 170810 50680 170840
rect 50740 170810 50800 170840
rect 50860 170810 50920 170840
rect 50980 170810 51040 170840
rect 51100 170810 51160 170840
rect 51220 170810 51280 170840
rect 51340 170810 51400 170840
rect 51460 170810 51520 170840
rect 51580 170810 51640 170840
rect 51700 170810 51760 170840
rect 51820 170810 51880 170840
rect 51940 170810 52000 170840
rect 52060 170810 52120 170840
rect 52180 170810 52240 170840
rect 52300 170810 52360 170840
rect 52420 170810 52480 170840
rect 52540 170810 52600 170840
rect 52660 170810 52720 170840
rect 52780 170810 52840 170840
rect 52900 170810 52960 170840
rect 53020 170810 53080 170840
rect 53140 170810 53200 170840
rect 53260 170810 53320 170840
rect 53380 170810 53440 170840
rect 53500 170810 53560 170840
rect 53620 170810 53680 170840
rect 53740 170810 53800 170840
rect 53860 170810 53920 170840
rect 53980 170810 54040 170840
rect 54100 170810 54160 170840
rect 54220 170810 54280 170840
rect 54340 170810 54400 170840
rect 54460 170810 54520 170840
rect 54580 170810 54640 170840
rect 54700 170810 54760 170840
rect 54820 170810 54880 170840
rect 54940 170810 55000 170840
rect 55060 170810 55120 170840
rect 55180 170810 55240 170840
rect 55300 170810 55360 170840
rect 55420 170810 55480 170840
rect 55540 170810 55600 170840
rect 55660 170810 55720 170840
rect 55780 170810 55840 170840
rect 55900 170810 55960 170840
rect 56020 170810 56080 170840
rect 56140 170810 56200 170840
rect 56260 170810 56320 170840
rect 56380 170810 56440 170840
rect 56500 170810 56560 170840
rect 56620 170810 56680 170840
rect 56740 170810 56800 170840
rect 56860 170810 56920 170840
rect 56980 170810 57040 170840
rect 57100 170810 57160 170840
rect 57220 170810 57280 170840
rect 57340 170810 57400 170840
rect 57460 170810 57520 170840
rect 57580 170810 57640 170840
rect 57700 170810 57760 170840
rect 57820 170810 57880 170840
rect 57940 170810 58000 170840
rect 58060 170810 58120 170840
rect 58180 170810 58240 170840
rect 58300 170810 58360 170840
rect 58420 170810 58480 170840
rect 58540 170810 58600 170840
rect 58660 170810 58720 170840
rect 58780 170810 58840 170840
rect 58900 170810 58960 170840
rect 59020 170810 59080 170840
rect 59140 170810 59200 170840
rect 59260 170810 59320 170840
rect 59380 170810 59440 170840
rect 59500 170810 59560 170840
rect 59620 170810 59680 170840
rect 59740 170810 59800 170840
rect 60140 170760 60150 170840
rect 60290 170760 60300 170840
rect 60440 170760 60450 170840
rect 60850 170789 60860 170869
rect 61170 170789 61180 170869
rect 61590 170789 61600 170869
rect 61910 170789 61920 170869
rect 62060 170840 62140 170850
rect 62210 170840 62290 170850
rect 62680 170840 62710 170870
rect 73245 170840 73270 170870
rect 74270 170869 74350 170879
rect 74590 170869 74670 170879
rect 75010 170869 75090 170879
rect 75330 170869 75410 170879
rect 73560 170840 73640 170850
rect 73710 170840 73790 170850
rect 73860 170840 73940 170850
rect 62140 170760 62150 170840
rect 62290 170760 62300 170840
rect 62560 170810 62620 170840
rect 62680 170810 62740 170840
rect 73245 170810 73300 170840
rect 73640 170760 73650 170840
rect 73790 170760 73800 170840
rect 73940 170760 73950 170840
rect 74350 170789 74360 170869
rect 74670 170789 74680 170869
rect 75090 170789 75100 170869
rect 75410 170789 75420 170869
rect 75560 170840 75640 170850
rect 75710 170840 75790 170850
rect 76180 170840 76210 170870
rect 86745 170840 86770 170870
rect 87770 170869 87850 170879
rect 88090 170869 88170 170879
rect 88510 170869 88590 170879
rect 88830 170869 88910 170879
rect 87060 170840 87140 170850
rect 87210 170840 87290 170850
rect 87360 170840 87440 170850
rect 75640 170760 75650 170840
rect 75790 170760 75800 170840
rect 76060 170810 76120 170840
rect 76180 170810 76240 170840
rect 86745 170810 86800 170840
rect 87140 170760 87150 170840
rect 87290 170760 87300 170840
rect 87440 170760 87450 170840
rect 87850 170789 87860 170869
rect 88170 170789 88180 170869
rect 88590 170789 88600 170869
rect 88910 170789 88920 170869
rect 89060 170840 89140 170850
rect 89210 170840 89290 170850
rect 89680 170840 89710 170870
rect 100245 170840 100270 170870
rect 101270 170869 101350 170879
rect 101590 170869 101670 170879
rect 102010 170869 102090 170879
rect 102330 170869 102410 170879
rect 114770 170869 114850 170879
rect 115090 170869 115170 170879
rect 115510 170869 115590 170879
rect 115830 170869 115910 170879
rect 100560 170840 100640 170850
rect 100710 170840 100790 170850
rect 100860 170840 100940 170850
rect 89140 170760 89150 170840
rect 89290 170760 89300 170840
rect 89560 170810 89620 170840
rect 89680 170810 89740 170840
rect 100245 170810 100300 170840
rect 100640 170760 100650 170840
rect 100790 170760 100800 170840
rect 100940 170760 100950 170840
rect 101350 170789 101360 170869
rect 101670 170789 101680 170869
rect 102090 170789 102100 170869
rect 102410 170789 102420 170869
rect 114850 170789 114860 170869
rect 115170 170789 115180 170869
rect 115590 170789 115600 170869
rect 115910 170789 115920 170869
rect 116060 170840 116140 170850
rect 116210 170840 116290 170850
rect 116680 170840 116710 170870
rect 127245 170840 127270 170870
rect 128270 170869 128350 170879
rect 128590 170869 128670 170879
rect 129010 170869 129090 170879
rect 129330 170869 129410 170879
rect 141665 170870 141745 170880
rect 141985 170870 142065 170880
rect 145200 170870 145265 170880
rect 145505 170870 145585 170880
rect 145825 170870 145905 170880
rect 127560 170840 127640 170850
rect 127710 170840 127790 170850
rect 127860 170840 127940 170850
rect 116140 170760 116150 170840
rect 116290 170760 116300 170840
rect 116560 170810 116620 170840
rect 116680 170810 116740 170840
rect 127245 170810 127300 170840
rect 127640 170760 127650 170840
rect 127790 170760 127800 170840
rect 127940 170760 127950 170840
rect 128350 170789 128360 170869
rect 128670 170789 128680 170869
rect 129090 170789 129100 170869
rect 129410 170789 129420 170869
rect 129560 170840 129640 170850
rect 129710 170840 129790 170850
rect 130180 170840 130210 170870
rect 140740 170840 140770 170870
rect 141060 170840 141140 170850
rect 141210 170840 141290 170850
rect 141360 170840 141440 170850
rect 129640 170760 129650 170840
rect 129790 170760 129800 170840
rect 130060 170810 130120 170840
rect 130180 170810 130240 170840
rect 140740 170810 140800 170840
rect 141140 170760 141150 170840
rect 141290 170760 141300 170840
rect 141440 170760 141450 170840
rect 141745 170790 141755 170870
rect 142065 170790 142075 170870
rect 145265 170790 145275 170870
rect 145585 170790 145595 170870
rect 145905 170790 145915 170870
rect 146620 170860 146630 170940
rect 146940 170860 146950 170940
rect 146700 170780 146780 170790
rect 49180 170690 49210 170750
rect 49300 170690 49330 170750
rect 49420 170690 49450 170750
rect 49540 170690 49570 170750
rect 49660 170690 49690 170750
rect 49780 170690 49810 170750
rect 49900 170690 49930 170750
rect 50020 170690 50050 170750
rect 50140 170690 50170 170750
rect 50260 170690 50290 170750
rect 50380 170690 50410 170750
rect 50500 170690 50530 170750
rect 50620 170690 50650 170750
rect 50740 170690 50770 170750
rect 50860 170690 50890 170750
rect 50980 170690 51010 170750
rect 51100 170690 51130 170750
rect 51220 170690 51250 170750
rect 51340 170690 51370 170750
rect 51460 170690 51490 170750
rect 51580 170690 51610 170750
rect 51700 170690 51730 170750
rect 51820 170690 51850 170750
rect 51940 170690 51970 170750
rect 52060 170690 52090 170750
rect 52180 170690 52210 170750
rect 52300 170690 52330 170750
rect 52420 170690 52450 170750
rect 52540 170690 52570 170750
rect 52660 170690 52690 170750
rect 52780 170690 52810 170750
rect 52900 170690 52930 170750
rect 53020 170690 53050 170750
rect 53140 170690 53170 170750
rect 53260 170690 53290 170750
rect 53380 170690 53410 170750
rect 53500 170690 53530 170750
rect 53620 170690 53650 170750
rect 53740 170690 53770 170750
rect 53860 170690 53890 170750
rect 53980 170690 54010 170750
rect 54100 170690 54130 170750
rect 54220 170690 54250 170750
rect 54340 170690 54370 170750
rect 54460 170690 54490 170750
rect 54580 170690 54610 170750
rect 54700 170690 54730 170750
rect 54820 170690 54850 170750
rect 54940 170690 54970 170750
rect 55060 170690 55090 170750
rect 55180 170690 55210 170750
rect 55300 170690 55330 170750
rect 55420 170690 55450 170750
rect 55540 170690 55570 170750
rect 55660 170690 55690 170750
rect 55780 170690 55810 170750
rect 55900 170690 55930 170750
rect 56020 170690 56050 170750
rect 56140 170690 56170 170750
rect 56260 170690 56290 170750
rect 56380 170690 56410 170750
rect 56500 170690 56530 170750
rect 56620 170690 56650 170750
rect 56740 170690 56770 170750
rect 56860 170690 56890 170750
rect 56980 170690 57010 170750
rect 57100 170690 57130 170750
rect 57220 170690 57250 170750
rect 57340 170690 57370 170750
rect 57460 170690 57490 170750
rect 57580 170690 57610 170750
rect 57700 170690 57730 170750
rect 57820 170690 57850 170750
rect 57940 170690 57970 170750
rect 58060 170690 58090 170750
rect 58180 170690 58210 170750
rect 58300 170690 58330 170750
rect 58420 170690 58450 170750
rect 58540 170690 58570 170750
rect 58660 170690 58690 170750
rect 58780 170690 58810 170750
rect 58900 170690 58930 170750
rect 59020 170690 59050 170750
rect 59140 170690 59170 170750
rect 59260 170690 59290 170750
rect 59380 170690 59410 170750
rect 59500 170690 59530 170750
rect 59620 170690 59650 170750
rect 59740 170690 59770 170750
rect 60610 170709 60690 170719
rect 60930 170709 61010 170719
rect 61350 170709 61430 170719
rect 61670 170709 61750 170719
rect 48500 170660 48640 170670
rect 48710 170660 48790 170670
rect 60060 170660 60140 170670
rect 60210 170660 60290 170670
rect 60360 170660 60440 170670
rect 43060 170620 43140 170630
rect 43380 170620 43460 170630
rect 43140 170540 43150 170620
rect 43460 170540 43470 170620
rect 43905 170550 43985 170560
rect 44225 170550 44305 170560
rect 44545 170550 44625 170560
rect 44865 170550 44945 170560
rect 45185 170550 45265 170560
rect 45505 170550 45585 170560
rect 45825 170550 45905 170560
rect 46145 170550 46225 170560
rect 46465 170550 46545 170560
rect 46785 170550 46865 170560
rect 47105 170550 47185 170560
rect 47425 170550 47505 170560
rect 47745 170550 47825 170560
rect 48065 170550 48145 170560
rect 43985 170470 43995 170550
rect 44305 170470 44315 170550
rect 44625 170470 44635 170550
rect 44945 170470 44955 170550
rect 45265 170470 45275 170550
rect 45585 170470 45595 170550
rect 45905 170470 45915 170550
rect 46225 170470 46235 170550
rect 46545 170470 46555 170550
rect 46865 170470 46875 170550
rect 47185 170470 47195 170550
rect 47505 170470 47515 170550
rect 47825 170470 47835 170550
rect 48145 170470 48155 170550
rect 48500 170490 48605 170660
rect 48640 170580 48650 170660
rect 48790 170580 48800 170660
rect 60140 170580 60150 170660
rect 60290 170580 60300 170660
rect 60440 170580 60450 170660
rect 60690 170629 60700 170709
rect 61010 170629 61020 170709
rect 61430 170629 61440 170709
rect 61750 170629 61760 170709
rect 62680 170690 62710 170750
rect 73245 170690 73270 170750
rect 74110 170709 74190 170719
rect 74430 170709 74510 170719
rect 74850 170709 74930 170719
rect 75170 170709 75250 170719
rect 62060 170660 62140 170670
rect 62210 170660 62290 170670
rect 73560 170660 73640 170670
rect 73710 170660 73790 170670
rect 73860 170660 73940 170670
rect 62140 170580 62150 170660
rect 62290 170580 62300 170660
rect 73640 170580 73650 170660
rect 73790 170580 73800 170660
rect 73940 170580 73950 170660
rect 74190 170629 74200 170709
rect 74510 170629 74520 170709
rect 74930 170629 74940 170709
rect 75250 170629 75260 170709
rect 76180 170690 76210 170750
rect 86745 170690 86770 170750
rect 87610 170709 87690 170719
rect 87930 170709 88010 170719
rect 88350 170709 88430 170719
rect 88670 170709 88750 170719
rect 75560 170660 75640 170670
rect 75710 170660 75790 170670
rect 87060 170660 87140 170670
rect 87210 170660 87290 170670
rect 87360 170660 87440 170670
rect 75640 170580 75650 170660
rect 75790 170580 75800 170660
rect 87140 170580 87150 170660
rect 87290 170580 87300 170660
rect 87440 170580 87450 170660
rect 87690 170629 87700 170709
rect 88010 170629 88020 170709
rect 88430 170629 88440 170709
rect 88750 170629 88760 170709
rect 89680 170690 89710 170750
rect 100245 170690 100270 170750
rect 101110 170709 101190 170719
rect 101430 170709 101510 170719
rect 101850 170709 101930 170719
rect 102170 170709 102250 170719
rect 114610 170709 114690 170719
rect 114930 170709 115010 170719
rect 115350 170709 115430 170719
rect 115670 170709 115750 170719
rect 89060 170660 89140 170670
rect 89210 170660 89290 170670
rect 100560 170660 100640 170670
rect 100710 170660 100790 170670
rect 100860 170660 100940 170670
rect 89140 170580 89150 170660
rect 89290 170580 89300 170660
rect 100640 170580 100650 170660
rect 100790 170580 100800 170660
rect 100940 170580 100950 170660
rect 101190 170629 101200 170709
rect 101510 170629 101520 170709
rect 101930 170629 101940 170709
rect 102250 170629 102260 170709
rect 114690 170629 114700 170709
rect 115010 170629 115020 170709
rect 115430 170629 115440 170709
rect 115750 170629 115760 170709
rect 116680 170690 116710 170750
rect 127245 170690 127270 170750
rect 128110 170709 128190 170719
rect 128430 170709 128510 170719
rect 128850 170709 128930 170719
rect 129170 170709 129250 170719
rect 116060 170660 116140 170670
rect 116210 170660 116290 170670
rect 127560 170660 127640 170670
rect 127710 170660 127790 170670
rect 127860 170660 127940 170670
rect 116140 170580 116150 170660
rect 116290 170580 116300 170660
rect 127640 170580 127650 170660
rect 127790 170580 127800 170660
rect 127940 170580 127950 170660
rect 128190 170629 128200 170709
rect 128510 170629 128520 170709
rect 128930 170629 128940 170709
rect 129250 170629 129260 170709
rect 130180 170690 130210 170750
rect 140740 170690 140770 170750
rect 141825 170710 141905 170720
rect 142145 170710 142200 170720
rect 145345 170710 145425 170720
rect 145665 170710 145745 170720
rect 145985 170710 146065 170720
rect 129560 170660 129640 170670
rect 129710 170660 129790 170670
rect 141060 170660 141140 170670
rect 141210 170660 141290 170670
rect 141360 170660 141440 170670
rect 129640 170580 129650 170660
rect 129790 170580 129800 170660
rect 141140 170580 141150 170660
rect 141290 170580 141300 170660
rect 141440 170580 141450 170660
rect 141905 170630 141915 170710
rect 145425 170630 145435 170710
rect 145745 170630 145755 170710
rect 146065 170630 146075 170710
rect 146780 170700 146790 170780
rect 146540 170620 146620 170630
rect 146860 170620 146940 170630
rect 60770 170549 60850 170559
rect 61090 170549 61170 170559
rect 61510 170549 61590 170559
rect 61830 170549 61910 170559
rect 74270 170549 74350 170559
rect 74590 170549 74670 170559
rect 75010 170549 75090 170559
rect 75330 170549 75410 170559
rect 87770 170549 87850 170559
rect 88090 170549 88170 170559
rect 88510 170549 88590 170559
rect 88830 170549 88910 170559
rect 101270 170549 101350 170559
rect 101590 170549 101670 170559
rect 102010 170549 102090 170559
rect 102330 170549 102410 170559
rect 114770 170549 114850 170559
rect 115090 170549 115170 170559
rect 115510 170549 115590 170559
rect 115830 170549 115910 170559
rect 128270 170549 128350 170559
rect 128590 170549 128670 170559
rect 129010 170549 129090 170559
rect 129330 170549 129410 170559
rect 141665 170550 141745 170560
rect 141985 170550 142065 170560
rect 145200 170550 145265 170560
rect 145505 170550 145585 170560
rect 145825 170550 145905 170560
rect 48500 170480 48640 170490
rect 48710 170480 48790 170490
rect 60060 170480 60140 170490
rect 60210 170480 60290 170490
rect 60360 170480 60440 170490
rect 42950 170460 42980 170470
rect 43220 170460 43300 170470
rect 42980 170380 42990 170460
rect 43300 170380 43310 170460
rect 44065 170390 44145 170400
rect 44385 170390 44465 170400
rect 44705 170390 44785 170400
rect 45025 170390 45105 170400
rect 45345 170390 45425 170400
rect 45665 170390 45745 170400
rect 45985 170390 46065 170400
rect 46305 170390 46385 170400
rect 46625 170390 46705 170400
rect 46945 170390 47025 170400
rect 47265 170390 47345 170400
rect 47585 170390 47665 170400
rect 47905 170390 47985 170400
rect 48225 170390 48305 170400
rect 44145 170310 44155 170390
rect 44465 170310 44475 170390
rect 44785 170310 44795 170390
rect 45105 170310 45115 170390
rect 45425 170310 45435 170390
rect 45745 170310 45755 170390
rect 46065 170310 46075 170390
rect 46385 170310 46395 170390
rect 46705 170310 46715 170390
rect 47025 170310 47035 170390
rect 47345 170310 47355 170390
rect 47665 170310 47675 170390
rect 47985 170310 47995 170390
rect 48305 170310 48315 170390
rect 48500 170310 48605 170480
rect 48640 170400 48650 170480
rect 48790 170400 48800 170480
rect 60140 170400 60150 170480
rect 60290 170400 60300 170480
rect 60440 170400 60450 170480
rect 60850 170469 60860 170549
rect 61170 170469 61180 170549
rect 61590 170469 61600 170549
rect 61910 170469 61920 170549
rect 62060 170480 62140 170490
rect 62210 170480 62290 170490
rect 73560 170480 73640 170490
rect 73710 170480 73790 170490
rect 73860 170480 73940 170490
rect 62140 170400 62150 170480
rect 62290 170400 62300 170480
rect 73640 170400 73650 170480
rect 73790 170400 73800 170480
rect 73940 170400 73950 170480
rect 74350 170469 74360 170549
rect 74670 170469 74680 170549
rect 75090 170469 75100 170549
rect 75410 170469 75420 170549
rect 75560 170480 75640 170490
rect 75710 170480 75790 170490
rect 87060 170480 87140 170490
rect 87210 170480 87290 170490
rect 87360 170480 87440 170490
rect 75640 170400 75650 170480
rect 75790 170400 75800 170480
rect 87140 170400 87150 170480
rect 87290 170400 87300 170480
rect 87440 170400 87450 170480
rect 87850 170469 87860 170549
rect 88170 170469 88180 170549
rect 88590 170469 88600 170549
rect 88910 170469 88920 170549
rect 89060 170480 89140 170490
rect 89210 170480 89290 170490
rect 100560 170480 100640 170490
rect 100710 170480 100790 170490
rect 100860 170480 100940 170490
rect 89140 170400 89150 170480
rect 89290 170400 89300 170480
rect 100640 170400 100650 170480
rect 100790 170400 100800 170480
rect 100940 170400 100950 170480
rect 101350 170469 101360 170549
rect 101670 170469 101680 170549
rect 102090 170469 102100 170549
rect 102410 170469 102420 170549
rect 114850 170469 114860 170549
rect 115170 170469 115180 170549
rect 115590 170469 115600 170549
rect 115910 170469 115920 170549
rect 116060 170480 116140 170490
rect 116210 170480 116290 170490
rect 127560 170480 127640 170490
rect 127710 170480 127790 170490
rect 127860 170480 127940 170490
rect 116140 170400 116150 170480
rect 116290 170400 116300 170480
rect 127640 170400 127650 170480
rect 127790 170400 127800 170480
rect 127940 170400 127950 170480
rect 128350 170469 128360 170549
rect 128670 170469 128680 170549
rect 129090 170469 129100 170549
rect 129410 170469 129420 170549
rect 129560 170480 129640 170490
rect 129710 170480 129790 170490
rect 141060 170480 141140 170490
rect 141210 170480 141290 170490
rect 141360 170480 141440 170490
rect 129640 170400 129650 170480
rect 129790 170400 129800 170480
rect 141140 170400 141150 170480
rect 141290 170400 141300 170480
rect 141440 170400 141450 170480
rect 141745 170470 141755 170550
rect 142065 170470 142075 170550
rect 145265 170470 145275 170550
rect 145585 170470 145595 170550
rect 145905 170470 145915 170550
rect 146620 170540 146630 170620
rect 146940 170540 146950 170620
rect 146700 170460 146780 170470
rect 60610 170389 60690 170399
rect 60930 170389 61010 170399
rect 61350 170389 61430 170399
rect 61670 170389 61750 170399
rect 74110 170389 74190 170399
rect 74430 170389 74510 170399
rect 74850 170389 74930 170399
rect 75170 170389 75250 170399
rect 87610 170389 87690 170399
rect 87930 170389 88010 170399
rect 88350 170389 88430 170399
rect 88670 170389 88750 170399
rect 101110 170389 101190 170399
rect 101430 170389 101510 170399
rect 101850 170389 101930 170399
rect 102170 170389 102250 170399
rect 114610 170389 114690 170399
rect 114930 170389 115010 170399
rect 115350 170389 115430 170399
rect 115670 170389 115750 170399
rect 128110 170389 128190 170399
rect 128430 170389 128510 170399
rect 128850 170389 128930 170399
rect 129170 170389 129250 170399
rect 141825 170390 141905 170400
rect 142145 170390 142200 170400
rect 145345 170390 145425 170400
rect 145665 170390 145745 170400
rect 145985 170390 146065 170400
rect 43060 170300 43140 170310
rect 43380 170300 43460 170310
rect 48500 170300 48640 170310
rect 48710 170300 48790 170310
rect 60060 170300 60140 170310
rect 60210 170300 60290 170310
rect 60360 170300 60440 170310
rect 60690 170309 60700 170389
rect 61010 170309 61020 170389
rect 61430 170309 61440 170389
rect 61750 170309 61760 170389
rect 62060 170300 62140 170310
rect 62210 170300 62290 170310
rect 73560 170300 73640 170310
rect 73710 170300 73790 170310
rect 73860 170300 73940 170310
rect 74190 170309 74200 170389
rect 74510 170309 74520 170389
rect 74930 170309 74940 170389
rect 75250 170309 75260 170389
rect 75560 170300 75640 170310
rect 75710 170300 75790 170310
rect 87060 170300 87140 170310
rect 87210 170300 87290 170310
rect 87360 170300 87440 170310
rect 87690 170309 87700 170389
rect 88010 170309 88020 170389
rect 88430 170309 88440 170389
rect 88750 170309 88760 170389
rect 89060 170300 89140 170310
rect 89210 170300 89290 170310
rect 100560 170300 100640 170310
rect 100710 170300 100790 170310
rect 100860 170300 100940 170310
rect 101190 170309 101200 170389
rect 101510 170309 101520 170389
rect 101930 170309 101940 170389
rect 102250 170309 102260 170389
rect 114690 170309 114700 170389
rect 115010 170309 115020 170389
rect 115430 170309 115440 170389
rect 115750 170309 115760 170389
rect 116060 170300 116140 170310
rect 116210 170300 116290 170310
rect 127560 170300 127640 170310
rect 127710 170300 127790 170310
rect 127860 170300 127940 170310
rect 128190 170309 128200 170389
rect 128510 170309 128520 170389
rect 128930 170309 128940 170389
rect 129250 170309 129260 170389
rect 141905 170310 141915 170390
rect 145425 170310 145435 170390
rect 145745 170310 145755 170390
rect 146065 170310 146075 170390
rect 146780 170380 146790 170460
rect 129560 170300 129640 170310
rect 129710 170300 129790 170310
rect 141060 170300 141140 170310
rect 141210 170300 141290 170310
rect 141360 170300 141440 170310
rect 146540 170300 146620 170310
rect 146860 170300 146940 170310
rect 43140 170220 43150 170300
rect 43460 170220 43470 170300
rect 43905 170230 43985 170240
rect 44225 170230 44305 170240
rect 44545 170230 44625 170240
rect 44865 170230 44945 170240
rect 45185 170230 45265 170240
rect 45505 170230 45585 170240
rect 45825 170230 45905 170240
rect 46145 170230 46225 170240
rect 46465 170230 46545 170240
rect 46785 170230 46865 170240
rect 47105 170230 47185 170240
rect 47425 170230 47505 170240
rect 47745 170230 47825 170240
rect 48065 170230 48145 170240
rect 43985 170150 43995 170230
rect 44305 170150 44315 170230
rect 44625 170150 44635 170230
rect 44945 170150 44955 170230
rect 45265 170150 45275 170230
rect 45585 170150 45595 170230
rect 45905 170150 45915 170230
rect 46225 170150 46235 170230
rect 46545 170150 46555 170230
rect 46865 170150 46875 170230
rect 47185 170150 47195 170230
rect 47505 170150 47515 170230
rect 47825 170150 47835 170230
rect 48145 170150 48155 170230
rect 42950 170140 42980 170150
rect 43220 170140 43300 170150
rect 42980 170060 42990 170140
rect 43300 170060 43310 170140
rect 48500 170130 48605 170300
rect 48640 170220 48650 170300
rect 48790 170220 48800 170300
rect 60140 170220 60150 170300
rect 60290 170220 60300 170300
rect 60440 170220 60450 170300
rect 60770 170229 60850 170239
rect 61090 170229 61170 170239
rect 61510 170229 61590 170239
rect 61830 170229 61910 170239
rect 48500 170120 48640 170130
rect 48710 170120 48790 170130
rect 49270 170120 49350 170130
rect 49420 170120 49500 170130
rect 49570 170120 49650 170130
rect 44065 170070 44145 170080
rect 44385 170070 44465 170080
rect 44705 170070 44785 170080
rect 45025 170070 45105 170080
rect 45345 170070 45425 170080
rect 45665 170070 45745 170080
rect 45985 170070 46065 170080
rect 46305 170070 46385 170080
rect 46625 170070 46705 170080
rect 46945 170070 47025 170080
rect 47265 170070 47345 170080
rect 47585 170070 47665 170080
rect 47905 170070 47985 170080
rect 48225 170070 48305 170080
rect 44145 169990 44155 170070
rect 44465 169990 44475 170070
rect 44785 169990 44795 170070
rect 45105 169990 45115 170070
rect 45425 169990 45435 170070
rect 45745 169990 45755 170070
rect 46065 169990 46075 170070
rect 46385 169990 46395 170070
rect 46705 169990 46715 170070
rect 47025 169990 47035 170070
rect 47345 169990 47355 170070
rect 47665 169990 47675 170070
rect 47985 169990 47995 170070
rect 48305 169990 48315 170070
rect 43060 169980 43140 169990
rect 43380 169980 43460 169990
rect 43140 169900 43150 169980
rect 43460 169900 43470 169980
rect 48500 169950 48605 170120
rect 48640 170040 48650 170120
rect 48790 170040 48800 170120
rect 49350 170040 49360 170120
rect 49500 170040 49510 170120
rect 49650 170040 49660 170120
rect 48500 169940 48640 169950
rect 48710 169940 48790 169950
rect 49270 169940 49350 169950
rect 49420 169940 49500 169950
rect 49570 169940 49650 169950
rect 43905 169910 43985 169920
rect 44225 169910 44305 169920
rect 44545 169910 44625 169920
rect 44865 169910 44945 169920
rect 45185 169910 45265 169920
rect 45505 169910 45585 169920
rect 45825 169910 45905 169920
rect 46145 169910 46225 169920
rect 46465 169910 46545 169920
rect 46785 169910 46865 169920
rect 47105 169910 47185 169920
rect 47425 169910 47505 169920
rect 47745 169910 47825 169920
rect 48065 169910 48145 169920
rect 43985 169830 43995 169910
rect 44305 169830 44315 169910
rect 44625 169830 44635 169910
rect 44945 169830 44955 169910
rect 45265 169830 45275 169910
rect 45585 169830 45595 169910
rect 45905 169830 45915 169910
rect 46225 169830 46235 169910
rect 46545 169830 46555 169910
rect 46865 169830 46875 169910
rect 47185 169830 47195 169910
rect 47505 169830 47515 169910
rect 47825 169830 47835 169910
rect 48145 169830 48155 169910
rect 42950 169820 42980 169830
rect 43220 169820 43300 169830
rect 42980 169740 42990 169820
rect 43300 169740 43310 169820
rect 48500 169770 48605 169940
rect 48640 169860 48650 169940
rect 48790 169860 48800 169940
rect 49350 169860 49360 169940
rect 49500 169860 49510 169940
rect 49650 169860 49660 169940
rect 48500 169760 48640 169770
rect 48710 169760 48790 169770
rect 49270 169760 49350 169770
rect 49420 169760 49500 169770
rect 49570 169760 49650 169770
rect 44065 169750 44145 169760
rect 44385 169750 44465 169760
rect 44705 169750 44785 169760
rect 45025 169750 45105 169760
rect 45345 169750 45425 169760
rect 45665 169750 45745 169760
rect 45985 169750 46065 169760
rect 46305 169750 46385 169760
rect 46625 169750 46705 169760
rect 46945 169750 47025 169760
rect 47265 169750 47345 169760
rect 47585 169750 47665 169760
rect 47905 169750 47985 169760
rect 48225 169750 48305 169760
rect 44145 169670 44155 169750
rect 44465 169670 44475 169750
rect 44785 169670 44795 169750
rect 45105 169670 45115 169750
rect 45425 169670 45435 169750
rect 45745 169670 45755 169750
rect 46065 169670 46075 169750
rect 46385 169670 46395 169750
rect 46705 169670 46715 169750
rect 47025 169670 47035 169750
rect 47345 169670 47355 169750
rect 47665 169670 47675 169750
rect 47985 169670 47995 169750
rect 48305 169670 48315 169750
rect 43060 169660 43140 169670
rect 43380 169660 43460 169670
rect 43140 169580 43150 169660
rect 43460 169580 43470 169660
rect 43905 169590 43985 169600
rect 44225 169590 44305 169600
rect 44545 169590 44625 169600
rect 44865 169590 44945 169600
rect 45185 169590 45265 169600
rect 45505 169590 45585 169600
rect 45825 169590 45905 169600
rect 46145 169590 46225 169600
rect 46465 169590 46545 169600
rect 46785 169590 46865 169600
rect 47105 169590 47185 169600
rect 47425 169590 47505 169600
rect 47745 169590 47825 169600
rect 48065 169590 48145 169600
rect 48500 169590 48605 169760
rect 48640 169680 48650 169760
rect 48790 169680 48800 169760
rect 49350 169680 49360 169760
rect 49500 169680 49510 169760
rect 49650 169680 49660 169760
rect 43985 169510 43995 169590
rect 44305 169510 44315 169590
rect 44625 169510 44635 169590
rect 44945 169510 44955 169590
rect 45265 169510 45275 169590
rect 45585 169510 45595 169590
rect 45905 169510 45915 169590
rect 46225 169510 46235 169590
rect 46545 169510 46555 169590
rect 46865 169510 46875 169590
rect 47185 169510 47195 169590
rect 47505 169510 47515 169590
rect 47825 169510 47835 169590
rect 48145 169510 48155 169590
rect 48500 169580 48640 169590
rect 48710 169580 48790 169590
rect 49270 169580 49350 169590
rect 49420 169580 49500 169590
rect 49570 169580 49650 169590
rect 42950 169500 42980 169510
rect 43220 169500 43300 169510
rect 42980 169420 42990 169500
rect 43300 169420 43310 169500
rect 44065 169430 44145 169440
rect 44385 169430 44465 169440
rect 44705 169430 44785 169440
rect 45025 169430 45105 169440
rect 45345 169430 45425 169440
rect 45665 169430 45745 169440
rect 45985 169430 46065 169440
rect 46305 169430 46385 169440
rect 46625 169430 46705 169440
rect 46945 169430 47025 169440
rect 47265 169430 47345 169440
rect 47585 169430 47665 169440
rect 47905 169430 47985 169440
rect 48225 169430 48305 169440
rect 44145 169350 44155 169430
rect 44465 169350 44475 169430
rect 44785 169350 44795 169430
rect 45105 169350 45115 169430
rect 45425 169350 45435 169430
rect 45745 169350 45755 169430
rect 46065 169350 46075 169430
rect 46385 169350 46395 169430
rect 46705 169350 46715 169430
rect 47025 169350 47035 169430
rect 47345 169350 47355 169430
rect 47665 169350 47675 169430
rect 47985 169350 47995 169430
rect 48305 169350 48315 169430
rect 48500 169410 48605 169580
rect 48640 169500 48650 169580
rect 48790 169500 48800 169580
rect 49350 169500 49360 169580
rect 49500 169500 49510 169580
rect 49650 169500 49660 169580
rect 48500 169400 48640 169410
rect 48710 169400 48790 169410
rect 49270 169400 49350 169410
rect 49420 169400 49500 169410
rect 49570 169400 49650 169410
rect 43060 169340 43140 169350
rect 43380 169340 43460 169350
rect 43140 169260 43150 169340
rect 43460 169260 43470 169340
rect 43905 169270 43985 169280
rect 44225 169270 44305 169280
rect 44545 169270 44625 169280
rect 44865 169270 44945 169280
rect 45185 169270 45265 169280
rect 45505 169270 45585 169280
rect 45825 169270 45905 169280
rect 46145 169270 46225 169280
rect 46465 169270 46545 169280
rect 46785 169270 46865 169280
rect 47105 169270 47185 169280
rect 47425 169270 47505 169280
rect 47745 169270 47825 169280
rect 48065 169270 48145 169280
rect 43985 169190 43995 169270
rect 44305 169190 44315 169270
rect 44625 169190 44635 169270
rect 44945 169190 44955 169270
rect 45265 169190 45275 169270
rect 45585 169190 45595 169270
rect 45905 169190 45915 169270
rect 46225 169190 46235 169270
rect 46545 169190 46555 169270
rect 46865 169190 46875 169270
rect 47185 169190 47195 169270
rect 47505 169190 47515 169270
rect 47825 169190 47835 169270
rect 48145 169190 48155 169270
rect 48500 169230 48605 169400
rect 48640 169320 48650 169400
rect 48790 169320 48800 169400
rect 49350 169320 49360 169400
rect 49500 169320 49510 169400
rect 49650 169320 49660 169400
rect 48500 169220 48640 169230
rect 48710 169220 48790 169230
rect 49270 169220 49350 169230
rect 49420 169220 49500 169230
rect 49570 169220 49650 169230
rect 42950 169180 42980 169190
rect 43220 169180 43300 169190
rect 42980 169100 42990 169180
rect 43300 169100 43310 169180
rect 44065 169110 44145 169120
rect 44385 169110 44465 169120
rect 44705 169110 44785 169120
rect 45025 169110 45105 169120
rect 45345 169110 45425 169120
rect 45665 169110 45745 169120
rect 45985 169110 46065 169120
rect 46305 169110 46385 169120
rect 46625 169110 46705 169120
rect 46945 169110 47025 169120
rect 47265 169110 47345 169120
rect 47585 169110 47665 169120
rect 47905 169110 47985 169120
rect 48225 169110 48305 169120
rect 44145 169030 44155 169110
rect 44465 169030 44475 169110
rect 44785 169030 44795 169110
rect 45105 169030 45115 169110
rect 45425 169030 45435 169110
rect 45745 169030 45755 169110
rect 46065 169030 46075 169110
rect 46385 169030 46395 169110
rect 46705 169030 46715 169110
rect 47025 169030 47035 169110
rect 47345 169030 47355 169110
rect 47665 169030 47675 169110
rect 47985 169030 47995 169110
rect 48305 169030 48315 169110
rect 48500 169050 48605 169220
rect 48640 169140 48650 169220
rect 48790 169140 48800 169220
rect 49350 169140 49360 169220
rect 49500 169140 49510 169220
rect 49650 169140 49660 169220
rect 48500 169040 48640 169050
rect 48710 169040 48790 169050
rect 49270 169040 49350 169050
rect 49420 169040 49500 169050
rect 49570 169040 49650 169050
rect 43060 169020 43140 169030
rect 43380 169020 43460 169030
rect 43140 168940 43150 169020
rect 43460 168940 43470 169020
rect 43905 168950 43985 168960
rect 44225 168950 44305 168960
rect 44545 168950 44625 168960
rect 44865 168950 44945 168960
rect 45185 168950 45265 168960
rect 45505 168950 45585 168960
rect 45825 168950 45905 168960
rect 46145 168950 46225 168960
rect 46465 168950 46545 168960
rect 46785 168950 46865 168960
rect 47105 168950 47185 168960
rect 47425 168950 47505 168960
rect 47745 168950 47825 168960
rect 48065 168950 48145 168960
rect 43985 168870 43995 168950
rect 44305 168870 44315 168950
rect 44625 168870 44635 168950
rect 44945 168870 44955 168950
rect 45265 168870 45275 168950
rect 45585 168870 45595 168950
rect 45905 168870 45915 168950
rect 46225 168870 46235 168950
rect 46545 168870 46555 168950
rect 46865 168870 46875 168950
rect 47185 168870 47195 168950
rect 47505 168870 47515 168950
rect 47825 168870 47835 168950
rect 48145 168870 48155 168950
rect 48500 168870 48605 169040
rect 48640 168960 48650 169040
rect 48790 168960 48800 169040
rect 49350 168960 49360 169040
rect 49500 168960 49510 169040
rect 49650 168960 49660 169040
rect 42950 168860 42980 168870
rect 43220 168860 43300 168870
rect 48500 168860 48640 168870
rect 48710 168860 48790 168870
rect 49270 168860 49350 168870
rect 49420 168860 49500 168870
rect 49570 168860 49650 168870
rect 42980 168780 42990 168860
rect 43300 168780 43310 168860
rect 44065 168790 44145 168800
rect 44385 168790 44465 168800
rect 44705 168790 44785 168800
rect 45025 168790 45105 168800
rect 45345 168790 45425 168800
rect 45665 168790 45745 168800
rect 45985 168790 46065 168800
rect 46305 168790 46385 168800
rect 46625 168790 46705 168800
rect 46945 168790 47025 168800
rect 47265 168790 47345 168800
rect 47585 168790 47665 168800
rect 47905 168790 47985 168800
rect 48225 168790 48305 168800
rect 44145 168710 44155 168790
rect 44465 168710 44475 168790
rect 44785 168710 44795 168790
rect 45105 168710 45115 168790
rect 45425 168710 45435 168790
rect 45745 168710 45755 168790
rect 46065 168710 46075 168790
rect 46385 168710 46395 168790
rect 46705 168710 46715 168790
rect 47025 168710 47035 168790
rect 47345 168710 47355 168790
rect 47665 168710 47675 168790
rect 47985 168710 47995 168790
rect 48305 168710 48315 168790
rect 43060 168700 43140 168710
rect 43380 168700 43460 168710
rect 43140 168620 43150 168700
rect 43460 168620 43470 168700
rect 48500 168690 48605 168860
rect 48640 168780 48650 168860
rect 48790 168780 48800 168860
rect 49350 168780 49360 168860
rect 49500 168780 49510 168860
rect 49650 168780 49660 168860
rect 48500 168680 48640 168690
rect 48710 168680 48790 168690
rect 49270 168680 49350 168690
rect 49420 168680 49500 168690
rect 49570 168680 49650 168690
rect 43905 168630 43985 168640
rect 44225 168630 44305 168640
rect 44545 168630 44625 168640
rect 44865 168630 44945 168640
rect 45185 168630 45265 168640
rect 45505 168630 45585 168640
rect 45825 168630 45905 168640
rect 46145 168630 46225 168640
rect 46465 168630 46545 168640
rect 46785 168630 46865 168640
rect 47105 168630 47185 168640
rect 47425 168630 47505 168640
rect 47745 168630 47825 168640
rect 48065 168630 48145 168640
rect 43985 168550 43995 168630
rect 44305 168550 44315 168630
rect 44625 168550 44635 168630
rect 44945 168550 44955 168630
rect 45265 168550 45275 168630
rect 45585 168550 45595 168630
rect 45905 168550 45915 168630
rect 46225 168550 46235 168630
rect 46545 168550 46555 168630
rect 46865 168550 46875 168630
rect 47185 168550 47195 168630
rect 47505 168550 47515 168630
rect 47825 168550 47835 168630
rect 48145 168550 48155 168630
rect 42950 168540 42980 168550
rect 43220 168540 43300 168550
rect 42980 168460 42990 168540
rect 43300 168460 43310 168540
rect 48500 168510 48605 168680
rect 48640 168600 48650 168680
rect 48790 168600 48800 168680
rect 49350 168600 49360 168680
rect 49500 168600 49510 168680
rect 49650 168600 49660 168680
rect 48500 168500 48640 168510
rect 48710 168500 48790 168510
rect 49270 168500 49350 168510
rect 49420 168500 49500 168510
rect 49570 168500 49650 168510
rect 44065 168470 44145 168480
rect 44385 168470 44465 168480
rect 44705 168470 44785 168480
rect 45025 168470 45105 168480
rect 45345 168470 45425 168480
rect 45665 168470 45745 168480
rect 45985 168470 46065 168480
rect 46305 168470 46385 168480
rect 46625 168470 46705 168480
rect 46945 168470 47025 168480
rect 47265 168470 47345 168480
rect 47585 168470 47665 168480
rect 47905 168470 47985 168480
rect 48225 168470 48305 168480
rect 44145 168390 44155 168470
rect 44465 168390 44475 168470
rect 44785 168390 44795 168470
rect 45105 168390 45115 168470
rect 45425 168390 45435 168470
rect 45745 168390 45755 168470
rect 46065 168390 46075 168470
rect 46385 168390 46395 168470
rect 46705 168390 46715 168470
rect 47025 168390 47035 168470
rect 47345 168390 47355 168470
rect 47665 168390 47675 168470
rect 47985 168390 47995 168470
rect 48305 168390 48315 168470
rect 43060 168380 43140 168390
rect 43380 168380 43460 168390
rect 43140 168300 43150 168380
rect 43460 168300 43470 168380
rect 48500 168330 48605 168500
rect 48640 168420 48650 168500
rect 48790 168420 48800 168500
rect 49350 168420 49360 168500
rect 49500 168420 49510 168500
rect 49650 168420 49660 168500
rect 48500 168320 48640 168330
rect 48710 168320 48790 168330
rect 49270 168320 49350 168330
rect 49420 168320 49500 168330
rect 49570 168320 49650 168330
rect 43905 168310 43985 168320
rect 44225 168310 44305 168320
rect 44545 168310 44625 168320
rect 44865 168310 44945 168320
rect 45185 168310 45265 168320
rect 45505 168310 45585 168320
rect 45825 168310 45905 168320
rect 46145 168310 46225 168320
rect 46465 168310 46545 168320
rect 46785 168310 46865 168320
rect 47105 168310 47185 168320
rect 47425 168310 47505 168320
rect 47745 168310 47825 168320
rect 48065 168310 48145 168320
rect 43985 168230 43995 168310
rect 44305 168230 44315 168310
rect 44625 168230 44635 168310
rect 44945 168230 44955 168310
rect 45265 168230 45275 168310
rect 45585 168230 45595 168310
rect 45905 168230 45915 168310
rect 46225 168230 46235 168310
rect 46545 168230 46555 168310
rect 46865 168230 46875 168310
rect 47185 168230 47195 168310
rect 47505 168230 47515 168310
rect 47825 168230 47835 168310
rect 48145 168230 48155 168310
rect 42950 168220 42980 168230
rect 43220 168220 43300 168230
rect 42980 168140 42990 168220
rect 43300 168140 43310 168220
rect 44065 168150 44145 168160
rect 44385 168150 44465 168160
rect 44705 168150 44785 168160
rect 45025 168150 45105 168160
rect 45345 168150 45425 168160
rect 45665 168150 45745 168160
rect 45985 168150 46065 168160
rect 46305 168150 46385 168160
rect 46625 168150 46705 168160
rect 46945 168150 47025 168160
rect 47265 168150 47345 168160
rect 47585 168150 47665 168160
rect 47905 168150 47985 168160
rect 48225 168150 48305 168160
rect 48500 168150 48605 168320
rect 48640 168240 48650 168320
rect 48790 168240 48800 168320
rect 49350 168240 49360 168320
rect 49500 168240 49510 168320
rect 49650 168240 49660 168320
rect 44145 168070 44155 168150
rect 44465 168070 44475 168150
rect 44785 168070 44795 168150
rect 45105 168070 45115 168150
rect 45425 168070 45435 168150
rect 45745 168070 45755 168150
rect 46065 168070 46075 168150
rect 46385 168070 46395 168150
rect 46705 168070 46715 168150
rect 47025 168070 47035 168150
rect 47345 168070 47355 168150
rect 47665 168070 47675 168150
rect 47985 168070 47995 168150
rect 48305 168070 48315 168150
rect 48500 168140 48640 168150
rect 48710 168140 48790 168150
rect 49270 168140 49350 168150
rect 49420 168140 49500 168150
rect 49570 168140 49650 168150
rect 43060 168060 43140 168070
rect 43380 168060 43460 168070
rect 43140 167980 43150 168060
rect 43460 167980 43470 168060
rect 43905 167990 43985 168000
rect 44225 167990 44305 168000
rect 44545 167990 44625 168000
rect 44865 167990 44945 168000
rect 45185 167990 45265 168000
rect 45505 167990 45585 168000
rect 45825 167990 45905 168000
rect 46145 167990 46225 168000
rect 46465 167990 46545 168000
rect 46785 167990 46865 168000
rect 47105 167990 47185 168000
rect 47425 167990 47505 168000
rect 47745 167990 47825 168000
rect 48065 167990 48145 168000
rect 43985 167910 43995 167990
rect 44305 167910 44315 167990
rect 44625 167910 44635 167990
rect 44945 167910 44955 167990
rect 45265 167910 45275 167990
rect 45585 167910 45595 167990
rect 45905 167910 45915 167990
rect 46225 167910 46235 167990
rect 46545 167910 46555 167990
rect 46865 167910 46875 167990
rect 47185 167910 47195 167990
rect 47505 167910 47515 167990
rect 47825 167910 47835 167990
rect 48145 167910 48155 167990
rect 48500 167970 48605 168140
rect 48640 168060 48650 168140
rect 48790 168060 48800 168140
rect 49350 168060 49360 168140
rect 49500 168060 49510 168140
rect 49650 168060 49660 168140
rect 48500 167960 48640 167970
rect 48710 167960 48790 167970
rect 49270 167960 49350 167970
rect 49420 167960 49500 167970
rect 49570 167960 49650 167970
rect 42950 167900 42980 167910
rect 43220 167900 43300 167910
rect 42980 167820 42990 167900
rect 43300 167820 43310 167900
rect 44065 167830 44145 167840
rect 44385 167830 44465 167840
rect 44705 167830 44785 167840
rect 45025 167830 45105 167840
rect 45345 167830 45425 167840
rect 45665 167830 45745 167840
rect 45985 167830 46065 167840
rect 46305 167830 46385 167840
rect 46625 167830 46705 167840
rect 46945 167830 47025 167840
rect 47265 167830 47345 167840
rect 47585 167830 47665 167840
rect 47905 167830 47985 167840
rect 48225 167830 48305 167840
rect 44145 167750 44155 167830
rect 44465 167750 44475 167830
rect 44785 167750 44795 167830
rect 45105 167750 45115 167830
rect 45425 167750 45435 167830
rect 45745 167750 45755 167830
rect 46065 167750 46075 167830
rect 46385 167750 46395 167830
rect 46705 167750 46715 167830
rect 47025 167750 47035 167830
rect 47345 167750 47355 167830
rect 47665 167750 47675 167830
rect 47985 167750 47995 167830
rect 48305 167750 48315 167830
rect 48500 167790 48605 167960
rect 48640 167880 48650 167960
rect 48790 167880 48800 167960
rect 49350 167880 49360 167960
rect 49500 167880 49510 167960
rect 49650 167880 49660 167960
rect 48500 167780 48640 167790
rect 48710 167780 48790 167790
rect 49270 167780 49350 167790
rect 49420 167780 49500 167790
rect 49570 167780 49650 167790
rect 43060 167740 43140 167750
rect 43380 167740 43460 167750
rect 43140 167660 43150 167740
rect 43460 167660 43470 167740
rect 43905 167670 43985 167680
rect 44225 167670 44305 167680
rect 44545 167670 44625 167680
rect 44865 167670 44945 167680
rect 45185 167670 45265 167680
rect 45505 167670 45585 167680
rect 45825 167670 45905 167680
rect 46145 167670 46225 167680
rect 46465 167670 46545 167680
rect 46785 167670 46865 167680
rect 47105 167670 47185 167680
rect 47425 167670 47505 167680
rect 47745 167670 47825 167680
rect 48065 167670 48145 167680
rect 43985 167590 43995 167670
rect 44305 167590 44315 167670
rect 44625 167590 44635 167670
rect 44945 167590 44955 167670
rect 45265 167590 45275 167670
rect 45585 167590 45595 167670
rect 45905 167590 45915 167670
rect 46225 167590 46235 167670
rect 46545 167590 46555 167670
rect 46865 167590 46875 167670
rect 47185 167590 47195 167670
rect 47505 167590 47515 167670
rect 47825 167590 47835 167670
rect 48145 167590 48155 167670
rect 48500 167610 48605 167780
rect 48640 167700 48650 167780
rect 48790 167700 48800 167780
rect 49350 167700 49360 167780
rect 49500 167700 49510 167780
rect 49650 167700 49660 167780
rect 48500 167600 48640 167610
rect 48710 167600 48790 167610
rect 49270 167600 49350 167610
rect 49420 167600 49500 167610
rect 49570 167600 49650 167610
rect 42950 167580 42980 167590
rect 43220 167580 43300 167590
rect 42980 167500 42990 167580
rect 43300 167500 43310 167580
rect 44065 167510 44145 167520
rect 44385 167510 44465 167520
rect 44705 167510 44785 167520
rect 45025 167510 45105 167520
rect 45345 167510 45425 167520
rect 45665 167510 45745 167520
rect 45985 167510 46065 167520
rect 46305 167510 46385 167520
rect 46625 167510 46705 167520
rect 46945 167510 47025 167520
rect 47265 167510 47345 167520
rect 47585 167510 47665 167520
rect 47905 167510 47985 167520
rect 48225 167510 48305 167520
rect 44145 167430 44155 167510
rect 44465 167430 44475 167510
rect 44785 167430 44795 167510
rect 45105 167430 45115 167510
rect 45425 167430 45435 167510
rect 45745 167430 45755 167510
rect 46065 167430 46075 167510
rect 46385 167430 46395 167510
rect 46705 167430 46715 167510
rect 47025 167430 47035 167510
rect 47345 167430 47355 167510
rect 47665 167430 47675 167510
rect 47985 167430 47995 167510
rect 48305 167430 48315 167510
rect 48500 167430 48605 167600
rect 48640 167520 48650 167600
rect 48790 167520 48800 167600
rect 49350 167520 49360 167600
rect 49500 167520 49510 167600
rect 49650 167520 49660 167600
rect 43060 167420 43140 167430
rect 43380 167420 43460 167430
rect 48500 167420 48640 167430
rect 48710 167420 48790 167430
rect 49270 167420 49350 167430
rect 49420 167420 49500 167430
rect 49570 167420 49650 167430
rect 43140 167340 43150 167420
rect 43460 167340 43470 167420
rect 43905 167350 43985 167360
rect 44225 167350 44305 167360
rect 44545 167350 44625 167360
rect 44865 167350 44945 167360
rect 45185 167350 45265 167360
rect 45505 167350 45585 167360
rect 45825 167350 45905 167360
rect 46145 167350 46225 167360
rect 46465 167350 46545 167360
rect 46785 167350 46865 167360
rect 47105 167350 47185 167360
rect 47425 167350 47505 167360
rect 47745 167350 47825 167360
rect 48065 167350 48145 167360
rect 43985 167270 43995 167350
rect 44305 167270 44315 167350
rect 44625 167270 44635 167350
rect 44945 167270 44955 167350
rect 45265 167270 45275 167350
rect 45585 167270 45595 167350
rect 45905 167270 45915 167350
rect 46225 167270 46235 167350
rect 46545 167270 46555 167350
rect 46865 167270 46875 167350
rect 47185 167270 47195 167350
rect 47505 167270 47515 167350
rect 47825 167270 47835 167350
rect 48145 167270 48155 167350
rect 42950 167260 42980 167270
rect 43220 167260 43300 167270
rect 42980 167180 42990 167260
rect 43300 167180 43310 167260
rect 48500 167250 48605 167420
rect 48640 167340 48650 167420
rect 48790 167340 48800 167420
rect 49350 167340 49360 167420
rect 49500 167340 49510 167420
rect 49650 167340 49660 167420
rect 48500 167240 48640 167250
rect 48710 167240 48790 167250
rect 49270 167240 49350 167250
rect 49420 167240 49500 167250
rect 49570 167240 49650 167250
rect 44065 167190 44145 167200
rect 44385 167190 44465 167200
rect 44705 167190 44785 167200
rect 45025 167190 45105 167200
rect 45345 167190 45425 167200
rect 45665 167190 45745 167200
rect 45985 167190 46065 167200
rect 46305 167190 46385 167200
rect 46625 167190 46705 167200
rect 46945 167190 47025 167200
rect 47265 167190 47345 167200
rect 47585 167190 47665 167200
rect 47905 167190 47985 167200
rect 48225 167190 48305 167200
rect 44145 167110 44155 167190
rect 44465 167110 44475 167190
rect 44785 167110 44795 167190
rect 45105 167110 45115 167190
rect 45425 167110 45435 167190
rect 45745 167110 45755 167190
rect 46065 167110 46075 167190
rect 46385 167110 46395 167190
rect 46705 167110 46715 167190
rect 47025 167110 47035 167190
rect 47345 167110 47355 167190
rect 47665 167110 47675 167190
rect 47985 167110 47995 167190
rect 48305 167110 48315 167190
rect 43060 167100 43140 167110
rect 43380 167100 43460 167110
rect 43140 167020 43150 167100
rect 43460 167020 43470 167100
rect 48500 167070 48605 167240
rect 48640 167160 48650 167240
rect 48790 167160 48800 167240
rect 49350 167160 49360 167240
rect 49500 167160 49510 167240
rect 49650 167160 49660 167240
rect 48500 167060 48640 167070
rect 48710 167060 48790 167070
rect 49270 167060 49350 167070
rect 49420 167060 49500 167070
rect 49570 167060 49650 167070
rect 43905 167030 43985 167040
rect 44225 167030 44305 167040
rect 44545 167030 44625 167040
rect 44865 167030 44945 167040
rect 45185 167030 45265 167040
rect 45505 167030 45585 167040
rect 45825 167030 45905 167040
rect 46145 167030 46225 167040
rect 46465 167030 46545 167040
rect 46785 167030 46865 167040
rect 47105 167030 47185 167040
rect 47425 167030 47505 167040
rect 47745 167030 47825 167040
rect 48065 167030 48145 167040
rect 43985 166950 43995 167030
rect 44305 166950 44315 167030
rect 44625 166950 44635 167030
rect 44945 166950 44955 167030
rect 45265 166950 45275 167030
rect 45585 166950 45595 167030
rect 45905 166950 45915 167030
rect 46225 166950 46235 167030
rect 46545 166950 46555 167030
rect 46865 166950 46875 167030
rect 47185 166950 47195 167030
rect 47505 166950 47515 167030
rect 47825 166950 47835 167030
rect 48145 166950 48155 167030
rect 42950 166940 42980 166950
rect 43220 166940 43300 166950
rect 42980 166860 42990 166940
rect 43300 166860 43310 166940
rect 48500 166890 48605 167060
rect 48640 166980 48650 167060
rect 48790 166980 48800 167060
rect 49350 166980 49360 167060
rect 49500 166980 49510 167060
rect 49650 166980 49660 167060
rect 48500 166880 48640 166890
rect 48710 166880 48790 166890
rect 49270 166880 49350 166890
rect 49420 166880 49500 166890
rect 49570 166880 49650 166890
rect 44065 166870 44145 166880
rect 44385 166870 44465 166880
rect 44705 166870 44785 166880
rect 45025 166870 45105 166880
rect 45345 166870 45425 166880
rect 45665 166870 45745 166880
rect 45985 166870 46065 166880
rect 46305 166870 46385 166880
rect 46625 166870 46705 166880
rect 46945 166870 47025 166880
rect 47265 166870 47345 166880
rect 47585 166870 47665 166880
rect 47905 166870 47985 166880
rect 48225 166870 48305 166880
rect 44145 166790 44155 166870
rect 44465 166790 44475 166870
rect 44785 166790 44795 166870
rect 45105 166790 45115 166870
rect 45425 166790 45435 166870
rect 45745 166790 45755 166870
rect 46065 166790 46075 166870
rect 46385 166790 46395 166870
rect 46705 166790 46715 166870
rect 47025 166790 47035 166870
rect 47345 166790 47355 166870
rect 47665 166790 47675 166870
rect 47985 166790 47995 166870
rect 48305 166790 48315 166870
rect 43060 166780 43140 166790
rect 43380 166780 43460 166790
rect 43140 166700 43150 166780
rect 43460 166700 43470 166780
rect 43905 166710 43985 166720
rect 44225 166710 44305 166720
rect 44545 166710 44625 166720
rect 44865 166710 44945 166720
rect 45185 166710 45265 166720
rect 45505 166710 45585 166720
rect 45825 166710 45905 166720
rect 46145 166710 46225 166720
rect 46465 166710 46545 166720
rect 46785 166710 46865 166720
rect 47105 166710 47185 166720
rect 47425 166710 47505 166720
rect 47745 166710 47825 166720
rect 48065 166710 48145 166720
rect 48500 166710 48605 166880
rect 48640 166800 48650 166880
rect 48790 166800 48800 166880
rect 49350 166800 49360 166880
rect 49500 166800 49510 166880
rect 49650 166800 49660 166880
rect 43985 166630 43995 166710
rect 44305 166630 44315 166710
rect 44625 166630 44635 166710
rect 44945 166630 44955 166710
rect 45265 166630 45275 166710
rect 45585 166630 45595 166710
rect 45905 166630 45915 166710
rect 46225 166630 46235 166710
rect 46545 166630 46555 166710
rect 46865 166630 46875 166710
rect 47185 166630 47195 166710
rect 47505 166630 47515 166710
rect 47825 166630 47835 166710
rect 48145 166630 48155 166710
rect 48500 166700 48640 166710
rect 48710 166700 48790 166710
rect 49270 166700 49350 166710
rect 49420 166700 49500 166710
rect 49570 166700 49650 166710
rect 42950 166620 42980 166630
rect 43220 166620 43300 166630
rect 42980 166540 42990 166620
rect 43300 166540 43310 166620
rect 44065 166550 44145 166560
rect 44385 166550 44465 166560
rect 44705 166550 44785 166560
rect 45025 166550 45105 166560
rect 45345 166550 45425 166560
rect 45665 166550 45745 166560
rect 45985 166550 46065 166560
rect 46305 166550 46385 166560
rect 46625 166550 46705 166560
rect 46945 166550 47025 166560
rect 47265 166550 47345 166560
rect 47585 166550 47665 166560
rect 47905 166550 47985 166560
rect 48225 166550 48305 166560
rect 44145 166470 44155 166550
rect 44465 166470 44475 166550
rect 44785 166470 44795 166550
rect 45105 166470 45115 166550
rect 45425 166470 45435 166550
rect 45745 166470 45755 166550
rect 46065 166470 46075 166550
rect 46385 166470 46395 166550
rect 46705 166470 46715 166550
rect 47025 166470 47035 166550
rect 47345 166470 47355 166550
rect 47665 166470 47675 166550
rect 47985 166470 47995 166550
rect 48305 166470 48315 166550
rect 48500 166530 48605 166700
rect 48640 166620 48650 166700
rect 48790 166620 48800 166700
rect 49350 166620 49360 166700
rect 49500 166620 49510 166700
rect 49650 166620 49660 166700
rect 48500 166520 48640 166530
rect 48710 166520 48790 166530
rect 49270 166520 49350 166530
rect 49420 166520 49500 166530
rect 49570 166520 49650 166530
rect 43060 166460 43140 166470
rect 43380 166460 43460 166470
rect 43140 166380 43150 166460
rect 43460 166380 43470 166460
rect 43905 166390 43985 166400
rect 44225 166390 44305 166400
rect 44545 166390 44625 166400
rect 44865 166390 44945 166400
rect 45185 166390 45265 166400
rect 45505 166390 45585 166400
rect 45825 166390 45905 166400
rect 46145 166390 46225 166400
rect 46465 166390 46545 166400
rect 46785 166390 46865 166400
rect 47105 166390 47185 166400
rect 47425 166390 47505 166400
rect 47745 166390 47825 166400
rect 48065 166390 48145 166400
rect 43985 166310 43995 166390
rect 44305 166310 44315 166390
rect 44625 166310 44635 166390
rect 44945 166310 44955 166390
rect 45265 166310 45275 166390
rect 45585 166310 45595 166390
rect 45905 166310 45915 166390
rect 46225 166310 46235 166390
rect 46545 166310 46555 166390
rect 46865 166310 46875 166390
rect 47185 166310 47195 166390
rect 47505 166310 47515 166390
rect 47825 166310 47835 166390
rect 48145 166310 48155 166390
rect 48500 166350 48605 166520
rect 48640 166440 48650 166520
rect 48790 166440 48800 166520
rect 49350 166440 49360 166520
rect 49500 166440 49510 166520
rect 49650 166440 49660 166520
rect 48500 166340 48640 166350
rect 48710 166340 48790 166350
rect 49270 166340 49350 166350
rect 49420 166340 49500 166350
rect 49570 166340 49650 166350
rect 42950 166300 42980 166310
rect 43220 166300 43300 166310
rect 42980 166220 42990 166300
rect 43300 166220 43310 166300
rect 44065 166230 44145 166240
rect 44385 166230 44465 166240
rect 44705 166230 44785 166240
rect 45025 166230 45105 166240
rect 45345 166230 45425 166240
rect 45665 166230 45745 166240
rect 45985 166230 46065 166240
rect 46305 166230 46385 166240
rect 46625 166230 46705 166240
rect 46945 166230 47025 166240
rect 47265 166230 47345 166240
rect 47585 166230 47665 166240
rect 47905 166230 47985 166240
rect 48225 166230 48305 166240
rect 44145 166150 44155 166230
rect 44465 166150 44475 166230
rect 44785 166150 44795 166230
rect 45105 166150 45115 166230
rect 45425 166150 45435 166230
rect 45745 166150 45755 166230
rect 46065 166150 46075 166230
rect 46385 166150 46395 166230
rect 46705 166150 46715 166230
rect 47025 166150 47035 166230
rect 47345 166150 47355 166230
rect 47665 166150 47675 166230
rect 47985 166150 47995 166230
rect 48305 166150 48315 166230
rect 48500 166170 48605 166340
rect 48640 166260 48650 166340
rect 48790 166260 48800 166340
rect 49350 166260 49360 166340
rect 49500 166260 49510 166340
rect 49650 166260 49660 166340
rect 48500 166160 48640 166170
rect 48710 166160 48790 166170
rect 49270 166160 49350 166170
rect 49420 166160 49500 166170
rect 49570 166160 49650 166170
rect 43060 166140 43140 166150
rect 43380 166140 43460 166150
rect 43140 166060 43150 166140
rect 43460 166060 43470 166140
rect 43905 166070 43985 166080
rect 44225 166070 44305 166080
rect 44545 166070 44625 166080
rect 44865 166070 44945 166080
rect 45185 166070 45265 166080
rect 45505 166070 45585 166080
rect 45825 166070 45905 166080
rect 46145 166070 46225 166080
rect 46465 166070 46545 166080
rect 46785 166070 46865 166080
rect 47105 166070 47185 166080
rect 47425 166070 47505 166080
rect 47745 166070 47825 166080
rect 48065 166070 48145 166080
rect 43985 165990 43995 166070
rect 44305 165990 44315 166070
rect 44625 165990 44635 166070
rect 44945 165990 44955 166070
rect 45265 165990 45275 166070
rect 45585 165990 45595 166070
rect 45905 165990 45915 166070
rect 46225 165990 46235 166070
rect 46545 165990 46555 166070
rect 46865 165990 46875 166070
rect 47185 165990 47195 166070
rect 47505 165990 47515 166070
rect 47825 165990 47835 166070
rect 48145 165990 48155 166070
rect 48500 165990 48605 166160
rect 48640 166080 48650 166160
rect 48790 166080 48800 166160
rect 49350 166080 49360 166160
rect 49500 166080 49510 166160
rect 49650 166080 49660 166160
rect 42950 165980 42980 165990
rect 43220 165980 43300 165990
rect 48500 165980 48640 165990
rect 48710 165980 48790 165990
rect 49270 165980 49350 165990
rect 49420 165980 49500 165990
rect 49570 165980 49650 165990
rect 42980 165900 42990 165980
rect 43300 165900 43310 165980
rect 44065 165910 44145 165920
rect 44385 165910 44465 165920
rect 44705 165910 44785 165920
rect 45025 165910 45105 165920
rect 45345 165910 45425 165920
rect 45665 165910 45745 165920
rect 45985 165910 46065 165920
rect 46305 165910 46385 165920
rect 46625 165910 46705 165920
rect 46945 165910 47025 165920
rect 47265 165910 47345 165920
rect 47585 165910 47665 165920
rect 47905 165910 47985 165920
rect 48225 165910 48305 165920
rect 44145 165830 44155 165910
rect 44465 165830 44475 165910
rect 44785 165830 44795 165910
rect 45105 165830 45115 165910
rect 45425 165830 45435 165910
rect 45745 165830 45755 165910
rect 46065 165830 46075 165910
rect 46385 165830 46395 165910
rect 46705 165830 46715 165910
rect 47025 165830 47035 165910
rect 47345 165830 47355 165910
rect 47665 165830 47675 165910
rect 47985 165830 47995 165910
rect 48305 165830 48315 165910
rect 43060 165820 43140 165830
rect 43380 165820 43460 165830
rect 43140 165740 43150 165820
rect 43460 165740 43470 165820
rect 48500 165810 48605 165980
rect 48640 165900 48650 165980
rect 48790 165900 48800 165980
rect 49350 165900 49360 165980
rect 49500 165900 49510 165980
rect 49650 165900 49660 165980
rect 48500 165800 48640 165810
rect 48710 165800 48790 165810
rect 49270 165800 49350 165810
rect 49420 165800 49500 165810
rect 49570 165800 49650 165810
rect 43905 165750 43985 165760
rect 44225 165750 44305 165760
rect 44545 165750 44625 165760
rect 44865 165750 44945 165760
rect 45185 165750 45265 165760
rect 45505 165750 45585 165760
rect 45825 165750 45905 165760
rect 46145 165750 46225 165760
rect 46465 165750 46545 165760
rect 46785 165750 46865 165760
rect 47105 165750 47185 165760
rect 47425 165750 47505 165760
rect 47745 165750 47825 165760
rect 48065 165750 48145 165760
rect 43985 165670 43995 165750
rect 44305 165670 44315 165750
rect 44625 165670 44635 165750
rect 44945 165670 44955 165750
rect 45265 165670 45275 165750
rect 45585 165670 45595 165750
rect 45905 165670 45915 165750
rect 46225 165670 46235 165750
rect 46545 165670 46555 165750
rect 46865 165670 46875 165750
rect 47185 165670 47195 165750
rect 47505 165670 47515 165750
rect 47825 165670 47835 165750
rect 48145 165670 48155 165750
rect 42950 165660 42980 165670
rect 43220 165660 43300 165670
rect 42980 165580 42990 165660
rect 43300 165580 43310 165660
rect 48500 165630 48605 165800
rect 48640 165720 48650 165800
rect 48790 165720 48800 165800
rect 49350 165720 49360 165800
rect 49500 165720 49510 165800
rect 49650 165720 49660 165800
rect 48500 165620 48640 165630
rect 48710 165620 48790 165630
rect 49270 165620 49350 165630
rect 49420 165620 49500 165630
rect 49570 165620 49650 165630
rect 44065 165590 44145 165600
rect 44385 165590 44465 165600
rect 44705 165590 44785 165600
rect 45025 165590 45105 165600
rect 45345 165590 45425 165600
rect 45665 165590 45745 165600
rect 45985 165590 46065 165600
rect 46305 165590 46385 165600
rect 46625 165590 46705 165600
rect 46945 165590 47025 165600
rect 47265 165590 47345 165600
rect 47585 165590 47665 165600
rect 47905 165590 47985 165600
rect 48225 165590 48305 165600
rect 44145 165510 44155 165590
rect 44465 165510 44475 165590
rect 44785 165510 44795 165590
rect 45105 165510 45115 165590
rect 45425 165510 45435 165590
rect 45745 165510 45755 165590
rect 46065 165510 46075 165590
rect 46385 165510 46395 165590
rect 46705 165510 46715 165590
rect 47025 165510 47035 165590
rect 47345 165510 47355 165590
rect 47665 165510 47675 165590
rect 47985 165510 47995 165590
rect 48305 165510 48315 165590
rect 43060 165500 43140 165510
rect 43380 165500 43460 165510
rect 43140 165420 43150 165500
rect 43460 165420 43470 165500
rect 48500 165450 48605 165620
rect 48640 165540 48650 165620
rect 48790 165540 48800 165620
rect 49350 165540 49360 165620
rect 49500 165540 49510 165620
rect 49650 165540 49660 165620
rect 48500 165440 48640 165450
rect 48710 165440 48790 165450
rect 49270 165440 49350 165450
rect 49420 165440 49500 165450
rect 49570 165440 49650 165450
rect 43905 165430 43985 165440
rect 44225 165430 44305 165440
rect 44545 165430 44625 165440
rect 44865 165430 44945 165440
rect 45185 165430 45265 165440
rect 45505 165430 45585 165440
rect 45825 165430 45905 165440
rect 46145 165430 46225 165440
rect 46465 165430 46545 165440
rect 46785 165430 46865 165440
rect 47105 165430 47185 165440
rect 47425 165430 47505 165440
rect 47745 165430 47825 165440
rect 48065 165430 48145 165440
rect 43985 165350 43995 165430
rect 44305 165350 44315 165430
rect 44625 165350 44635 165430
rect 44945 165350 44955 165430
rect 45265 165350 45275 165430
rect 45585 165350 45595 165430
rect 45905 165350 45915 165430
rect 46225 165350 46235 165430
rect 46545 165350 46555 165430
rect 46865 165350 46875 165430
rect 47185 165350 47195 165430
rect 47505 165350 47515 165430
rect 47825 165350 47835 165430
rect 48145 165350 48155 165430
rect 42950 165340 42980 165350
rect 43220 165340 43300 165350
rect 42980 165260 42990 165340
rect 43300 165260 43310 165340
rect 44065 165270 44145 165280
rect 44385 165270 44465 165280
rect 44705 165270 44785 165280
rect 45025 165270 45105 165280
rect 45345 165270 45425 165280
rect 45665 165270 45745 165280
rect 45985 165270 46065 165280
rect 46305 165270 46385 165280
rect 46625 165270 46705 165280
rect 46945 165270 47025 165280
rect 47265 165270 47345 165280
rect 47585 165270 47665 165280
rect 47905 165270 47985 165280
rect 48225 165270 48305 165280
rect 48500 165270 48605 165440
rect 48640 165360 48650 165440
rect 48790 165360 48800 165440
rect 49350 165360 49360 165440
rect 49500 165360 49510 165440
rect 49650 165360 49660 165440
rect 44145 165190 44155 165270
rect 44465 165190 44475 165270
rect 44785 165190 44795 165270
rect 45105 165190 45115 165270
rect 45425 165190 45435 165270
rect 45745 165190 45755 165270
rect 46065 165190 46075 165270
rect 46385 165190 46395 165270
rect 46705 165190 46715 165270
rect 47025 165190 47035 165270
rect 47345 165190 47355 165270
rect 47665 165190 47675 165270
rect 47985 165190 47995 165270
rect 48305 165190 48315 165270
rect 48500 165260 48640 165270
rect 48710 165260 48790 165270
rect 49270 165260 49350 165270
rect 49420 165260 49500 165270
rect 49570 165260 49650 165270
rect 43060 165180 43140 165190
rect 43380 165180 43460 165190
rect 43140 165100 43150 165180
rect 43460 165100 43470 165180
rect 43905 165110 43985 165120
rect 44225 165110 44305 165120
rect 44545 165110 44625 165120
rect 44865 165110 44945 165120
rect 45185 165110 45265 165120
rect 45505 165110 45585 165120
rect 45825 165110 45905 165120
rect 46145 165110 46225 165120
rect 46465 165110 46545 165120
rect 46785 165110 46865 165120
rect 47105 165110 47185 165120
rect 47425 165110 47505 165120
rect 47745 165110 47825 165120
rect 48065 165110 48145 165120
rect 43985 165030 43995 165110
rect 44305 165030 44315 165110
rect 44625 165030 44635 165110
rect 44945 165030 44955 165110
rect 45265 165030 45275 165110
rect 45585 165030 45595 165110
rect 45905 165030 45915 165110
rect 46225 165030 46235 165110
rect 46545 165030 46555 165110
rect 46865 165030 46875 165110
rect 47185 165030 47195 165110
rect 47505 165030 47515 165110
rect 47825 165030 47835 165110
rect 48145 165030 48155 165110
rect 48500 165090 48605 165260
rect 48640 165180 48650 165260
rect 48790 165180 48800 165260
rect 49350 165180 49360 165260
rect 49500 165180 49510 165260
rect 49650 165180 49660 165260
rect 48500 165080 48640 165090
rect 48710 165080 48790 165090
rect 49270 165080 49350 165090
rect 49420 165080 49500 165090
rect 49570 165080 49650 165090
rect 42950 165020 42980 165030
rect 43220 165020 43300 165030
rect 42980 164940 42990 165020
rect 43300 164940 43310 165020
rect 44065 164950 44145 164960
rect 44385 164950 44465 164960
rect 44705 164950 44785 164960
rect 45025 164950 45105 164960
rect 45345 164950 45425 164960
rect 45665 164950 45745 164960
rect 45985 164950 46065 164960
rect 46305 164950 46385 164960
rect 46625 164950 46705 164960
rect 46945 164950 47025 164960
rect 47265 164950 47345 164960
rect 47585 164950 47665 164960
rect 47905 164950 47985 164960
rect 48225 164950 48305 164960
rect 44145 164870 44155 164950
rect 44465 164870 44475 164950
rect 44785 164870 44795 164950
rect 45105 164870 45115 164950
rect 45425 164870 45435 164950
rect 45745 164870 45755 164950
rect 46065 164870 46075 164950
rect 46385 164870 46395 164950
rect 46705 164870 46715 164950
rect 47025 164870 47035 164950
rect 47345 164870 47355 164950
rect 47665 164870 47675 164950
rect 47985 164870 47995 164950
rect 48305 164870 48315 164950
rect 48500 164910 48605 165080
rect 48640 165000 48650 165080
rect 48790 165000 48800 165080
rect 49350 165000 49360 165080
rect 49500 165000 49510 165080
rect 49650 165000 49660 165080
rect 48500 164900 48640 164910
rect 48710 164900 48790 164910
rect 49270 164900 49350 164910
rect 49420 164900 49500 164910
rect 49570 164900 49650 164910
rect 43060 164860 43140 164870
rect 43380 164860 43460 164870
rect 43140 164780 43150 164860
rect 43460 164780 43470 164860
rect 43905 164790 43985 164800
rect 44225 164790 44305 164800
rect 44545 164790 44625 164800
rect 44865 164790 44945 164800
rect 45185 164790 45265 164800
rect 45505 164790 45585 164800
rect 45825 164790 45905 164800
rect 46145 164790 46225 164800
rect 46465 164790 46545 164800
rect 46785 164790 46865 164800
rect 47105 164790 47185 164800
rect 47425 164790 47505 164800
rect 47745 164790 47825 164800
rect 48065 164790 48145 164800
rect 43985 164710 43995 164790
rect 44305 164710 44315 164790
rect 44625 164710 44635 164790
rect 44945 164710 44955 164790
rect 45265 164710 45275 164790
rect 45585 164710 45595 164790
rect 45905 164710 45915 164790
rect 46225 164710 46235 164790
rect 46545 164710 46555 164790
rect 46865 164710 46875 164790
rect 47185 164710 47195 164790
rect 47505 164710 47515 164790
rect 47825 164710 47835 164790
rect 48145 164710 48155 164790
rect 48500 164730 48605 164900
rect 48640 164820 48650 164900
rect 48790 164820 48800 164900
rect 49350 164820 49360 164900
rect 49500 164820 49510 164900
rect 49650 164820 49660 164900
rect 48500 164720 48640 164730
rect 48710 164720 48790 164730
rect 49270 164720 49350 164730
rect 49420 164720 49500 164730
rect 49570 164720 49650 164730
rect 42950 164700 42980 164710
rect 43220 164700 43300 164710
rect 42980 164620 42990 164700
rect 43300 164620 43310 164700
rect 44065 164630 44145 164640
rect 44385 164630 44465 164640
rect 44705 164630 44785 164640
rect 45025 164630 45105 164640
rect 45345 164630 45425 164640
rect 45665 164630 45745 164640
rect 45985 164630 46065 164640
rect 46305 164630 46385 164640
rect 46625 164630 46705 164640
rect 46945 164630 47025 164640
rect 47265 164630 47345 164640
rect 47585 164630 47665 164640
rect 47905 164630 47985 164640
rect 48225 164630 48305 164640
rect 44145 164550 44155 164630
rect 44465 164550 44475 164630
rect 44785 164550 44795 164630
rect 45105 164550 45115 164630
rect 45425 164550 45435 164630
rect 45745 164550 45755 164630
rect 46065 164550 46075 164630
rect 46385 164550 46395 164630
rect 46705 164550 46715 164630
rect 47025 164550 47035 164630
rect 47345 164550 47355 164630
rect 47665 164550 47675 164630
rect 47985 164550 47995 164630
rect 48305 164550 48315 164630
rect 48500 164550 48605 164720
rect 48640 164640 48650 164720
rect 48790 164640 48800 164720
rect 49350 164640 49360 164720
rect 49500 164640 49510 164720
rect 49650 164640 49660 164720
rect 43060 164540 43140 164550
rect 43380 164540 43460 164550
rect 48500 164540 48640 164550
rect 48710 164540 48790 164550
rect 49270 164540 49350 164550
rect 49420 164540 49500 164550
rect 49570 164540 49650 164550
rect 43140 164460 43150 164540
rect 43460 164460 43470 164540
rect 43905 164470 43985 164480
rect 44225 164470 44305 164480
rect 44545 164470 44625 164480
rect 44865 164470 44945 164480
rect 45185 164470 45265 164480
rect 45505 164470 45585 164480
rect 45825 164470 45905 164480
rect 46145 164470 46225 164480
rect 46465 164470 46545 164480
rect 46785 164470 46865 164480
rect 47105 164470 47185 164480
rect 47425 164470 47505 164480
rect 47745 164470 47825 164480
rect 48065 164470 48145 164480
rect 43985 164390 43995 164470
rect 44305 164390 44315 164470
rect 44625 164390 44635 164470
rect 44945 164390 44955 164470
rect 45265 164390 45275 164470
rect 45585 164390 45595 164470
rect 45905 164390 45915 164470
rect 46225 164390 46235 164470
rect 46545 164390 46555 164470
rect 46865 164390 46875 164470
rect 47185 164390 47195 164470
rect 47505 164390 47515 164470
rect 47825 164390 47835 164470
rect 48145 164390 48155 164470
rect 42950 164380 42980 164390
rect 43220 164380 43300 164390
rect 42980 164300 42990 164380
rect 43300 164300 43310 164380
rect 48500 164370 48605 164540
rect 48640 164460 48650 164540
rect 48790 164460 48800 164540
rect 49350 164460 49360 164540
rect 49500 164460 49510 164540
rect 49650 164460 49660 164540
rect 48500 164360 48640 164370
rect 48710 164360 48790 164370
rect 49270 164360 49350 164370
rect 49420 164360 49500 164370
rect 49570 164360 49650 164370
rect 44065 164310 44145 164320
rect 44385 164310 44465 164320
rect 44705 164310 44785 164320
rect 45025 164310 45105 164320
rect 45345 164310 45425 164320
rect 45665 164310 45745 164320
rect 45985 164310 46065 164320
rect 46305 164310 46385 164320
rect 46625 164310 46705 164320
rect 46945 164310 47025 164320
rect 47265 164310 47345 164320
rect 47585 164310 47665 164320
rect 47905 164310 47985 164320
rect 48225 164310 48305 164320
rect 44145 164230 44155 164310
rect 44465 164230 44475 164310
rect 44785 164230 44795 164310
rect 45105 164230 45115 164310
rect 45425 164230 45435 164310
rect 45745 164230 45755 164310
rect 46065 164230 46075 164310
rect 46385 164230 46395 164310
rect 46705 164230 46715 164310
rect 47025 164230 47035 164310
rect 47345 164230 47355 164310
rect 47665 164230 47675 164310
rect 47985 164230 47995 164310
rect 48305 164230 48315 164310
rect 43060 164220 43140 164230
rect 43380 164220 43460 164230
rect 43140 164140 43150 164220
rect 43460 164140 43470 164220
rect 48500 164190 48605 164360
rect 48640 164280 48650 164360
rect 48790 164280 48800 164360
rect 49350 164280 49360 164360
rect 49500 164280 49510 164360
rect 49650 164280 49660 164360
rect 49790 164200 49800 170200
rect 49910 170120 49990 170130
rect 50210 170120 50290 170130
rect 49990 170040 50000 170120
rect 50290 170040 50300 170120
rect 49910 169940 49990 169950
rect 50210 169940 50290 169950
rect 49990 169860 50000 169940
rect 50290 169860 50300 169940
rect 49910 169760 49990 169770
rect 50210 169760 50290 169770
rect 49990 169680 50000 169760
rect 50290 169680 50300 169760
rect 49910 169580 49990 169590
rect 50210 169580 50290 169590
rect 49990 169500 50000 169580
rect 50290 169500 50300 169580
rect 49910 169400 49990 169410
rect 50210 169400 50290 169410
rect 49990 169320 50000 169400
rect 50290 169320 50300 169400
rect 49910 169220 49990 169230
rect 50210 169220 50290 169230
rect 49990 169140 50000 169220
rect 50290 169140 50300 169220
rect 49910 169040 49990 169050
rect 50210 169040 50290 169050
rect 49990 168960 50000 169040
rect 50290 168960 50300 169040
rect 49910 168860 49990 168870
rect 50210 168860 50290 168870
rect 49990 168780 50000 168860
rect 50290 168780 50300 168860
rect 49910 168680 49990 168690
rect 50210 168680 50290 168690
rect 49990 168600 50000 168680
rect 50290 168600 50300 168680
rect 49910 168500 49990 168510
rect 50210 168500 50290 168510
rect 49990 168420 50000 168500
rect 50290 168420 50300 168500
rect 49910 168320 49990 168330
rect 50210 168320 50290 168330
rect 49990 168240 50000 168320
rect 50290 168240 50300 168320
rect 49910 168140 49990 168150
rect 50210 168140 50290 168150
rect 49990 168060 50000 168140
rect 50290 168060 50300 168140
rect 49910 167960 49990 167970
rect 50210 167960 50290 167970
rect 49990 167880 50000 167960
rect 50290 167880 50300 167960
rect 49910 167780 49990 167790
rect 50210 167780 50290 167790
rect 49990 167700 50000 167780
rect 50290 167700 50300 167780
rect 49910 167600 49990 167610
rect 50210 167600 50290 167610
rect 49990 167520 50000 167600
rect 50290 167520 50300 167600
rect 49910 167420 49990 167430
rect 50210 167420 50290 167430
rect 49990 167340 50000 167420
rect 50290 167340 50300 167420
rect 49910 167240 49990 167250
rect 50210 167240 50290 167250
rect 49990 167160 50000 167240
rect 50290 167160 50300 167240
rect 49910 167060 49990 167070
rect 50210 167060 50290 167070
rect 49990 166980 50000 167060
rect 50290 166980 50300 167060
rect 49910 166880 49990 166890
rect 50210 166880 50290 166890
rect 49990 166800 50000 166880
rect 50290 166800 50300 166880
rect 49910 166700 49990 166710
rect 50210 166700 50290 166710
rect 49990 166620 50000 166700
rect 50290 166620 50300 166700
rect 49910 166520 49990 166530
rect 50210 166520 50290 166530
rect 49990 166440 50000 166520
rect 50290 166440 50300 166520
rect 49910 166340 49990 166350
rect 50210 166340 50290 166350
rect 49990 166260 50000 166340
rect 50290 166260 50300 166340
rect 49910 166160 49990 166170
rect 50210 166160 50290 166170
rect 49990 166080 50000 166160
rect 50290 166080 50300 166160
rect 49910 165980 49990 165990
rect 50210 165980 50290 165990
rect 49990 165900 50000 165980
rect 50290 165900 50300 165980
rect 49910 165800 49990 165810
rect 50210 165800 50290 165810
rect 49990 165720 50000 165800
rect 50290 165720 50300 165800
rect 49910 165620 49990 165630
rect 50210 165620 50290 165630
rect 49990 165540 50000 165620
rect 50290 165540 50300 165620
rect 49910 165440 49990 165450
rect 50210 165440 50290 165450
rect 49990 165360 50000 165440
rect 50290 165360 50300 165440
rect 49910 165260 49990 165270
rect 50210 165260 50290 165270
rect 49990 165180 50000 165260
rect 50290 165180 50300 165260
rect 49910 165080 49990 165090
rect 50210 165080 50290 165090
rect 49990 165000 50000 165080
rect 50290 165000 50300 165080
rect 49910 164900 49990 164910
rect 50210 164900 50290 164910
rect 49990 164820 50000 164900
rect 50290 164820 50300 164900
rect 49910 164720 49990 164730
rect 50210 164720 50290 164730
rect 49990 164640 50000 164720
rect 50290 164640 50300 164720
rect 49910 164540 49990 164550
rect 50210 164540 50290 164550
rect 49990 164460 50000 164540
rect 50290 164460 50300 164540
rect 49910 164360 49990 164370
rect 50210 164360 50290 164370
rect 49990 164280 50000 164360
rect 50290 164280 50300 164360
rect 50470 164200 50480 170200
rect 50530 170120 50610 170130
rect 50680 170120 50760 170130
rect 50830 170120 50910 170130
rect 50610 170040 50620 170120
rect 50760 170040 50770 170120
rect 50910 170040 50920 170120
rect 50530 169940 50610 169950
rect 50680 169940 50760 169950
rect 50830 169940 50910 169950
rect 50610 169860 50620 169940
rect 50760 169860 50770 169940
rect 50910 169860 50920 169940
rect 50530 169760 50610 169770
rect 50680 169760 50760 169770
rect 50830 169760 50910 169770
rect 50610 169680 50620 169760
rect 50760 169680 50770 169760
rect 50910 169680 50920 169760
rect 50530 169580 50610 169590
rect 50680 169580 50760 169590
rect 50830 169580 50910 169590
rect 50610 169500 50620 169580
rect 50760 169500 50770 169580
rect 50910 169500 50920 169580
rect 50530 169400 50610 169410
rect 50680 169400 50760 169410
rect 50830 169400 50910 169410
rect 50610 169320 50620 169400
rect 50760 169320 50770 169400
rect 50910 169320 50920 169400
rect 50530 169220 50610 169230
rect 50680 169220 50760 169230
rect 50830 169220 50910 169230
rect 50610 169140 50620 169220
rect 50760 169140 50770 169220
rect 50910 169140 50920 169220
rect 50530 169040 50610 169050
rect 50680 169040 50760 169050
rect 50830 169040 50910 169050
rect 50610 168960 50620 169040
rect 50760 168960 50770 169040
rect 50910 168960 50920 169040
rect 50530 168860 50610 168870
rect 50680 168860 50760 168870
rect 50830 168860 50910 168870
rect 50610 168780 50620 168860
rect 50760 168780 50770 168860
rect 50910 168780 50920 168860
rect 50530 168680 50610 168690
rect 50680 168680 50760 168690
rect 50830 168680 50910 168690
rect 50610 168600 50620 168680
rect 50760 168600 50770 168680
rect 50910 168600 50920 168680
rect 50530 168500 50610 168510
rect 50680 168500 50760 168510
rect 50830 168500 50910 168510
rect 50610 168420 50620 168500
rect 50760 168420 50770 168500
rect 50910 168420 50920 168500
rect 50530 168320 50610 168330
rect 50680 168320 50760 168330
rect 50830 168320 50910 168330
rect 50610 168240 50620 168320
rect 50760 168240 50770 168320
rect 50910 168240 50920 168320
rect 50530 168140 50610 168150
rect 50680 168140 50760 168150
rect 50830 168140 50910 168150
rect 50610 168060 50620 168140
rect 50760 168060 50770 168140
rect 50910 168060 50920 168140
rect 50530 167960 50610 167970
rect 50680 167960 50760 167970
rect 50830 167960 50910 167970
rect 50610 167880 50620 167960
rect 50760 167880 50770 167960
rect 50910 167880 50920 167960
rect 50530 167780 50610 167790
rect 50680 167780 50760 167790
rect 50830 167780 50910 167790
rect 50610 167700 50620 167780
rect 50760 167700 50770 167780
rect 50910 167700 50920 167780
rect 50530 167600 50610 167610
rect 50680 167600 50760 167610
rect 50830 167600 50910 167610
rect 50610 167520 50620 167600
rect 50760 167520 50770 167600
rect 50910 167520 50920 167600
rect 50530 167420 50610 167430
rect 50680 167420 50760 167430
rect 50830 167420 50910 167430
rect 50610 167340 50620 167420
rect 50760 167340 50770 167420
rect 50910 167340 50920 167420
rect 50530 167240 50610 167250
rect 50680 167240 50760 167250
rect 50830 167240 50910 167250
rect 50610 167160 50620 167240
rect 50760 167160 50770 167240
rect 50910 167160 50920 167240
rect 50530 167060 50610 167070
rect 50680 167060 50760 167070
rect 50830 167060 50910 167070
rect 50610 166980 50620 167060
rect 50760 166980 50770 167060
rect 50910 166980 50920 167060
rect 50530 166880 50610 166890
rect 50680 166880 50760 166890
rect 50830 166880 50910 166890
rect 50610 166800 50620 166880
rect 50760 166800 50770 166880
rect 50910 166800 50920 166880
rect 50530 166700 50610 166710
rect 50680 166700 50760 166710
rect 50830 166700 50910 166710
rect 50610 166620 50620 166700
rect 50760 166620 50770 166700
rect 50910 166620 50920 166700
rect 50530 166520 50610 166530
rect 50680 166520 50760 166530
rect 50830 166520 50910 166530
rect 50610 166440 50620 166520
rect 50760 166440 50770 166520
rect 50910 166440 50920 166520
rect 50530 166340 50610 166350
rect 50680 166340 50760 166350
rect 50830 166340 50910 166350
rect 50610 166260 50620 166340
rect 50760 166260 50770 166340
rect 50910 166260 50920 166340
rect 50530 166160 50610 166170
rect 50680 166160 50760 166170
rect 50830 166160 50910 166170
rect 50610 166080 50620 166160
rect 50760 166080 50770 166160
rect 50910 166080 50920 166160
rect 50530 165980 50610 165990
rect 50680 165980 50760 165990
rect 50830 165980 50910 165990
rect 50610 165900 50620 165980
rect 50760 165900 50770 165980
rect 50910 165900 50920 165980
rect 50530 165800 50610 165810
rect 50680 165800 50760 165810
rect 50830 165800 50910 165810
rect 50610 165720 50620 165800
rect 50760 165720 50770 165800
rect 50910 165720 50920 165800
rect 50530 165620 50610 165630
rect 50680 165620 50760 165630
rect 50830 165620 50910 165630
rect 50610 165540 50620 165620
rect 50760 165540 50770 165620
rect 50910 165540 50920 165620
rect 50530 165440 50610 165450
rect 50680 165440 50760 165450
rect 50830 165440 50910 165450
rect 50610 165360 50620 165440
rect 50760 165360 50770 165440
rect 50910 165360 50920 165440
rect 50530 165260 50610 165270
rect 50680 165260 50760 165270
rect 50830 165260 50910 165270
rect 50610 165180 50620 165260
rect 50760 165180 50770 165260
rect 50910 165180 50920 165260
rect 50530 165080 50610 165090
rect 50680 165080 50760 165090
rect 50830 165080 50910 165090
rect 50610 165000 50620 165080
rect 50760 165000 50770 165080
rect 50910 165000 50920 165080
rect 50530 164900 50610 164910
rect 50680 164900 50760 164910
rect 50830 164900 50910 164910
rect 50610 164820 50620 164900
rect 50760 164820 50770 164900
rect 50910 164820 50920 164900
rect 50530 164720 50610 164730
rect 50680 164720 50760 164730
rect 50830 164720 50910 164730
rect 50610 164640 50620 164720
rect 50760 164640 50770 164720
rect 50910 164640 50920 164720
rect 50530 164540 50610 164550
rect 50680 164540 50760 164550
rect 50830 164540 50910 164550
rect 50610 164460 50620 164540
rect 50760 164460 50770 164540
rect 50910 164460 50920 164540
rect 50530 164360 50610 164370
rect 50680 164360 50760 164370
rect 50830 164360 50910 164370
rect 50610 164280 50620 164360
rect 50760 164280 50770 164360
rect 50910 164280 50920 164360
rect 51050 164200 51060 170200
rect 51170 170120 51250 170130
rect 51470 170120 51550 170130
rect 51250 170040 51260 170120
rect 51550 170040 51560 170120
rect 51170 169940 51250 169950
rect 51470 169940 51550 169950
rect 51250 169860 51260 169940
rect 51550 169860 51560 169940
rect 51170 169760 51250 169770
rect 51470 169760 51550 169770
rect 51250 169680 51260 169760
rect 51550 169680 51560 169760
rect 51170 169580 51250 169590
rect 51470 169580 51550 169590
rect 51250 169500 51260 169580
rect 51550 169500 51560 169580
rect 51170 169400 51250 169410
rect 51470 169400 51550 169410
rect 51250 169320 51260 169400
rect 51550 169320 51560 169400
rect 51170 169220 51250 169230
rect 51470 169220 51550 169230
rect 51250 169140 51260 169220
rect 51550 169140 51560 169220
rect 51170 169040 51250 169050
rect 51470 169040 51550 169050
rect 51250 168960 51260 169040
rect 51550 168960 51560 169040
rect 51170 168860 51250 168870
rect 51470 168860 51550 168870
rect 51250 168780 51260 168860
rect 51550 168780 51560 168860
rect 51170 168680 51250 168690
rect 51470 168680 51550 168690
rect 51250 168600 51260 168680
rect 51550 168600 51560 168680
rect 51170 168500 51250 168510
rect 51470 168500 51550 168510
rect 51250 168420 51260 168500
rect 51550 168420 51560 168500
rect 51170 168320 51250 168330
rect 51470 168320 51550 168330
rect 51250 168240 51260 168320
rect 51550 168240 51560 168320
rect 51170 168140 51250 168150
rect 51470 168140 51550 168150
rect 51250 168060 51260 168140
rect 51550 168060 51560 168140
rect 51170 167960 51250 167970
rect 51470 167960 51550 167970
rect 51250 167880 51260 167960
rect 51550 167880 51560 167960
rect 51170 167780 51250 167790
rect 51470 167780 51550 167790
rect 51250 167700 51260 167780
rect 51550 167700 51560 167780
rect 51170 167600 51250 167610
rect 51470 167600 51550 167610
rect 51250 167520 51260 167600
rect 51550 167520 51560 167600
rect 51170 167420 51250 167430
rect 51470 167420 51550 167430
rect 51250 167340 51260 167420
rect 51550 167340 51560 167420
rect 51170 167240 51250 167250
rect 51470 167240 51550 167250
rect 51250 167160 51260 167240
rect 51550 167160 51560 167240
rect 51170 167060 51250 167070
rect 51470 167060 51550 167070
rect 51250 166980 51260 167060
rect 51550 166980 51560 167060
rect 51170 166880 51250 166890
rect 51470 166880 51550 166890
rect 51250 166800 51260 166880
rect 51550 166800 51560 166880
rect 51170 166700 51250 166710
rect 51470 166700 51550 166710
rect 51250 166620 51260 166700
rect 51550 166620 51560 166700
rect 51170 166520 51250 166530
rect 51470 166520 51550 166530
rect 51250 166440 51260 166520
rect 51550 166440 51560 166520
rect 51170 166340 51250 166350
rect 51470 166340 51550 166350
rect 51250 166260 51260 166340
rect 51550 166260 51560 166340
rect 51170 166160 51250 166170
rect 51470 166160 51550 166170
rect 51250 166080 51260 166160
rect 51550 166080 51560 166160
rect 51170 165980 51250 165990
rect 51470 165980 51550 165990
rect 51250 165900 51260 165980
rect 51550 165900 51560 165980
rect 51170 165800 51250 165810
rect 51470 165800 51550 165810
rect 51250 165720 51260 165800
rect 51550 165720 51560 165800
rect 51170 165620 51250 165630
rect 51470 165620 51550 165630
rect 51250 165540 51260 165620
rect 51550 165540 51560 165620
rect 51170 165440 51250 165450
rect 51470 165440 51550 165450
rect 51250 165360 51260 165440
rect 51550 165360 51560 165440
rect 51170 165260 51250 165270
rect 51470 165260 51550 165270
rect 51250 165180 51260 165260
rect 51550 165180 51560 165260
rect 51170 165080 51250 165090
rect 51470 165080 51550 165090
rect 51250 165000 51260 165080
rect 51550 165000 51560 165080
rect 51170 164900 51250 164910
rect 51470 164900 51550 164910
rect 51250 164820 51260 164900
rect 51550 164820 51560 164900
rect 51170 164720 51250 164730
rect 51470 164720 51550 164730
rect 51250 164640 51260 164720
rect 51550 164640 51560 164720
rect 51170 164540 51250 164550
rect 51470 164540 51550 164550
rect 51250 164460 51260 164540
rect 51550 164460 51560 164540
rect 51170 164360 51250 164370
rect 51470 164360 51550 164370
rect 51250 164280 51260 164360
rect 51550 164280 51560 164360
rect 51730 164200 51740 170200
rect 51790 170120 51870 170130
rect 51940 170120 52020 170130
rect 52090 170120 52170 170130
rect 51870 170040 51880 170120
rect 52020 170040 52030 170120
rect 52170 170040 52180 170120
rect 51790 169940 51870 169950
rect 51940 169940 52020 169950
rect 52090 169940 52170 169950
rect 51870 169860 51880 169940
rect 52020 169860 52030 169940
rect 52170 169860 52180 169940
rect 51790 169760 51870 169770
rect 51940 169760 52020 169770
rect 52090 169760 52170 169770
rect 51870 169680 51880 169760
rect 52020 169680 52030 169760
rect 52170 169680 52180 169760
rect 51790 169580 51870 169590
rect 51940 169580 52020 169590
rect 52090 169580 52170 169590
rect 51870 169500 51880 169580
rect 52020 169500 52030 169580
rect 52170 169500 52180 169580
rect 51790 169400 51870 169410
rect 51940 169400 52020 169410
rect 52090 169400 52170 169410
rect 51870 169320 51880 169400
rect 52020 169320 52030 169400
rect 52170 169320 52180 169400
rect 51790 169220 51870 169230
rect 51940 169220 52020 169230
rect 52090 169220 52170 169230
rect 51870 169140 51880 169220
rect 52020 169140 52030 169220
rect 52170 169140 52180 169220
rect 51790 169040 51870 169050
rect 51940 169040 52020 169050
rect 52090 169040 52170 169050
rect 51870 168960 51880 169040
rect 52020 168960 52030 169040
rect 52170 168960 52180 169040
rect 51790 168860 51870 168870
rect 51940 168860 52020 168870
rect 52090 168860 52170 168870
rect 51870 168780 51880 168860
rect 52020 168780 52030 168860
rect 52170 168780 52180 168860
rect 51790 168680 51870 168690
rect 51940 168680 52020 168690
rect 52090 168680 52170 168690
rect 51870 168600 51880 168680
rect 52020 168600 52030 168680
rect 52170 168600 52180 168680
rect 51790 168500 51870 168510
rect 51940 168500 52020 168510
rect 52090 168500 52170 168510
rect 51870 168420 51880 168500
rect 52020 168420 52030 168500
rect 52170 168420 52180 168500
rect 51790 168320 51870 168330
rect 51940 168320 52020 168330
rect 52090 168320 52170 168330
rect 51870 168240 51880 168320
rect 52020 168240 52030 168320
rect 52170 168240 52180 168320
rect 51790 168140 51870 168150
rect 51940 168140 52020 168150
rect 52090 168140 52170 168150
rect 51870 168060 51880 168140
rect 52020 168060 52030 168140
rect 52170 168060 52180 168140
rect 51790 167960 51870 167970
rect 51940 167960 52020 167970
rect 52090 167960 52170 167970
rect 51870 167880 51880 167960
rect 52020 167880 52030 167960
rect 52170 167880 52180 167960
rect 51790 167780 51870 167790
rect 51940 167780 52020 167790
rect 52090 167780 52170 167790
rect 51870 167700 51880 167780
rect 52020 167700 52030 167780
rect 52170 167700 52180 167780
rect 51790 167600 51870 167610
rect 51940 167600 52020 167610
rect 52090 167600 52170 167610
rect 51870 167520 51880 167600
rect 52020 167520 52030 167600
rect 52170 167520 52180 167600
rect 51790 167420 51870 167430
rect 51940 167420 52020 167430
rect 52090 167420 52170 167430
rect 51870 167340 51880 167420
rect 52020 167340 52030 167420
rect 52170 167340 52180 167420
rect 51790 167240 51870 167250
rect 51940 167240 52020 167250
rect 52090 167240 52170 167250
rect 51870 167160 51880 167240
rect 52020 167160 52030 167240
rect 52170 167160 52180 167240
rect 51790 167060 51870 167070
rect 51940 167060 52020 167070
rect 52090 167060 52170 167070
rect 51870 166980 51880 167060
rect 52020 166980 52030 167060
rect 52170 166980 52180 167060
rect 51790 166880 51870 166890
rect 51940 166880 52020 166890
rect 52090 166880 52170 166890
rect 51870 166800 51880 166880
rect 52020 166800 52030 166880
rect 52170 166800 52180 166880
rect 51790 166700 51870 166710
rect 51940 166700 52020 166710
rect 52090 166700 52170 166710
rect 51870 166620 51880 166700
rect 52020 166620 52030 166700
rect 52170 166620 52180 166700
rect 51790 166520 51870 166530
rect 51940 166520 52020 166530
rect 52090 166520 52170 166530
rect 51870 166440 51880 166520
rect 52020 166440 52030 166520
rect 52170 166440 52180 166520
rect 51790 166340 51870 166350
rect 51940 166340 52020 166350
rect 52090 166340 52170 166350
rect 51870 166260 51880 166340
rect 52020 166260 52030 166340
rect 52170 166260 52180 166340
rect 51790 166160 51870 166170
rect 51940 166160 52020 166170
rect 52090 166160 52170 166170
rect 51870 166080 51880 166160
rect 52020 166080 52030 166160
rect 52170 166080 52180 166160
rect 51790 165980 51870 165990
rect 51940 165980 52020 165990
rect 52090 165980 52170 165990
rect 51870 165900 51880 165980
rect 52020 165900 52030 165980
rect 52170 165900 52180 165980
rect 51790 165800 51870 165810
rect 51940 165800 52020 165810
rect 52090 165800 52170 165810
rect 51870 165720 51880 165800
rect 52020 165720 52030 165800
rect 52170 165720 52180 165800
rect 51790 165620 51870 165630
rect 51940 165620 52020 165630
rect 52090 165620 52170 165630
rect 51870 165540 51880 165620
rect 52020 165540 52030 165620
rect 52170 165540 52180 165620
rect 51790 165440 51870 165450
rect 51940 165440 52020 165450
rect 52090 165440 52170 165450
rect 51870 165360 51880 165440
rect 52020 165360 52030 165440
rect 52170 165360 52180 165440
rect 51790 165260 51870 165270
rect 51940 165260 52020 165270
rect 52090 165260 52170 165270
rect 51870 165180 51880 165260
rect 52020 165180 52030 165260
rect 52170 165180 52180 165260
rect 51790 165080 51870 165090
rect 51940 165080 52020 165090
rect 52090 165080 52170 165090
rect 51870 165000 51880 165080
rect 52020 165000 52030 165080
rect 52170 165000 52180 165080
rect 51790 164900 51870 164910
rect 51940 164900 52020 164910
rect 52090 164900 52170 164910
rect 51870 164820 51880 164900
rect 52020 164820 52030 164900
rect 52170 164820 52180 164900
rect 51790 164720 51870 164730
rect 51940 164720 52020 164730
rect 52090 164720 52170 164730
rect 51870 164640 51880 164720
rect 52020 164640 52030 164720
rect 52170 164640 52180 164720
rect 51790 164540 51870 164550
rect 51940 164540 52020 164550
rect 52090 164540 52170 164550
rect 51870 164460 51880 164540
rect 52020 164460 52030 164540
rect 52170 164460 52180 164540
rect 51790 164360 51870 164370
rect 51940 164360 52020 164370
rect 52090 164360 52170 164370
rect 51870 164280 51880 164360
rect 52020 164280 52030 164360
rect 52170 164280 52180 164360
rect 52310 164200 52320 170200
rect 52430 170120 52510 170130
rect 52730 170120 52810 170130
rect 52510 170040 52520 170120
rect 52810 170040 52820 170120
rect 52430 169940 52510 169950
rect 52730 169940 52810 169950
rect 52510 169860 52520 169940
rect 52810 169860 52820 169940
rect 52430 169760 52510 169770
rect 52730 169760 52810 169770
rect 52510 169680 52520 169760
rect 52810 169680 52820 169760
rect 52430 169580 52510 169590
rect 52730 169580 52810 169590
rect 52510 169500 52520 169580
rect 52810 169500 52820 169580
rect 52430 169400 52510 169410
rect 52730 169400 52810 169410
rect 52510 169320 52520 169400
rect 52810 169320 52820 169400
rect 52430 169220 52510 169230
rect 52730 169220 52810 169230
rect 52510 169140 52520 169220
rect 52810 169140 52820 169220
rect 52430 169040 52510 169050
rect 52730 169040 52810 169050
rect 52510 168960 52520 169040
rect 52810 168960 52820 169040
rect 52430 168860 52510 168870
rect 52730 168860 52810 168870
rect 52510 168780 52520 168860
rect 52810 168780 52820 168860
rect 52430 168680 52510 168690
rect 52730 168680 52810 168690
rect 52510 168600 52520 168680
rect 52810 168600 52820 168680
rect 52430 168500 52510 168510
rect 52730 168500 52810 168510
rect 52510 168420 52520 168500
rect 52810 168420 52820 168500
rect 52430 168320 52510 168330
rect 52730 168320 52810 168330
rect 52510 168240 52520 168320
rect 52810 168240 52820 168320
rect 52430 168140 52510 168150
rect 52730 168140 52810 168150
rect 52510 168060 52520 168140
rect 52810 168060 52820 168140
rect 52430 167960 52510 167970
rect 52730 167960 52810 167970
rect 52510 167880 52520 167960
rect 52810 167880 52820 167960
rect 52430 167780 52510 167790
rect 52730 167780 52810 167790
rect 52510 167700 52520 167780
rect 52810 167700 52820 167780
rect 52430 167600 52510 167610
rect 52730 167600 52810 167610
rect 52510 167520 52520 167600
rect 52810 167520 52820 167600
rect 52430 167420 52510 167430
rect 52730 167420 52810 167430
rect 52510 167340 52520 167420
rect 52810 167340 52820 167420
rect 52430 167240 52510 167250
rect 52730 167240 52810 167250
rect 52510 167160 52520 167240
rect 52810 167160 52820 167240
rect 52430 167060 52510 167070
rect 52730 167060 52810 167070
rect 52510 166980 52520 167060
rect 52810 166980 52820 167060
rect 52430 166880 52510 166890
rect 52730 166880 52810 166890
rect 52510 166800 52520 166880
rect 52810 166800 52820 166880
rect 52430 166700 52510 166710
rect 52730 166700 52810 166710
rect 52510 166620 52520 166700
rect 52810 166620 52820 166700
rect 52430 166520 52510 166530
rect 52730 166520 52810 166530
rect 52510 166440 52520 166520
rect 52810 166440 52820 166520
rect 52430 166340 52510 166350
rect 52730 166340 52810 166350
rect 52510 166260 52520 166340
rect 52810 166260 52820 166340
rect 52430 166160 52510 166170
rect 52730 166160 52810 166170
rect 52510 166080 52520 166160
rect 52810 166080 52820 166160
rect 52430 165980 52510 165990
rect 52730 165980 52810 165990
rect 52510 165900 52520 165980
rect 52810 165900 52820 165980
rect 52430 165800 52510 165810
rect 52730 165800 52810 165810
rect 52510 165720 52520 165800
rect 52810 165720 52820 165800
rect 52430 165620 52510 165630
rect 52730 165620 52810 165630
rect 52510 165540 52520 165620
rect 52810 165540 52820 165620
rect 52430 165440 52510 165450
rect 52730 165440 52810 165450
rect 52510 165360 52520 165440
rect 52810 165360 52820 165440
rect 52430 165260 52510 165270
rect 52730 165260 52810 165270
rect 52510 165180 52520 165260
rect 52810 165180 52820 165260
rect 52430 165080 52510 165090
rect 52730 165080 52810 165090
rect 52510 165000 52520 165080
rect 52810 165000 52820 165080
rect 52430 164900 52510 164910
rect 52730 164900 52810 164910
rect 52510 164820 52520 164900
rect 52810 164820 52820 164900
rect 52430 164720 52510 164730
rect 52730 164720 52810 164730
rect 52510 164640 52520 164720
rect 52810 164640 52820 164720
rect 52430 164540 52510 164550
rect 52730 164540 52810 164550
rect 52510 164460 52520 164540
rect 52810 164460 52820 164540
rect 52430 164360 52510 164370
rect 52730 164360 52810 164370
rect 52510 164280 52520 164360
rect 52810 164280 52820 164360
rect 52990 164200 53000 170200
rect 53050 170120 53130 170130
rect 53200 170120 53280 170130
rect 53350 170120 53430 170130
rect 53130 170040 53140 170120
rect 53280 170040 53290 170120
rect 53430 170040 53440 170120
rect 53050 169940 53130 169950
rect 53200 169940 53280 169950
rect 53350 169940 53430 169950
rect 53130 169860 53140 169940
rect 53280 169860 53290 169940
rect 53430 169860 53440 169940
rect 53050 169760 53130 169770
rect 53200 169760 53280 169770
rect 53350 169760 53430 169770
rect 53130 169680 53140 169760
rect 53280 169680 53290 169760
rect 53430 169680 53440 169760
rect 53050 169580 53130 169590
rect 53200 169580 53280 169590
rect 53350 169580 53430 169590
rect 53130 169500 53140 169580
rect 53280 169500 53290 169580
rect 53430 169500 53440 169580
rect 53050 169400 53130 169410
rect 53200 169400 53280 169410
rect 53350 169400 53430 169410
rect 53130 169320 53140 169400
rect 53280 169320 53290 169400
rect 53430 169320 53440 169400
rect 53050 169220 53130 169230
rect 53200 169220 53280 169230
rect 53350 169220 53430 169230
rect 53130 169140 53140 169220
rect 53280 169140 53290 169220
rect 53430 169140 53440 169220
rect 53050 169040 53130 169050
rect 53200 169040 53280 169050
rect 53350 169040 53430 169050
rect 53130 168960 53140 169040
rect 53280 168960 53290 169040
rect 53430 168960 53440 169040
rect 53050 168860 53130 168870
rect 53200 168860 53280 168870
rect 53350 168860 53430 168870
rect 53130 168780 53140 168860
rect 53280 168780 53290 168860
rect 53430 168780 53440 168860
rect 53050 168680 53130 168690
rect 53200 168680 53280 168690
rect 53350 168680 53430 168690
rect 53130 168600 53140 168680
rect 53280 168600 53290 168680
rect 53430 168600 53440 168680
rect 53050 168500 53130 168510
rect 53200 168500 53280 168510
rect 53350 168500 53430 168510
rect 53130 168420 53140 168500
rect 53280 168420 53290 168500
rect 53430 168420 53440 168500
rect 53050 168320 53130 168330
rect 53200 168320 53280 168330
rect 53350 168320 53430 168330
rect 53130 168240 53140 168320
rect 53280 168240 53290 168320
rect 53430 168240 53440 168320
rect 53050 168140 53130 168150
rect 53200 168140 53280 168150
rect 53350 168140 53430 168150
rect 53130 168060 53140 168140
rect 53280 168060 53290 168140
rect 53430 168060 53440 168140
rect 53050 167960 53130 167970
rect 53200 167960 53280 167970
rect 53350 167960 53430 167970
rect 53130 167880 53140 167960
rect 53280 167880 53290 167960
rect 53430 167880 53440 167960
rect 53050 167780 53130 167790
rect 53200 167780 53280 167790
rect 53350 167780 53430 167790
rect 53130 167700 53140 167780
rect 53280 167700 53290 167780
rect 53430 167700 53440 167780
rect 53050 167600 53130 167610
rect 53200 167600 53280 167610
rect 53350 167600 53430 167610
rect 53130 167520 53140 167600
rect 53280 167520 53290 167600
rect 53430 167520 53440 167600
rect 53050 167420 53130 167430
rect 53200 167420 53280 167430
rect 53350 167420 53430 167430
rect 53130 167340 53140 167420
rect 53280 167340 53290 167420
rect 53430 167340 53440 167420
rect 53050 167240 53130 167250
rect 53200 167240 53280 167250
rect 53350 167240 53430 167250
rect 53130 167160 53140 167240
rect 53280 167160 53290 167240
rect 53430 167160 53440 167240
rect 53050 167060 53130 167070
rect 53200 167060 53280 167070
rect 53350 167060 53430 167070
rect 53130 166980 53140 167060
rect 53280 166980 53290 167060
rect 53430 166980 53440 167060
rect 53050 166880 53130 166890
rect 53200 166880 53280 166890
rect 53350 166880 53430 166890
rect 53130 166800 53140 166880
rect 53280 166800 53290 166880
rect 53430 166800 53440 166880
rect 53050 166700 53130 166710
rect 53200 166700 53280 166710
rect 53350 166700 53430 166710
rect 53130 166620 53140 166700
rect 53280 166620 53290 166700
rect 53430 166620 53440 166700
rect 53050 166520 53130 166530
rect 53200 166520 53280 166530
rect 53350 166520 53430 166530
rect 53130 166440 53140 166520
rect 53280 166440 53290 166520
rect 53430 166440 53440 166520
rect 53050 166340 53130 166350
rect 53200 166340 53280 166350
rect 53350 166340 53430 166350
rect 53130 166260 53140 166340
rect 53280 166260 53290 166340
rect 53430 166260 53440 166340
rect 53050 166160 53130 166170
rect 53200 166160 53280 166170
rect 53350 166160 53430 166170
rect 53130 166080 53140 166160
rect 53280 166080 53290 166160
rect 53430 166080 53440 166160
rect 53050 165980 53130 165990
rect 53200 165980 53280 165990
rect 53350 165980 53430 165990
rect 53130 165900 53140 165980
rect 53280 165900 53290 165980
rect 53430 165900 53440 165980
rect 53050 165800 53130 165810
rect 53200 165800 53280 165810
rect 53350 165800 53430 165810
rect 53130 165720 53140 165800
rect 53280 165720 53290 165800
rect 53430 165720 53440 165800
rect 53050 165620 53130 165630
rect 53200 165620 53280 165630
rect 53350 165620 53430 165630
rect 53130 165540 53140 165620
rect 53280 165540 53290 165620
rect 53430 165540 53440 165620
rect 53050 165440 53130 165450
rect 53200 165440 53280 165450
rect 53350 165440 53430 165450
rect 53130 165360 53140 165440
rect 53280 165360 53290 165440
rect 53430 165360 53440 165440
rect 53050 165260 53130 165270
rect 53200 165260 53280 165270
rect 53350 165260 53430 165270
rect 53130 165180 53140 165260
rect 53280 165180 53290 165260
rect 53430 165180 53440 165260
rect 53050 165080 53130 165090
rect 53200 165080 53280 165090
rect 53350 165080 53430 165090
rect 53130 165000 53140 165080
rect 53280 165000 53290 165080
rect 53430 165000 53440 165080
rect 53050 164900 53130 164910
rect 53200 164900 53280 164910
rect 53350 164900 53430 164910
rect 53130 164820 53140 164900
rect 53280 164820 53290 164900
rect 53430 164820 53440 164900
rect 53050 164720 53130 164730
rect 53200 164720 53280 164730
rect 53350 164720 53430 164730
rect 53130 164640 53140 164720
rect 53280 164640 53290 164720
rect 53430 164640 53440 164720
rect 53050 164540 53130 164550
rect 53200 164540 53280 164550
rect 53350 164540 53430 164550
rect 53130 164460 53140 164540
rect 53280 164460 53290 164540
rect 53430 164460 53440 164540
rect 53050 164360 53130 164370
rect 53200 164360 53280 164370
rect 53350 164360 53430 164370
rect 53130 164280 53140 164360
rect 53280 164280 53290 164360
rect 53430 164280 53440 164360
rect 53570 164200 53580 170200
rect 53690 170120 53770 170130
rect 53990 170120 54070 170130
rect 53770 170040 53780 170120
rect 54070 170040 54080 170120
rect 53690 169940 53770 169950
rect 53990 169940 54070 169950
rect 53770 169860 53780 169940
rect 54070 169860 54080 169940
rect 53690 169760 53770 169770
rect 53990 169760 54070 169770
rect 53770 169680 53780 169760
rect 54070 169680 54080 169760
rect 53690 169580 53770 169590
rect 53990 169580 54070 169590
rect 53770 169500 53780 169580
rect 54070 169500 54080 169580
rect 53690 169400 53770 169410
rect 53990 169400 54070 169410
rect 53770 169320 53780 169400
rect 54070 169320 54080 169400
rect 53690 169220 53770 169230
rect 53990 169220 54070 169230
rect 53770 169140 53780 169220
rect 54070 169140 54080 169220
rect 53690 169040 53770 169050
rect 53990 169040 54070 169050
rect 53770 168960 53780 169040
rect 54070 168960 54080 169040
rect 53690 168860 53770 168870
rect 53990 168860 54070 168870
rect 53770 168780 53780 168860
rect 54070 168780 54080 168860
rect 53690 168680 53770 168690
rect 53990 168680 54070 168690
rect 53770 168600 53780 168680
rect 54070 168600 54080 168680
rect 53690 168500 53770 168510
rect 53990 168500 54070 168510
rect 53770 168420 53780 168500
rect 54070 168420 54080 168500
rect 53690 168320 53770 168330
rect 53990 168320 54070 168330
rect 53770 168240 53780 168320
rect 54070 168240 54080 168320
rect 53690 168140 53770 168150
rect 53990 168140 54070 168150
rect 53770 168060 53780 168140
rect 54070 168060 54080 168140
rect 53690 167960 53770 167970
rect 53990 167960 54070 167970
rect 53770 167880 53780 167960
rect 54070 167880 54080 167960
rect 53690 167780 53770 167790
rect 53990 167780 54070 167790
rect 53770 167700 53780 167780
rect 54070 167700 54080 167780
rect 53690 167600 53770 167610
rect 53990 167600 54070 167610
rect 53770 167520 53780 167600
rect 54070 167520 54080 167600
rect 53690 167420 53770 167430
rect 53990 167420 54070 167430
rect 53770 167340 53780 167420
rect 54070 167340 54080 167420
rect 53690 167240 53770 167250
rect 53990 167240 54070 167250
rect 53770 167160 53780 167240
rect 54070 167160 54080 167240
rect 53690 167060 53770 167070
rect 53990 167060 54070 167070
rect 53770 166980 53780 167060
rect 54070 166980 54080 167060
rect 53690 166880 53770 166890
rect 53990 166880 54070 166890
rect 53770 166800 53780 166880
rect 54070 166800 54080 166880
rect 53690 166700 53770 166710
rect 53990 166700 54070 166710
rect 53770 166620 53780 166700
rect 54070 166620 54080 166700
rect 53690 166520 53770 166530
rect 53990 166520 54070 166530
rect 53770 166440 53780 166520
rect 54070 166440 54080 166520
rect 53690 166340 53770 166350
rect 53990 166340 54070 166350
rect 53770 166260 53780 166340
rect 54070 166260 54080 166340
rect 53690 166160 53770 166170
rect 53990 166160 54070 166170
rect 53770 166080 53780 166160
rect 54070 166080 54080 166160
rect 53690 165980 53770 165990
rect 53990 165980 54070 165990
rect 53770 165900 53780 165980
rect 54070 165900 54080 165980
rect 53690 165800 53770 165810
rect 53990 165800 54070 165810
rect 53770 165720 53780 165800
rect 54070 165720 54080 165800
rect 53690 165620 53770 165630
rect 53990 165620 54070 165630
rect 53770 165540 53780 165620
rect 54070 165540 54080 165620
rect 53690 165440 53770 165450
rect 53990 165440 54070 165450
rect 53770 165360 53780 165440
rect 54070 165360 54080 165440
rect 53690 165260 53770 165270
rect 53990 165260 54070 165270
rect 53770 165180 53780 165260
rect 54070 165180 54080 165260
rect 53690 165080 53770 165090
rect 53990 165080 54070 165090
rect 53770 165000 53780 165080
rect 54070 165000 54080 165080
rect 53690 164900 53770 164910
rect 53990 164900 54070 164910
rect 53770 164820 53780 164900
rect 54070 164820 54080 164900
rect 53690 164720 53770 164730
rect 53990 164720 54070 164730
rect 53770 164640 53780 164720
rect 54070 164640 54080 164720
rect 53690 164540 53770 164550
rect 53990 164540 54070 164550
rect 53770 164460 53780 164540
rect 54070 164460 54080 164540
rect 53690 164360 53770 164370
rect 53990 164360 54070 164370
rect 53770 164280 53780 164360
rect 54070 164280 54080 164360
rect 54250 164200 54260 170200
rect 54310 170120 54390 170130
rect 54460 170120 54540 170130
rect 54610 170120 54690 170130
rect 54390 170040 54400 170120
rect 54540 170040 54550 170120
rect 54690 170040 54700 170120
rect 54310 169940 54390 169950
rect 54460 169940 54540 169950
rect 54610 169940 54690 169950
rect 54390 169860 54400 169940
rect 54540 169860 54550 169940
rect 54690 169860 54700 169940
rect 54310 169760 54390 169770
rect 54460 169760 54540 169770
rect 54610 169760 54690 169770
rect 54390 169680 54400 169760
rect 54540 169680 54550 169760
rect 54690 169680 54700 169760
rect 54310 169580 54390 169590
rect 54460 169580 54540 169590
rect 54610 169580 54690 169590
rect 54390 169500 54400 169580
rect 54540 169500 54550 169580
rect 54690 169500 54700 169580
rect 54310 169400 54390 169410
rect 54460 169400 54540 169410
rect 54610 169400 54690 169410
rect 54390 169320 54400 169400
rect 54540 169320 54550 169400
rect 54690 169320 54700 169400
rect 54310 169220 54390 169230
rect 54460 169220 54540 169230
rect 54610 169220 54690 169230
rect 54390 169140 54400 169220
rect 54540 169140 54550 169220
rect 54690 169140 54700 169220
rect 54310 169040 54390 169050
rect 54460 169040 54540 169050
rect 54610 169040 54690 169050
rect 54390 168960 54400 169040
rect 54540 168960 54550 169040
rect 54690 168960 54700 169040
rect 54310 168860 54390 168870
rect 54460 168860 54540 168870
rect 54610 168860 54690 168870
rect 54390 168780 54400 168860
rect 54540 168780 54550 168860
rect 54690 168780 54700 168860
rect 54310 168680 54390 168690
rect 54460 168680 54540 168690
rect 54610 168680 54690 168690
rect 54390 168600 54400 168680
rect 54540 168600 54550 168680
rect 54690 168600 54700 168680
rect 54310 168500 54390 168510
rect 54460 168500 54540 168510
rect 54610 168500 54690 168510
rect 54390 168420 54400 168500
rect 54540 168420 54550 168500
rect 54690 168420 54700 168500
rect 54310 168320 54390 168330
rect 54460 168320 54540 168330
rect 54610 168320 54690 168330
rect 54390 168240 54400 168320
rect 54540 168240 54550 168320
rect 54690 168240 54700 168320
rect 54310 168140 54390 168150
rect 54460 168140 54540 168150
rect 54610 168140 54690 168150
rect 54390 168060 54400 168140
rect 54540 168060 54550 168140
rect 54690 168060 54700 168140
rect 54310 167960 54390 167970
rect 54460 167960 54540 167970
rect 54610 167960 54690 167970
rect 54390 167880 54400 167960
rect 54540 167880 54550 167960
rect 54690 167880 54700 167960
rect 54310 167780 54390 167790
rect 54460 167780 54540 167790
rect 54610 167780 54690 167790
rect 54390 167700 54400 167780
rect 54540 167700 54550 167780
rect 54690 167700 54700 167780
rect 54310 167600 54390 167610
rect 54460 167600 54540 167610
rect 54610 167600 54690 167610
rect 54390 167520 54400 167600
rect 54540 167520 54550 167600
rect 54690 167520 54700 167600
rect 54310 167420 54390 167430
rect 54460 167420 54540 167430
rect 54610 167420 54690 167430
rect 54390 167340 54400 167420
rect 54540 167340 54550 167420
rect 54690 167340 54700 167420
rect 54310 167240 54390 167250
rect 54460 167240 54540 167250
rect 54610 167240 54690 167250
rect 54390 167160 54400 167240
rect 54540 167160 54550 167240
rect 54690 167160 54700 167240
rect 54310 167060 54390 167070
rect 54460 167060 54540 167070
rect 54610 167060 54690 167070
rect 54390 166980 54400 167060
rect 54540 166980 54550 167060
rect 54690 166980 54700 167060
rect 54310 166880 54390 166890
rect 54460 166880 54540 166890
rect 54610 166880 54690 166890
rect 54390 166800 54400 166880
rect 54540 166800 54550 166880
rect 54690 166800 54700 166880
rect 54310 166700 54390 166710
rect 54460 166700 54540 166710
rect 54610 166700 54690 166710
rect 54390 166620 54400 166700
rect 54540 166620 54550 166700
rect 54690 166620 54700 166700
rect 54310 166520 54390 166530
rect 54460 166520 54540 166530
rect 54610 166520 54690 166530
rect 54390 166440 54400 166520
rect 54540 166440 54550 166520
rect 54690 166440 54700 166520
rect 54310 166340 54390 166350
rect 54460 166340 54540 166350
rect 54610 166340 54690 166350
rect 54390 166260 54400 166340
rect 54540 166260 54550 166340
rect 54690 166260 54700 166340
rect 54310 166160 54390 166170
rect 54460 166160 54540 166170
rect 54610 166160 54690 166170
rect 54390 166080 54400 166160
rect 54540 166080 54550 166160
rect 54690 166080 54700 166160
rect 54310 165980 54390 165990
rect 54460 165980 54540 165990
rect 54610 165980 54690 165990
rect 54390 165900 54400 165980
rect 54540 165900 54550 165980
rect 54690 165900 54700 165980
rect 54310 165800 54390 165810
rect 54460 165800 54540 165810
rect 54610 165800 54690 165810
rect 54390 165720 54400 165800
rect 54540 165720 54550 165800
rect 54690 165720 54700 165800
rect 54310 165620 54390 165630
rect 54460 165620 54540 165630
rect 54610 165620 54690 165630
rect 54390 165540 54400 165620
rect 54540 165540 54550 165620
rect 54690 165540 54700 165620
rect 54310 165440 54390 165450
rect 54460 165440 54540 165450
rect 54610 165440 54690 165450
rect 54390 165360 54400 165440
rect 54540 165360 54550 165440
rect 54690 165360 54700 165440
rect 54310 165260 54390 165270
rect 54460 165260 54540 165270
rect 54610 165260 54690 165270
rect 54390 165180 54400 165260
rect 54540 165180 54550 165260
rect 54690 165180 54700 165260
rect 54310 165080 54390 165090
rect 54460 165080 54540 165090
rect 54610 165080 54690 165090
rect 54390 165000 54400 165080
rect 54540 165000 54550 165080
rect 54690 165000 54700 165080
rect 54310 164900 54390 164910
rect 54460 164900 54540 164910
rect 54610 164900 54690 164910
rect 54390 164820 54400 164900
rect 54540 164820 54550 164900
rect 54690 164820 54700 164900
rect 54310 164720 54390 164730
rect 54460 164720 54540 164730
rect 54610 164720 54690 164730
rect 54390 164640 54400 164720
rect 54540 164640 54550 164720
rect 54690 164640 54700 164720
rect 54310 164540 54390 164550
rect 54460 164540 54540 164550
rect 54610 164540 54690 164550
rect 54390 164460 54400 164540
rect 54540 164460 54550 164540
rect 54690 164460 54700 164540
rect 54310 164360 54390 164370
rect 54460 164360 54540 164370
rect 54610 164360 54690 164370
rect 54390 164280 54400 164360
rect 54540 164280 54550 164360
rect 54690 164280 54700 164360
rect 54830 164200 54840 170200
rect 54950 170120 55030 170130
rect 55250 170120 55330 170130
rect 55030 170040 55040 170120
rect 55330 170040 55340 170120
rect 54950 169940 55030 169950
rect 55250 169940 55330 169950
rect 55030 169860 55040 169940
rect 55330 169860 55340 169940
rect 54950 169760 55030 169770
rect 55250 169760 55330 169770
rect 55030 169680 55040 169760
rect 55330 169680 55340 169760
rect 54950 169580 55030 169590
rect 55250 169580 55330 169590
rect 55030 169500 55040 169580
rect 55330 169500 55340 169580
rect 54950 169400 55030 169410
rect 55250 169400 55330 169410
rect 55030 169320 55040 169400
rect 55330 169320 55340 169400
rect 54950 169220 55030 169230
rect 55250 169220 55330 169230
rect 55030 169140 55040 169220
rect 55330 169140 55340 169220
rect 54950 169040 55030 169050
rect 55250 169040 55330 169050
rect 55030 168960 55040 169040
rect 55330 168960 55340 169040
rect 54950 168860 55030 168870
rect 55250 168860 55330 168870
rect 55030 168780 55040 168860
rect 55330 168780 55340 168860
rect 54950 168680 55030 168690
rect 55250 168680 55330 168690
rect 55030 168600 55040 168680
rect 55330 168600 55340 168680
rect 54950 168500 55030 168510
rect 55250 168500 55330 168510
rect 55030 168420 55040 168500
rect 55330 168420 55340 168500
rect 54950 168320 55030 168330
rect 55250 168320 55330 168330
rect 55030 168240 55040 168320
rect 55330 168240 55340 168320
rect 54950 168140 55030 168150
rect 55250 168140 55330 168150
rect 55030 168060 55040 168140
rect 55330 168060 55340 168140
rect 54950 167960 55030 167970
rect 55250 167960 55330 167970
rect 55030 167880 55040 167960
rect 55330 167880 55340 167960
rect 54950 167780 55030 167790
rect 55250 167780 55330 167790
rect 55030 167700 55040 167780
rect 55330 167700 55340 167780
rect 54950 167600 55030 167610
rect 55250 167600 55330 167610
rect 55030 167520 55040 167600
rect 55330 167520 55340 167600
rect 54950 167420 55030 167430
rect 55250 167420 55330 167430
rect 55030 167340 55040 167420
rect 55330 167340 55340 167420
rect 54950 167240 55030 167250
rect 55250 167240 55330 167250
rect 55030 167160 55040 167240
rect 55330 167160 55340 167240
rect 54950 167060 55030 167070
rect 55250 167060 55330 167070
rect 55030 166980 55040 167060
rect 55330 166980 55340 167060
rect 54950 166880 55030 166890
rect 55250 166880 55330 166890
rect 55030 166800 55040 166880
rect 55330 166800 55340 166880
rect 54950 166700 55030 166710
rect 55250 166700 55330 166710
rect 55030 166620 55040 166700
rect 55330 166620 55340 166700
rect 54950 166520 55030 166530
rect 55250 166520 55330 166530
rect 55030 166440 55040 166520
rect 55330 166440 55340 166520
rect 54950 166340 55030 166350
rect 55250 166340 55330 166350
rect 55030 166260 55040 166340
rect 55330 166260 55340 166340
rect 54950 166160 55030 166170
rect 55250 166160 55330 166170
rect 55030 166080 55040 166160
rect 55330 166080 55340 166160
rect 54950 165980 55030 165990
rect 55250 165980 55330 165990
rect 55030 165900 55040 165980
rect 55330 165900 55340 165980
rect 54950 165800 55030 165810
rect 55250 165800 55330 165810
rect 55030 165720 55040 165800
rect 55330 165720 55340 165800
rect 54950 165620 55030 165630
rect 55250 165620 55330 165630
rect 55030 165540 55040 165620
rect 55330 165540 55340 165620
rect 54950 165440 55030 165450
rect 55250 165440 55330 165450
rect 55030 165360 55040 165440
rect 55330 165360 55340 165440
rect 54950 165260 55030 165270
rect 55250 165260 55330 165270
rect 55030 165180 55040 165260
rect 55330 165180 55340 165260
rect 54950 165080 55030 165090
rect 55250 165080 55330 165090
rect 55030 165000 55040 165080
rect 55330 165000 55340 165080
rect 54950 164900 55030 164910
rect 55250 164900 55330 164910
rect 55030 164820 55040 164900
rect 55330 164820 55340 164900
rect 54950 164720 55030 164730
rect 55250 164720 55330 164730
rect 55030 164640 55040 164720
rect 55330 164640 55340 164720
rect 54950 164540 55030 164550
rect 55250 164540 55330 164550
rect 55030 164460 55040 164540
rect 55330 164460 55340 164540
rect 54950 164360 55030 164370
rect 55250 164360 55330 164370
rect 55030 164280 55040 164360
rect 55330 164280 55340 164360
rect 55510 164200 55520 170200
rect 55570 170120 55650 170130
rect 55720 170120 55800 170130
rect 55870 170120 55950 170130
rect 55650 170040 55660 170120
rect 55800 170040 55810 170120
rect 55950 170040 55960 170120
rect 55570 169940 55650 169950
rect 55720 169940 55800 169950
rect 55870 169940 55950 169950
rect 55650 169860 55660 169940
rect 55800 169860 55810 169940
rect 55950 169860 55960 169940
rect 55570 169760 55650 169770
rect 55720 169760 55800 169770
rect 55870 169760 55950 169770
rect 55650 169680 55660 169760
rect 55800 169680 55810 169760
rect 55950 169680 55960 169760
rect 55570 169580 55650 169590
rect 55720 169580 55800 169590
rect 55870 169580 55950 169590
rect 55650 169500 55660 169580
rect 55800 169500 55810 169580
rect 55950 169500 55960 169580
rect 55570 169400 55650 169410
rect 55720 169400 55800 169410
rect 55870 169400 55950 169410
rect 55650 169320 55660 169400
rect 55800 169320 55810 169400
rect 55950 169320 55960 169400
rect 55570 169220 55650 169230
rect 55720 169220 55800 169230
rect 55870 169220 55950 169230
rect 55650 169140 55660 169220
rect 55800 169140 55810 169220
rect 55950 169140 55960 169220
rect 55570 169040 55650 169050
rect 55720 169040 55800 169050
rect 55870 169040 55950 169050
rect 55650 168960 55660 169040
rect 55800 168960 55810 169040
rect 55950 168960 55960 169040
rect 55570 168860 55650 168870
rect 55720 168860 55800 168870
rect 55870 168860 55950 168870
rect 55650 168780 55660 168860
rect 55800 168780 55810 168860
rect 55950 168780 55960 168860
rect 55570 168680 55650 168690
rect 55720 168680 55800 168690
rect 55870 168680 55950 168690
rect 55650 168600 55660 168680
rect 55800 168600 55810 168680
rect 55950 168600 55960 168680
rect 55570 168500 55650 168510
rect 55720 168500 55800 168510
rect 55870 168500 55950 168510
rect 55650 168420 55660 168500
rect 55800 168420 55810 168500
rect 55950 168420 55960 168500
rect 55570 168320 55650 168330
rect 55720 168320 55800 168330
rect 55870 168320 55950 168330
rect 55650 168240 55660 168320
rect 55800 168240 55810 168320
rect 55950 168240 55960 168320
rect 55570 168140 55650 168150
rect 55720 168140 55800 168150
rect 55870 168140 55950 168150
rect 55650 168060 55660 168140
rect 55800 168060 55810 168140
rect 55950 168060 55960 168140
rect 55570 167960 55650 167970
rect 55720 167960 55800 167970
rect 55870 167960 55950 167970
rect 55650 167880 55660 167960
rect 55800 167880 55810 167960
rect 55950 167880 55960 167960
rect 55570 167780 55650 167790
rect 55720 167780 55800 167790
rect 55870 167780 55950 167790
rect 55650 167700 55660 167780
rect 55800 167700 55810 167780
rect 55950 167700 55960 167780
rect 55570 167600 55650 167610
rect 55720 167600 55800 167610
rect 55870 167600 55950 167610
rect 55650 167520 55660 167600
rect 55800 167520 55810 167600
rect 55950 167520 55960 167600
rect 55570 167420 55650 167430
rect 55720 167420 55800 167430
rect 55870 167420 55950 167430
rect 55650 167340 55660 167420
rect 55800 167340 55810 167420
rect 55950 167340 55960 167420
rect 55570 167240 55650 167250
rect 55720 167240 55800 167250
rect 55870 167240 55950 167250
rect 55650 167160 55660 167240
rect 55800 167160 55810 167240
rect 55950 167160 55960 167240
rect 55570 167060 55650 167070
rect 55720 167060 55800 167070
rect 55870 167060 55950 167070
rect 55650 166980 55660 167060
rect 55800 166980 55810 167060
rect 55950 166980 55960 167060
rect 55570 166880 55650 166890
rect 55720 166880 55800 166890
rect 55870 166880 55950 166890
rect 55650 166800 55660 166880
rect 55800 166800 55810 166880
rect 55950 166800 55960 166880
rect 55570 166700 55650 166710
rect 55720 166700 55800 166710
rect 55870 166700 55950 166710
rect 55650 166620 55660 166700
rect 55800 166620 55810 166700
rect 55950 166620 55960 166700
rect 55570 166520 55650 166530
rect 55720 166520 55800 166530
rect 55870 166520 55950 166530
rect 55650 166440 55660 166520
rect 55800 166440 55810 166520
rect 55950 166440 55960 166520
rect 55570 166340 55650 166350
rect 55720 166340 55800 166350
rect 55870 166340 55950 166350
rect 55650 166260 55660 166340
rect 55800 166260 55810 166340
rect 55950 166260 55960 166340
rect 55570 166160 55650 166170
rect 55720 166160 55800 166170
rect 55870 166160 55950 166170
rect 55650 166080 55660 166160
rect 55800 166080 55810 166160
rect 55950 166080 55960 166160
rect 55570 165980 55650 165990
rect 55720 165980 55800 165990
rect 55870 165980 55950 165990
rect 55650 165900 55660 165980
rect 55800 165900 55810 165980
rect 55950 165900 55960 165980
rect 55570 165800 55650 165810
rect 55720 165800 55800 165810
rect 55870 165800 55950 165810
rect 55650 165720 55660 165800
rect 55800 165720 55810 165800
rect 55950 165720 55960 165800
rect 55570 165620 55650 165630
rect 55720 165620 55800 165630
rect 55870 165620 55950 165630
rect 55650 165540 55660 165620
rect 55800 165540 55810 165620
rect 55950 165540 55960 165620
rect 55570 165440 55650 165450
rect 55720 165440 55800 165450
rect 55870 165440 55950 165450
rect 55650 165360 55660 165440
rect 55800 165360 55810 165440
rect 55950 165360 55960 165440
rect 55570 165260 55650 165270
rect 55720 165260 55800 165270
rect 55870 165260 55950 165270
rect 55650 165180 55660 165260
rect 55800 165180 55810 165260
rect 55950 165180 55960 165260
rect 55570 165080 55650 165090
rect 55720 165080 55800 165090
rect 55870 165080 55950 165090
rect 55650 165000 55660 165080
rect 55800 165000 55810 165080
rect 55950 165000 55960 165080
rect 55570 164900 55650 164910
rect 55720 164900 55800 164910
rect 55870 164900 55950 164910
rect 55650 164820 55660 164900
rect 55800 164820 55810 164900
rect 55950 164820 55960 164900
rect 55570 164720 55650 164730
rect 55720 164720 55800 164730
rect 55870 164720 55950 164730
rect 55650 164640 55660 164720
rect 55800 164640 55810 164720
rect 55950 164640 55960 164720
rect 55570 164540 55650 164550
rect 55720 164540 55800 164550
rect 55870 164540 55950 164550
rect 55650 164460 55660 164540
rect 55800 164460 55810 164540
rect 55950 164460 55960 164540
rect 55570 164360 55650 164370
rect 55720 164360 55800 164370
rect 55870 164360 55950 164370
rect 55650 164280 55660 164360
rect 55800 164280 55810 164360
rect 55950 164280 55960 164360
rect 56090 164200 56100 170200
rect 56210 170120 56290 170130
rect 56510 170120 56590 170130
rect 56290 170040 56300 170120
rect 56590 170040 56600 170120
rect 56210 169940 56290 169950
rect 56510 169940 56590 169950
rect 56290 169860 56300 169940
rect 56590 169860 56600 169940
rect 56210 169760 56290 169770
rect 56510 169760 56590 169770
rect 56290 169680 56300 169760
rect 56590 169680 56600 169760
rect 56210 169580 56290 169590
rect 56510 169580 56590 169590
rect 56290 169500 56300 169580
rect 56590 169500 56600 169580
rect 56210 169400 56290 169410
rect 56510 169400 56590 169410
rect 56290 169320 56300 169400
rect 56590 169320 56600 169400
rect 56210 169220 56290 169230
rect 56510 169220 56590 169230
rect 56290 169140 56300 169220
rect 56590 169140 56600 169220
rect 56210 169040 56290 169050
rect 56510 169040 56590 169050
rect 56290 168960 56300 169040
rect 56590 168960 56600 169040
rect 56210 168860 56290 168870
rect 56510 168860 56590 168870
rect 56290 168780 56300 168860
rect 56590 168780 56600 168860
rect 56210 168680 56290 168690
rect 56510 168680 56590 168690
rect 56290 168600 56300 168680
rect 56590 168600 56600 168680
rect 56210 168500 56290 168510
rect 56510 168500 56590 168510
rect 56290 168420 56300 168500
rect 56590 168420 56600 168500
rect 56210 168320 56290 168330
rect 56510 168320 56590 168330
rect 56290 168240 56300 168320
rect 56590 168240 56600 168320
rect 56210 168140 56290 168150
rect 56510 168140 56590 168150
rect 56290 168060 56300 168140
rect 56590 168060 56600 168140
rect 56210 167960 56290 167970
rect 56510 167960 56590 167970
rect 56290 167880 56300 167960
rect 56590 167880 56600 167960
rect 56210 167780 56290 167790
rect 56510 167780 56590 167790
rect 56290 167700 56300 167780
rect 56590 167700 56600 167780
rect 56210 167600 56290 167610
rect 56510 167600 56590 167610
rect 56290 167520 56300 167600
rect 56590 167520 56600 167600
rect 56210 167420 56290 167430
rect 56510 167420 56590 167430
rect 56290 167340 56300 167420
rect 56590 167340 56600 167420
rect 56210 167240 56290 167250
rect 56510 167240 56590 167250
rect 56290 167160 56300 167240
rect 56590 167160 56600 167240
rect 56210 167060 56290 167070
rect 56510 167060 56590 167070
rect 56290 166980 56300 167060
rect 56590 166980 56600 167060
rect 56210 166880 56290 166890
rect 56510 166880 56590 166890
rect 56290 166800 56300 166880
rect 56590 166800 56600 166880
rect 56210 166700 56290 166710
rect 56510 166700 56590 166710
rect 56290 166620 56300 166700
rect 56590 166620 56600 166700
rect 56210 166520 56290 166530
rect 56510 166520 56590 166530
rect 56290 166440 56300 166520
rect 56590 166440 56600 166520
rect 56210 166340 56290 166350
rect 56510 166340 56590 166350
rect 56290 166260 56300 166340
rect 56590 166260 56600 166340
rect 56210 166160 56290 166170
rect 56510 166160 56590 166170
rect 56290 166080 56300 166160
rect 56590 166080 56600 166160
rect 56210 165980 56290 165990
rect 56510 165980 56590 165990
rect 56290 165900 56300 165980
rect 56590 165900 56600 165980
rect 56210 165800 56290 165810
rect 56510 165800 56590 165810
rect 56290 165720 56300 165800
rect 56590 165720 56600 165800
rect 56210 165620 56290 165630
rect 56510 165620 56590 165630
rect 56290 165540 56300 165620
rect 56590 165540 56600 165620
rect 56210 165440 56290 165450
rect 56510 165440 56590 165450
rect 56290 165360 56300 165440
rect 56590 165360 56600 165440
rect 56210 165260 56290 165270
rect 56510 165260 56590 165270
rect 56290 165180 56300 165260
rect 56590 165180 56600 165260
rect 56210 165080 56290 165090
rect 56510 165080 56590 165090
rect 56290 165000 56300 165080
rect 56590 165000 56600 165080
rect 56210 164900 56290 164910
rect 56510 164900 56590 164910
rect 56290 164820 56300 164900
rect 56590 164820 56600 164900
rect 56210 164720 56290 164730
rect 56510 164720 56590 164730
rect 56290 164640 56300 164720
rect 56590 164640 56600 164720
rect 56210 164540 56290 164550
rect 56510 164540 56590 164550
rect 56290 164460 56300 164540
rect 56590 164460 56600 164540
rect 56210 164360 56290 164370
rect 56510 164360 56590 164370
rect 56290 164280 56300 164360
rect 56590 164280 56600 164360
rect 56770 164200 56780 170200
rect 56830 170120 56910 170130
rect 56980 170120 57060 170130
rect 57130 170120 57210 170130
rect 56910 170040 56920 170120
rect 57060 170040 57070 170120
rect 57210 170040 57220 170120
rect 56830 169940 56910 169950
rect 56980 169940 57060 169950
rect 57130 169940 57210 169950
rect 56910 169860 56920 169940
rect 57060 169860 57070 169940
rect 57210 169860 57220 169940
rect 56830 169760 56910 169770
rect 56980 169760 57060 169770
rect 57130 169760 57210 169770
rect 56910 169680 56920 169760
rect 57060 169680 57070 169760
rect 57210 169680 57220 169760
rect 56830 169580 56910 169590
rect 56980 169580 57060 169590
rect 57130 169580 57210 169590
rect 56910 169500 56920 169580
rect 57060 169500 57070 169580
rect 57210 169500 57220 169580
rect 56830 169400 56910 169410
rect 56980 169400 57060 169410
rect 57130 169400 57210 169410
rect 56910 169320 56920 169400
rect 57060 169320 57070 169400
rect 57210 169320 57220 169400
rect 56830 169220 56910 169230
rect 56980 169220 57060 169230
rect 57130 169220 57210 169230
rect 56910 169140 56920 169220
rect 57060 169140 57070 169220
rect 57210 169140 57220 169220
rect 56830 169040 56910 169050
rect 56980 169040 57060 169050
rect 57130 169040 57210 169050
rect 56910 168960 56920 169040
rect 57060 168960 57070 169040
rect 57210 168960 57220 169040
rect 56830 168860 56910 168870
rect 56980 168860 57060 168870
rect 57130 168860 57210 168870
rect 56910 168780 56920 168860
rect 57060 168780 57070 168860
rect 57210 168780 57220 168860
rect 56830 168680 56910 168690
rect 56980 168680 57060 168690
rect 57130 168680 57210 168690
rect 56910 168600 56920 168680
rect 57060 168600 57070 168680
rect 57210 168600 57220 168680
rect 56830 168500 56910 168510
rect 56980 168500 57060 168510
rect 57130 168500 57210 168510
rect 56910 168420 56920 168500
rect 57060 168420 57070 168500
rect 57210 168420 57220 168500
rect 56830 168320 56910 168330
rect 56980 168320 57060 168330
rect 57130 168320 57210 168330
rect 56910 168240 56920 168320
rect 57060 168240 57070 168320
rect 57210 168240 57220 168320
rect 56830 168140 56910 168150
rect 56980 168140 57060 168150
rect 57130 168140 57210 168150
rect 56910 168060 56920 168140
rect 57060 168060 57070 168140
rect 57210 168060 57220 168140
rect 56830 167960 56910 167970
rect 56980 167960 57060 167970
rect 57130 167960 57210 167970
rect 56910 167880 56920 167960
rect 57060 167880 57070 167960
rect 57210 167880 57220 167960
rect 56830 167780 56910 167790
rect 56980 167780 57060 167790
rect 57130 167780 57210 167790
rect 56910 167700 56920 167780
rect 57060 167700 57070 167780
rect 57210 167700 57220 167780
rect 56830 167600 56910 167610
rect 56980 167600 57060 167610
rect 57130 167600 57210 167610
rect 56910 167520 56920 167600
rect 57060 167520 57070 167600
rect 57210 167520 57220 167600
rect 56830 167420 56910 167430
rect 56980 167420 57060 167430
rect 57130 167420 57210 167430
rect 56910 167340 56920 167420
rect 57060 167340 57070 167420
rect 57210 167340 57220 167420
rect 56830 167240 56910 167250
rect 56980 167240 57060 167250
rect 57130 167240 57210 167250
rect 56910 167160 56920 167240
rect 57060 167160 57070 167240
rect 57210 167160 57220 167240
rect 56830 167060 56910 167070
rect 56980 167060 57060 167070
rect 57130 167060 57210 167070
rect 56910 166980 56920 167060
rect 57060 166980 57070 167060
rect 57210 166980 57220 167060
rect 56830 166880 56910 166890
rect 56980 166880 57060 166890
rect 57130 166880 57210 166890
rect 56910 166800 56920 166880
rect 57060 166800 57070 166880
rect 57210 166800 57220 166880
rect 56830 166700 56910 166710
rect 56980 166700 57060 166710
rect 57130 166700 57210 166710
rect 56910 166620 56920 166700
rect 57060 166620 57070 166700
rect 57210 166620 57220 166700
rect 56830 166520 56910 166530
rect 56980 166520 57060 166530
rect 57130 166520 57210 166530
rect 56910 166440 56920 166520
rect 57060 166440 57070 166520
rect 57210 166440 57220 166520
rect 56830 166340 56910 166350
rect 56980 166340 57060 166350
rect 57130 166340 57210 166350
rect 56910 166260 56920 166340
rect 57060 166260 57070 166340
rect 57210 166260 57220 166340
rect 56830 166160 56910 166170
rect 56980 166160 57060 166170
rect 57130 166160 57210 166170
rect 56910 166080 56920 166160
rect 57060 166080 57070 166160
rect 57210 166080 57220 166160
rect 56830 165980 56910 165990
rect 56980 165980 57060 165990
rect 57130 165980 57210 165990
rect 56910 165900 56920 165980
rect 57060 165900 57070 165980
rect 57210 165900 57220 165980
rect 56830 165800 56910 165810
rect 56980 165800 57060 165810
rect 57130 165800 57210 165810
rect 56910 165720 56920 165800
rect 57060 165720 57070 165800
rect 57210 165720 57220 165800
rect 56830 165620 56910 165630
rect 56980 165620 57060 165630
rect 57130 165620 57210 165630
rect 56910 165540 56920 165620
rect 57060 165540 57070 165620
rect 57210 165540 57220 165620
rect 56830 165440 56910 165450
rect 56980 165440 57060 165450
rect 57130 165440 57210 165450
rect 56910 165360 56920 165440
rect 57060 165360 57070 165440
rect 57210 165360 57220 165440
rect 56830 165260 56910 165270
rect 56980 165260 57060 165270
rect 57130 165260 57210 165270
rect 56910 165180 56920 165260
rect 57060 165180 57070 165260
rect 57210 165180 57220 165260
rect 56830 165080 56910 165090
rect 56980 165080 57060 165090
rect 57130 165080 57210 165090
rect 56910 165000 56920 165080
rect 57060 165000 57070 165080
rect 57210 165000 57220 165080
rect 56830 164900 56910 164910
rect 56980 164900 57060 164910
rect 57130 164900 57210 164910
rect 56910 164820 56920 164900
rect 57060 164820 57070 164900
rect 57210 164820 57220 164900
rect 56830 164720 56910 164730
rect 56980 164720 57060 164730
rect 57130 164720 57210 164730
rect 56910 164640 56920 164720
rect 57060 164640 57070 164720
rect 57210 164640 57220 164720
rect 56830 164540 56910 164550
rect 56980 164540 57060 164550
rect 57130 164540 57210 164550
rect 56910 164460 56920 164540
rect 57060 164460 57070 164540
rect 57210 164460 57220 164540
rect 56830 164360 56910 164370
rect 56980 164360 57060 164370
rect 57130 164360 57210 164370
rect 56910 164280 56920 164360
rect 57060 164280 57070 164360
rect 57210 164280 57220 164360
rect 57350 164200 57360 170200
rect 57470 170120 57550 170130
rect 57770 170120 57850 170130
rect 57550 170040 57560 170120
rect 57850 170040 57860 170120
rect 57470 169940 57550 169950
rect 57770 169940 57850 169950
rect 57550 169860 57560 169940
rect 57850 169860 57860 169940
rect 57470 169760 57550 169770
rect 57770 169760 57850 169770
rect 57550 169680 57560 169760
rect 57850 169680 57860 169760
rect 57470 169580 57550 169590
rect 57770 169580 57850 169590
rect 57550 169500 57560 169580
rect 57850 169500 57860 169580
rect 57470 169400 57550 169410
rect 57770 169400 57850 169410
rect 57550 169320 57560 169400
rect 57850 169320 57860 169400
rect 57470 169220 57550 169230
rect 57770 169220 57850 169230
rect 57550 169140 57560 169220
rect 57850 169140 57860 169220
rect 57470 169040 57550 169050
rect 57770 169040 57850 169050
rect 57550 168960 57560 169040
rect 57850 168960 57860 169040
rect 57470 168860 57550 168870
rect 57770 168860 57850 168870
rect 57550 168780 57560 168860
rect 57850 168780 57860 168860
rect 57470 168680 57550 168690
rect 57770 168680 57850 168690
rect 57550 168600 57560 168680
rect 57850 168600 57860 168680
rect 57470 168500 57550 168510
rect 57770 168500 57850 168510
rect 57550 168420 57560 168500
rect 57850 168420 57860 168500
rect 57470 168320 57550 168330
rect 57770 168320 57850 168330
rect 57550 168240 57560 168320
rect 57850 168240 57860 168320
rect 57470 168140 57550 168150
rect 57770 168140 57850 168150
rect 57550 168060 57560 168140
rect 57850 168060 57860 168140
rect 57470 167960 57550 167970
rect 57770 167960 57850 167970
rect 57550 167880 57560 167960
rect 57850 167880 57860 167960
rect 57470 167780 57550 167790
rect 57770 167780 57850 167790
rect 57550 167700 57560 167780
rect 57850 167700 57860 167780
rect 57470 167600 57550 167610
rect 57770 167600 57850 167610
rect 57550 167520 57560 167600
rect 57850 167520 57860 167600
rect 57470 167420 57550 167430
rect 57770 167420 57850 167430
rect 57550 167340 57560 167420
rect 57850 167340 57860 167420
rect 57470 167240 57550 167250
rect 57770 167240 57850 167250
rect 57550 167160 57560 167240
rect 57850 167160 57860 167240
rect 57470 167060 57550 167070
rect 57770 167060 57850 167070
rect 57550 166980 57560 167060
rect 57850 166980 57860 167060
rect 57470 166880 57550 166890
rect 57770 166880 57850 166890
rect 57550 166800 57560 166880
rect 57850 166800 57860 166880
rect 57470 166700 57550 166710
rect 57770 166700 57850 166710
rect 57550 166620 57560 166700
rect 57850 166620 57860 166700
rect 57470 166520 57550 166530
rect 57770 166520 57850 166530
rect 57550 166440 57560 166520
rect 57850 166440 57860 166520
rect 57470 166340 57550 166350
rect 57770 166340 57850 166350
rect 57550 166260 57560 166340
rect 57850 166260 57860 166340
rect 57470 166160 57550 166170
rect 57770 166160 57850 166170
rect 57550 166080 57560 166160
rect 57850 166080 57860 166160
rect 57470 165980 57550 165990
rect 57770 165980 57850 165990
rect 57550 165900 57560 165980
rect 57850 165900 57860 165980
rect 57470 165800 57550 165810
rect 57770 165800 57850 165810
rect 57550 165720 57560 165800
rect 57850 165720 57860 165800
rect 57470 165620 57550 165630
rect 57770 165620 57850 165630
rect 57550 165540 57560 165620
rect 57850 165540 57860 165620
rect 57470 165440 57550 165450
rect 57770 165440 57850 165450
rect 57550 165360 57560 165440
rect 57850 165360 57860 165440
rect 57470 165260 57550 165270
rect 57770 165260 57850 165270
rect 57550 165180 57560 165260
rect 57850 165180 57860 165260
rect 57470 165080 57550 165090
rect 57770 165080 57850 165090
rect 57550 165000 57560 165080
rect 57850 165000 57860 165080
rect 57470 164900 57550 164910
rect 57770 164900 57850 164910
rect 57550 164820 57560 164900
rect 57850 164820 57860 164900
rect 57470 164720 57550 164730
rect 57770 164720 57850 164730
rect 57550 164640 57560 164720
rect 57850 164640 57860 164720
rect 57470 164540 57550 164550
rect 57770 164540 57850 164550
rect 57550 164460 57560 164540
rect 57850 164460 57860 164540
rect 57470 164360 57550 164370
rect 57770 164360 57850 164370
rect 57550 164280 57560 164360
rect 57850 164280 57860 164360
rect 58030 164200 58040 170200
rect 58090 170120 58170 170130
rect 58240 170120 58320 170130
rect 58390 170120 58470 170130
rect 58170 170040 58180 170120
rect 58320 170040 58330 170120
rect 58470 170040 58480 170120
rect 58090 169940 58170 169950
rect 58240 169940 58320 169950
rect 58390 169940 58470 169950
rect 58170 169860 58180 169940
rect 58320 169860 58330 169940
rect 58470 169860 58480 169940
rect 58090 169760 58170 169770
rect 58240 169760 58320 169770
rect 58390 169760 58470 169770
rect 58170 169680 58180 169760
rect 58320 169680 58330 169760
rect 58470 169680 58480 169760
rect 58090 169580 58170 169590
rect 58240 169580 58320 169590
rect 58390 169580 58470 169590
rect 58170 169500 58180 169580
rect 58320 169500 58330 169580
rect 58470 169500 58480 169580
rect 58090 169400 58170 169410
rect 58240 169400 58320 169410
rect 58390 169400 58470 169410
rect 58170 169320 58180 169400
rect 58320 169320 58330 169400
rect 58470 169320 58480 169400
rect 58090 169220 58170 169230
rect 58240 169220 58320 169230
rect 58390 169220 58470 169230
rect 58170 169140 58180 169220
rect 58320 169140 58330 169220
rect 58470 169140 58480 169220
rect 58090 169040 58170 169050
rect 58240 169040 58320 169050
rect 58390 169040 58470 169050
rect 58170 168960 58180 169040
rect 58320 168960 58330 169040
rect 58470 168960 58480 169040
rect 58090 168860 58170 168870
rect 58240 168860 58320 168870
rect 58390 168860 58470 168870
rect 58170 168780 58180 168860
rect 58320 168780 58330 168860
rect 58470 168780 58480 168860
rect 58090 168680 58170 168690
rect 58240 168680 58320 168690
rect 58390 168680 58470 168690
rect 58170 168600 58180 168680
rect 58320 168600 58330 168680
rect 58470 168600 58480 168680
rect 58090 168500 58170 168510
rect 58240 168500 58320 168510
rect 58390 168500 58470 168510
rect 58170 168420 58180 168500
rect 58320 168420 58330 168500
rect 58470 168420 58480 168500
rect 58090 168320 58170 168330
rect 58240 168320 58320 168330
rect 58390 168320 58470 168330
rect 58170 168240 58180 168320
rect 58320 168240 58330 168320
rect 58470 168240 58480 168320
rect 58090 168140 58170 168150
rect 58240 168140 58320 168150
rect 58390 168140 58470 168150
rect 58170 168060 58180 168140
rect 58320 168060 58330 168140
rect 58470 168060 58480 168140
rect 58090 167960 58170 167970
rect 58240 167960 58320 167970
rect 58390 167960 58470 167970
rect 58170 167880 58180 167960
rect 58320 167880 58330 167960
rect 58470 167880 58480 167960
rect 58090 167780 58170 167790
rect 58240 167780 58320 167790
rect 58390 167780 58470 167790
rect 58170 167700 58180 167780
rect 58320 167700 58330 167780
rect 58470 167700 58480 167780
rect 58090 167600 58170 167610
rect 58240 167600 58320 167610
rect 58390 167600 58470 167610
rect 58170 167520 58180 167600
rect 58320 167520 58330 167600
rect 58470 167520 58480 167600
rect 58090 167420 58170 167430
rect 58240 167420 58320 167430
rect 58390 167420 58470 167430
rect 58170 167340 58180 167420
rect 58320 167340 58330 167420
rect 58470 167340 58480 167420
rect 58090 167240 58170 167250
rect 58240 167240 58320 167250
rect 58390 167240 58470 167250
rect 58170 167160 58180 167240
rect 58320 167160 58330 167240
rect 58470 167160 58480 167240
rect 58090 167060 58170 167070
rect 58240 167060 58320 167070
rect 58390 167060 58470 167070
rect 58170 166980 58180 167060
rect 58320 166980 58330 167060
rect 58470 166980 58480 167060
rect 58090 166880 58170 166890
rect 58240 166880 58320 166890
rect 58390 166880 58470 166890
rect 58170 166800 58180 166880
rect 58320 166800 58330 166880
rect 58470 166800 58480 166880
rect 58090 166700 58170 166710
rect 58240 166700 58320 166710
rect 58390 166700 58470 166710
rect 58170 166620 58180 166700
rect 58320 166620 58330 166700
rect 58470 166620 58480 166700
rect 58090 166520 58170 166530
rect 58240 166520 58320 166530
rect 58390 166520 58470 166530
rect 58170 166440 58180 166520
rect 58320 166440 58330 166520
rect 58470 166440 58480 166520
rect 58090 166340 58170 166350
rect 58240 166340 58320 166350
rect 58390 166340 58470 166350
rect 58170 166260 58180 166340
rect 58320 166260 58330 166340
rect 58470 166260 58480 166340
rect 58090 166160 58170 166170
rect 58240 166160 58320 166170
rect 58390 166160 58470 166170
rect 58170 166080 58180 166160
rect 58320 166080 58330 166160
rect 58470 166080 58480 166160
rect 58090 165980 58170 165990
rect 58240 165980 58320 165990
rect 58390 165980 58470 165990
rect 58170 165900 58180 165980
rect 58320 165900 58330 165980
rect 58470 165900 58480 165980
rect 58090 165800 58170 165810
rect 58240 165800 58320 165810
rect 58390 165800 58470 165810
rect 58170 165720 58180 165800
rect 58320 165720 58330 165800
rect 58470 165720 58480 165800
rect 58090 165620 58170 165630
rect 58240 165620 58320 165630
rect 58390 165620 58470 165630
rect 58170 165540 58180 165620
rect 58320 165540 58330 165620
rect 58470 165540 58480 165620
rect 58090 165440 58170 165450
rect 58240 165440 58320 165450
rect 58390 165440 58470 165450
rect 58170 165360 58180 165440
rect 58320 165360 58330 165440
rect 58470 165360 58480 165440
rect 58090 165260 58170 165270
rect 58240 165260 58320 165270
rect 58390 165260 58470 165270
rect 58170 165180 58180 165260
rect 58320 165180 58330 165260
rect 58470 165180 58480 165260
rect 58090 165080 58170 165090
rect 58240 165080 58320 165090
rect 58390 165080 58470 165090
rect 58170 165000 58180 165080
rect 58320 165000 58330 165080
rect 58470 165000 58480 165080
rect 58090 164900 58170 164910
rect 58240 164900 58320 164910
rect 58390 164900 58470 164910
rect 58170 164820 58180 164900
rect 58320 164820 58330 164900
rect 58470 164820 58480 164900
rect 58090 164720 58170 164730
rect 58240 164720 58320 164730
rect 58390 164720 58470 164730
rect 58170 164640 58180 164720
rect 58320 164640 58330 164720
rect 58470 164640 58480 164720
rect 58090 164540 58170 164550
rect 58240 164540 58320 164550
rect 58390 164540 58470 164550
rect 58170 164460 58180 164540
rect 58320 164460 58330 164540
rect 58470 164460 58480 164540
rect 58090 164360 58170 164370
rect 58240 164360 58320 164370
rect 58390 164360 58470 164370
rect 58170 164280 58180 164360
rect 58320 164280 58330 164360
rect 58470 164280 58480 164360
rect 58610 164200 58620 170200
rect 58730 170120 58810 170130
rect 59030 170120 59110 170130
rect 58810 170040 58820 170120
rect 59110 170040 59120 170120
rect 58730 169940 58810 169950
rect 59030 169940 59110 169950
rect 58810 169860 58820 169940
rect 59110 169860 59120 169940
rect 58730 169760 58810 169770
rect 59030 169760 59110 169770
rect 58810 169680 58820 169760
rect 59110 169680 59120 169760
rect 58730 169580 58810 169590
rect 59030 169580 59110 169590
rect 58810 169500 58820 169580
rect 59110 169500 59120 169580
rect 58730 169400 58810 169410
rect 59030 169400 59110 169410
rect 58810 169320 58820 169400
rect 59110 169320 59120 169400
rect 58730 169220 58810 169230
rect 59030 169220 59110 169230
rect 58810 169140 58820 169220
rect 59110 169140 59120 169220
rect 58730 169040 58810 169050
rect 59030 169040 59110 169050
rect 58810 168960 58820 169040
rect 59110 168960 59120 169040
rect 58730 168860 58810 168870
rect 59030 168860 59110 168870
rect 58810 168780 58820 168860
rect 59110 168780 59120 168860
rect 58730 168680 58810 168690
rect 59030 168680 59110 168690
rect 58810 168600 58820 168680
rect 59110 168600 59120 168680
rect 58730 168500 58810 168510
rect 59030 168500 59110 168510
rect 58810 168420 58820 168500
rect 59110 168420 59120 168500
rect 58730 168320 58810 168330
rect 59030 168320 59110 168330
rect 58810 168240 58820 168320
rect 59110 168240 59120 168320
rect 58730 168140 58810 168150
rect 59030 168140 59110 168150
rect 58810 168060 58820 168140
rect 59110 168060 59120 168140
rect 58730 167960 58810 167970
rect 59030 167960 59110 167970
rect 58810 167880 58820 167960
rect 59110 167880 59120 167960
rect 58730 167780 58810 167790
rect 59030 167780 59110 167790
rect 58810 167700 58820 167780
rect 59110 167700 59120 167780
rect 58730 167600 58810 167610
rect 59030 167600 59110 167610
rect 58810 167520 58820 167600
rect 59110 167520 59120 167600
rect 58730 167420 58810 167430
rect 59030 167420 59110 167430
rect 58810 167340 58820 167420
rect 59110 167340 59120 167420
rect 58730 167240 58810 167250
rect 59030 167240 59110 167250
rect 58810 167160 58820 167240
rect 59110 167160 59120 167240
rect 58730 167060 58810 167070
rect 59030 167060 59110 167070
rect 58810 166980 58820 167060
rect 59110 166980 59120 167060
rect 58730 166880 58810 166890
rect 59030 166880 59110 166890
rect 58810 166800 58820 166880
rect 59110 166800 59120 166880
rect 58730 166700 58810 166710
rect 59030 166700 59110 166710
rect 58810 166620 58820 166700
rect 59110 166620 59120 166700
rect 58730 166520 58810 166530
rect 59030 166520 59110 166530
rect 58810 166440 58820 166520
rect 59110 166440 59120 166520
rect 58730 166340 58810 166350
rect 59030 166340 59110 166350
rect 58810 166260 58820 166340
rect 59110 166260 59120 166340
rect 58730 166160 58810 166170
rect 59030 166160 59110 166170
rect 58810 166080 58820 166160
rect 59110 166080 59120 166160
rect 58730 165980 58810 165990
rect 59030 165980 59110 165990
rect 58810 165900 58820 165980
rect 59110 165900 59120 165980
rect 58730 165800 58810 165810
rect 59030 165800 59110 165810
rect 58810 165720 58820 165800
rect 59110 165720 59120 165800
rect 58730 165620 58810 165630
rect 59030 165620 59110 165630
rect 58810 165540 58820 165620
rect 59110 165540 59120 165620
rect 58730 165440 58810 165450
rect 59030 165440 59110 165450
rect 58810 165360 58820 165440
rect 59110 165360 59120 165440
rect 58730 165260 58810 165270
rect 59030 165260 59110 165270
rect 58810 165180 58820 165260
rect 59110 165180 59120 165260
rect 58730 165080 58810 165090
rect 59030 165080 59110 165090
rect 58810 165000 58820 165080
rect 59110 165000 59120 165080
rect 58730 164900 58810 164910
rect 59030 164900 59110 164910
rect 58810 164820 58820 164900
rect 59110 164820 59120 164900
rect 58730 164720 58810 164730
rect 59030 164720 59110 164730
rect 58810 164640 58820 164720
rect 59110 164640 59120 164720
rect 58730 164540 58810 164550
rect 59030 164540 59110 164550
rect 58810 164460 58820 164540
rect 59110 164460 59120 164540
rect 58730 164360 58810 164370
rect 59030 164360 59110 164370
rect 58810 164280 58820 164360
rect 59110 164280 59120 164360
rect 59290 164200 59300 170200
rect 60850 170149 60860 170229
rect 61170 170149 61180 170229
rect 61590 170149 61600 170229
rect 61910 170149 61920 170229
rect 62140 170220 62150 170300
rect 62290 170220 62300 170300
rect 73640 170220 73650 170300
rect 73790 170220 73800 170300
rect 73940 170220 73950 170300
rect 74270 170229 74350 170239
rect 74590 170229 74670 170239
rect 75010 170229 75090 170239
rect 75330 170229 75410 170239
rect 74350 170149 74360 170229
rect 74670 170149 74680 170229
rect 75090 170149 75100 170229
rect 75410 170149 75420 170229
rect 75640 170220 75650 170300
rect 75790 170220 75800 170300
rect 87140 170220 87150 170300
rect 87290 170220 87300 170300
rect 87440 170220 87450 170300
rect 87770 170229 87850 170239
rect 88090 170229 88170 170239
rect 88510 170229 88590 170239
rect 88830 170229 88910 170239
rect 87850 170149 87860 170229
rect 88170 170149 88180 170229
rect 88590 170149 88600 170229
rect 88910 170149 88920 170229
rect 89140 170220 89150 170300
rect 89290 170220 89300 170300
rect 100640 170220 100650 170300
rect 100790 170220 100800 170300
rect 100940 170220 100950 170300
rect 101270 170229 101350 170239
rect 101590 170229 101670 170239
rect 102010 170229 102090 170239
rect 102330 170229 102410 170239
rect 114770 170229 114850 170239
rect 115090 170229 115170 170239
rect 115510 170229 115590 170239
rect 115830 170229 115910 170239
rect 101350 170149 101360 170229
rect 101670 170149 101680 170229
rect 102090 170149 102100 170229
rect 102410 170149 102420 170229
rect 114850 170149 114860 170229
rect 115170 170149 115180 170229
rect 115590 170149 115600 170229
rect 115910 170149 115920 170229
rect 116140 170220 116150 170300
rect 116290 170220 116300 170300
rect 127640 170220 127650 170300
rect 127790 170220 127800 170300
rect 127940 170220 127950 170300
rect 128270 170229 128350 170239
rect 128590 170229 128670 170239
rect 129010 170229 129090 170239
rect 129330 170229 129410 170239
rect 128350 170149 128360 170229
rect 128670 170149 128680 170229
rect 129090 170149 129100 170229
rect 129410 170149 129420 170229
rect 129640 170220 129650 170300
rect 129790 170220 129800 170300
rect 141140 170220 141150 170300
rect 141290 170220 141300 170300
rect 141440 170220 141450 170300
rect 141665 170230 141745 170240
rect 141985 170230 142065 170240
rect 145200 170230 145265 170240
rect 145505 170230 145585 170240
rect 145825 170230 145905 170240
rect 141745 170150 141755 170230
rect 142065 170150 142075 170230
rect 145265 170150 145275 170230
rect 145585 170150 145595 170230
rect 145905 170150 145915 170230
rect 146620 170220 146630 170300
rect 146940 170220 146950 170300
rect 146700 170140 146780 170150
rect 59350 170120 59430 170130
rect 59500 170120 59580 170130
rect 59650 170120 59730 170130
rect 60060 170120 60140 170130
rect 60210 170120 60290 170130
rect 60360 170120 60440 170130
rect 62060 170120 62140 170130
rect 62210 170120 62290 170130
rect 73560 170120 73640 170130
rect 73710 170120 73790 170130
rect 73860 170120 73940 170130
rect 75560 170120 75640 170130
rect 75710 170120 75790 170130
rect 87060 170120 87140 170130
rect 87210 170120 87290 170130
rect 87360 170120 87440 170130
rect 89060 170120 89140 170130
rect 89210 170120 89290 170130
rect 100560 170120 100640 170130
rect 100710 170120 100790 170130
rect 100860 170120 100940 170130
rect 116060 170120 116140 170130
rect 116210 170120 116290 170130
rect 127560 170120 127640 170130
rect 127710 170120 127790 170130
rect 127860 170120 127940 170130
rect 129560 170120 129640 170130
rect 129710 170120 129790 170130
rect 140710 170120 140730 170130
rect 141060 170120 141140 170130
rect 141210 170120 141290 170130
rect 141360 170120 141440 170130
rect 59430 170040 59440 170120
rect 59580 170040 59590 170120
rect 59730 170040 59740 170120
rect 60140 170040 60150 170120
rect 60290 170040 60300 170120
rect 60440 170040 60450 170120
rect 60610 170069 60690 170079
rect 60930 170069 61010 170079
rect 61350 170069 61430 170079
rect 61670 170069 61750 170079
rect 60690 169989 60700 170069
rect 61010 169989 61020 170069
rect 61430 169989 61440 170069
rect 61750 169989 61760 170069
rect 62140 170040 62150 170120
rect 62290 170040 62300 170120
rect 73640 170040 73650 170120
rect 73790 170040 73800 170120
rect 73940 170040 73950 170120
rect 74110 170069 74190 170079
rect 74430 170069 74510 170079
rect 74850 170069 74930 170079
rect 75170 170069 75250 170079
rect 74190 169989 74200 170069
rect 74510 169989 74520 170069
rect 74930 169989 74940 170069
rect 75250 169989 75260 170069
rect 75640 170040 75650 170120
rect 75790 170040 75800 170120
rect 87140 170040 87150 170120
rect 87290 170040 87300 170120
rect 87440 170040 87450 170120
rect 87610 170069 87690 170079
rect 87930 170069 88010 170079
rect 88350 170069 88430 170079
rect 88670 170069 88750 170079
rect 87690 169989 87700 170069
rect 88010 169989 88020 170069
rect 88430 169989 88440 170069
rect 88750 169989 88760 170069
rect 89140 170040 89150 170120
rect 89290 170040 89300 170120
rect 100640 170040 100650 170120
rect 100790 170040 100800 170120
rect 100940 170040 100950 170120
rect 101110 170069 101190 170079
rect 101430 170069 101510 170079
rect 101850 170069 101930 170079
rect 102170 170069 102250 170079
rect 114610 170069 114690 170079
rect 114930 170069 115010 170079
rect 115350 170069 115430 170079
rect 115670 170069 115750 170079
rect 101190 169989 101200 170069
rect 101510 169989 101520 170069
rect 101930 169989 101940 170069
rect 102250 169989 102260 170069
rect 114690 169989 114700 170069
rect 115010 169989 115020 170069
rect 115430 169989 115440 170069
rect 115750 169989 115760 170069
rect 116140 170040 116150 170120
rect 116290 170040 116300 170120
rect 127640 170040 127650 170120
rect 127790 170040 127800 170120
rect 127940 170040 127950 170120
rect 128110 170069 128190 170079
rect 128430 170069 128510 170079
rect 128850 170069 128930 170079
rect 129170 170069 129250 170079
rect 128190 169989 128200 170069
rect 128510 169989 128520 170069
rect 128930 169989 128940 170069
rect 129250 169989 129260 170069
rect 129640 170040 129650 170120
rect 129790 170040 129800 170120
rect 140730 170040 140740 170120
rect 141140 170040 141150 170120
rect 141290 170040 141300 170120
rect 141440 170040 141450 170120
rect 141825 170070 141905 170080
rect 142145 170070 142200 170080
rect 145345 170070 145425 170080
rect 145665 170070 145745 170080
rect 145985 170070 146065 170080
rect 141905 169990 141915 170070
rect 145425 169990 145435 170070
rect 145745 169990 145755 170070
rect 146065 169990 146075 170070
rect 146780 170060 146790 170140
rect 146540 169980 146620 169990
rect 146860 169980 146940 169990
rect 59350 169940 59430 169950
rect 59500 169940 59580 169950
rect 59650 169940 59730 169950
rect 60060 169940 60140 169950
rect 60210 169940 60290 169950
rect 60360 169940 60440 169950
rect 62060 169940 62140 169950
rect 62210 169940 62290 169950
rect 73560 169940 73640 169950
rect 73710 169940 73790 169950
rect 73860 169940 73940 169950
rect 75560 169940 75640 169950
rect 75710 169940 75790 169950
rect 87060 169940 87140 169950
rect 87210 169940 87290 169950
rect 87360 169940 87440 169950
rect 89060 169940 89140 169950
rect 89210 169940 89290 169950
rect 100560 169940 100640 169950
rect 100710 169940 100790 169950
rect 100860 169940 100940 169950
rect 116060 169940 116140 169950
rect 116210 169940 116290 169950
rect 127560 169940 127640 169950
rect 127710 169940 127790 169950
rect 127860 169940 127940 169950
rect 129560 169940 129640 169950
rect 129710 169940 129790 169950
rect 140710 169940 140730 169950
rect 141060 169940 141140 169950
rect 141210 169940 141290 169950
rect 141360 169940 141440 169950
rect 59430 169860 59440 169940
rect 59580 169860 59590 169940
rect 59730 169860 59740 169940
rect 60140 169860 60150 169940
rect 60290 169860 60300 169940
rect 60440 169860 60450 169940
rect 60770 169909 60850 169919
rect 61090 169909 61170 169919
rect 61510 169909 61590 169919
rect 61830 169909 61910 169919
rect 60850 169829 60860 169909
rect 61170 169829 61180 169909
rect 61590 169829 61600 169909
rect 61910 169829 61920 169909
rect 62140 169860 62150 169940
rect 62290 169860 62300 169940
rect 73640 169860 73650 169940
rect 73790 169860 73800 169940
rect 73940 169860 73950 169940
rect 74270 169909 74350 169919
rect 74590 169909 74670 169919
rect 75010 169909 75090 169919
rect 75330 169909 75410 169919
rect 74350 169829 74360 169909
rect 74670 169829 74680 169909
rect 75090 169829 75100 169909
rect 75410 169829 75420 169909
rect 75640 169860 75650 169940
rect 75790 169860 75800 169940
rect 87140 169860 87150 169940
rect 87290 169860 87300 169940
rect 87440 169860 87450 169940
rect 87770 169909 87850 169919
rect 88090 169909 88170 169919
rect 88510 169909 88590 169919
rect 88830 169909 88910 169919
rect 87850 169829 87860 169909
rect 88170 169829 88180 169909
rect 88590 169829 88600 169909
rect 88910 169829 88920 169909
rect 89140 169860 89150 169940
rect 89290 169860 89300 169940
rect 100640 169860 100650 169940
rect 100790 169860 100800 169940
rect 100940 169860 100950 169940
rect 101270 169909 101350 169919
rect 101590 169909 101670 169919
rect 102010 169909 102090 169919
rect 102330 169909 102410 169919
rect 114770 169909 114850 169919
rect 115090 169909 115170 169919
rect 115510 169909 115590 169919
rect 115830 169909 115910 169919
rect 101350 169829 101360 169909
rect 101670 169829 101680 169909
rect 102090 169829 102100 169909
rect 102410 169829 102420 169909
rect 114850 169829 114860 169909
rect 115170 169829 115180 169909
rect 115590 169829 115600 169909
rect 115910 169829 115920 169909
rect 116140 169860 116150 169940
rect 116290 169860 116300 169940
rect 127640 169860 127650 169940
rect 127790 169860 127800 169940
rect 127940 169860 127950 169940
rect 128270 169909 128350 169919
rect 128590 169909 128670 169919
rect 129010 169909 129090 169919
rect 129330 169909 129410 169919
rect 128350 169829 128360 169909
rect 128670 169829 128680 169909
rect 129090 169829 129100 169909
rect 129410 169829 129420 169909
rect 129640 169860 129650 169940
rect 129790 169860 129800 169940
rect 140730 169860 140740 169940
rect 141140 169860 141150 169940
rect 141290 169860 141300 169940
rect 141440 169860 141450 169940
rect 141665 169910 141745 169920
rect 141985 169910 142065 169920
rect 145200 169910 145265 169920
rect 145505 169910 145585 169920
rect 145825 169910 145905 169920
rect 141745 169830 141755 169910
rect 142065 169830 142075 169910
rect 145265 169830 145275 169910
rect 145585 169830 145595 169910
rect 145905 169830 145915 169910
rect 146620 169900 146630 169980
rect 146940 169900 146950 169980
rect 146700 169820 146780 169830
rect 59350 169760 59430 169770
rect 59500 169760 59580 169770
rect 59650 169760 59730 169770
rect 60060 169760 60140 169770
rect 60210 169760 60290 169770
rect 60360 169760 60440 169770
rect 62060 169760 62140 169770
rect 62210 169760 62290 169770
rect 73560 169760 73640 169770
rect 73710 169760 73790 169770
rect 73860 169760 73940 169770
rect 75560 169760 75640 169770
rect 75710 169760 75790 169770
rect 87060 169760 87140 169770
rect 87210 169760 87290 169770
rect 87360 169760 87440 169770
rect 89060 169760 89140 169770
rect 89210 169760 89290 169770
rect 100560 169760 100640 169770
rect 100710 169760 100790 169770
rect 100860 169760 100940 169770
rect 116060 169760 116140 169770
rect 116210 169760 116290 169770
rect 127560 169760 127640 169770
rect 127710 169760 127790 169770
rect 127860 169760 127940 169770
rect 129560 169760 129640 169770
rect 129710 169760 129790 169770
rect 140710 169760 140730 169770
rect 141060 169760 141140 169770
rect 141210 169760 141290 169770
rect 141360 169760 141440 169770
rect 59430 169680 59440 169760
rect 59580 169680 59590 169760
rect 59730 169680 59740 169760
rect 60140 169680 60150 169760
rect 60290 169680 60300 169760
rect 60440 169680 60450 169760
rect 60610 169749 60690 169759
rect 60930 169749 61010 169759
rect 61350 169749 61430 169759
rect 61670 169749 61750 169759
rect 60690 169669 60700 169749
rect 61010 169669 61020 169749
rect 61430 169669 61440 169749
rect 61750 169669 61760 169749
rect 62140 169680 62150 169760
rect 62290 169680 62300 169760
rect 73640 169680 73650 169760
rect 73790 169680 73800 169760
rect 73940 169680 73950 169760
rect 74110 169749 74190 169759
rect 74430 169749 74510 169759
rect 74850 169749 74930 169759
rect 75170 169749 75250 169759
rect 74190 169669 74200 169749
rect 74510 169669 74520 169749
rect 74930 169669 74940 169749
rect 75250 169669 75260 169749
rect 75640 169680 75650 169760
rect 75790 169680 75800 169760
rect 87140 169680 87150 169760
rect 87290 169680 87300 169760
rect 87440 169680 87450 169760
rect 87610 169749 87690 169759
rect 87930 169749 88010 169759
rect 88350 169749 88430 169759
rect 88670 169749 88750 169759
rect 87690 169669 87700 169749
rect 88010 169669 88020 169749
rect 88430 169669 88440 169749
rect 88750 169669 88760 169749
rect 89140 169680 89150 169760
rect 89290 169680 89300 169760
rect 100640 169680 100650 169760
rect 100790 169680 100800 169760
rect 100940 169680 100950 169760
rect 101110 169749 101190 169759
rect 101430 169749 101510 169759
rect 101850 169749 101930 169759
rect 102170 169749 102250 169759
rect 114610 169749 114690 169759
rect 114930 169749 115010 169759
rect 115350 169749 115430 169759
rect 115670 169749 115750 169759
rect 101190 169669 101200 169749
rect 101510 169669 101520 169749
rect 101930 169669 101940 169749
rect 102250 169669 102260 169749
rect 114690 169669 114700 169749
rect 115010 169669 115020 169749
rect 115430 169669 115440 169749
rect 115750 169669 115760 169749
rect 116140 169680 116150 169760
rect 116290 169680 116300 169760
rect 127640 169680 127650 169760
rect 127790 169680 127800 169760
rect 127940 169680 127950 169760
rect 128110 169749 128190 169759
rect 128430 169749 128510 169759
rect 128850 169749 128930 169759
rect 129170 169749 129250 169759
rect 128190 169669 128200 169749
rect 128510 169669 128520 169749
rect 128930 169669 128940 169749
rect 129250 169669 129260 169749
rect 129640 169680 129650 169760
rect 129790 169680 129800 169760
rect 140730 169680 140740 169760
rect 141140 169680 141150 169760
rect 141290 169680 141300 169760
rect 141440 169680 141450 169760
rect 141825 169750 141905 169760
rect 142145 169750 142200 169760
rect 145345 169750 145425 169760
rect 145665 169750 145745 169760
rect 145985 169750 146065 169760
rect 141905 169670 141915 169750
rect 145425 169670 145435 169750
rect 145745 169670 145755 169750
rect 146065 169670 146075 169750
rect 146780 169740 146790 169820
rect 146540 169660 146620 169670
rect 146860 169660 146940 169670
rect 59350 169580 59430 169590
rect 59500 169580 59580 169590
rect 59650 169580 59730 169590
rect 60060 169580 60140 169590
rect 60210 169580 60290 169590
rect 60360 169580 60440 169590
rect 60770 169589 60850 169599
rect 61090 169589 61170 169599
rect 61510 169589 61590 169599
rect 61830 169589 61910 169599
rect 59430 169500 59440 169580
rect 59580 169500 59590 169580
rect 59730 169500 59740 169580
rect 60140 169500 60150 169580
rect 60290 169500 60300 169580
rect 60440 169500 60450 169580
rect 60850 169509 60860 169589
rect 61170 169509 61180 169589
rect 61590 169509 61600 169589
rect 61910 169509 61920 169589
rect 62060 169580 62140 169590
rect 62210 169580 62290 169590
rect 73560 169580 73640 169590
rect 73710 169580 73790 169590
rect 73860 169580 73940 169590
rect 74270 169589 74350 169599
rect 74590 169589 74670 169599
rect 75010 169589 75090 169599
rect 75330 169589 75410 169599
rect 62140 169500 62150 169580
rect 62290 169500 62300 169580
rect 73640 169500 73650 169580
rect 73790 169500 73800 169580
rect 73940 169500 73950 169580
rect 74350 169509 74360 169589
rect 74670 169509 74680 169589
rect 75090 169509 75100 169589
rect 75410 169509 75420 169589
rect 75560 169580 75640 169590
rect 75710 169580 75790 169590
rect 87060 169580 87140 169590
rect 87210 169580 87290 169590
rect 87360 169580 87440 169590
rect 87770 169589 87850 169599
rect 88090 169589 88170 169599
rect 88510 169589 88590 169599
rect 88830 169589 88910 169599
rect 75640 169500 75650 169580
rect 75790 169500 75800 169580
rect 87140 169500 87150 169580
rect 87290 169500 87300 169580
rect 87440 169500 87450 169580
rect 87850 169509 87860 169589
rect 88170 169509 88180 169589
rect 88590 169509 88600 169589
rect 88910 169509 88920 169589
rect 89060 169580 89140 169590
rect 89210 169580 89290 169590
rect 100560 169580 100640 169590
rect 100710 169580 100790 169590
rect 100860 169580 100940 169590
rect 101270 169589 101350 169599
rect 101590 169589 101670 169599
rect 102010 169589 102090 169599
rect 102330 169589 102410 169599
rect 114770 169589 114850 169599
rect 115090 169589 115170 169599
rect 115510 169589 115590 169599
rect 115830 169589 115910 169599
rect 89140 169500 89150 169580
rect 89290 169500 89300 169580
rect 100640 169500 100650 169580
rect 100790 169500 100800 169580
rect 100940 169500 100950 169580
rect 101350 169509 101360 169589
rect 101670 169509 101680 169589
rect 102090 169509 102100 169589
rect 102410 169509 102420 169589
rect 114850 169509 114860 169589
rect 115170 169509 115180 169589
rect 115590 169509 115600 169589
rect 115910 169509 115920 169589
rect 116060 169580 116140 169590
rect 116210 169580 116290 169590
rect 127560 169580 127640 169590
rect 127710 169580 127790 169590
rect 127860 169580 127940 169590
rect 128270 169589 128350 169599
rect 128590 169589 128670 169599
rect 129010 169589 129090 169599
rect 129330 169589 129410 169599
rect 141665 169590 141745 169600
rect 141985 169590 142065 169600
rect 145200 169590 145265 169600
rect 145505 169590 145585 169600
rect 145825 169590 145905 169600
rect 116140 169500 116150 169580
rect 116290 169500 116300 169580
rect 127640 169500 127650 169580
rect 127790 169500 127800 169580
rect 127940 169500 127950 169580
rect 128350 169509 128360 169589
rect 128670 169509 128680 169589
rect 129090 169509 129100 169589
rect 129410 169509 129420 169589
rect 129560 169580 129640 169590
rect 129710 169580 129790 169590
rect 140710 169580 140730 169590
rect 141060 169580 141140 169590
rect 141210 169580 141290 169590
rect 141360 169580 141440 169590
rect 129640 169500 129650 169580
rect 129790 169500 129800 169580
rect 140730 169500 140740 169580
rect 141140 169500 141150 169580
rect 141290 169500 141300 169580
rect 141440 169500 141450 169580
rect 141745 169510 141755 169590
rect 142065 169510 142075 169590
rect 145265 169510 145275 169590
rect 145585 169510 145595 169590
rect 145905 169510 145915 169590
rect 146620 169580 146630 169660
rect 146940 169580 146950 169660
rect 146700 169500 146780 169510
rect 60610 169429 60690 169439
rect 60930 169429 61010 169439
rect 61350 169429 61430 169439
rect 61670 169429 61750 169439
rect 74110 169429 74190 169439
rect 74430 169429 74510 169439
rect 74850 169429 74930 169439
rect 75170 169429 75250 169439
rect 87610 169429 87690 169439
rect 87930 169429 88010 169439
rect 88350 169429 88430 169439
rect 88670 169429 88750 169439
rect 101110 169429 101190 169439
rect 101430 169429 101510 169439
rect 101850 169429 101930 169439
rect 102170 169429 102250 169439
rect 114610 169429 114690 169439
rect 114930 169429 115010 169439
rect 115350 169429 115430 169439
rect 115670 169429 115750 169439
rect 128110 169429 128190 169439
rect 128430 169429 128510 169439
rect 128850 169429 128930 169439
rect 129170 169429 129250 169439
rect 141825 169430 141905 169440
rect 142145 169430 142200 169440
rect 145345 169430 145425 169440
rect 145665 169430 145745 169440
rect 145985 169430 146065 169440
rect 59350 169400 59430 169410
rect 59500 169400 59580 169410
rect 59650 169400 59730 169410
rect 60060 169400 60140 169410
rect 60210 169400 60290 169410
rect 60360 169400 60440 169410
rect 59430 169320 59440 169400
rect 59580 169320 59590 169400
rect 59730 169320 59740 169400
rect 60140 169320 60150 169400
rect 60290 169320 60300 169400
rect 60440 169320 60450 169400
rect 60690 169349 60700 169429
rect 61010 169349 61020 169429
rect 61430 169349 61440 169429
rect 61750 169349 61760 169429
rect 62060 169400 62140 169410
rect 62210 169400 62290 169410
rect 73560 169400 73640 169410
rect 73710 169400 73790 169410
rect 73860 169400 73940 169410
rect 62140 169320 62150 169400
rect 62290 169320 62300 169400
rect 73640 169320 73650 169400
rect 73790 169320 73800 169400
rect 73940 169320 73950 169400
rect 74190 169349 74200 169429
rect 74510 169349 74520 169429
rect 74930 169349 74940 169429
rect 75250 169349 75260 169429
rect 75560 169400 75640 169410
rect 75710 169400 75790 169410
rect 87060 169400 87140 169410
rect 87210 169400 87290 169410
rect 87360 169400 87440 169410
rect 75640 169320 75650 169400
rect 75790 169320 75800 169400
rect 87140 169320 87150 169400
rect 87290 169320 87300 169400
rect 87440 169320 87450 169400
rect 87690 169349 87700 169429
rect 88010 169349 88020 169429
rect 88430 169349 88440 169429
rect 88750 169349 88760 169429
rect 89060 169400 89140 169410
rect 89210 169400 89290 169410
rect 100560 169400 100640 169410
rect 100710 169400 100790 169410
rect 100860 169400 100940 169410
rect 89140 169320 89150 169400
rect 89290 169320 89300 169400
rect 100640 169320 100650 169400
rect 100790 169320 100800 169400
rect 100940 169320 100950 169400
rect 101190 169349 101200 169429
rect 101510 169349 101520 169429
rect 101930 169349 101940 169429
rect 102250 169349 102260 169429
rect 114690 169349 114700 169429
rect 115010 169349 115020 169429
rect 115430 169349 115440 169429
rect 115750 169349 115760 169429
rect 116060 169400 116140 169410
rect 116210 169400 116290 169410
rect 127560 169400 127640 169410
rect 127710 169400 127790 169410
rect 127860 169400 127940 169410
rect 116140 169320 116150 169400
rect 116290 169320 116300 169400
rect 127640 169320 127650 169400
rect 127790 169320 127800 169400
rect 127940 169320 127950 169400
rect 128190 169349 128200 169429
rect 128510 169349 128520 169429
rect 128930 169349 128940 169429
rect 129250 169349 129260 169429
rect 129560 169400 129640 169410
rect 129710 169400 129790 169410
rect 140710 169400 140730 169410
rect 141060 169400 141140 169410
rect 141210 169400 141290 169410
rect 141360 169400 141440 169410
rect 129640 169320 129650 169400
rect 129790 169320 129800 169400
rect 140730 169320 140740 169400
rect 141140 169320 141150 169400
rect 141290 169320 141300 169400
rect 141440 169320 141450 169400
rect 141905 169350 141915 169430
rect 145425 169350 145435 169430
rect 145745 169350 145755 169430
rect 146065 169350 146075 169430
rect 146780 169420 146790 169500
rect 146540 169340 146620 169350
rect 146860 169340 146940 169350
rect 60770 169269 60850 169279
rect 61090 169269 61170 169279
rect 61510 169269 61590 169279
rect 61830 169269 61910 169279
rect 74270 169269 74350 169279
rect 74590 169269 74670 169279
rect 75010 169269 75090 169279
rect 75330 169269 75410 169279
rect 87770 169269 87850 169279
rect 88090 169269 88170 169279
rect 88510 169269 88590 169279
rect 88830 169269 88910 169279
rect 101270 169269 101350 169279
rect 101590 169269 101670 169279
rect 102010 169269 102090 169279
rect 102330 169269 102410 169279
rect 114770 169269 114850 169279
rect 115090 169269 115170 169279
rect 115510 169269 115590 169279
rect 115830 169269 115910 169279
rect 128270 169269 128350 169279
rect 128590 169269 128670 169279
rect 129010 169269 129090 169279
rect 129330 169269 129410 169279
rect 141665 169270 141745 169280
rect 141985 169270 142065 169280
rect 145200 169270 145265 169280
rect 145505 169270 145585 169280
rect 145825 169270 145905 169280
rect 59350 169220 59430 169230
rect 59500 169220 59580 169230
rect 59650 169220 59730 169230
rect 60060 169220 60140 169230
rect 60210 169220 60290 169230
rect 60360 169220 60440 169230
rect 59430 169140 59440 169220
rect 59580 169140 59590 169220
rect 59730 169140 59740 169220
rect 60140 169140 60150 169220
rect 60290 169140 60300 169220
rect 60440 169140 60450 169220
rect 60850 169189 60860 169269
rect 61170 169189 61180 169269
rect 61590 169189 61600 169269
rect 61910 169189 61920 169269
rect 62060 169220 62140 169230
rect 62210 169220 62290 169230
rect 73560 169220 73640 169230
rect 73710 169220 73790 169230
rect 73860 169220 73940 169230
rect 62140 169140 62150 169220
rect 62290 169140 62300 169220
rect 73640 169140 73650 169220
rect 73790 169140 73800 169220
rect 73940 169140 73950 169220
rect 74350 169189 74360 169269
rect 74670 169189 74680 169269
rect 75090 169189 75100 169269
rect 75410 169189 75420 169269
rect 75560 169220 75640 169230
rect 75710 169220 75790 169230
rect 87060 169220 87140 169230
rect 87210 169220 87290 169230
rect 87360 169220 87440 169230
rect 75640 169140 75650 169220
rect 75790 169140 75800 169220
rect 87140 169140 87150 169220
rect 87290 169140 87300 169220
rect 87440 169140 87450 169220
rect 87850 169189 87860 169269
rect 88170 169189 88180 169269
rect 88590 169189 88600 169269
rect 88910 169189 88920 169269
rect 89060 169220 89140 169230
rect 89210 169220 89290 169230
rect 100560 169220 100640 169230
rect 100710 169220 100790 169230
rect 100860 169220 100940 169230
rect 89140 169140 89150 169220
rect 89290 169140 89300 169220
rect 100640 169140 100650 169220
rect 100790 169140 100800 169220
rect 100940 169140 100950 169220
rect 101350 169189 101360 169269
rect 101670 169189 101680 169269
rect 102090 169189 102100 169269
rect 102410 169189 102420 169269
rect 114850 169189 114860 169269
rect 115170 169189 115180 169269
rect 115590 169189 115600 169269
rect 115910 169189 115920 169269
rect 116060 169220 116140 169230
rect 116210 169220 116290 169230
rect 127560 169220 127640 169230
rect 127710 169220 127790 169230
rect 127860 169220 127940 169230
rect 116140 169140 116150 169220
rect 116290 169140 116300 169220
rect 127640 169140 127650 169220
rect 127790 169140 127800 169220
rect 127940 169140 127950 169220
rect 128350 169189 128360 169269
rect 128670 169189 128680 169269
rect 129090 169189 129100 169269
rect 129410 169189 129420 169269
rect 129560 169220 129640 169230
rect 129710 169220 129790 169230
rect 140710 169220 140730 169230
rect 141060 169220 141140 169230
rect 141210 169220 141290 169230
rect 141360 169220 141440 169230
rect 129640 169140 129650 169220
rect 129790 169140 129800 169220
rect 140730 169140 140740 169220
rect 141140 169140 141150 169220
rect 141290 169140 141300 169220
rect 141440 169140 141450 169220
rect 141745 169190 141755 169270
rect 142065 169190 142075 169270
rect 145265 169190 145275 169270
rect 145585 169190 145595 169270
rect 145905 169190 145915 169270
rect 146620 169260 146630 169340
rect 146940 169260 146950 169340
rect 146700 169180 146780 169190
rect 60610 169109 60690 169119
rect 60930 169109 61010 169119
rect 61350 169109 61430 169119
rect 61670 169109 61750 169119
rect 74110 169109 74190 169119
rect 74430 169109 74510 169119
rect 74850 169109 74930 169119
rect 75170 169109 75250 169119
rect 87610 169109 87690 169119
rect 87930 169109 88010 169119
rect 88350 169109 88430 169119
rect 88670 169109 88750 169119
rect 101110 169109 101190 169119
rect 101430 169109 101510 169119
rect 101850 169109 101930 169119
rect 102170 169109 102250 169119
rect 114610 169109 114690 169119
rect 114930 169109 115010 169119
rect 115350 169109 115430 169119
rect 115670 169109 115750 169119
rect 128110 169109 128190 169119
rect 128430 169109 128510 169119
rect 128850 169109 128930 169119
rect 129170 169109 129250 169119
rect 141825 169110 141905 169120
rect 142145 169110 142200 169120
rect 145345 169110 145425 169120
rect 145665 169110 145745 169120
rect 145985 169110 146065 169120
rect 59350 169040 59430 169050
rect 59500 169040 59580 169050
rect 59650 169040 59730 169050
rect 60060 169040 60140 169050
rect 60210 169040 60290 169050
rect 60360 169040 60440 169050
rect 59430 168960 59440 169040
rect 59580 168960 59590 169040
rect 59730 168960 59740 169040
rect 60140 168960 60150 169040
rect 60290 168960 60300 169040
rect 60440 168960 60450 169040
rect 60690 169029 60700 169109
rect 61010 169029 61020 169109
rect 61430 169029 61440 169109
rect 61750 169029 61760 169109
rect 62060 169040 62140 169050
rect 62210 169040 62290 169050
rect 73560 169040 73640 169050
rect 73710 169040 73790 169050
rect 73860 169040 73940 169050
rect 62140 168960 62150 169040
rect 62290 168960 62300 169040
rect 73640 168960 73650 169040
rect 73790 168960 73800 169040
rect 73940 168960 73950 169040
rect 74190 169029 74200 169109
rect 74510 169029 74520 169109
rect 74930 169029 74940 169109
rect 75250 169029 75260 169109
rect 75560 169040 75640 169050
rect 75710 169040 75790 169050
rect 87060 169040 87140 169050
rect 87210 169040 87290 169050
rect 87360 169040 87440 169050
rect 75640 168960 75650 169040
rect 75790 168960 75800 169040
rect 87140 168960 87150 169040
rect 87290 168960 87300 169040
rect 87440 168960 87450 169040
rect 87690 169029 87700 169109
rect 88010 169029 88020 169109
rect 88430 169029 88440 169109
rect 88750 169029 88760 169109
rect 89060 169040 89140 169050
rect 89210 169040 89290 169050
rect 100560 169040 100640 169050
rect 100710 169040 100790 169050
rect 100860 169040 100940 169050
rect 89140 168960 89150 169040
rect 89290 168960 89300 169040
rect 100640 168960 100650 169040
rect 100790 168960 100800 169040
rect 100940 168960 100950 169040
rect 101190 169029 101200 169109
rect 101510 169029 101520 169109
rect 101930 169029 101940 169109
rect 102250 169029 102260 169109
rect 114690 169029 114700 169109
rect 115010 169029 115020 169109
rect 115430 169029 115440 169109
rect 115750 169029 115760 169109
rect 116060 169040 116140 169050
rect 116210 169040 116290 169050
rect 127560 169040 127640 169050
rect 127710 169040 127790 169050
rect 127860 169040 127940 169050
rect 116140 168960 116150 169040
rect 116290 168960 116300 169040
rect 127640 168960 127650 169040
rect 127790 168960 127800 169040
rect 127940 168960 127950 169040
rect 128190 169029 128200 169109
rect 128510 169029 128520 169109
rect 128930 169029 128940 169109
rect 129250 169029 129260 169109
rect 129560 169040 129640 169050
rect 129710 169040 129790 169050
rect 140710 169040 140730 169050
rect 141060 169040 141140 169050
rect 141210 169040 141290 169050
rect 141360 169040 141440 169050
rect 129640 168960 129650 169040
rect 129790 168960 129800 169040
rect 140730 168960 140740 169040
rect 141140 168960 141150 169040
rect 141290 168960 141300 169040
rect 141440 168960 141450 169040
rect 141905 169030 141915 169110
rect 145425 169030 145435 169110
rect 145745 169030 145755 169110
rect 146065 169030 146075 169110
rect 146780 169100 146790 169180
rect 146540 169020 146620 169030
rect 146860 169020 146940 169030
rect 60770 168949 60850 168959
rect 61090 168949 61170 168959
rect 61510 168949 61590 168959
rect 61830 168949 61910 168959
rect 74270 168949 74350 168959
rect 74590 168949 74670 168959
rect 75010 168949 75090 168959
rect 75330 168949 75410 168959
rect 87770 168949 87850 168959
rect 88090 168949 88170 168959
rect 88510 168949 88590 168959
rect 88830 168949 88910 168959
rect 101270 168949 101350 168959
rect 101590 168949 101670 168959
rect 102010 168949 102090 168959
rect 102330 168949 102410 168959
rect 114770 168949 114850 168959
rect 115090 168949 115170 168959
rect 115510 168949 115590 168959
rect 115830 168949 115910 168959
rect 128270 168949 128350 168959
rect 128590 168949 128670 168959
rect 129010 168949 129090 168959
rect 129330 168949 129410 168959
rect 141665 168950 141745 168960
rect 141985 168950 142065 168960
rect 145200 168950 145265 168960
rect 145505 168950 145585 168960
rect 145825 168950 145905 168960
rect 59350 168860 59430 168870
rect 59500 168860 59580 168870
rect 59650 168860 59730 168870
rect 60060 168860 60140 168870
rect 60210 168860 60290 168870
rect 60360 168860 60440 168870
rect 60850 168869 60860 168949
rect 61170 168869 61180 168949
rect 61590 168869 61600 168949
rect 61910 168869 61920 168949
rect 62060 168860 62140 168870
rect 62210 168860 62290 168870
rect 73560 168860 73640 168870
rect 73710 168860 73790 168870
rect 73860 168860 73940 168870
rect 74350 168869 74360 168949
rect 74670 168869 74680 168949
rect 75090 168869 75100 168949
rect 75410 168869 75420 168949
rect 75560 168860 75640 168870
rect 75710 168860 75790 168870
rect 87060 168860 87140 168870
rect 87210 168860 87290 168870
rect 87360 168860 87440 168870
rect 87850 168869 87860 168949
rect 88170 168869 88180 168949
rect 88590 168869 88600 168949
rect 88910 168869 88920 168949
rect 89060 168860 89140 168870
rect 89210 168860 89290 168870
rect 100560 168860 100640 168870
rect 100710 168860 100790 168870
rect 100860 168860 100940 168870
rect 101350 168869 101360 168949
rect 101670 168869 101680 168949
rect 102090 168869 102100 168949
rect 102410 168869 102420 168949
rect 114850 168869 114860 168949
rect 115170 168869 115180 168949
rect 115590 168869 115600 168949
rect 115910 168869 115920 168949
rect 116060 168860 116140 168870
rect 116210 168860 116290 168870
rect 127560 168860 127640 168870
rect 127710 168860 127790 168870
rect 127860 168860 127940 168870
rect 128350 168869 128360 168949
rect 128670 168869 128680 168949
rect 129090 168869 129100 168949
rect 129410 168869 129420 168949
rect 141745 168870 141755 168950
rect 142065 168870 142075 168950
rect 145265 168870 145275 168950
rect 145585 168870 145595 168950
rect 145905 168870 145915 168950
rect 146620 168940 146630 169020
rect 146940 168940 146950 169020
rect 129560 168860 129640 168870
rect 129710 168860 129790 168870
rect 140710 168860 140730 168870
rect 141060 168860 141140 168870
rect 141210 168860 141290 168870
rect 141360 168860 141440 168870
rect 146700 168860 146780 168870
rect 59430 168780 59440 168860
rect 59580 168780 59590 168860
rect 59730 168780 59740 168860
rect 60140 168780 60150 168860
rect 60290 168780 60300 168860
rect 60440 168780 60450 168860
rect 60610 168789 60690 168799
rect 60930 168789 61010 168799
rect 61350 168789 61430 168799
rect 61670 168789 61750 168799
rect 60690 168709 60700 168789
rect 61010 168709 61020 168789
rect 61430 168709 61440 168789
rect 61750 168709 61760 168789
rect 62140 168780 62150 168860
rect 62290 168780 62300 168860
rect 73640 168780 73650 168860
rect 73790 168780 73800 168860
rect 73940 168780 73950 168860
rect 74110 168789 74190 168799
rect 74430 168789 74510 168799
rect 74850 168789 74930 168799
rect 75170 168789 75250 168799
rect 74190 168709 74200 168789
rect 74510 168709 74520 168789
rect 74930 168709 74940 168789
rect 75250 168709 75260 168789
rect 75640 168780 75650 168860
rect 75790 168780 75800 168860
rect 87140 168780 87150 168860
rect 87290 168780 87300 168860
rect 87440 168780 87450 168860
rect 87610 168789 87690 168799
rect 87930 168789 88010 168799
rect 88350 168789 88430 168799
rect 88670 168789 88750 168799
rect 87690 168709 87700 168789
rect 88010 168709 88020 168789
rect 88430 168709 88440 168789
rect 88750 168709 88760 168789
rect 89140 168780 89150 168860
rect 89290 168780 89300 168860
rect 100640 168780 100650 168860
rect 100790 168780 100800 168860
rect 100940 168780 100950 168860
rect 101110 168789 101190 168799
rect 101430 168789 101510 168799
rect 101850 168789 101930 168799
rect 102170 168789 102250 168799
rect 114610 168789 114690 168799
rect 114930 168789 115010 168799
rect 115350 168789 115430 168799
rect 115670 168789 115750 168799
rect 101190 168709 101200 168789
rect 101510 168709 101520 168789
rect 101930 168709 101940 168789
rect 102250 168709 102260 168789
rect 114690 168709 114700 168789
rect 115010 168709 115020 168789
rect 115430 168709 115440 168789
rect 115750 168709 115760 168789
rect 116140 168780 116150 168860
rect 116290 168780 116300 168860
rect 127640 168780 127650 168860
rect 127790 168780 127800 168860
rect 127940 168780 127950 168860
rect 128110 168789 128190 168799
rect 128430 168789 128510 168799
rect 128850 168789 128930 168799
rect 129170 168789 129250 168799
rect 128190 168709 128200 168789
rect 128510 168709 128520 168789
rect 128930 168709 128940 168789
rect 129250 168709 129260 168789
rect 129640 168780 129650 168860
rect 129790 168780 129800 168860
rect 140730 168780 140740 168860
rect 141140 168780 141150 168860
rect 141290 168780 141300 168860
rect 141440 168780 141450 168860
rect 141825 168790 141905 168800
rect 142145 168790 142200 168800
rect 145345 168790 145425 168800
rect 145665 168790 145745 168800
rect 145985 168790 146065 168800
rect 141905 168710 141915 168790
rect 145425 168710 145435 168790
rect 145745 168710 145755 168790
rect 146065 168710 146075 168790
rect 146780 168780 146790 168860
rect 146540 168700 146620 168710
rect 146860 168700 146940 168710
rect 59350 168680 59430 168690
rect 59500 168680 59580 168690
rect 59650 168680 59730 168690
rect 60060 168680 60140 168690
rect 60210 168680 60290 168690
rect 60360 168680 60440 168690
rect 62060 168680 62140 168690
rect 62210 168680 62290 168690
rect 73560 168680 73640 168690
rect 73710 168680 73790 168690
rect 73860 168680 73940 168690
rect 75560 168680 75640 168690
rect 75710 168680 75790 168690
rect 87060 168680 87140 168690
rect 87210 168680 87290 168690
rect 87360 168680 87440 168690
rect 89060 168680 89140 168690
rect 89210 168680 89290 168690
rect 100560 168680 100640 168690
rect 100710 168680 100790 168690
rect 100860 168680 100940 168690
rect 116060 168680 116140 168690
rect 116210 168680 116290 168690
rect 127560 168680 127640 168690
rect 127710 168680 127790 168690
rect 127860 168680 127940 168690
rect 129560 168680 129640 168690
rect 129710 168680 129790 168690
rect 140710 168680 140730 168690
rect 141060 168680 141140 168690
rect 141210 168680 141290 168690
rect 141360 168680 141440 168690
rect 59430 168600 59440 168680
rect 59580 168600 59590 168680
rect 59730 168600 59740 168680
rect 60140 168600 60150 168680
rect 60290 168600 60300 168680
rect 60440 168600 60450 168680
rect 60770 168629 60850 168639
rect 61090 168629 61170 168639
rect 61510 168629 61590 168639
rect 61830 168629 61910 168639
rect 60850 168549 60860 168629
rect 61170 168549 61180 168629
rect 61590 168549 61600 168629
rect 61910 168549 61920 168629
rect 62140 168600 62150 168680
rect 62290 168600 62300 168680
rect 73640 168600 73650 168680
rect 73790 168600 73800 168680
rect 73940 168600 73950 168680
rect 74270 168629 74350 168639
rect 74590 168629 74670 168639
rect 75010 168629 75090 168639
rect 75330 168629 75410 168639
rect 74350 168549 74360 168629
rect 74670 168549 74680 168629
rect 75090 168549 75100 168629
rect 75410 168549 75420 168629
rect 75640 168600 75650 168680
rect 75790 168600 75800 168680
rect 87140 168600 87150 168680
rect 87290 168600 87300 168680
rect 87440 168600 87450 168680
rect 87770 168629 87850 168639
rect 88090 168629 88170 168639
rect 88510 168629 88590 168639
rect 88830 168629 88910 168639
rect 87850 168549 87860 168629
rect 88170 168549 88180 168629
rect 88590 168549 88600 168629
rect 88910 168549 88920 168629
rect 89140 168600 89150 168680
rect 89290 168600 89300 168680
rect 100640 168600 100650 168680
rect 100790 168600 100800 168680
rect 100940 168600 100950 168680
rect 101270 168629 101350 168639
rect 101590 168629 101670 168639
rect 102010 168629 102090 168639
rect 102330 168629 102410 168639
rect 114770 168629 114850 168639
rect 115090 168629 115170 168639
rect 115510 168629 115590 168639
rect 115830 168629 115910 168639
rect 101350 168549 101360 168629
rect 101670 168549 101680 168629
rect 102090 168549 102100 168629
rect 102410 168549 102420 168629
rect 114850 168549 114860 168629
rect 115170 168549 115180 168629
rect 115590 168549 115600 168629
rect 115910 168549 115920 168629
rect 116140 168600 116150 168680
rect 116290 168600 116300 168680
rect 127640 168600 127650 168680
rect 127790 168600 127800 168680
rect 127940 168600 127950 168680
rect 128270 168629 128350 168639
rect 128590 168629 128670 168639
rect 129010 168629 129090 168639
rect 129330 168629 129410 168639
rect 128350 168549 128360 168629
rect 128670 168549 128680 168629
rect 129090 168549 129100 168629
rect 129410 168549 129420 168629
rect 129640 168600 129650 168680
rect 129790 168600 129800 168680
rect 140730 168600 140740 168680
rect 141140 168600 141150 168680
rect 141290 168600 141300 168680
rect 141440 168600 141450 168680
rect 141665 168630 141745 168640
rect 141985 168630 142065 168640
rect 145200 168630 145265 168640
rect 145505 168630 145585 168640
rect 145825 168630 145905 168640
rect 141745 168550 141755 168630
rect 142065 168550 142075 168630
rect 145265 168550 145275 168630
rect 145585 168550 145595 168630
rect 145905 168550 145915 168630
rect 146620 168620 146630 168700
rect 146940 168620 146950 168700
rect 146700 168540 146780 168550
rect 59350 168500 59430 168510
rect 59500 168500 59580 168510
rect 59650 168500 59730 168510
rect 60060 168500 60140 168510
rect 60210 168500 60290 168510
rect 60360 168500 60440 168510
rect 62060 168500 62140 168510
rect 62210 168500 62290 168510
rect 73560 168500 73640 168510
rect 73710 168500 73790 168510
rect 73860 168500 73940 168510
rect 75560 168500 75640 168510
rect 75710 168500 75790 168510
rect 87060 168500 87140 168510
rect 87210 168500 87290 168510
rect 87360 168500 87440 168510
rect 89060 168500 89140 168510
rect 89210 168500 89290 168510
rect 100560 168500 100640 168510
rect 100710 168500 100790 168510
rect 100860 168500 100940 168510
rect 116060 168500 116140 168510
rect 116210 168500 116290 168510
rect 127560 168500 127640 168510
rect 127710 168500 127790 168510
rect 127860 168500 127940 168510
rect 129560 168500 129640 168510
rect 129710 168500 129790 168510
rect 140710 168500 140730 168510
rect 141060 168500 141140 168510
rect 141210 168500 141290 168510
rect 141360 168500 141440 168510
rect 59430 168420 59440 168500
rect 59580 168420 59590 168500
rect 59730 168420 59740 168500
rect 60140 168420 60150 168500
rect 60290 168420 60300 168500
rect 60440 168420 60450 168500
rect 60610 168469 60690 168479
rect 60930 168469 61010 168479
rect 61350 168469 61430 168479
rect 61670 168469 61750 168479
rect 60690 168389 60700 168469
rect 61010 168389 61020 168469
rect 61430 168389 61440 168469
rect 61750 168389 61760 168469
rect 62140 168420 62150 168500
rect 62290 168420 62300 168500
rect 73640 168420 73650 168500
rect 73790 168420 73800 168500
rect 73940 168420 73950 168500
rect 74110 168469 74190 168479
rect 74430 168469 74510 168479
rect 74850 168469 74930 168479
rect 75170 168469 75250 168479
rect 74190 168389 74200 168469
rect 74510 168389 74520 168469
rect 74930 168389 74940 168469
rect 75250 168389 75260 168469
rect 75640 168420 75650 168500
rect 75790 168420 75800 168500
rect 87140 168420 87150 168500
rect 87290 168420 87300 168500
rect 87440 168420 87450 168500
rect 87610 168469 87690 168479
rect 87930 168469 88010 168479
rect 88350 168469 88430 168479
rect 88670 168469 88750 168479
rect 87690 168389 87700 168469
rect 88010 168389 88020 168469
rect 88430 168389 88440 168469
rect 88750 168389 88760 168469
rect 89140 168420 89150 168500
rect 89290 168420 89300 168500
rect 100640 168420 100650 168500
rect 100790 168420 100800 168500
rect 100940 168420 100950 168500
rect 101110 168469 101190 168479
rect 101430 168469 101510 168479
rect 101850 168469 101930 168479
rect 102170 168469 102250 168479
rect 114610 168469 114690 168479
rect 114930 168469 115010 168479
rect 115350 168469 115430 168479
rect 115670 168469 115750 168479
rect 101190 168389 101200 168469
rect 101510 168389 101520 168469
rect 101930 168389 101940 168469
rect 102250 168389 102260 168469
rect 114690 168389 114700 168469
rect 115010 168389 115020 168469
rect 115430 168389 115440 168469
rect 115750 168389 115760 168469
rect 116140 168420 116150 168500
rect 116290 168420 116300 168500
rect 127640 168420 127650 168500
rect 127790 168420 127800 168500
rect 127940 168420 127950 168500
rect 128110 168469 128190 168479
rect 128430 168469 128510 168479
rect 128850 168469 128930 168479
rect 129170 168469 129250 168479
rect 128190 168389 128200 168469
rect 128510 168389 128520 168469
rect 128930 168389 128940 168469
rect 129250 168389 129260 168469
rect 129640 168420 129650 168500
rect 129790 168420 129800 168500
rect 140730 168420 140740 168500
rect 141140 168420 141150 168500
rect 141290 168420 141300 168500
rect 141440 168420 141450 168500
rect 141825 168470 141905 168480
rect 142145 168470 142200 168480
rect 145345 168470 145425 168480
rect 145665 168470 145745 168480
rect 145985 168470 146065 168480
rect 141905 168390 141915 168470
rect 145425 168390 145435 168470
rect 145745 168390 145755 168470
rect 146065 168390 146075 168470
rect 146780 168460 146790 168540
rect 146540 168380 146620 168390
rect 146860 168380 146940 168390
rect 59350 168320 59430 168330
rect 59500 168320 59580 168330
rect 59650 168320 59730 168330
rect 60060 168320 60140 168330
rect 60210 168320 60290 168330
rect 60360 168320 60440 168330
rect 62060 168320 62140 168330
rect 62210 168320 62290 168330
rect 73560 168320 73640 168330
rect 73710 168320 73790 168330
rect 73860 168320 73940 168330
rect 75560 168320 75640 168330
rect 75710 168320 75790 168330
rect 87060 168320 87140 168330
rect 87210 168320 87290 168330
rect 87360 168320 87440 168330
rect 89060 168320 89140 168330
rect 89210 168320 89290 168330
rect 100560 168320 100640 168330
rect 100710 168320 100790 168330
rect 100860 168320 100940 168330
rect 116060 168320 116140 168330
rect 116210 168320 116290 168330
rect 127560 168320 127640 168330
rect 127710 168320 127790 168330
rect 127860 168320 127940 168330
rect 129560 168320 129640 168330
rect 129710 168320 129790 168330
rect 140710 168320 140730 168330
rect 141060 168320 141140 168330
rect 141210 168320 141290 168330
rect 141360 168320 141440 168330
rect 59430 168240 59440 168320
rect 59580 168240 59590 168320
rect 59730 168240 59740 168320
rect 60140 168240 60150 168320
rect 60290 168240 60300 168320
rect 60440 168240 60450 168320
rect 60770 168309 60850 168319
rect 61090 168309 61170 168319
rect 61510 168309 61590 168319
rect 61830 168309 61910 168319
rect 60850 168229 60860 168309
rect 61170 168229 61180 168309
rect 61590 168229 61600 168309
rect 61910 168229 61920 168309
rect 62140 168240 62150 168320
rect 62290 168240 62300 168320
rect 73640 168240 73650 168320
rect 73790 168240 73800 168320
rect 73940 168240 73950 168320
rect 74270 168309 74350 168319
rect 74590 168309 74670 168319
rect 75010 168309 75090 168319
rect 75330 168309 75410 168319
rect 74350 168229 74360 168309
rect 74670 168229 74680 168309
rect 75090 168229 75100 168309
rect 75410 168229 75420 168309
rect 75640 168240 75650 168320
rect 75790 168240 75800 168320
rect 87140 168240 87150 168320
rect 87290 168240 87300 168320
rect 87440 168240 87450 168320
rect 87770 168309 87850 168319
rect 88090 168309 88170 168319
rect 88510 168309 88590 168319
rect 88830 168309 88910 168319
rect 87850 168229 87860 168309
rect 88170 168229 88180 168309
rect 88590 168229 88600 168309
rect 88910 168229 88920 168309
rect 89140 168240 89150 168320
rect 89290 168240 89300 168320
rect 100640 168240 100650 168320
rect 100790 168240 100800 168320
rect 100940 168240 100950 168320
rect 101270 168309 101350 168319
rect 101590 168309 101670 168319
rect 102010 168309 102090 168319
rect 102330 168309 102410 168319
rect 114770 168309 114850 168319
rect 115090 168309 115170 168319
rect 115510 168309 115590 168319
rect 115830 168309 115910 168319
rect 101350 168229 101360 168309
rect 101670 168229 101680 168309
rect 102090 168229 102100 168309
rect 102410 168229 102420 168309
rect 114850 168229 114860 168309
rect 115170 168229 115180 168309
rect 115590 168229 115600 168309
rect 115910 168229 115920 168309
rect 116140 168240 116150 168320
rect 116290 168240 116300 168320
rect 127640 168240 127650 168320
rect 127790 168240 127800 168320
rect 127940 168240 127950 168320
rect 128270 168309 128350 168319
rect 128590 168309 128670 168319
rect 129010 168309 129090 168319
rect 129330 168309 129410 168319
rect 128350 168229 128360 168309
rect 128670 168229 128680 168309
rect 129090 168229 129100 168309
rect 129410 168229 129420 168309
rect 129640 168240 129650 168320
rect 129790 168240 129800 168320
rect 140730 168240 140740 168320
rect 141140 168240 141150 168320
rect 141290 168240 141300 168320
rect 141440 168240 141450 168320
rect 141665 168310 141745 168320
rect 141985 168310 142065 168320
rect 145200 168310 145265 168320
rect 145505 168310 145585 168320
rect 145825 168310 145905 168320
rect 141745 168230 141755 168310
rect 142065 168230 142075 168310
rect 145265 168230 145275 168310
rect 145585 168230 145595 168310
rect 145905 168230 145915 168310
rect 146620 168300 146630 168380
rect 146940 168300 146950 168380
rect 146700 168220 146780 168230
rect 59350 168140 59430 168150
rect 59500 168140 59580 168150
rect 59650 168140 59730 168150
rect 60060 168140 60140 168150
rect 60210 168140 60290 168150
rect 60360 168140 60440 168150
rect 60610 168149 60690 168159
rect 60930 168149 61010 168159
rect 61350 168149 61430 168159
rect 61670 168149 61750 168159
rect 59430 168060 59440 168140
rect 59580 168060 59590 168140
rect 59730 168060 59740 168140
rect 60140 168060 60150 168140
rect 60290 168060 60300 168140
rect 60440 168060 60450 168140
rect 60690 168069 60700 168149
rect 61010 168069 61020 168149
rect 61430 168069 61440 168149
rect 61750 168069 61760 168149
rect 62060 168140 62140 168150
rect 62210 168140 62290 168150
rect 73560 168140 73640 168150
rect 73710 168140 73790 168150
rect 73860 168140 73940 168150
rect 74110 168149 74190 168159
rect 74430 168149 74510 168159
rect 74850 168149 74930 168159
rect 75170 168149 75250 168159
rect 62140 168060 62150 168140
rect 62290 168060 62300 168140
rect 73640 168060 73650 168140
rect 73790 168060 73800 168140
rect 73940 168060 73950 168140
rect 74190 168069 74200 168149
rect 74510 168069 74520 168149
rect 74930 168069 74940 168149
rect 75250 168069 75260 168149
rect 75560 168140 75640 168150
rect 75710 168140 75790 168150
rect 87060 168140 87140 168150
rect 87210 168140 87290 168150
rect 87360 168140 87440 168150
rect 87610 168149 87690 168159
rect 87930 168149 88010 168159
rect 88350 168149 88430 168159
rect 88670 168149 88750 168159
rect 75640 168060 75650 168140
rect 75790 168060 75800 168140
rect 87140 168060 87150 168140
rect 87290 168060 87300 168140
rect 87440 168060 87450 168140
rect 87690 168069 87700 168149
rect 88010 168069 88020 168149
rect 88430 168069 88440 168149
rect 88750 168069 88760 168149
rect 89060 168140 89140 168150
rect 89210 168140 89290 168150
rect 100560 168140 100640 168150
rect 100710 168140 100790 168150
rect 100860 168140 100940 168150
rect 101110 168149 101190 168159
rect 101430 168149 101510 168159
rect 101850 168149 101930 168159
rect 102170 168149 102250 168159
rect 114610 168149 114690 168159
rect 114930 168149 115010 168159
rect 115350 168149 115430 168159
rect 115670 168149 115750 168159
rect 89140 168060 89150 168140
rect 89290 168060 89300 168140
rect 100640 168060 100650 168140
rect 100790 168060 100800 168140
rect 100940 168060 100950 168140
rect 101190 168069 101200 168149
rect 101510 168069 101520 168149
rect 101930 168069 101940 168149
rect 102250 168069 102260 168149
rect 114690 168069 114700 168149
rect 115010 168069 115020 168149
rect 115430 168069 115440 168149
rect 115750 168069 115760 168149
rect 116060 168140 116140 168150
rect 116210 168140 116290 168150
rect 127560 168140 127640 168150
rect 127710 168140 127790 168150
rect 127860 168140 127940 168150
rect 128110 168149 128190 168159
rect 128430 168149 128510 168159
rect 128850 168149 128930 168159
rect 129170 168149 129250 168159
rect 141825 168150 141905 168160
rect 142145 168150 142200 168160
rect 145345 168150 145425 168160
rect 145665 168150 145745 168160
rect 145985 168150 146065 168160
rect 116140 168060 116150 168140
rect 116290 168060 116300 168140
rect 127640 168060 127650 168140
rect 127790 168060 127800 168140
rect 127940 168060 127950 168140
rect 128190 168069 128200 168149
rect 128510 168069 128520 168149
rect 128930 168069 128940 168149
rect 129250 168069 129260 168149
rect 129560 168140 129640 168150
rect 129710 168140 129790 168150
rect 140710 168140 140730 168150
rect 141060 168140 141140 168150
rect 141210 168140 141290 168150
rect 141360 168140 141440 168150
rect 129640 168060 129650 168140
rect 129790 168060 129800 168140
rect 140730 168060 140740 168140
rect 141140 168060 141150 168140
rect 141290 168060 141300 168140
rect 141440 168060 141450 168140
rect 141905 168070 141915 168150
rect 145425 168070 145435 168150
rect 145745 168070 145755 168150
rect 146065 168070 146075 168150
rect 146780 168140 146790 168220
rect 146540 168060 146620 168070
rect 146860 168060 146940 168070
rect 60770 167989 60850 167999
rect 61090 167989 61170 167999
rect 61510 167989 61590 167999
rect 61830 167989 61910 167999
rect 74270 167989 74350 167999
rect 74590 167989 74670 167999
rect 75010 167989 75090 167999
rect 75330 167989 75410 167999
rect 87770 167989 87850 167999
rect 88090 167989 88170 167999
rect 88510 167989 88590 167999
rect 88830 167989 88910 167999
rect 101270 167989 101350 167999
rect 101590 167989 101670 167999
rect 102010 167989 102090 167999
rect 102330 167989 102410 167999
rect 114770 167989 114850 167999
rect 115090 167989 115170 167999
rect 115510 167989 115590 167999
rect 115830 167989 115910 167999
rect 128270 167989 128350 167999
rect 128590 167989 128670 167999
rect 129010 167989 129090 167999
rect 129330 167989 129410 167999
rect 141665 167990 141745 168000
rect 141985 167990 142065 168000
rect 145200 167990 145265 168000
rect 145505 167990 145585 168000
rect 145825 167990 145905 168000
rect 59350 167960 59430 167970
rect 59500 167960 59580 167970
rect 59650 167960 59730 167970
rect 60060 167960 60140 167970
rect 60210 167960 60290 167970
rect 60360 167960 60440 167970
rect 59430 167880 59440 167960
rect 59580 167880 59590 167960
rect 59730 167880 59740 167960
rect 60140 167880 60150 167960
rect 60290 167880 60300 167960
rect 60440 167880 60450 167960
rect 60850 167909 60860 167989
rect 61170 167909 61180 167989
rect 61590 167909 61600 167989
rect 61910 167909 61920 167989
rect 62060 167960 62140 167970
rect 62210 167960 62290 167970
rect 73560 167960 73640 167970
rect 73710 167960 73790 167970
rect 73860 167960 73940 167970
rect 62140 167880 62150 167960
rect 62290 167880 62300 167960
rect 73640 167880 73650 167960
rect 73790 167880 73800 167960
rect 73940 167880 73950 167960
rect 74350 167909 74360 167989
rect 74670 167909 74680 167989
rect 75090 167909 75100 167989
rect 75410 167909 75420 167989
rect 75560 167960 75640 167970
rect 75710 167960 75790 167970
rect 87060 167960 87140 167970
rect 87210 167960 87290 167970
rect 87360 167960 87440 167970
rect 75640 167880 75650 167960
rect 75790 167880 75800 167960
rect 87140 167880 87150 167960
rect 87290 167880 87300 167960
rect 87440 167880 87450 167960
rect 87850 167909 87860 167989
rect 88170 167909 88180 167989
rect 88590 167909 88600 167989
rect 88910 167909 88920 167989
rect 89060 167960 89140 167970
rect 89210 167960 89290 167970
rect 100560 167960 100640 167970
rect 100710 167960 100790 167970
rect 100860 167960 100940 167970
rect 89140 167880 89150 167960
rect 89290 167880 89300 167960
rect 100640 167880 100650 167960
rect 100790 167880 100800 167960
rect 100940 167880 100950 167960
rect 101350 167909 101360 167989
rect 101670 167909 101680 167989
rect 102090 167909 102100 167989
rect 102410 167909 102420 167989
rect 114850 167909 114860 167989
rect 115170 167909 115180 167989
rect 115590 167909 115600 167989
rect 115910 167909 115920 167989
rect 116060 167960 116140 167970
rect 116210 167960 116290 167970
rect 127560 167960 127640 167970
rect 127710 167960 127790 167970
rect 127860 167960 127940 167970
rect 116140 167880 116150 167960
rect 116290 167880 116300 167960
rect 127640 167880 127650 167960
rect 127790 167880 127800 167960
rect 127940 167880 127950 167960
rect 128350 167909 128360 167989
rect 128670 167909 128680 167989
rect 129090 167909 129100 167989
rect 129410 167909 129420 167989
rect 129560 167960 129640 167970
rect 129710 167960 129790 167970
rect 140710 167960 140730 167970
rect 141060 167960 141140 167970
rect 141210 167960 141290 167970
rect 141360 167960 141440 167970
rect 129640 167880 129650 167960
rect 129790 167880 129800 167960
rect 140730 167880 140740 167960
rect 141140 167880 141150 167960
rect 141290 167880 141300 167960
rect 141440 167880 141450 167960
rect 141745 167910 141755 167990
rect 142065 167910 142075 167990
rect 145265 167910 145275 167990
rect 145585 167910 145595 167990
rect 145905 167910 145915 167990
rect 146620 167980 146630 168060
rect 146940 167980 146950 168060
rect 146700 167900 146780 167910
rect 60610 167829 60690 167839
rect 60930 167829 61010 167839
rect 61350 167829 61430 167839
rect 61670 167829 61750 167839
rect 74110 167829 74190 167839
rect 74430 167829 74510 167839
rect 74850 167829 74930 167839
rect 75170 167829 75250 167839
rect 87610 167829 87690 167839
rect 87930 167829 88010 167839
rect 88350 167829 88430 167839
rect 88670 167829 88750 167839
rect 101110 167829 101190 167839
rect 101430 167829 101510 167839
rect 101850 167829 101930 167839
rect 102170 167829 102250 167839
rect 114610 167829 114690 167839
rect 114930 167829 115010 167839
rect 115350 167829 115430 167839
rect 115670 167829 115750 167839
rect 128110 167829 128190 167839
rect 128430 167829 128510 167839
rect 128850 167829 128930 167839
rect 129170 167829 129250 167839
rect 141825 167830 141905 167840
rect 142145 167830 142200 167840
rect 145345 167830 145425 167840
rect 145665 167830 145745 167840
rect 145985 167830 146065 167840
rect 59350 167780 59430 167790
rect 59500 167780 59580 167790
rect 59650 167780 59730 167790
rect 60060 167780 60140 167790
rect 60210 167780 60290 167790
rect 60360 167780 60440 167790
rect 59430 167700 59440 167780
rect 59580 167700 59590 167780
rect 59730 167700 59740 167780
rect 60140 167700 60150 167780
rect 60290 167700 60300 167780
rect 60440 167700 60450 167780
rect 60690 167749 60700 167829
rect 61010 167749 61020 167829
rect 61430 167749 61440 167829
rect 61750 167749 61760 167829
rect 62060 167780 62140 167790
rect 62210 167780 62290 167790
rect 73560 167780 73640 167790
rect 73710 167780 73790 167790
rect 73860 167780 73940 167790
rect 62140 167700 62150 167780
rect 62290 167700 62300 167780
rect 73640 167700 73650 167780
rect 73790 167700 73800 167780
rect 73940 167700 73950 167780
rect 74190 167749 74200 167829
rect 74510 167749 74520 167829
rect 74930 167749 74940 167829
rect 75250 167749 75260 167829
rect 75560 167780 75640 167790
rect 75710 167780 75790 167790
rect 87060 167780 87140 167790
rect 87210 167780 87290 167790
rect 87360 167780 87440 167790
rect 75640 167700 75650 167780
rect 75790 167700 75800 167780
rect 87140 167700 87150 167780
rect 87290 167700 87300 167780
rect 87440 167700 87450 167780
rect 87690 167749 87700 167829
rect 88010 167749 88020 167829
rect 88430 167749 88440 167829
rect 88750 167749 88760 167829
rect 89060 167780 89140 167790
rect 89210 167780 89290 167790
rect 100560 167780 100640 167790
rect 100710 167780 100790 167790
rect 100860 167780 100940 167790
rect 89140 167700 89150 167780
rect 89290 167700 89300 167780
rect 100640 167700 100650 167780
rect 100790 167700 100800 167780
rect 100940 167700 100950 167780
rect 101190 167749 101200 167829
rect 101510 167749 101520 167829
rect 101930 167749 101940 167829
rect 102250 167749 102260 167829
rect 114690 167749 114700 167829
rect 115010 167749 115020 167829
rect 115430 167749 115440 167829
rect 115750 167749 115760 167829
rect 116060 167780 116140 167790
rect 116210 167780 116290 167790
rect 127560 167780 127640 167790
rect 127710 167780 127790 167790
rect 127860 167780 127940 167790
rect 116140 167700 116150 167780
rect 116290 167700 116300 167780
rect 127640 167700 127650 167780
rect 127790 167700 127800 167780
rect 127940 167700 127950 167780
rect 128190 167749 128200 167829
rect 128510 167749 128520 167829
rect 128930 167749 128940 167829
rect 129250 167749 129260 167829
rect 129560 167780 129640 167790
rect 129710 167780 129790 167790
rect 140710 167780 140730 167790
rect 141060 167780 141140 167790
rect 141210 167780 141290 167790
rect 141360 167780 141440 167790
rect 129640 167700 129650 167780
rect 129790 167700 129800 167780
rect 140730 167700 140740 167780
rect 141140 167700 141150 167780
rect 141290 167700 141300 167780
rect 141440 167700 141450 167780
rect 141905 167750 141915 167830
rect 145425 167750 145435 167830
rect 145745 167750 145755 167830
rect 146065 167750 146075 167830
rect 146780 167820 146790 167900
rect 146540 167740 146620 167750
rect 146860 167740 146940 167750
rect 60770 167669 60850 167679
rect 61090 167669 61170 167679
rect 61510 167669 61590 167679
rect 61830 167669 61910 167679
rect 74270 167669 74350 167679
rect 74590 167669 74670 167679
rect 75010 167669 75090 167679
rect 75330 167669 75410 167679
rect 87770 167669 87850 167679
rect 88090 167669 88170 167679
rect 88510 167669 88590 167679
rect 88830 167669 88910 167679
rect 101270 167669 101350 167679
rect 101590 167669 101670 167679
rect 102010 167669 102090 167679
rect 102330 167669 102410 167679
rect 114770 167669 114850 167679
rect 115090 167669 115170 167679
rect 115510 167669 115590 167679
rect 115830 167669 115910 167679
rect 128270 167669 128350 167679
rect 128590 167669 128670 167679
rect 129010 167669 129090 167679
rect 129330 167669 129410 167679
rect 141665 167670 141745 167680
rect 141985 167670 142065 167680
rect 145200 167670 145265 167680
rect 145505 167670 145585 167680
rect 145825 167670 145905 167680
rect 59350 167600 59430 167610
rect 59500 167600 59580 167610
rect 59650 167600 59730 167610
rect 60060 167600 60140 167610
rect 60210 167600 60290 167610
rect 60360 167600 60440 167610
rect 59430 167520 59440 167600
rect 59580 167520 59590 167600
rect 59730 167520 59740 167600
rect 60140 167520 60150 167600
rect 60290 167520 60300 167600
rect 60440 167520 60450 167600
rect 60850 167589 60860 167669
rect 61170 167589 61180 167669
rect 61590 167589 61600 167669
rect 61910 167589 61920 167669
rect 62060 167600 62140 167610
rect 62210 167600 62290 167610
rect 73560 167600 73640 167610
rect 73710 167600 73790 167610
rect 73860 167600 73940 167610
rect 62140 167520 62150 167600
rect 62290 167520 62300 167600
rect 73640 167520 73650 167600
rect 73790 167520 73800 167600
rect 73940 167520 73950 167600
rect 74350 167589 74360 167669
rect 74670 167589 74680 167669
rect 75090 167589 75100 167669
rect 75410 167589 75420 167669
rect 75560 167600 75640 167610
rect 75710 167600 75790 167610
rect 87060 167600 87140 167610
rect 87210 167600 87290 167610
rect 87360 167600 87440 167610
rect 75640 167520 75650 167600
rect 75790 167520 75800 167600
rect 87140 167520 87150 167600
rect 87290 167520 87300 167600
rect 87440 167520 87450 167600
rect 87850 167589 87860 167669
rect 88170 167589 88180 167669
rect 88590 167589 88600 167669
rect 88910 167589 88920 167669
rect 89060 167600 89140 167610
rect 89210 167600 89290 167610
rect 100560 167600 100640 167610
rect 100710 167600 100790 167610
rect 100860 167600 100940 167610
rect 89140 167520 89150 167600
rect 89290 167520 89300 167600
rect 100640 167520 100650 167600
rect 100790 167520 100800 167600
rect 100940 167520 100950 167600
rect 101350 167589 101360 167669
rect 101670 167589 101680 167669
rect 102090 167589 102100 167669
rect 102410 167589 102420 167669
rect 114850 167589 114860 167669
rect 115170 167589 115180 167669
rect 115590 167589 115600 167669
rect 115910 167589 115920 167669
rect 116060 167600 116140 167610
rect 116210 167600 116290 167610
rect 127560 167600 127640 167610
rect 127710 167600 127790 167610
rect 127860 167600 127940 167610
rect 116140 167520 116150 167600
rect 116290 167520 116300 167600
rect 127640 167520 127650 167600
rect 127790 167520 127800 167600
rect 127940 167520 127950 167600
rect 128350 167589 128360 167669
rect 128670 167589 128680 167669
rect 129090 167589 129100 167669
rect 129410 167589 129420 167669
rect 129560 167600 129640 167610
rect 129710 167600 129790 167610
rect 140710 167600 140730 167610
rect 141060 167600 141140 167610
rect 141210 167600 141290 167610
rect 141360 167600 141440 167610
rect 129640 167520 129650 167600
rect 129790 167520 129800 167600
rect 140730 167520 140740 167600
rect 141140 167520 141150 167600
rect 141290 167520 141300 167600
rect 141440 167520 141450 167600
rect 141745 167590 141755 167670
rect 142065 167590 142075 167670
rect 145265 167590 145275 167670
rect 145585 167590 145595 167670
rect 145905 167590 145915 167670
rect 146620 167660 146630 167740
rect 146940 167660 146950 167740
rect 146700 167580 146780 167590
rect 60610 167509 60690 167519
rect 60930 167509 61010 167519
rect 61350 167509 61430 167519
rect 61670 167509 61750 167519
rect 74110 167509 74190 167519
rect 74430 167509 74510 167519
rect 74850 167509 74930 167519
rect 75170 167509 75250 167519
rect 87610 167509 87690 167519
rect 87930 167509 88010 167519
rect 88350 167509 88430 167519
rect 88670 167509 88750 167519
rect 101110 167509 101190 167519
rect 101430 167509 101510 167519
rect 101850 167509 101930 167519
rect 102170 167509 102250 167519
rect 114610 167509 114690 167519
rect 114930 167509 115010 167519
rect 115350 167509 115430 167519
rect 115670 167509 115750 167519
rect 128110 167509 128190 167519
rect 128430 167509 128510 167519
rect 128850 167509 128930 167519
rect 129170 167509 129250 167519
rect 141825 167510 141905 167520
rect 142145 167510 142200 167520
rect 145345 167510 145425 167520
rect 145665 167510 145745 167520
rect 145985 167510 146065 167520
rect 59350 167420 59430 167430
rect 59500 167420 59580 167430
rect 59650 167420 59730 167430
rect 60060 167420 60140 167430
rect 60210 167420 60290 167430
rect 60360 167420 60440 167430
rect 60690 167429 60700 167509
rect 61010 167429 61020 167509
rect 61430 167429 61440 167509
rect 61750 167429 61760 167509
rect 62060 167420 62140 167430
rect 62210 167420 62290 167430
rect 73560 167420 73640 167430
rect 73710 167420 73790 167430
rect 73860 167420 73940 167430
rect 74190 167429 74200 167509
rect 74510 167429 74520 167509
rect 74930 167429 74940 167509
rect 75250 167429 75260 167509
rect 75560 167420 75640 167430
rect 75710 167420 75790 167430
rect 87060 167420 87140 167430
rect 87210 167420 87290 167430
rect 87360 167420 87440 167430
rect 87690 167429 87700 167509
rect 88010 167429 88020 167509
rect 88430 167429 88440 167509
rect 88750 167429 88760 167509
rect 89060 167420 89140 167430
rect 89210 167420 89290 167430
rect 100560 167420 100640 167430
rect 100710 167420 100790 167430
rect 100860 167420 100940 167430
rect 101190 167429 101200 167509
rect 101510 167429 101520 167509
rect 101930 167429 101940 167509
rect 102250 167429 102260 167509
rect 114690 167429 114700 167509
rect 115010 167429 115020 167509
rect 115430 167429 115440 167509
rect 115750 167429 115760 167509
rect 116060 167420 116140 167430
rect 116210 167420 116290 167430
rect 127560 167420 127640 167430
rect 127710 167420 127790 167430
rect 127860 167420 127940 167430
rect 128190 167429 128200 167509
rect 128510 167429 128520 167509
rect 128930 167429 128940 167509
rect 129250 167429 129260 167509
rect 141905 167430 141915 167510
rect 145425 167430 145435 167510
rect 145745 167430 145755 167510
rect 146065 167430 146075 167510
rect 146780 167500 146790 167580
rect 129560 167420 129640 167430
rect 129710 167420 129790 167430
rect 140710 167420 140730 167430
rect 141060 167420 141140 167430
rect 141210 167420 141290 167430
rect 141360 167420 141440 167430
rect 146540 167420 146620 167430
rect 146860 167420 146940 167430
rect 59430 167340 59440 167420
rect 59580 167340 59590 167420
rect 59730 167340 59740 167420
rect 60140 167340 60150 167420
rect 60290 167340 60300 167420
rect 60440 167340 60450 167420
rect 60770 167349 60850 167359
rect 61090 167349 61170 167359
rect 61510 167349 61590 167359
rect 61830 167349 61910 167359
rect 60850 167269 60860 167349
rect 61170 167269 61180 167349
rect 61590 167269 61600 167349
rect 61910 167269 61920 167349
rect 62140 167340 62150 167420
rect 62290 167340 62300 167420
rect 73640 167340 73650 167420
rect 73790 167340 73800 167420
rect 73940 167340 73950 167420
rect 74270 167349 74350 167359
rect 74590 167349 74670 167359
rect 75010 167349 75090 167359
rect 75330 167349 75410 167359
rect 74350 167269 74360 167349
rect 74670 167269 74680 167349
rect 75090 167269 75100 167349
rect 75410 167269 75420 167349
rect 75640 167340 75650 167420
rect 75790 167340 75800 167420
rect 87140 167340 87150 167420
rect 87290 167340 87300 167420
rect 87440 167340 87450 167420
rect 87770 167349 87850 167359
rect 88090 167349 88170 167359
rect 88510 167349 88590 167359
rect 88830 167349 88910 167359
rect 87850 167269 87860 167349
rect 88170 167269 88180 167349
rect 88590 167269 88600 167349
rect 88910 167269 88920 167349
rect 89140 167340 89150 167420
rect 89290 167340 89300 167420
rect 100640 167340 100650 167420
rect 100790 167340 100800 167420
rect 100940 167340 100950 167420
rect 101270 167349 101350 167359
rect 101590 167349 101670 167359
rect 102010 167349 102090 167359
rect 102330 167349 102410 167359
rect 114770 167349 114850 167359
rect 115090 167349 115170 167359
rect 115510 167349 115590 167359
rect 115830 167349 115910 167359
rect 101350 167269 101360 167349
rect 101670 167269 101680 167349
rect 102090 167269 102100 167349
rect 102410 167269 102420 167349
rect 114850 167269 114860 167349
rect 115170 167269 115180 167349
rect 115590 167269 115600 167349
rect 115910 167269 115920 167349
rect 116140 167340 116150 167420
rect 116290 167340 116300 167420
rect 127640 167340 127650 167420
rect 127790 167340 127800 167420
rect 127940 167340 127950 167420
rect 128270 167349 128350 167359
rect 128590 167349 128670 167359
rect 129010 167349 129090 167359
rect 129330 167349 129410 167359
rect 128350 167269 128360 167349
rect 128670 167269 128680 167349
rect 129090 167269 129100 167349
rect 129410 167269 129420 167349
rect 129640 167340 129650 167420
rect 129790 167340 129800 167420
rect 140730 167340 140740 167420
rect 141140 167340 141150 167420
rect 141290 167340 141300 167420
rect 141440 167340 141450 167420
rect 141665 167350 141745 167360
rect 141985 167350 142065 167360
rect 145200 167350 145265 167360
rect 145505 167350 145585 167360
rect 145825 167350 145905 167360
rect 141745 167270 141755 167350
rect 142065 167270 142075 167350
rect 145265 167270 145275 167350
rect 145585 167270 145595 167350
rect 145905 167270 145915 167350
rect 146620 167340 146630 167420
rect 146940 167340 146950 167420
rect 146700 167260 146780 167270
rect 59350 167240 59430 167250
rect 59500 167240 59580 167250
rect 59650 167240 59730 167250
rect 60060 167240 60140 167250
rect 60210 167240 60290 167250
rect 60360 167240 60440 167250
rect 62060 167240 62140 167250
rect 62210 167240 62290 167250
rect 73560 167240 73640 167250
rect 73710 167240 73790 167250
rect 73860 167240 73940 167250
rect 75560 167240 75640 167250
rect 75710 167240 75790 167250
rect 87060 167240 87140 167250
rect 87210 167240 87290 167250
rect 87360 167240 87440 167250
rect 89060 167240 89140 167250
rect 89210 167240 89290 167250
rect 100560 167240 100640 167250
rect 100710 167240 100790 167250
rect 100860 167240 100940 167250
rect 116060 167240 116140 167250
rect 116210 167240 116290 167250
rect 127560 167240 127640 167250
rect 127710 167240 127790 167250
rect 127860 167240 127940 167250
rect 129560 167240 129640 167250
rect 129710 167240 129790 167250
rect 140710 167240 140730 167250
rect 141060 167240 141140 167250
rect 141210 167240 141290 167250
rect 141360 167240 141440 167250
rect 59430 167160 59440 167240
rect 59580 167160 59590 167240
rect 59730 167160 59740 167240
rect 60140 167160 60150 167240
rect 60290 167160 60300 167240
rect 60440 167160 60450 167240
rect 60610 167189 60690 167199
rect 60930 167189 61010 167199
rect 61350 167189 61430 167199
rect 61670 167189 61750 167199
rect 60690 167109 60700 167189
rect 61010 167109 61020 167189
rect 61430 167109 61440 167189
rect 61750 167109 61760 167189
rect 62140 167160 62150 167240
rect 62290 167160 62300 167240
rect 73640 167160 73650 167240
rect 73790 167160 73800 167240
rect 73940 167160 73950 167240
rect 74110 167189 74190 167199
rect 74430 167189 74510 167199
rect 74850 167189 74930 167199
rect 75170 167189 75250 167199
rect 74190 167109 74200 167189
rect 74510 167109 74520 167189
rect 74930 167109 74940 167189
rect 75250 167109 75260 167189
rect 75640 167160 75650 167240
rect 75790 167160 75800 167240
rect 87140 167160 87150 167240
rect 87290 167160 87300 167240
rect 87440 167160 87450 167240
rect 87610 167189 87690 167199
rect 87930 167189 88010 167199
rect 88350 167189 88430 167199
rect 88670 167189 88750 167199
rect 87690 167109 87700 167189
rect 88010 167109 88020 167189
rect 88430 167109 88440 167189
rect 88750 167109 88760 167189
rect 89140 167160 89150 167240
rect 89290 167160 89300 167240
rect 100640 167160 100650 167240
rect 100790 167160 100800 167240
rect 100940 167160 100950 167240
rect 101110 167189 101190 167199
rect 101430 167189 101510 167199
rect 101850 167189 101930 167199
rect 102170 167189 102250 167199
rect 114610 167189 114690 167199
rect 114930 167189 115010 167199
rect 115350 167189 115430 167199
rect 115670 167189 115750 167199
rect 101190 167109 101200 167189
rect 101510 167109 101520 167189
rect 101930 167109 101940 167189
rect 102250 167109 102260 167189
rect 114690 167109 114700 167189
rect 115010 167109 115020 167189
rect 115430 167109 115440 167189
rect 115750 167109 115760 167189
rect 116140 167160 116150 167240
rect 116290 167160 116300 167240
rect 127640 167160 127650 167240
rect 127790 167160 127800 167240
rect 127940 167160 127950 167240
rect 128110 167189 128190 167199
rect 128430 167189 128510 167199
rect 128850 167189 128930 167199
rect 129170 167189 129250 167199
rect 128190 167109 128200 167189
rect 128510 167109 128520 167189
rect 128930 167109 128940 167189
rect 129250 167109 129260 167189
rect 129640 167160 129650 167240
rect 129790 167160 129800 167240
rect 140730 167160 140740 167240
rect 141140 167160 141150 167240
rect 141290 167160 141300 167240
rect 141440 167160 141450 167240
rect 141825 167190 141905 167200
rect 142145 167190 142200 167200
rect 145345 167190 145425 167200
rect 145665 167190 145745 167200
rect 145985 167190 146065 167200
rect 141905 167110 141915 167190
rect 145425 167110 145435 167190
rect 145745 167110 145755 167190
rect 146065 167110 146075 167190
rect 146780 167180 146790 167260
rect 146540 167100 146620 167110
rect 146860 167100 146940 167110
rect 59350 167060 59430 167070
rect 59500 167060 59580 167070
rect 59650 167060 59730 167070
rect 60060 167060 60140 167070
rect 60210 167060 60290 167070
rect 60360 167060 60440 167070
rect 62060 167060 62140 167070
rect 62210 167060 62290 167070
rect 73560 167060 73640 167070
rect 73710 167060 73790 167070
rect 73860 167060 73940 167070
rect 75560 167060 75640 167070
rect 75710 167060 75790 167070
rect 87060 167060 87140 167070
rect 87210 167060 87290 167070
rect 87360 167060 87440 167070
rect 89060 167060 89140 167070
rect 89210 167060 89290 167070
rect 100560 167060 100640 167070
rect 100710 167060 100790 167070
rect 100860 167060 100940 167070
rect 116060 167060 116140 167070
rect 116210 167060 116290 167070
rect 127560 167060 127640 167070
rect 127710 167060 127790 167070
rect 127860 167060 127940 167070
rect 129560 167060 129640 167070
rect 129710 167060 129790 167070
rect 140710 167060 140730 167070
rect 141060 167060 141140 167070
rect 141210 167060 141290 167070
rect 141360 167060 141440 167070
rect 59430 166980 59440 167060
rect 59580 166980 59590 167060
rect 59730 166980 59740 167060
rect 60140 166980 60150 167060
rect 60290 166980 60300 167060
rect 60440 166980 60450 167060
rect 60770 167029 60850 167039
rect 61090 167029 61170 167039
rect 61510 167029 61590 167039
rect 61830 167029 61910 167039
rect 60850 166949 60860 167029
rect 61170 166949 61180 167029
rect 61590 166949 61600 167029
rect 61910 166949 61920 167029
rect 62140 166980 62150 167060
rect 62290 166980 62300 167060
rect 73640 166980 73650 167060
rect 73790 166980 73800 167060
rect 73940 166980 73950 167060
rect 74270 167029 74350 167039
rect 74590 167029 74670 167039
rect 75010 167029 75090 167039
rect 75330 167029 75410 167039
rect 74350 166949 74360 167029
rect 74670 166949 74680 167029
rect 75090 166949 75100 167029
rect 75410 166949 75420 167029
rect 75640 166980 75650 167060
rect 75790 166980 75800 167060
rect 87140 166980 87150 167060
rect 87290 166980 87300 167060
rect 87440 166980 87450 167060
rect 87770 167029 87850 167039
rect 88090 167029 88170 167039
rect 88510 167029 88590 167039
rect 88830 167029 88910 167039
rect 87850 166949 87860 167029
rect 88170 166949 88180 167029
rect 88590 166949 88600 167029
rect 88910 166949 88920 167029
rect 89140 166980 89150 167060
rect 89290 166980 89300 167060
rect 100640 166980 100650 167060
rect 100790 166980 100800 167060
rect 100940 166980 100950 167060
rect 101270 167029 101350 167039
rect 101590 167029 101670 167039
rect 102010 167029 102090 167039
rect 102330 167029 102410 167039
rect 114770 167029 114850 167039
rect 115090 167029 115170 167039
rect 115510 167029 115590 167039
rect 115830 167029 115910 167039
rect 101350 166949 101360 167029
rect 101670 166949 101680 167029
rect 102090 166949 102100 167029
rect 102410 166949 102420 167029
rect 114850 166949 114860 167029
rect 115170 166949 115180 167029
rect 115590 166949 115600 167029
rect 115910 166949 115920 167029
rect 116140 166980 116150 167060
rect 116290 166980 116300 167060
rect 127640 166980 127650 167060
rect 127790 166980 127800 167060
rect 127940 166980 127950 167060
rect 128270 167029 128350 167039
rect 128590 167029 128670 167039
rect 129010 167029 129090 167039
rect 129330 167029 129410 167039
rect 128350 166949 128360 167029
rect 128670 166949 128680 167029
rect 129090 166949 129100 167029
rect 129410 166949 129420 167029
rect 129640 166980 129650 167060
rect 129790 166980 129800 167060
rect 140730 166980 140740 167060
rect 141140 166980 141150 167060
rect 141290 166980 141300 167060
rect 141440 166980 141450 167060
rect 141665 167030 141745 167040
rect 141985 167030 142065 167040
rect 145200 167030 145265 167040
rect 145505 167030 145585 167040
rect 145825 167030 145905 167040
rect 141745 166950 141755 167030
rect 142065 166950 142075 167030
rect 145265 166950 145275 167030
rect 145585 166950 145595 167030
rect 145905 166950 145915 167030
rect 146620 167020 146630 167100
rect 146940 167020 146950 167100
rect 146700 166940 146780 166950
rect 59350 166880 59430 166890
rect 59500 166880 59580 166890
rect 59650 166880 59730 166890
rect 60060 166880 60140 166890
rect 60210 166880 60290 166890
rect 60360 166880 60440 166890
rect 62060 166880 62140 166890
rect 62210 166880 62290 166890
rect 73560 166880 73640 166890
rect 73710 166880 73790 166890
rect 73860 166880 73940 166890
rect 75560 166880 75640 166890
rect 75710 166880 75790 166890
rect 87060 166880 87140 166890
rect 87210 166880 87290 166890
rect 87360 166880 87440 166890
rect 89060 166880 89140 166890
rect 89210 166880 89290 166890
rect 100560 166880 100640 166890
rect 100710 166880 100790 166890
rect 100860 166880 100940 166890
rect 116060 166880 116140 166890
rect 116210 166880 116290 166890
rect 127560 166880 127640 166890
rect 127710 166880 127790 166890
rect 127860 166880 127940 166890
rect 129560 166880 129640 166890
rect 129710 166880 129790 166890
rect 140710 166880 140730 166890
rect 141060 166880 141140 166890
rect 141210 166880 141290 166890
rect 141360 166880 141440 166890
rect 59430 166800 59440 166880
rect 59580 166800 59590 166880
rect 59730 166800 59740 166880
rect 60140 166800 60150 166880
rect 60290 166800 60300 166880
rect 60440 166800 60450 166880
rect 60610 166869 60690 166879
rect 60930 166869 61010 166879
rect 61350 166869 61430 166879
rect 61670 166869 61750 166879
rect 60690 166789 60700 166869
rect 61010 166789 61020 166869
rect 61430 166789 61440 166869
rect 61750 166789 61760 166869
rect 62140 166800 62150 166880
rect 62290 166800 62300 166880
rect 73640 166800 73650 166880
rect 73790 166800 73800 166880
rect 73940 166800 73950 166880
rect 74110 166869 74190 166879
rect 74430 166869 74510 166879
rect 74850 166869 74930 166879
rect 75170 166869 75250 166879
rect 74190 166789 74200 166869
rect 74510 166789 74520 166869
rect 74930 166789 74940 166869
rect 75250 166789 75260 166869
rect 75640 166800 75650 166880
rect 75790 166800 75800 166880
rect 87140 166800 87150 166880
rect 87290 166800 87300 166880
rect 87440 166800 87450 166880
rect 87610 166869 87690 166879
rect 87930 166869 88010 166879
rect 88350 166869 88430 166879
rect 88670 166869 88750 166879
rect 87690 166789 87700 166869
rect 88010 166789 88020 166869
rect 88430 166789 88440 166869
rect 88750 166789 88760 166869
rect 89140 166800 89150 166880
rect 89290 166800 89300 166880
rect 100640 166800 100650 166880
rect 100790 166800 100800 166880
rect 100940 166800 100950 166880
rect 101110 166869 101190 166879
rect 101430 166869 101510 166879
rect 101850 166869 101930 166879
rect 102170 166869 102250 166879
rect 114610 166869 114690 166879
rect 114930 166869 115010 166879
rect 115350 166869 115430 166879
rect 115670 166869 115750 166879
rect 101190 166789 101200 166869
rect 101510 166789 101520 166869
rect 101930 166789 101940 166869
rect 102250 166789 102260 166869
rect 114690 166789 114700 166869
rect 115010 166789 115020 166869
rect 115430 166789 115440 166869
rect 115750 166789 115760 166869
rect 116140 166800 116150 166880
rect 116290 166800 116300 166880
rect 127640 166800 127650 166880
rect 127790 166800 127800 166880
rect 127940 166800 127950 166880
rect 128110 166869 128190 166879
rect 128430 166869 128510 166879
rect 128850 166869 128930 166879
rect 129170 166869 129250 166879
rect 128190 166789 128200 166869
rect 128510 166789 128520 166869
rect 128930 166789 128940 166869
rect 129250 166789 129260 166869
rect 129640 166800 129650 166880
rect 129790 166800 129800 166880
rect 140730 166800 140740 166880
rect 141140 166800 141150 166880
rect 141290 166800 141300 166880
rect 141440 166800 141450 166880
rect 141825 166870 141905 166880
rect 142145 166870 142200 166880
rect 145345 166870 145425 166880
rect 145665 166870 145745 166880
rect 145985 166870 146065 166880
rect 141905 166790 141915 166870
rect 145425 166790 145435 166870
rect 145745 166790 145755 166870
rect 146065 166790 146075 166870
rect 146780 166860 146790 166940
rect 146540 166780 146620 166790
rect 146860 166780 146940 166790
rect 59350 166700 59430 166710
rect 59500 166700 59580 166710
rect 59650 166700 59730 166710
rect 60060 166700 60140 166710
rect 60210 166700 60290 166710
rect 60360 166700 60440 166710
rect 60770 166709 60850 166719
rect 61090 166709 61170 166719
rect 61510 166709 61590 166719
rect 61830 166709 61910 166719
rect 59430 166620 59440 166700
rect 59580 166620 59590 166700
rect 59730 166620 59740 166700
rect 60140 166620 60150 166700
rect 60290 166620 60300 166700
rect 60440 166620 60450 166700
rect 60850 166629 60860 166709
rect 61170 166629 61180 166709
rect 61590 166629 61600 166709
rect 61910 166629 61920 166709
rect 62060 166700 62140 166710
rect 62210 166700 62290 166710
rect 73560 166700 73640 166710
rect 73710 166700 73790 166710
rect 73860 166700 73940 166710
rect 74270 166709 74350 166719
rect 74590 166709 74670 166719
rect 75010 166709 75090 166719
rect 75330 166709 75410 166719
rect 62140 166620 62150 166700
rect 62290 166620 62300 166700
rect 73640 166620 73650 166700
rect 73790 166620 73800 166700
rect 73940 166620 73950 166700
rect 74350 166629 74360 166709
rect 74670 166629 74680 166709
rect 75090 166629 75100 166709
rect 75410 166629 75420 166709
rect 75560 166700 75640 166710
rect 75710 166700 75790 166710
rect 87060 166700 87140 166710
rect 87210 166700 87290 166710
rect 87360 166700 87440 166710
rect 87770 166709 87850 166719
rect 88090 166709 88170 166719
rect 88510 166709 88590 166719
rect 88830 166709 88910 166719
rect 75640 166620 75650 166700
rect 75790 166620 75800 166700
rect 87140 166620 87150 166700
rect 87290 166620 87300 166700
rect 87440 166620 87450 166700
rect 87850 166629 87860 166709
rect 88170 166629 88180 166709
rect 88590 166629 88600 166709
rect 88910 166629 88920 166709
rect 89060 166700 89140 166710
rect 89210 166700 89290 166710
rect 100560 166700 100640 166710
rect 100710 166700 100790 166710
rect 100860 166700 100940 166710
rect 101270 166709 101350 166719
rect 101590 166709 101670 166719
rect 102010 166709 102090 166719
rect 102330 166709 102410 166719
rect 114770 166709 114850 166719
rect 115090 166709 115170 166719
rect 115510 166709 115590 166719
rect 115830 166709 115910 166719
rect 89140 166620 89150 166700
rect 89290 166620 89300 166700
rect 100640 166620 100650 166700
rect 100790 166620 100800 166700
rect 100940 166620 100950 166700
rect 101350 166629 101360 166709
rect 101670 166629 101680 166709
rect 102090 166629 102100 166709
rect 102410 166629 102420 166709
rect 114850 166629 114860 166709
rect 115170 166629 115180 166709
rect 115590 166629 115600 166709
rect 115910 166629 115920 166709
rect 116060 166700 116140 166710
rect 116210 166700 116290 166710
rect 127560 166700 127640 166710
rect 127710 166700 127790 166710
rect 127860 166700 127940 166710
rect 128270 166709 128350 166719
rect 128590 166709 128670 166719
rect 129010 166709 129090 166719
rect 129330 166709 129410 166719
rect 141665 166710 141745 166720
rect 141985 166710 142065 166720
rect 145200 166710 145265 166720
rect 145505 166710 145585 166720
rect 145825 166710 145905 166720
rect 116140 166620 116150 166700
rect 116290 166620 116300 166700
rect 127640 166620 127650 166700
rect 127790 166620 127800 166700
rect 127940 166620 127950 166700
rect 128350 166629 128360 166709
rect 128670 166629 128680 166709
rect 129090 166629 129100 166709
rect 129410 166629 129420 166709
rect 129560 166700 129640 166710
rect 129710 166700 129790 166710
rect 140710 166700 140730 166710
rect 141060 166700 141140 166710
rect 141210 166700 141290 166710
rect 141360 166700 141440 166710
rect 129640 166620 129650 166700
rect 129790 166620 129800 166700
rect 140730 166620 140740 166700
rect 141140 166620 141150 166700
rect 141290 166620 141300 166700
rect 141440 166620 141450 166700
rect 141745 166630 141755 166710
rect 142065 166630 142075 166710
rect 145265 166630 145275 166710
rect 145585 166630 145595 166710
rect 145905 166630 145915 166710
rect 146620 166700 146630 166780
rect 146940 166700 146950 166780
rect 146700 166620 146780 166630
rect 60610 166549 60690 166559
rect 60930 166549 61010 166559
rect 61350 166549 61430 166559
rect 61670 166549 61750 166559
rect 74110 166549 74190 166559
rect 74430 166549 74510 166559
rect 74850 166549 74930 166559
rect 75170 166549 75250 166559
rect 87610 166549 87690 166559
rect 87930 166549 88010 166559
rect 88350 166549 88430 166559
rect 88670 166549 88750 166559
rect 101110 166549 101190 166559
rect 101430 166549 101510 166559
rect 101850 166549 101930 166559
rect 102170 166549 102250 166559
rect 114610 166549 114690 166559
rect 114930 166549 115010 166559
rect 115350 166549 115430 166559
rect 115670 166549 115750 166559
rect 128110 166549 128190 166559
rect 128430 166549 128510 166559
rect 128850 166549 128930 166559
rect 129170 166549 129250 166559
rect 141825 166550 141905 166560
rect 142145 166550 142200 166560
rect 145345 166550 145425 166560
rect 145665 166550 145745 166560
rect 145985 166550 146065 166560
rect 59350 166520 59430 166530
rect 59500 166520 59580 166530
rect 59650 166520 59730 166530
rect 60060 166520 60140 166530
rect 60210 166520 60290 166530
rect 60360 166520 60440 166530
rect 59430 166440 59440 166520
rect 59580 166440 59590 166520
rect 59730 166440 59740 166520
rect 60140 166440 60150 166520
rect 60290 166440 60300 166520
rect 60440 166440 60450 166520
rect 60690 166469 60700 166549
rect 61010 166469 61020 166549
rect 61430 166469 61440 166549
rect 61750 166469 61760 166549
rect 62060 166520 62140 166530
rect 62210 166520 62290 166530
rect 73560 166520 73640 166530
rect 73710 166520 73790 166530
rect 73860 166520 73940 166530
rect 62140 166440 62150 166520
rect 62290 166440 62300 166520
rect 73640 166440 73650 166520
rect 73790 166440 73800 166520
rect 73940 166440 73950 166520
rect 74190 166469 74200 166549
rect 74510 166469 74520 166549
rect 74930 166469 74940 166549
rect 75250 166469 75260 166549
rect 75560 166520 75640 166530
rect 75710 166520 75790 166530
rect 87060 166520 87140 166530
rect 87210 166520 87290 166530
rect 87360 166520 87440 166530
rect 75640 166440 75650 166520
rect 75790 166440 75800 166520
rect 87140 166440 87150 166520
rect 87290 166440 87300 166520
rect 87440 166440 87450 166520
rect 87690 166469 87700 166549
rect 88010 166469 88020 166549
rect 88430 166469 88440 166549
rect 88750 166469 88760 166549
rect 89060 166520 89140 166530
rect 89210 166520 89290 166530
rect 100560 166520 100640 166530
rect 100710 166520 100790 166530
rect 100860 166520 100940 166530
rect 89140 166440 89150 166520
rect 89290 166440 89300 166520
rect 100640 166440 100650 166520
rect 100790 166440 100800 166520
rect 100940 166440 100950 166520
rect 101190 166469 101200 166549
rect 101510 166469 101520 166549
rect 101930 166469 101940 166549
rect 102250 166469 102260 166549
rect 114690 166469 114700 166549
rect 115010 166469 115020 166549
rect 115430 166469 115440 166549
rect 115750 166469 115760 166549
rect 116060 166520 116140 166530
rect 116210 166520 116290 166530
rect 127560 166520 127640 166530
rect 127710 166520 127790 166530
rect 127860 166520 127940 166530
rect 116140 166440 116150 166520
rect 116290 166440 116300 166520
rect 127640 166440 127650 166520
rect 127790 166440 127800 166520
rect 127940 166440 127950 166520
rect 128190 166469 128200 166549
rect 128510 166469 128520 166549
rect 128930 166469 128940 166549
rect 129250 166469 129260 166549
rect 129560 166520 129640 166530
rect 129710 166520 129790 166530
rect 140710 166520 140730 166530
rect 141060 166520 141140 166530
rect 141210 166520 141290 166530
rect 141360 166520 141440 166530
rect 129640 166440 129650 166520
rect 129790 166440 129800 166520
rect 140730 166440 140740 166520
rect 141140 166440 141150 166520
rect 141290 166440 141300 166520
rect 141440 166440 141450 166520
rect 141905 166470 141915 166550
rect 145425 166470 145435 166550
rect 145745 166470 145755 166550
rect 146065 166470 146075 166550
rect 146780 166540 146790 166620
rect 146540 166460 146620 166470
rect 146860 166460 146940 166470
rect 60770 166389 60850 166399
rect 61090 166389 61170 166399
rect 61510 166389 61590 166399
rect 61830 166389 61910 166399
rect 74270 166389 74350 166399
rect 74590 166389 74670 166399
rect 75010 166389 75090 166399
rect 75330 166389 75410 166399
rect 87770 166389 87850 166399
rect 88090 166389 88170 166399
rect 88510 166389 88590 166399
rect 88830 166389 88910 166399
rect 101270 166389 101350 166399
rect 101590 166389 101670 166399
rect 102010 166389 102090 166399
rect 102330 166389 102410 166399
rect 114770 166389 114850 166399
rect 115090 166389 115170 166399
rect 115510 166389 115590 166399
rect 115830 166389 115910 166399
rect 128270 166389 128350 166399
rect 128590 166389 128670 166399
rect 129010 166389 129090 166399
rect 129330 166389 129410 166399
rect 141665 166390 141745 166400
rect 141985 166390 142065 166400
rect 145200 166390 145265 166400
rect 145505 166390 145585 166400
rect 145825 166390 145905 166400
rect 59350 166340 59430 166350
rect 59500 166340 59580 166350
rect 59650 166340 59730 166350
rect 60060 166340 60140 166350
rect 60210 166340 60290 166350
rect 60360 166340 60440 166350
rect 59430 166260 59440 166340
rect 59580 166260 59590 166340
rect 59730 166260 59740 166340
rect 60140 166260 60150 166340
rect 60290 166260 60300 166340
rect 60440 166260 60450 166340
rect 60850 166309 60860 166389
rect 61170 166309 61180 166389
rect 61590 166309 61600 166389
rect 61910 166309 61920 166389
rect 62060 166340 62140 166350
rect 62210 166340 62290 166350
rect 73560 166340 73640 166350
rect 73710 166340 73790 166350
rect 73860 166340 73940 166350
rect 62140 166260 62150 166340
rect 62290 166260 62300 166340
rect 73640 166260 73650 166340
rect 73790 166260 73800 166340
rect 73940 166260 73950 166340
rect 74350 166309 74360 166389
rect 74670 166309 74680 166389
rect 75090 166309 75100 166389
rect 75410 166309 75420 166389
rect 75560 166340 75640 166350
rect 75710 166340 75790 166350
rect 87060 166340 87140 166350
rect 87210 166340 87290 166350
rect 87360 166340 87440 166350
rect 75640 166260 75650 166340
rect 75790 166260 75800 166340
rect 87140 166260 87150 166340
rect 87290 166260 87300 166340
rect 87440 166260 87450 166340
rect 87850 166309 87860 166389
rect 88170 166309 88180 166389
rect 88590 166309 88600 166389
rect 88910 166309 88920 166389
rect 89060 166340 89140 166350
rect 89210 166340 89290 166350
rect 100560 166340 100640 166350
rect 100710 166340 100790 166350
rect 100860 166340 100940 166350
rect 89140 166260 89150 166340
rect 89290 166260 89300 166340
rect 100640 166260 100650 166340
rect 100790 166260 100800 166340
rect 100940 166260 100950 166340
rect 101350 166309 101360 166389
rect 101670 166309 101680 166389
rect 102090 166309 102100 166389
rect 102410 166309 102420 166389
rect 114850 166309 114860 166389
rect 115170 166309 115180 166389
rect 115590 166309 115600 166389
rect 115910 166309 115920 166389
rect 116060 166340 116140 166350
rect 116210 166340 116290 166350
rect 127560 166340 127640 166350
rect 127710 166340 127790 166350
rect 127860 166340 127940 166350
rect 116140 166260 116150 166340
rect 116290 166260 116300 166340
rect 127640 166260 127650 166340
rect 127790 166260 127800 166340
rect 127940 166260 127950 166340
rect 128350 166309 128360 166389
rect 128670 166309 128680 166389
rect 129090 166309 129100 166389
rect 129410 166309 129420 166389
rect 129560 166340 129640 166350
rect 129710 166340 129790 166350
rect 140710 166340 140730 166350
rect 141060 166340 141140 166350
rect 141210 166340 141290 166350
rect 141360 166340 141440 166350
rect 129640 166260 129650 166340
rect 129790 166260 129800 166340
rect 140730 166260 140740 166340
rect 141140 166260 141150 166340
rect 141290 166260 141300 166340
rect 141440 166260 141450 166340
rect 141745 166310 141755 166390
rect 142065 166310 142075 166390
rect 145265 166310 145275 166390
rect 145585 166310 145595 166390
rect 145905 166310 145915 166390
rect 146620 166380 146630 166460
rect 146940 166380 146950 166460
rect 146700 166300 146780 166310
rect 60610 166229 60690 166239
rect 60930 166229 61010 166239
rect 61350 166229 61430 166239
rect 61670 166229 61750 166239
rect 74110 166229 74190 166239
rect 74430 166229 74510 166239
rect 74850 166229 74930 166239
rect 75170 166229 75250 166239
rect 87610 166229 87690 166239
rect 87930 166229 88010 166239
rect 88350 166229 88430 166239
rect 88670 166229 88750 166239
rect 101110 166229 101190 166239
rect 101430 166229 101510 166239
rect 101850 166229 101930 166239
rect 102170 166229 102250 166239
rect 114610 166229 114690 166239
rect 114930 166229 115010 166239
rect 115350 166229 115430 166239
rect 115670 166229 115750 166239
rect 128110 166229 128190 166239
rect 128430 166229 128510 166239
rect 128850 166229 128930 166239
rect 129170 166229 129250 166239
rect 141825 166230 141905 166240
rect 142145 166230 142200 166240
rect 145345 166230 145425 166240
rect 145665 166230 145745 166240
rect 145985 166230 146065 166240
rect 59350 166160 59430 166170
rect 59500 166160 59580 166170
rect 59650 166160 59730 166170
rect 60060 166160 60140 166170
rect 60210 166160 60290 166170
rect 60360 166160 60440 166170
rect 59430 166080 59440 166160
rect 59580 166080 59590 166160
rect 59730 166080 59740 166160
rect 60140 166080 60150 166160
rect 60290 166080 60300 166160
rect 60440 166080 60450 166160
rect 60690 166149 60700 166229
rect 61010 166149 61020 166229
rect 61430 166149 61440 166229
rect 61750 166149 61760 166229
rect 62060 166160 62140 166170
rect 62210 166160 62290 166170
rect 73560 166160 73640 166170
rect 73710 166160 73790 166170
rect 73860 166160 73940 166170
rect 62140 166080 62150 166160
rect 62290 166080 62300 166160
rect 73640 166080 73650 166160
rect 73790 166080 73800 166160
rect 73940 166080 73950 166160
rect 74190 166149 74200 166229
rect 74510 166149 74520 166229
rect 74930 166149 74940 166229
rect 75250 166149 75260 166229
rect 75560 166160 75640 166170
rect 75710 166160 75790 166170
rect 87060 166160 87140 166170
rect 87210 166160 87290 166170
rect 87360 166160 87440 166170
rect 75640 166080 75650 166160
rect 75790 166080 75800 166160
rect 87140 166080 87150 166160
rect 87290 166080 87300 166160
rect 87440 166080 87450 166160
rect 87690 166149 87700 166229
rect 88010 166149 88020 166229
rect 88430 166149 88440 166229
rect 88750 166149 88760 166229
rect 89060 166160 89140 166170
rect 89210 166160 89290 166170
rect 100560 166160 100640 166170
rect 100710 166160 100790 166170
rect 100860 166160 100940 166170
rect 89140 166080 89150 166160
rect 89290 166080 89300 166160
rect 100640 166080 100650 166160
rect 100790 166080 100800 166160
rect 100940 166080 100950 166160
rect 101190 166149 101200 166229
rect 101510 166149 101520 166229
rect 101930 166149 101940 166229
rect 102250 166149 102260 166229
rect 114690 166149 114700 166229
rect 115010 166149 115020 166229
rect 115430 166149 115440 166229
rect 115750 166149 115760 166229
rect 116060 166160 116140 166170
rect 116210 166160 116290 166170
rect 127560 166160 127640 166170
rect 127710 166160 127790 166170
rect 127860 166160 127940 166170
rect 116140 166080 116150 166160
rect 116290 166080 116300 166160
rect 127640 166080 127650 166160
rect 127790 166080 127800 166160
rect 127940 166080 127950 166160
rect 128190 166149 128200 166229
rect 128510 166149 128520 166229
rect 128930 166149 128940 166229
rect 129250 166149 129260 166229
rect 129560 166160 129640 166170
rect 129710 166160 129790 166170
rect 140710 166160 140730 166170
rect 141060 166160 141140 166170
rect 141210 166160 141290 166170
rect 141360 166160 141440 166170
rect 129640 166080 129650 166160
rect 129790 166080 129800 166160
rect 140730 166080 140740 166160
rect 141140 166080 141150 166160
rect 141290 166080 141300 166160
rect 141440 166080 141450 166160
rect 141905 166150 141915 166230
rect 145425 166150 145435 166230
rect 145745 166150 145755 166230
rect 146065 166150 146075 166230
rect 146780 166220 146790 166300
rect 146540 166140 146620 166150
rect 146860 166140 146940 166150
rect 60770 166069 60850 166079
rect 61090 166069 61170 166079
rect 61510 166069 61590 166079
rect 61830 166069 61910 166079
rect 74270 166069 74350 166079
rect 74590 166069 74670 166079
rect 75010 166069 75090 166079
rect 75330 166069 75410 166079
rect 87770 166069 87850 166079
rect 88090 166069 88170 166079
rect 88510 166069 88590 166079
rect 88830 166069 88910 166079
rect 101270 166069 101350 166079
rect 101590 166069 101670 166079
rect 102010 166069 102090 166079
rect 102330 166069 102410 166079
rect 114770 166069 114850 166079
rect 115090 166069 115170 166079
rect 115510 166069 115590 166079
rect 115830 166069 115910 166079
rect 128270 166069 128350 166079
rect 128590 166069 128670 166079
rect 129010 166069 129090 166079
rect 129330 166069 129410 166079
rect 141665 166070 141745 166080
rect 141985 166070 142065 166080
rect 145200 166070 145265 166080
rect 145505 166070 145585 166080
rect 145825 166070 145905 166080
rect 59350 165980 59430 165990
rect 59500 165980 59580 165990
rect 59650 165980 59730 165990
rect 60060 165980 60140 165990
rect 60210 165980 60290 165990
rect 60360 165980 60440 165990
rect 60850 165989 60860 166069
rect 61170 165989 61180 166069
rect 61590 165989 61600 166069
rect 61910 165989 61920 166069
rect 62060 165980 62140 165990
rect 62210 165980 62290 165990
rect 73560 165980 73640 165990
rect 73710 165980 73790 165990
rect 73860 165980 73940 165990
rect 74350 165989 74360 166069
rect 74670 165989 74680 166069
rect 75090 165989 75100 166069
rect 75410 165989 75420 166069
rect 75560 165980 75640 165990
rect 75710 165980 75790 165990
rect 87060 165980 87140 165990
rect 87210 165980 87290 165990
rect 87360 165980 87440 165990
rect 87850 165989 87860 166069
rect 88170 165989 88180 166069
rect 88590 165989 88600 166069
rect 88910 165989 88920 166069
rect 89060 165980 89140 165990
rect 89210 165980 89290 165990
rect 100560 165980 100640 165990
rect 100710 165980 100790 165990
rect 100860 165980 100940 165990
rect 101350 165989 101360 166069
rect 101670 165989 101680 166069
rect 102090 165989 102100 166069
rect 102410 165989 102420 166069
rect 114850 165989 114860 166069
rect 115170 165989 115180 166069
rect 115590 165989 115600 166069
rect 115910 165989 115920 166069
rect 116060 165980 116140 165990
rect 116210 165980 116290 165990
rect 127560 165980 127640 165990
rect 127710 165980 127790 165990
rect 127860 165980 127940 165990
rect 128350 165989 128360 166069
rect 128670 165989 128680 166069
rect 129090 165989 129100 166069
rect 129410 165989 129420 166069
rect 141745 165990 141755 166070
rect 142065 165990 142075 166070
rect 145265 165990 145275 166070
rect 145585 165990 145595 166070
rect 145905 165990 145915 166070
rect 146620 166060 146630 166140
rect 146940 166060 146950 166140
rect 129560 165980 129640 165990
rect 129710 165980 129790 165990
rect 140710 165980 140730 165990
rect 141060 165980 141140 165990
rect 141210 165980 141290 165990
rect 141360 165980 141440 165990
rect 146700 165980 146780 165990
rect 59430 165900 59440 165980
rect 59580 165900 59590 165980
rect 59730 165900 59740 165980
rect 60140 165900 60150 165980
rect 60290 165900 60300 165980
rect 60440 165900 60450 165980
rect 60610 165909 60690 165919
rect 60930 165909 61010 165919
rect 61350 165909 61430 165919
rect 61670 165909 61750 165919
rect 60690 165829 60700 165909
rect 61010 165829 61020 165909
rect 61430 165829 61440 165909
rect 61750 165829 61760 165909
rect 62140 165900 62150 165980
rect 62290 165900 62300 165980
rect 73640 165900 73650 165980
rect 73790 165900 73800 165980
rect 73940 165900 73950 165980
rect 74110 165909 74190 165919
rect 74430 165909 74510 165919
rect 74850 165909 74930 165919
rect 75170 165909 75250 165919
rect 74190 165829 74200 165909
rect 74510 165829 74520 165909
rect 74930 165829 74940 165909
rect 75250 165829 75260 165909
rect 75640 165900 75650 165980
rect 75790 165900 75800 165980
rect 87140 165900 87150 165980
rect 87290 165900 87300 165980
rect 87440 165900 87450 165980
rect 87610 165909 87690 165919
rect 87930 165909 88010 165919
rect 88350 165909 88430 165919
rect 88670 165909 88750 165919
rect 87690 165829 87700 165909
rect 88010 165829 88020 165909
rect 88430 165829 88440 165909
rect 88750 165829 88760 165909
rect 89140 165900 89150 165980
rect 89290 165900 89300 165980
rect 100640 165900 100650 165980
rect 100790 165900 100800 165980
rect 100940 165900 100950 165980
rect 101110 165909 101190 165919
rect 101430 165909 101510 165919
rect 101850 165909 101930 165919
rect 102170 165909 102250 165919
rect 114610 165909 114690 165919
rect 114930 165909 115010 165919
rect 115350 165909 115430 165919
rect 115670 165909 115750 165919
rect 101190 165829 101200 165909
rect 101510 165829 101520 165909
rect 101930 165829 101940 165909
rect 102250 165829 102260 165909
rect 114690 165829 114700 165909
rect 115010 165829 115020 165909
rect 115430 165829 115440 165909
rect 115750 165829 115760 165909
rect 116140 165900 116150 165980
rect 116290 165900 116300 165980
rect 127640 165900 127650 165980
rect 127790 165900 127800 165980
rect 127940 165900 127950 165980
rect 128110 165909 128190 165919
rect 128430 165909 128510 165919
rect 128850 165909 128930 165919
rect 129170 165909 129250 165919
rect 128190 165829 128200 165909
rect 128510 165829 128520 165909
rect 128930 165829 128940 165909
rect 129250 165829 129260 165909
rect 129640 165900 129650 165980
rect 129790 165900 129800 165980
rect 140730 165900 140740 165980
rect 141140 165900 141150 165980
rect 141290 165900 141300 165980
rect 141440 165900 141450 165980
rect 141825 165910 141905 165920
rect 142145 165910 142200 165920
rect 145345 165910 145425 165920
rect 145665 165910 145745 165920
rect 145985 165910 146065 165920
rect 141905 165830 141915 165910
rect 145425 165830 145435 165910
rect 145745 165830 145755 165910
rect 146065 165830 146075 165910
rect 146780 165900 146790 165980
rect 146540 165820 146620 165830
rect 146860 165820 146940 165830
rect 59350 165800 59430 165810
rect 59500 165800 59580 165810
rect 59650 165800 59730 165810
rect 60060 165800 60140 165810
rect 60210 165800 60290 165810
rect 60360 165800 60440 165810
rect 62060 165800 62140 165810
rect 62210 165800 62290 165810
rect 73560 165800 73640 165810
rect 73710 165800 73790 165810
rect 73860 165800 73940 165810
rect 75560 165800 75640 165810
rect 75710 165800 75790 165810
rect 87060 165800 87140 165810
rect 87210 165800 87290 165810
rect 87360 165800 87440 165810
rect 89060 165800 89140 165810
rect 89210 165800 89290 165810
rect 100560 165800 100640 165810
rect 100710 165800 100790 165810
rect 100860 165800 100940 165810
rect 116060 165800 116140 165810
rect 116210 165800 116290 165810
rect 127560 165800 127640 165810
rect 127710 165800 127790 165810
rect 127860 165800 127940 165810
rect 129560 165800 129640 165810
rect 129710 165800 129790 165810
rect 140710 165800 140730 165810
rect 141060 165800 141140 165810
rect 141210 165800 141290 165810
rect 141360 165800 141440 165810
rect 59430 165720 59440 165800
rect 59580 165720 59590 165800
rect 59730 165720 59740 165800
rect 60140 165720 60150 165800
rect 60290 165720 60300 165800
rect 60440 165720 60450 165800
rect 60770 165749 60850 165759
rect 61090 165749 61170 165759
rect 61510 165749 61590 165759
rect 61830 165749 61910 165759
rect 60850 165669 60860 165749
rect 61170 165669 61180 165749
rect 61590 165669 61600 165749
rect 61910 165669 61920 165749
rect 62140 165720 62150 165800
rect 62290 165720 62300 165800
rect 73640 165720 73650 165800
rect 73790 165720 73800 165800
rect 73940 165720 73950 165800
rect 74270 165749 74350 165759
rect 74590 165749 74670 165759
rect 75010 165749 75090 165759
rect 75330 165749 75410 165759
rect 74350 165669 74360 165749
rect 74670 165669 74680 165749
rect 75090 165669 75100 165749
rect 75410 165669 75420 165749
rect 75640 165720 75650 165800
rect 75790 165720 75800 165800
rect 87140 165720 87150 165800
rect 87290 165720 87300 165800
rect 87440 165720 87450 165800
rect 87770 165749 87850 165759
rect 88090 165749 88170 165759
rect 88510 165749 88590 165759
rect 88830 165749 88910 165759
rect 87850 165669 87860 165749
rect 88170 165669 88180 165749
rect 88590 165669 88600 165749
rect 88910 165669 88920 165749
rect 89140 165720 89150 165800
rect 89290 165720 89300 165800
rect 100640 165720 100650 165800
rect 100790 165720 100800 165800
rect 100940 165720 100950 165800
rect 101270 165749 101350 165759
rect 101590 165749 101670 165759
rect 102010 165749 102090 165759
rect 102330 165749 102410 165759
rect 114770 165749 114850 165759
rect 115090 165749 115170 165759
rect 115510 165749 115590 165759
rect 115830 165749 115910 165759
rect 101350 165669 101360 165749
rect 101670 165669 101680 165749
rect 102090 165669 102100 165749
rect 102410 165669 102420 165749
rect 114850 165669 114860 165749
rect 115170 165669 115180 165749
rect 115590 165669 115600 165749
rect 115910 165669 115920 165749
rect 116140 165720 116150 165800
rect 116290 165720 116300 165800
rect 127640 165720 127650 165800
rect 127790 165720 127800 165800
rect 127940 165720 127950 165800
rect 128270 165749 128350 165759
rect 128590 165749 128670 165759
rect 129010 165749 129090 165759
rect 129330 165749 129410 165759
rect 128350 165669 128360 165749
rect 128670 165669 128680 165749
rect 129090 165669 129100 165749
rect 129410 165669 129420 165749
rect 129640 165720 129650 165800
rect 129790 165720 129800 165800
rect 140730 165720 140740 165800
rect 141140 165720 141150 165800
rect 141290 165720 141300 165800
rect 141440 165720 141450 165800
rect 141665 165750 141745 165760
rect 141985 165750 142065 165760
rect 145200 165750 145265 165760
rect 145505 165750 145585 165760
rect 145825 165750 145905 165760
rect 141745 165670 141755 165750
rect 142065 165670 142075 165750
rect 145265 165670 145275 165750
rect 145585 165670 145595 165750
rect 145905 165670 145915 165750
rect 146620 165740 146630 165820
rect 146940 165740 146950 165820
rect 146700 165660 146780 165670
rect 59350 165620 59430 165630
rect 59500 165620 59580 165630
rect 59650 165620 59730 165630
rect 60060 165620 60140 165630
rect 60210 165620 60290 165630
rect 60360 165620 60440 165630
rect 62060 165620 62140 165630
rect 62210 165620 62290 165630
rect 73560 165620 73640 165630
rect 73710 165620 73790 165630
rect 73860 165620 73940 165630
rect 75560 165620 75640 165630
rect 75710 165620 75790 165630
rect 87060 165620 87140 165630
rect 87210 165620 87290 165630
rect 87360 165620 87440 165630
rect 89060 165620 89140 165630
rect 89210 165620 89290 165630
rect 100560 165620 100640 165630
rect 100710 165620 100790 165630
rect 100860 165620 100940 165630
rect 116060 165620 116140 165630
rect 116210 165620 116290 165630
rect 127560 165620 127640 165630
rect 127710 165620 127790 165630
rect 127860 165620 127940 165630
rect 129560 165620 129640 165630
rect 129710 165620 129790 165630
rect 140710 165620 140730 165630
rect 141060 165620 141140 165630
rect 141210 165620 141290 165630
rect 141360 165620 141440 165630
rect 59430 165540 59440 165620
rect 59580 165540 59590 165620
rect 59730 165540 59740 165620
rect 60140 165540 60150 165620
rect 60290 165540 60300 165620
rect 60440 165540 60450 165620
rect 60610 165589 60690 165599
rect 60930 165589 61010 165599
rect 61350 165589 61430 165599
rect 61670 165589 61750 165599
rect 60690 165509 60700 165589
rect 61010 165509 61020 165589
rect 61430 165509 61440 165589
rect 61750 165509 61760 165589
rect 62140 165540 62150 165620
rect 62290 165540 62300 165620
rect 73640 165540 73650 165620
rect 73790 165540 73800 165620
rect 73940 165540 73950 165620
rect 74110 165589 74190 165599
rect 74430 165589 74510 165599
rect 74850 165589 74930 165599
rect 75170 165589 75250 165599
rect 74190 165509 74200 165589
rect 74510 165509 74520 165589
rect 74930 165509 74940 165589
rect 75250 165509 75260 165589
rect 75640 165540 75650 165620
rect 75790 165540 75800 165620
rect 87140 165540 87150 165620
rect 87290 165540 87300 165620
rect 87440 165540 87450 165620
rect 87610 165589 87690 165599
rect 87930 165589 88010 165599
rect 88350 165589 88430 165599
rect 88670 165589 88750 165599
rect 87690 165509 87700 165589
rect 88010 165509 88020 165589
rect 88430 165509 88440 165589
rect 88750 165509 88760 165589
rect 89140 165540 89150 165620
rect 89290 165540 89300 165620
rect 100640 165540 100650 165620
rect 100790 165540 100800 165620
rect 100940 165540 100950 165620
rect 101110 165589 101190 165599
rect 101430 165589 101510 165599
rect 101850 165589 101930 165599
rect 102170 165589 102250 165599
rect 114610 165589 114690 165599
rect 114930 165589 115010 165599
rect 115350 165589 115430 165599
rect 115670 165589 115750 165599
rect 101190 165509 101200 165589
rect 101510 165509 101520 165589
rect 101930 165509 101940 165589
rect 102250 165509 102260 165589
rect 114690 165509 114700 165589
rect 115010 165509 115020 165589
rect 115430 165509 115440 165589
rect 115750 165509 115760 165589
rect 116140 165540 116150 165620
rect 116290 165540 116300 165620
rect 127640 165540 127650 165620
rect 127790 165540 127800 165620
rect 127940 165540 127950 165620
rect 128110 165589 128190 165599
rect 128430 165589 128510 165599
rect 128850 165589 128930 165599
rect 129170 165589 129250 165599
rect 128190 165509 128200 165589
rect 128510 165509 128520 165589
rect 128930 165509 128940 165589
rect 129250 165509 129260 165589
rect 129640 165540 129650 165620
rect 129790 165540 129800 165620
rect 140730 165540 140740 165620
rect 141140 165540 141150 165620
rect 141290 165540 141300 165620
rect 141440 165540 141450 165620
rect 141825 165590 141905 165600
rect 142145 165590 142200 165600
rect 145345 165590 145425 165600
rect 145665 165590 145745 165600
rect 145985 165590 146065 165600
rect 141905 165510 141915 165590
rect 145425 165510 145435 165590
rect 145745 165510 145755 165590
rect 146065 165510 146075 165590
rect 146780 165580 146790 165660
rect 146540 165500 146620 165510
rect 146860 165500 146940 165510
rect 59350 165440 59430 165450
rect 59500 165440 59580 165450
rect 59650 165440 59730 165450
rect 60060 165440 60140 165450
rect 60210 165440 60290 165450
rect 60360 165440 60440 165450
rect 62060 165440 62140 165450
rect 62210 165440 62290 165450
rect 73560 165440 73640 165450
rect 73710 165440 73790 165450
rect 73860 165440 73940 165450
rect 75560 165440 75640 165450
rect 75710 165440 75790 165450
rect 87060 165440 87140 165450
rect 87210 165440 87290 165450
rect 87360 165440 87440 165450
rect 89060 165440 89140 165450
rect 89210 165440 89290 165450
rect 100560 165440 100640 165450
rect 100710 165440 100790 165450
rect 100860 165440 100940 165450
rect 116060 165440 116140 165450
rect 116210 165440 116290 165450
rect 127560 165440 127640 165450
rect 127710 165440 127790 165450
rect 127860 165440 127940 165450
rect 129560 165440 129640 165450
rect 129710 165440 129790 165450
rect 140710 165440 140730 165450
rect 141060 165440 141140 165450
rect 141210 165440 141290 165450
rect 141360 165440 141440 165450
rect 59430 165360 59440 165440
rect 59580 165360 59590 165440
rect 59730 165360 59740 165440
rect 60140 165360 60150 165440
rect 60290 165360 60300 165440
rect 60440 165360 60450 165440
rect 60770 165429 60850 165439
rect 61090 165429 61170 165439
rect 61510 165429 61590 165439
rect 61830 165429 61910 165439
rect 60850 165349 60860 165429
rect 61170 165349 61180 165429
rect 61590 165349 61600 165429
rect 61910 165349 61920 165429
rect 62140 165360 62150 165440
rect 62290 165360 62300 165440
rect 73640 165360 73650 165440
rect 73790 165360 73800 165440
rect 73940 165360 73950 165440
rect 74270 165429 74350 165439
rect 74590 165429 74670 165439
rect 75010 165429 75090 165439
rect 75330 165429 75410 165439
rect 74350 165349 74360 165429
rect 74670 165349 74680 165429
rect 75090 165349 75100 165429
rect 75410 165349 75420 165429
rect 75640 165360 75650 165440
rect 75790 165360 75800 165440
rect 87140 165360 87150 165440
rect 87290 165360 87300 165440
rect 87440 165360 87450 165440
rect 87770 165429 87850 165439
rect 88090 165429 88170 165439
rect 88510 165429 88590 165439
rect 88830 165429 88910 165439
rect 87850 165349 87860 165429
rect 88170 165349 88180 165429
rect 88590 165349 88600 165429
rect 88910 165349 88920 165429
rect 89140 165360 89150 165440
rect 89290 165360 89300 165440
rect 100640 165360 100650 165440
rect 100790 165360 100800 165440
rect 100940 165360 100950 165440
rect 101270 165429 101350 165439
rect 101590 165429 101670 165439
rect 102010 165429 102090 165439
rect 102330 165429 102410 165439
rect 114770 165429 114850 165439
rect 115090 165429 115170 165439
rect 115510 165429 115590 165439
rect 115830 165429 115910 165439
rect 101350 165349 101360 165429
rect 101670 165349 101680 165429
rect 102090 165349 102100 165429
rect 102410 165349 102420 165429
rect 114850 165349 114860 165429
rect 115170 165349 115180 165429
rect 115590 165349 115600 165429
rect 115910 165349 115920 165429
rect 116140 165360 116150 165440
rect 116290 165360 116300 165440
rect 127640 165360 127650 165440
rect 127790 165360 127800 165440
rect 127940 165360 127950 165440
rect 128270 165429 128350 165439
rect 128590 165429 128670 165439
rect 129010 165429 129090 165439
rect 129330 165429 129410 165439
rect 128350 165349 128360 165429
rect 128670 165349 128680 165429
rect 129090 165349 129100 165429
rect 129410 165349 129420 165429
rect 129640 165360 129650 165440
rect 129790 165360 129800 165440
rect 140730 165360 140740 165440
rect 141140 165360 141150 165440
rect 141290 165360 141300 165440
rect 141440 165360 141450 165440
rect 141665 165430 141745 165440
rect 141985 165430 142065 165440
rect 145200 165430 145265 165440
rect 145505 165430 145585 165440
rect 145825 165430 145905 165440
rect 141745 165350 141755 165430
rect 142065 165350 142075 165430
rect 145265 165350 145275 165430
rect 145585 165350 145595 165430
rect 145905 165350 145915 165430
rect 146620 165420 146630 165500
rect 146940 165420 146950 165500
rect 146700 165340 146780 165350
rect 59350 165260 59430 165270
rect 59500 165260 59580 165270
rect 59650 165260 59730 165270
rect 60060 165260 60140 165270
rect 60210 165260 60290 165270
rect 60360 165260 60440 165270
rect 60610 165269 60690 165279
rect 60930 165269 61010 165279
rect 61350 165269 61430 165279
rect 61670 165269 61750 165279
rect 59430 165180 59440 165260
rect 59580 165180 59590 165260
rect 59730 165180 59740 165260
rect 60140 165180 60150 165260
rect 60290 165180 60300 165260
rect 60440 165180 60450 165260
rect 60690 165189 60700 165269
rect 61010 165189 61020 165269
rect 61430 165189 61440 165269
rect 61750 165189 61760 165269
rect 62060 165260 62140 165270
rect 62210 165260 62290 165270
rect 73560 165260 73640 165270
rect 73710 165260 73790 165270
rect 73860 165260 73940 165270
rect 74110 165269 74190 165279
rect 74430 165269 74510 165279
rect 74850 165269 74930 165279
rect 75170 165269 75250 165279
rect 62140 165180 62150 165260
rect 62290 165180 62300 165260
rect 73640 165180 73650 165260
rect 73790 165180 73800 165260
rect 73940 165180 73950 165260
rect 74190 165189 74200 165269
rect 74510 165189 74520 165269
rect 74930 165189 74940 165269
rect 75250 165189 75260 165269
rect 75560 165260 75640 165270
rect 75710 165260 75790 165270
rect 87060 165260 87140 165270
rect 87210 165260 87290 165270
rect 87360 165260 87440 165270
rect 87610 165269 87690 165279
rect 87930 165269 88010 165279
rect 88350 165269 88430 165279
rect 88670 165269 88750 165279
rect 75640 165180 75650 165260
rect 75790 165180 75800 165260
rect 87140 165180 87150 165260
rect 87290 165180 87300 165260
rect 87440 165180 87450 165260
rect 87690 165189 87700 165269
rect 88010 165189 88020 165269
rect 88430 165189 88440 165269
rect 88750 165189 88760 165269
rect 89060 165260 89140 165270
rect 89210 165260 89290 165270
rect 100560 165260 100640 165270
rect 100710 165260 100790 165270
rect 100860 165260 100940 165270
rect 101110 165269 101190 165279
rect 101430 165269 101510 165279
rect 101850 165269 101930 165279
rect 102170 165269 102250 165279
rect 114610 165269 114690 165279
rect 114930 165269 115010 165279
rect 115350 165269 115430 165279
rect 115670 165269 115750 165279
rect 89140 165180 89150 165260
rect 89290 165180 89300 165260
rect 100640 165180 100650 165260
rect 100790 165180 100800 165260
rect 100940 165180 100950 165260
rect 101190 165189 101200 165269
rect 101510 165189 101520 165269
rect 101930 165189 101940 165269
rect 102250 165189 102260 165269
rect 114690 165189 114700 165269
rect 115010 165189 115020 165269
rect 115430 165189 115440 165269
rect 115750 165189 115760 165269
rect 116060 165260 116140 165270
rect 116210 165260 116290 165270
rect 127560 165260 127640 165270
rect 127710 165260 127790 165270
rect 127860 165260 127940 165270
rect 128110 165269 128190 165279
rect 128430 165269 128510 165279
rect 128850 165269 128930 165279
rect 129170 165269 129250 165279
rect 141825 165270 141905 165280
rect 142145 165270 142200 165280
rect 145345 165270 145425 165280
rect 145665 165270 145745 165280
rect 145985 165270 146065 165280
rect 116140 165180 116150 165260
rect 116290 165180 116300 165260
rect 127640 165180 127650 165260
rect 127790 165180 127800 165260
rect 127940 165180 127950 165260
rect 128190 165189 128200 165269
rect 128510 165189 128520 165269
rect 128930 165189 128940 165269
rect 129250 165189 129260 165269
rect 129560 165260 129640 165270
rect 129710 165260 129790 165270
rect 140710 165260 140730 165270
rect 141060 165260 141140 165270
rect 141210 165260 141290 165270
rect 141360 165260 141440 165270
rect 129640 165180 129650 165260
rect 129790 165180 129800 165260
rect 140730 165180 140740 165260
rect 141140 165180 141150 165260
rect 141290 165180 141300 165260
rect 141440 165180 141450 165260
rect 141905 165190 141915 165270
rect 145425 165190 145435 165270
rect 145745 165190 145755 165270
rect 146065 165190 146075 165270
rect 146780 165260 146790 165340
rect 146540 165180 146620 165190
rect 146860 165180 146940 165190
rect 60770 165109 60850 165119
rect 61090 165109 61170 165119
rect 61510 165109 61590 165119
rect 61830 165109 61910 165119
rect 74270 165109 74350 165119
rect 74590 165109 74670 165119
rect 75010 165109 75090 165119
rect 75330 165109 75410 165119
rect 87770 165109 87850 165119
rect 88090 165109 88170 165119
rect 88510 165109 88590 165119
rect 88830 165109 88910 165119
rect 101270 165109 101350 165119
rect 101590 165109 101670 165119
rect 102010 165109 102090 165119
rect 102330 165109 102410 165119
rect 114770 165109 114850 165119
rect 115090 165109 115170 165119
rect 115510 165109 115590 165119
rect 115830 165109 115910 165119
rect 128270 165109 128350 165119
rect 128590 165109 128670 165119
rect 129010 165109 129090 165119
rect 129330 165109 129410 165119
rect 141665 165110 141745 165120
rect 141985 165110 142065 165120
rect 145200 165110 145265 165120
rect 145505 165110 145585 165120
rect 145825 165110 145905 165120
rect 59350 165080 59430 165090
rect 59500 165080 59580 165090
rect 59650 165080 59730 165090
rect 60060 165080 60140 165090
rect 60210 165080 60290 165090
rect 60360 165080 60440 165090
rect 59430 165000 59440 165080
rect 59580 165000 59590 165080
rect 59730 165000 59740 165080
rect 60140 165000 60150 165080
rect 60290 165000 60300 165080
rect 60440 165000 60450 165080
rect 60850 165029 60860 165109
rect 61170 165029 61180 165109
rect 61590 165029 61600 165109
rect 61910 165029 61920 165109
rect 62060 165080 62140 165090
rect 62210 165080 62290 165090
rect 73560 165080 73640 165090
rect 73710 165080 73790 165090
rect 73860 165080 73940 165090
rect 62140 165000 62150 165080
rect 62290 165000 62300 165080
rect 73640 165000 73650 165080
rect 73790 165000 73800 165080
rect 73940 165000 73950 165080
rect 74350 165029 74360 165109
rect 74670 165029 74680 165109
rect 75090 165029 75100 165109
rect 75410 165029 75420 165109
rect 75560 165080 75640 165090
rect 75710 165080 75790 165090
rect 87060 165080 87140 165090
rect 87210 165080 87290 165090
rect 87360 165080 87440 165090
rect 75640 165000 75650 165080
rect 75790 165000 75800 165080
rect 87140 165000 87150 165080
rect 87290 165000 87300 165080
rect 87440 165000 87450 165080
rect 87850 165029 87860 165109
rect 88170 165029 88180 165109
rect 88590 165029 88600 165109
rect 88910 165029 88920 165109
rect 89060 165080 89140 165090
rect 89210 165080 89290 165090
rect 100560 165080 100640 165090
rect 100710 165080 100790 165090
rect 100860 165080 100940 165090
rect 89140 165000 89150 165080
rect 89290 165000 89300 165080
rect 100640 165000 100650 165080
rect 100790 165000 100800 165080
rect 100940 165000 100950 165080
rect 101350 165029 101360 165109
rect 101670 165029 101680 165109
rect 102090 165029 102100 165109
rect 102410 165029 102420 165109
rect 114850 165029 114860 165109
rect 115170 165029 115180 165109
rect 115590 165029 115600 165109
rect 115910 165029 115920 165109
rect 116060 165080 116140 165090
rect 116210 165080 116290 165090
rect 127560 165080 127640 165090
rect 127710 165080 127790 165090
rect 127860 165080 127940 165090
rect 116140 165000 116150 165080
rect 116290 165000 116300 165080
rect 127640 165000 127650 165080
rect 127790 165000 127800 165080
rect 127940 165000 127950 165080
rect 128350 165029 128360 165109
rect 128670 165029 128680 165109
rect 129090 165029 129100 165109
rect 129410 165029 129420 165109
rect 129560 165080 129640 165090
rect 129710 165080 129790 165090
rect 140710 165080 140730 165090
rect 141060 165080 141140 165090
rect 141210 165080 141290 165090
rect 141360 165080 141440 165090
rect 129640 165000 129650 165080
rect 129790 165000 129800 165080
rect 140730 165000 140740 165080
rect 141140 165000 141150 165080
rect 141290 165000 141300 165080
rect 141440 165000 141450 165080
rect 141745 165030 141755 165110
rect 142065 165030 142075 165110
rect 145265 165030 145275 165110
rect 145585 165030 145595 165110
rect 145905 165030 145915 165110
rect 146620 165100 146630 165180
rect 146940 165100 146950 165180
rect 146700 165020 146780 165030
rect 60610 164949 60690 164959
rect 60930 164949 61010 164959
rect 61350 164949 61430 164959
rect 61670 164949 61750 164959
rect 74110 164949 74190 164959
rect 74430 164949 74510 164959
rect 74850 164949 74930 164959
rect 75170 164949 75250 164959
rect 87610 164949 87690 164959
rect 87930 164949 88010 164959
rect 88350 164949 88430 164959
rect 88670 164949 88750 164959
rect 101110 164949 101190 164959
rect 101430 164949 101510 164959
rect 101850 164949 101930 164959
rect 102170 164949 102250 164959
rect 114610 164949 114690 164959
rect 114930 164949 115010 164959
rect 115350 164949 115430 164959
rect 115670 164949 115750 164959
rect 128110 164949 128190 164959
rect 128430 164949 128510 164959
rect 128850 164949 128930 164959
rect 129170 164949 129250 164959
rect 141825 164950 141905 164960
rect 142145 164950 142200 164960
rect 145345 164950 145425 164960
rect 145665 164950 145745 164960
rect 145985 164950 146065 164960
rect 59350 164900 59430 164910
rect 59500 164900 59580 164910
rect 59650 164900 59730 164910
rect 60060 164900 60140 164910
rect 60210 164900 60290 164910
rect 60360 164900 60440 164910
rect 59430 164820 59440 164900
rect 59580 164820 59590 164900
rect 59730 164820 59740 164900
rect 60140 164820 60150 164900
rect 60290 164820 60300 164900
rect 60440 164820 60450 164900
rect 60690 164869 60700 164949
rect 61010 164869 61020 164949
rect 61430 164869 61440 164949
rect 61750 164869 61760 164949
rect 62060 164900 62140 164910
rect 62210 164900 62290 164910
rect 73560 164900 73640 164910
rect 73710 164900 73790 164910
rect 73860 164900 73940 164910
rect 62140 164820 62150 164900
rect 62290 164820 62300 164900
rect 73640 164820 73650 164900
rect 73790 164820 73800 164900
rect 73940 164820 73950 164900
rect 74190 164869 74200 164949
rect 74510 164869 74520 164949
rect 74930 164869 74940 164949
rect 75250 164869 75260 164949
rect 75560 164900 75640 164910
rect 75710 164900 75790 164910
rect 87060 164900 87140 164910
rect 87210 164900 87290 164910
rect 87360 164900 87440 164910
rect 75640 164820 75650 164900
rect 75790 164820 75800 164900
rect 87140 164820 87150 164900
rect 87290 164820 87300 164900
rect 87440 164820 87450 164900
rect 87690 164869 87700 164949
rect 88010 164869 88020 164949
rect 88430 164869 88440 164949
rect 88750 164869 88760 164949
rect 89060 164900 89140 164910
rect 89210 164900 89290 164910
rect 100560 164900 100640 164910
rect 100710 164900 100790 164910
rect 100860 164900 100940 164910
rect 89140 164820 89150 164900
rect 89290 164820 89300 164900
rect 100640 164820 100650 164900
rect 100790 164820 100800 164900
rect 100940 164820 100950 164900
rect 101190 164869 101200 164949
rect 101510 164869 101520 164949
rect 101930 164869 101940 164949
rect 102250 164869 102260 164949
rect 114690 164869 114700 164949
rect 115010 164869 115020 164949
rect 115430 164869 115440 164949
rect 115750 164869 115760 164949
rect 116060 164900 116140 164910
rect 116210 164900 116290 164910
rect 127560 164900 127640 164910
rect 127710 164900 127790 164910
rect 127860 164900 127940 164910
rect 116140 164820 116150 164900
rect 116290 164820 116300 164900
rect 127640 164820 127650 164900
rect 127790 164820 127800 164900
rect 127940 164820 127950 164900
rect 128190 164869 128200 164949
rect 128510 164869 128520 164949
rect 128930 164869 128940 164949
rect 129250 164869 129260 164949
rect 129560 164900 129640 164910
rect 129710 164900 129790 164910
rect 140710 164900 140730 164910
rect 141060 164900 141140 164910
rect 141210 164900 141290 164910
rect 141360 164900 141440 164910
rect 129640 164820 129650 164900
rect 129790 164820 129800 164900
rect 140730 164820 140740 164900
rect 141140 164820 141150 164900
rect 141290 164820 141300 164900
rect 141440 164820 141450 164900
rect 141905 164870 141915 164950
rect 145425 164870 145435 164950
rect 145745 164870 145755 164950
rect 146065 164870 146075 164950
rect 146780 164940 146790 165020
rect 146540 164860 146620 164870
rect 146860 164860 146940 164870
rect 60770 164789 60850 164799
rect 61090 164789 61170 164799
rect 61510 164789 61590 164799
rect 61830 164789 61910 164799
rect 74270 164789 74350 164799
rect 74590 164789 74670 164799
rect 75010 164789 75090 164799
rect 75330 164789 75410 164799
rect 87770 164789 87850 164799
rect 88090 164789 88170 164799
rect 88510 164789 88590 164799
rect 88830 164789 88910 164799
rect 101270 164789 101350 164799
rect 101590 164789 101670 164799
rect 102010 164789 102090 164799
rect 102330 164789 102410 164799
rect 114770 164789 114850 164799
rect 115090 164789 115170 164799
rect 115510 164789 115590 164799
rect 115830 164789 115910 164799
rect 128270 164789 128350 164799
rect 128590 164789 128670 164799
rect 129010 164789 129090 164799
rect 129330 164789 129410 164799
rect 141665 164790 141745 164800
rect 141985 164790 142065 164800
rect 145200 164790 145265 164800
rect 145505 164790 145585 164800
rect 145825 164790 145905 164800
rect 59350 164720 59430 164730
rect 59500 164720 59580 164730
rect 59650 164720 59730 164730
rect 60060 164720 60140 164730
rect 60210 164720 60290 164730
rect 60360 164720 60440 164730
rect 59430 164640 59440 164720
rect 59580 164640 59590 164720
rect 59730 164640 59740 164720
rect 60140 164640 60150 164720
rect 60290 164640 60300 164720
rect 60440 164640 60450 164720
rect 60850 164709 60860 164789
rect 61170 164709 61180 164789
rect 61590 164709 61600 164789
rect 61910 164709 61920 164789
rect 62060 164720 62140 164730
rect 62210 164720 62290 164730
rect 73560 164720 73640 164730
rect 73710 164720 73790 164730
rect 73860 164720 73940 164730
rect 62140 164640 62150 164720
rect 62290 164640 62300 164720
rect 73640 164640 73650 164720
rect 73790 164640 73800 164720
rect 73940 164640 73950 164720
rect 74350 164709 74360 164789
rect 74670 164709 74680 164789
rect 75090 164709 75100 164789
rect 75410 164709 75420 164789
rect 75560 164720 75640 164730
rect 75710 164720 75790 164730
rect 87060 164720 87140 164730
rect 87210 164720 87290 164730
rect 87360 164720 87440 164730
rect 75640 164640 75650 164720
rect 75790 164640 75800 164720
rect 87140 164640 87150 164720
rect 87290 164640 87300 164720
rect 87440 164640 87450 164720
rect 87850 164709 87860 164789
rect 88170 164709 88180 164789
rect 88590 164709 88600 164789
rect 88910 164709 88920 164789
rect 89060 164720 89140 164730
rect 89210 164720 89290 164730
rect 100560 164720 100640 164730
rect 100710 164720 100790 164730
rect 100860 164720 100940 164730
rect 89140 164640 89150 164720
rect 89290 164640 89300 164720
rect 100640 164640 100650 164720
rect 100790 164640 100800 164720
rect 100940 164640 100950 164720
rect 101350 164709 101360 164789
rect 101670 164709 101680 164789
rect 102090 164709 102100 164789
rect 102410 164709 102420 164789
rect 114850 164709 114860 164789
rect 115170 164709 115180 164789
rect 115590 164709 115600 164789
rect 115910 164709 115920 164789
rect 116060 164720 116140 164730
rect 116210 164720 116290 164730
rect 127560 164720 127640 164730
rect 127710 164720 127790 164730
rect 127860 164720 127940 164730
rect 116140 164640 116150 164720
rect 116290 164640 116300 164720
rect 127640 164640 127650 164720
rect 127790 164640 127800 164720
rect 127940 164640 127950 164720
rect 128350 164709 128360 164789
rect 128670 164709 128680 164789
rect 129090 164709 129100 164789
rect 129410 164709 129420 164789
rect 129560 164720 129640 164730
rect 129710 164720 129790 164730
rect 140710 164720 140730 164730
rect 141060 164720 141140 164730
rect 141210 164720 141290 164730
rect 141360 164720 141440 164730
rect 129640 164640 129650 164720
rect 129790 164640 129800 164720
rect 140730 164640 140740 164720
rect 141140 164640 141150 164720
rect 141290 164640 141300 164720
rect 141440 164640 141450 164720
rect 141745 164710 141755 164790
rect 142065 164710 142075 164790
rect 145265 164710 145275 164790
rect 145585 164710 145595 164790
rect 145905 164710 145915 164790
rect 146620 164780 146630 164860
rect 146940 164780 146950 164860
rect 146700 164700 146780 164710
rect 60610 164629 60690 164639
rect 60930 164629 61010 164639
rect 61350 164629 61430 164639
rect 61670 164629 61750 164639
rect 74110 164629 74190 164639
rect 74430 164629 74510 164639
rect 74850 164629 74930 164639
rect 75170 164629 75250 164639
rect 87610 164629 87690 164639
rect 87930 164629 88010 164639
rect 88350 164629 88430 164639
rect 88670 164629 88750 164639
rect 101110 164629 101190 164639
rect 101430 164629 101510 164639
rect 101850 164629 101930 164639
rect 102170 164629 102250 164639
rect 114610 164629 114690 164639
rect 114930 164629 115010 164639
rect 115350 164629 115430 164639
rect 115670 164629 115750 164639
rect 128110 164629 128190 164639
rect 128430 164629 128510 164639
rect 128850 164629 128930 164639
rect 129170 164629 129250 164639
rect 141825 164630 141905 164640
rect 142145 164630 142200 164640
rect 145345 164630 145425 164640
rect 145665 164630 145745 164640
rect 145985 164630 146065 164640
rect 59350 164540 59430 164550
rect 59500 164540 59580 164550
rect 59650 164540 59730 164550
rect 60060 164540 60140 164550
rect 60210 164540 60290 164550
rect 60360 164540 60440 164550
rect 60690 164549 60700 164629
rect 61010 164549 61020 164629
rect 61430 164549 61440 164629
rect 61750 164549 61760 164629
rect 62060 164540 62140 164550
rect 62210 164540 62290 164550
rect 73560 164540 73640 164550
rect 73710 164540 73790 164550
rect 73860 164540 73940 164550
rect 74190 164549 74200 164629
rect 74510 164549 74520 164629
rect 74930 164549 74940 164629
rect 75250 164549 75260 164629
rect 75560 164540 75640 164550
rect 75710 164540 75790 164550
rect 87060 164540 87140 164550
rect 87210 164540 87290 164550
rect 87360 164540 87440 164550
rect 87690 164549 87700 164629
rect 88010 164549 88020 164629
rect 88430 164549 88440 164629
rect 88750 164549 88760 164629
rect 89060 164540 89140 164550
rect 89210 164540 89290 164550
rect 100560 164540 100640 164550
rect 100710 164540 100790 164550
rect 100860 164540 100940 164550
rect 101190 164549 101200 164629
rect 101510 164549 101520 164629
rect 101930 164549 101940 164629
rect 102250 164549 102260 164629
rect 114690 164549 114700 164629
rect 115010 164549 115020 164629
rect 115430 164549 115440 164629
rect 115750 164549 115760 164629
rect 116060 164540 116140 164550
rect 116210 164540 116290 164550
rect 127560 164540 127640 164550
rect 127710 164540 127790 164550
rect 127860 164540 127940 164550
rect 128190 164549 128200 164629
rect 128510 164549 128520 164629
rect 128930 164549 128940 164629
rect 129250 164549 129260 164629
rect 141905 164550 141915 164630
rect 145425 164550 145435 164630
rect 145745 164550 145755 164630
rect 146065 164550 146075 164630
rect 146780 164620 146790 164700
rect 129560 164540 129640 164550
rect 129710 164540 129790 164550
rect 140710 164540 140730 164550
rect 141060 164540 141140 164550
rect 141210 164540 141290 164550
rect 141360 164540 141440 164550
rect 146540 164540 146620 164550
rect 146860 164540 146940 164550
rect 59430 164460 59440 164540
rect 59580 164460 59590 164540
rect 59730 164460 59740 164540
rect 60140 164460 60150 164540
rect 60290 164460 60300 164540
rect 60440 164460 60450 164540
rect 60770 164469 60850 164479
rect 61090 164469 61170 164479
rect 61510 164469 61590 164479
rect 61830 164469 61910 164479
rect 60850 164389 60860 164469
rect 61170 164389 61180 164469
rect 61590 164389 61600 164469
rect 61910 164389 61920 164469
rect 62140 164460 62150 164540
rect 62290 164460 62300 164540
rect 73640 164460 73650 164540
rect 73790 164460 73800 164540
rect 73940 164460 73950 164540
rect 74270 164469 74350 164479
rect 74590 164469 74670 164479
rect 75010 164469 75090 164479
rect 75330 164469 75410 164479
rect 74350 164389 74360 164469
rect 74670 164389 74680 164469
rect 75090 164389 75100 164469
rect 75410 164389 75420 164469
rect 75640 164460 75650 164540
rect 75790 164460 75800 164540
rect 87140 164460 87150 164540
rect 87290 164460 87300 164540
rect 87440 164460 87450 164540
rect 87770 164469 87850 164479
rect 88090 164469 88170 164479
rect 88510 164469 88590 164479
rect 88830 164469 88910 164479
rect 87850 164389 87860 164469
rect 88170 164389 88180 164469
rect 88590 164389 88600 164469
rect 88910 164389 88920 164469
rect 89140 164460 89150 164540
rect 89290 164460 89300 164540
rect 100640 164460 100650 164540
rect 100790 164460 100800 164540
rect 100940 164460 100950 164540
rect 101270 164469 101350 164479
rect 101590 164469 101670 164479
rect 102010 164469 102090 164479
rect 102330 164469 102410 164479
rect 114770 164469 114850 164479
rect 115090 164469 115170 164479
rect 115510 164469 115590 164479
rect 115830 164469 115910 164479
rect 101350 164389 101360 164469
rect 101670 164389 101680 164469
rect 102090 164389 102100 164469
rect 102410 164389 102420 164469
rect 114850 164389 114860 164469
rect 115170 164389 115180 164469
rect 115590 164389 115600 164469
rect 115910 164389 115920 164469
rect 116140 164460 116150 164540
rect 116290 164460 116300 164540
rect 127640 164460 127650 164540
rect 127790 164460 127800 164540
rect 127940 164460 127950 164540
rect 128270 164469 128350 164479
rect 128590 164469 128670 164479
rect 129010 164469 129090 164479
rect 129330 164469 129410 164479
rect 128350 164389 128360 164469
rect 128670 164389 128680 164469
rect 129090 164389 129100 164469
rect 129410 164389 129420 164469
rect 129640 164460 129650 164540
rect 129790 164460 129800 164540
rect 140730 164460 140740 164540
rect 141140 164460 141150 164540
rect 141290 164460 141300 164540
rect 141440 164460 141450 164540
rect 141665 164470 141745 164480
rect 141985 164470 142065 164480
rect 145200 164470 145265 164480
rect 145505 164470 145585 164480
rect 145825 164470 145905 164480
rect 141745 164390 141755 164470
rect 142065 164390 142075 164470
rect 145265 164390 145275 164470
rect 145585 164390 145595 164470
rect 145905 164390 145915 164470
rect 146620 164460 146630 164540
rect 146940 164460 146950 164540
rect 146700 164380 146780 164390
rect 59350 164360 59430 164370
rect 59500 164360 59580 164370
rect 59650 164360 59730 164370
rect 60060 164360 60140 164370
rect 60210 164360 60290 164370
rect 60360 164360 60440 164370
rect 62060 164360 62140 164370
rect 62210 164360 62290 164370
rect 73560 164360 73640 164370
rect 73710 164360 73790 164370
rect 73860 164360 73940 164370
rect 75560 164360 75640 164370
rect 75710 164360 75790 164370
rect 87060 164360 87140 164370
rect 87210 164360 87290 164370
rect 87360 164360 87440 164370
rect 89060 164360 89140 164370
rect 89210 164360 89290 164370
rect 100560 164360 100640 164370
rect 100710 164360 100790 164370
rect 100860 164360 100940 164370
rect 116060 164360 116140 164370
rect 116210 164360 116290 164370
rect 127560 164360 127640 164370
rect 127710 164360 127790 164370
rect 127860 164360 127940 164370
rect 129560 164360 129640 164370
rect 129710 164360 129790 164370
rect 140710 164360 140730 164370
rect 141060 164360 141140 164370
rect 141210 164360 141290 164370
rect 141360 164360 141440 164370
rect 59430 164280 59440 164360
rect 59580 164280 59590 164360
rect 59730 164280 59740 164360
rect 60140 164280 60150 164360
rect 60290 164280 60300 164360
rect 60440 164280 60450 164360
rect 60610 164309 60690 164319
rect 60930 164309 61010 164319
rect 61350 164309 61430 164319
rect 61670 164309 61750 164319
rect 60690 164229 60700 164309
rect 61010 164229 61020 164309
rect 61430 164229 61440 164309
rect 61750 164229 61760 164309
rect 62140 164280 62150 164360
rect 62290 164280 62300 164360
rect 73640 164280 73650 164360
rect 73790 164280 73800 164360
rect 73940 164280 73950 164360
rect 74110 164309 74190 164319
rect 74430 164309 74510 164319
rect 74850 164309 74930 164319
rect 75170 164309 75250 164319
rect 74190 164229 74200 164309
rect 74510 164229 74520 164309
rect 74930 164229 74940 164309
rect 75250 164229 75260 164309
rect 75640 164280 75650 164360
rect 75790 164280 75800 164360
rect 87140 164280 87150 164360
rect 87290 164280 87300 164360
rect 87440 164280 87450 164360
rect 87610 164309 87690 164319
rect 87930 164309 88010 164319
rect 88350 164309 88430 164319
rect 88670 164309 88750 164319
rect 87690 164229 87700 164309
rect 88010 164229 88020 164309
rect 88430 164229 88440 164309
rect 88750 164229 88760 164309
rect 89140 164280 89150 164360
rect 89290 164280 89300 164360
rect 100640 164280 100650 164360
rect 100790 164280 100800 164360
rect 100940 164280 100950 164360
rect 101110 164309 101190 164319
rect 101430 164309 101510 164319
rect 101850 164309 101930 164319
rect 102170 164309 102250 164319
rect 114610 164309 114690 164319
rect 114930 164309 115010 164319
rect 115350 164309 115430 164319
rect 115670 164309 115750 164319
rect 101190 164229 101200 164309
rect 101510 164229 101520 164309
rect 101930 164229 101940 164309
rect 102250 164229 102260 164309
rect 114690 164229 114700 164309
rect 115010 164229 115020 164309
rect 115430 164229 115440 164309
rect 115750 164229 115760 164309
rect 116140 164280 116150 164360
rect 116290 164280 116300 164360
rect 127640 164280 127650 164360
rect 127790 164280 127800 164360
rect 127940 164280 127950 164360
rect 128110 164309 128190 164319
rect 128430 164309 128510 164319
rect 128850 164309 128930 164319
rect 129170 164309 129250 164319
rect 128190 164229 128200 164309
rect 128510 164229 128520 164309
rect 128930 164229 128940 164309
rect 129250 164229 129260 164309
rect 129640 164280 129650 164360
rect 129790 164280 129800 164360
rect 140730 164280 140740 164360
rect 141140 164280 141150 164360
rect 141290 164280 141300 164360
rect 141440 164280 141450 164360
rect 141825 164310 141905 164320
rect 142145 164310 142200 164320
rect 145345 164310 145425 164320
rect 145665 164310 145745 164320
rect 145985 164310 146065 164320
rect 141905 164230 141915 164310
rect 145425 164230 145435 164310
rect 145745 164230 145755 164310
rect 146065 164230 146075 164310
rect 146780 164300 146790 164380
rect 146540 164220 146620 164230
rect 146860 164220 146940 164230
rect 48500 164180 48640 164190
rect 48710 164180 48790 164190
rect 60060 164180 60140 164190
rect 60210 164180 60290 164190
rect 60360 164180 60440 164190
rect 62060 164180 62140 164190
rect 62210 164180 62290 164190
rect 73560 164180 73640 164190
rect 73710 164180 73790 164190
rect 73860 164180 73940 164190
rect 75560 164180 75640 164190
rect 75710 164180 75790 164190
rect 87060 164180 87140 164190
rect 87210 164180 87290 164190
rect 87360 164180 87440 164190
rect 89060 164180 89140 164190
rect 89210 164180 89290 164190
rect 100560 164180 100640 164190
rect 100710 164180 100790 164190
rect 100860 164180 100940 164190
rect 116060 164180 116140 164190
rect 116210 164180 116290 164190
rect 127560 164180 127640 164190
rect 127710 164180 127790 164190
rect 127860 164180 127940 164190
rect 129560 164180 129640 164190
rect 129710 164180 129790 164190
rect 141060 164180 141140 164190
rect 141210 164180 141290 164190
rect 141360 164180 141440 164190
rect 43905 164150 43985 164160
rect 44225 164150 44305 164160
rect 44545 164150 44625 164160
rect 44865 164150 44945 164160
rect 45185 164150 45265 164160
rect 45505 164150 45585 164160
rect 45825 164150 45905 164160
rect 46145 164150 46225 164160
rect 46465 164150 46545 164160
rect 46785 164150 46865 164160
rect 47105 164150 47185 164160
rect 47425 164150 47505 164160
rect 47745 164150 47825 164160
rect 48065 164150 48145 164160
rect 43985 164070 43995 164150
rect 44305 164070 44315 164150
rect 44625 164070 44635 164150
rect 44945 164070 44955 164150
rect 45265 164070 45275 164150
rect 45585 164070 45595 164150
rect 45905 164070 45915 164150
rect 46225 164070 46235 164150
rect 46545 164070 46555 164150
rect 46865 164070 46875 164150
rect 47185 164070 47195 164150
rect 47505 164070 47515 164150
rect 47825 164070 47835 164150
rect 48145 164070 48155 164150
rect 42950 164060 42980 164070
rect 43220 164060 43300 164070
rect 42980 163980 42990 164060
rect 43300 163980 43310 164060
rect 48500 164010 48605 164180
rect 48640 164100 48650 164180
rect 48790 164100 48800 164180
rect 60140 164100 60150 164180
rect 60290 164100 60300 164180
rect 60440 164100 60450 164180
rect 60770 164149 60850 164159
rect 61090 164149 61170 164159
rect 61510 164149 61590 164159
rect 61830 164149 61910 164159
rect 60850 164069 60860 164149
rect 61170 164069 61180 164149
rect 61590 164069 61600 164149
rect 61910 164069 61920 164149
rect 62140 164100 62150 164180
rect 62290 164100 62300 164180
rect 73640 164100 73650 164180
rect 73790 164100 73800 164180
rect 73940 164100 73950 164180
rect 74270 164149 74350 164159
rect 74590 164149 74670 164159
rect 75010 164149 75090 164159
rect 75330 164149 75410 164159
rect 74350 164069 74360 164149
rect 74670 164069 74680 164149
rect 75090 164069 75100 164149
rect 75410 164069 75420 164149
rect 75640 164100 75650 164180
rect 75790 164100 75800 164180
rect 87140 164100 87150 164180
rect 87290 164100 87300 164180
rect 87440 164100 87450 164180
rect 87770 164149 87850 164159
rect 88090 164149 88170 164159
rect 88510 164149 88590 164159
rect 88830 164149 88910 164159
rect 87850 164069 87860 164149
rect 88170 164069 88180 164149
rect 88590 164069 88600 164149
rect 88910 164069 88920 164149
rect 89140 164100 89150 164180
rect 89290 164100 89300 164180
rect 100640 164100 100650 164180
rect 100790 164100 100800 164180
rect 100940 164100 100950 164180
rect 101270 164149 101350 164159
rect 101590 164149 101670 164159
rect 102010 164149 102090 164159
rect 102330 164149 102410 164159
rect 114770 164149 114850 164159
rect 115090 164149 115170 164159
rect 115510 164149 115590 164159
rect 115830 164149 115910 164159
rect 101350 164069 101360 164149
rect 101670 164069 101680 164149
rect 102090 164069 102100 164149
rect 102410 164069 102420 164149
rect 114850 164069 114860 164149
rect 115170 164069 115180 164149
rect 115590 164069 115600 164149
rect 115910 164069 115920 164149
rect 116140 164100 116150 164180
rect 116290 164100 116300 164180
rect 127640 164100 127650 164180
rect 127790 164100 127800 164180
rect 127940 164100 127950 164180
rect 128270 164149 128350 164159
rect 128590 164149 128670 164159
rect 129010 164149 129090 164159
rect 129330 164149 129410 164159
rect 128350 164069 128360 164149
rect 128670 164069 128680 164149
rect 129090 164069 129100 164149
rect 129410 164069 129420 164149
rect 129640 164100 129650 164180
rect 129790 164100 129800 164180
rect 141140 164100 141150 164180
rect 141290 164100 141300 164180
rect 141440 164100 141450 164180
rect 141665 164150 141745 164160
rect 141985 164150 142065 164160
rect 145200 164150 145265 164160
rect 145505 164150 145585 164160
rect 145825 164150 145905 164160
rect 141745 164070 141755 164150
rect 142065 164070 142075 164150
rect 145265 164070 145275 164150
rect 145585 164070 145595 164150
rect 145905 164070 145915 164150
rect 146620 164140 146630 164220
rect 146940 164140 146950 164220
rect 146700 164060 146780 164070
rect 49155 164040 49235 164050
rect 49315 164040 49395 164050
rect 62655 164040 62735 164050
rect 76155 164040 76235 164050
rect 89655 164040 89735 164050
rect 116655 164040 116735 164050
rect 130155 164040 130235 164050
rect 48500 164000 48640 164010
rect 48710 164000 48790 164010
rect 44065 163990 44145 164000
rect 44385 163990 44465 164000
rect 44705 163990 44785 164000
rect 45025 163990 45105 164000
rect 45345 163990 45425 164000
rect 45665 163990 45745 164000
rect 45985 163990 46065 164000
rect 46305 163990 46385 164000
rect 46625 163990 46705 164000
rect 46945 163990 47025 164000
rect 47265 163990 47345 164000
rect 47585 163990 47665 164000
rect 47905 163990 47985 164000
rect 48225 163990 48305 164000
rect 44145 163910 44155 163990
rect 44465 163910 44475 163990
rect 44785 163910 44795 163990
rect 45105 163910 45115 163990
rect 45425 163910 45435 163990
rect 45745 163910 45755 163990
rect 46065 163910 46075 163990
rect 46385 163910 46395 163990
rect 46705 163910 46715 163990
rect 47025 163910 47035 163990
rect 47345 163910 47355 163990
rect 47665 163910 47675 163990
rect 47985 163910 47995 163990
rect 48305 163910 48315 163990
rect 43060 163900 43140 163910
rect 43380 163900 43460 163910
rect 43140 163820 43150 163900
rect 43460 163820 43470 163900
rect 43905 163830 43985 163840
rect 44225 163830 44305 163840
rect 44545 163830 44625 163840
rect 44865 163830 44945 163840
rect 45185 163830 45265 163840
rect 45505 163830 45585 163840
rect 45825 163830 45905 163840
rect 46145 163830 46225 163840
rect 46465 163830 46545 163840
rect 46785 163830 46865 163840
rect 47105 163830 47185 163840
rect 47425 163830 47505 163840
rect 47745 163830 47825 163840
rect 48065 163830 48145 163840
rect 48500 163830 48605 164000
rect 48640 163920 48650 164000
rect 48790 163920 48800 164000
rect 49235 163960 49245 164040
rect 49315 163960 49325 164040
rect 49395 163960 49405 164040
rect 60060 164000 60140 164010
rect 60210 164000 60290 164010
rect 60360 164000 60440 164010
rect 62060 164000 62140 164010
rect 62210 164000 62290 164010
rect 60140 163920 60150 164000
rect 60290 163920 60300 164000
rect 60440 163920 60450 164000
rect 60610 163989 60690 163999
rect 60930 163989 61010 163999
rect 61350 163989 61430 163999
rect 61670 163989 61750 163999
rect 60690 163909 60700 163989
rect 61010 163909 61020 163989
rect 61430 163909 61440 163989
rect 61750 163909 61760 163989
rect 62140 163920 62150 164000
rect 62290 163920 62300 164000
rect 62735 163960 62745 164040
rect 73560 164000 73640 164010
rect 73710 164000 73790 164010
rect 73860 164000 73940 164010
rect 75560 164000 75640 164010
rect 75710 164000 75790 164010
rect 73640 163920 73650 164000
rect 73790 163920 73800 164000
rect 73940 163920 73950 164000
rect 74110 163989 74190 163999
rect 74430 163989 74510 163999
rect 74850 163989 74930 163999
rect 75170 163989 75250 163999
rect 74190 163909 74200 163989
rect 74510 163909 74520 163989
rect 74930 163909 74940 163989
rect 75250 163909 75260 163989
rect 75640 163920 75650 164000
rect 75790 163920 75800 164000
rect 76235 163960 76245 164040
rect 87060 164000 87140 164010
rect 87210 164000 87290 164010
rect 87360 164000 87440 164010
rect 89060 164000 89140 164010
rect 89210 164000 89290 164010
rect 87140 163920 87150 164000
rect 87290 163920 87300 164000
rect 87440 163920 87450 164000
rect 87610 163989 87690 163999
rect 87930 163989 88010 163999
rect 88350 163989 88430 163999
rect 88670 163989 88750 163999
rect 87690 163909 87700 163989
rect 88010 163909 88020 163989
rect 88430 163909 88440 163989
rect 88750 163909 88760 163989
rect 89140 163920 89150 164000
rect 89290 163920 89300 164000
rect 89735 163960 89745 164040
rect 100560 164000 100640 164010
rect 100710 164000 100790 164010
rect 100860 164000 100940 164010
rect 116060 164000 116140 164010
rect 116210 164000 116290 164010
rect 100640 163920 100650 164000
rect 100790 163920 100800 164000
rect 100940 163920 100950 164000
rect 101110 163989 101190 163999
rect 101430 163989 101510 163999
rect 101850 163989 101930 163999
rect 102170 163989 102250 163999
rect 114610 163989 114690 163999
rect 114930 163989 115010 163999
rect 115350 163989 115430 163999
rect 115670 163989 115750 163999
rect 101190 163909 101200 163989
rect 101510 163909 101520 163989
rect 101930 163909 101940 163989
rect 102250 163909 102260 163989
rect 114690 163909 114700 163989
rect 115010 163909 115020 163989
rect 115430 163909 115440 163989
rect 115750 163909 115760 163989
rect 116140 163920 116150 164000
rect 116290 163920 116300 164000
rect 116735 163960 116745 164040
rect 127560 164000 127640 164010
rect 127710 164000 127790 164010
rect 127860 164000 127940 164010
rect 129560 164000 129640 164010
rect 129710 164000 129790 164010
rect 127640 163920 127650 164000
rect 127790 163920 127800 164000
rect 127940 163920 127950 164000
rect 128110 163989 128190 163999
rect 128430 163989 128510 163999
rect 128850 163989 128930 163999
rect 129170 163989 129250 163999
rect 128190 163909 128200 163989
rect 128510 163909 128520 163989
rect 128930 163909 128940 163989
rect 129250 163909 129260 163989
rect 129640 163920 129650 164000
rect 129790 163920 129800 164000
rect 130235 163960 130245 164040
rect 141060 164000 141140 164010
rect 141210 164000 141290 164010
rect 141360 164000 141440 164010
rect 141140 163920 141150 164000
rect 141290 163920 141300 164000
rect 141440 163920 141450 164000
rect 141825 163990 141905 164000
rect 142145 163990 142200 164000
rect 145345 163990 145425 164000
rect 145665 163990 145745 164000
rect 145985 163990 146065 164000
rect 141905 163910 141915 163990
rect 145425 163910 145435 163990
rect 145745 163910 145755 163990
rect 146065 163910 146075 163990
rect 146780 163980 146790 164060
rect 146540 163900 146620 163910
rect 146860 163900 146940 163910
rect 43985 163750 43995 163830
rect 44305 163750 44315 163830
rect 44625 163750 44635 163830
rect 44945 163750 44955 163830
rect 45265 163750 45275 163830
rect 45585 163750 45595 163830
rect 45905 163750 45915 163830
rect 46225 163750 46235 163830
rect 46545 163750 46555 163830
rect 46865 163750 46875 163830
rect 47185 163750 47195 163830
rect 47505 163750 47515 163830
rect 47825 163750 47835 163830
rect 48145 163750 48155 163830
rect 48500 163820 48640 163830
rect 48710 163820 48790 163830
rect 60060 163820 60140 163830
rect 60210 163820 60290 163830
rect 60360 163820 60440 163830
rect 60770 163829 60850 163839
rect 61090 163829 61170 163839
rect 61510 163829 61590 163839
rect 61830 163829 61910 163839
rect 42950 163740 42980 163750
rect 43220 163740 43300 163750
rect 42980 163660 42990 163740
rect 43300 163660 43310 163740
rect 44065 163670 44145 163680
rect 44385 163670 44465 163680
rect 44705 163670 44785 163680
rect 45025 163670 45105 163680
rect 45345 163670 45425 163680
rect 45665 163670 45745 163680
rect 45985 163670 46065 163680
rect 46305 163670 46385 163680
rect 46625 163670 46705 163680
rect 46945 163670 47025 163680
rect 47265 163670 47345 163680
rect 47585 163670 47665 163680
rect 47905 163670 47985 163680
rect 48225 163670 48305 163680
rect 44145 163590 44155 163670
rect 44465 163590 44475 163670
rect 44785 163590 44795 163670
rect 45105 163590 45115 163670
rect 45425 163590 45435 163670
rect 45745 163590 45755 163670
rect 46065 163590 46075 163670
rect 46385 163590 46395 163670
rect 46705 163590 46715 163670
rect 47025 163590 47035 163670
rect 47345 163590 47355 163670
rect 47665 163590 47675 163670
rect 47985 163590 47995 163670
rect 48305 163590 48315 163670
rect 48500 163650 48605 163820
rect 48640 163740 48650 163820
rect 48790 163740 48800 163820
rect 60140 163740 60150 163820
rect 60290 163740 60300 163820
rect 60440 163740 60450 163820
rect 60850 163749 60860 163829
rect 61170 163749 61180 163829
rect 61590 163749 61600 163829
rect 61910 163749 61920 163829
rect 62060 163820 62140 163830
rect 62210 163820 62290 163830
rect 73560 163820 73640 163830
rect 73710 163820 73790 163830
rect 73860 163820 73940 163830
rect 74270 163829 74350 163839
rect 74590 163829 74670 163839
rect 75010 163829 75090 163839
rect 75330 163829 75410 163839
rect 62140 163740 62150 163820
rect 62290 163740 62300 163820
rect 73640 163740 73650 163820
rect 73790 163740 73800 163820
rect 73940 163740 73950 163820
rect 74350 163749 74360 163829
rect 74670 163749 74680 163829
rect 75090 163749 75100 163829
rect 75410 163749 75420 163829
rect 75560 163820 75640 163830
rect 75710 163820 75790 163830
rect 87060 163820 87140 163830
rect 87210 163820 87290 163830
rect 87360 163820 87440 163830
rect 87770 163829 87850 163839
rect 88090 163829 88170 163839
rect 88510 163829 88590 163839
rect 88830 163829 88910 163839
rect 75640 163740 75650 163820
rect 75790 163740 75800 163820
rect 87140 163740 87150 163820
rect 87290 163740 87300 163820
rect 87440 163740 87450 163820
rect 87850 163749 87860 163829
rect 88170 163749 88180 163829
rect 88590 163749 88600 163829
rect 88910 163749 88920 163829
rect 89060 163820 89140 163830
rect 89210 163820 89290 163830
rect 100560 163820 100640 163830
rect 100710 163820 100790 163830
rect 100860 163820 100940 163830
rect 101270 163829 101350 163839
rect 101590 163829 101670 163839
rect 102010 163829 102090 163839
rect 102330 163829 102410 163839
rect 114770 163829 114850 163839
rect 115090 163829 115170 163839
rect 115510 163829 115590 163839
rect 115830 163829 115910 163839
rect 89140 163740 89150 163820
rect 89290 163740 89300 163820
rect 100640 163740 100650 163820
rect 100790 163740 100800 163820
rect 100940 163740 100950 163820
rect 101350 163749 101360 163829
rect 101670 163749 101680 163829
rect 102090 163749 102100 163829
rect 102410 163749 102420 163829
rect 114850 163749 114860 163829
rect 115170 163749 115180 163829
rect 115590 163749 115600 163829
rect 115910 163749 115920 163829
rect 116060 163820 116140 163830
rect 116210 163820 116290 163830
rect 127560 163820 127640 163830
rect 127710 163820 127790 163830
rect 127860 163820 127940 163830
rect 128270 163829 128350 163839
rect 128590 163829 128670 163839
rect 129010 163829 129090 163839
rect 129330 163829 129410 163839
rect 141665 163830 141745 163840
rect 141985 163830 142065 163840
rect 145200 163830 145265 163840
rect 145505 163830 145585 163840
rect 145825 163830 145905 163840
rect 116140 163740 116150 163820
rect 116290 163740 116300 163820
rect 127640 163740 127650 163820
rect 127790 163740 127800 163820
rect 127940 163740 127950 163820
rect 128350 163749 128360 163829
rect 128670 163749 128680 163829
rect 129090 163749 129100 163829
rect 129410 163749 129420 163829
rect 129560 163820 129640 163830
rect 129710 163820 129790 163830
rect 141060 163820 141140 163830
rect 141210 163820 141290 163830
rect 141360 163820 141440 163830
rect 129640 163740 129650 163820
rect 129790 163740 129800 163820
rect 141140 163740 141150 163820
rect 141290 163740 141300 163820
rect 141440 163740 141450 163820
rect 141745 163750 141755 163830
rect 142065 163750 142075 163830
rect 145265 163750 145275 163830
rect 145585 163750 145595 163830
rect 145905 163750 145915 163830
rect 146620 163820 146630 163900
rect 146940 163820 146950 163900
rect 146700 163740 146780 163750
rect 49180 163670 49210 163700
rect 49300 163670 49330 163700
rect 49420 163670 49450 163700
rect 49540 163670 49570 163700
rect 49660 163670 49690 163700
rect 49780 163670 49810 163700
rect 49900 163670 49930 163700
rect 50020 163670 50050 163700
rect 50140 163670 50170 163700
rect 50260 163670 50290 163700
rect 50380 163670 50410 163700
rect 50500 163670 50530 163700
rect 50620 163670 50650 163700
rect 50740 163670 50770 163700
rect 50860 163670 50890 163700
rect 50980 163670 51010 163700
rect 51100 163670 51130 163700
rect 51220 163670 51250 163700
rect 51340 163670 51370 163700
rect 51460 163670 51490 163700
rect 51580 163670 51610 163700
rect 51700 163670 51730 163700
rect 51820 163670 51850 163700
rect 51940 163670 51970 163700
rect 52060 163670 52090 163700
rect 52180 163670 52210 163700
rect 52300 163670 52330 163700
rect 52420 163670 52450 163700
rect 52540 163670 52570 163700
rect 52660 163670 52690 163700
rect 52780 163670 52810 163700
rect 52900 163670 52930 163700
rect 53020 163670 53050 163700
rect 53140 163670 53170 163700
rect 53260 163670 53290 163700
rect 53380 163670 53410 163700
rect 53500 163670 53530 163700
rect 53620 163670 53650 163700
rect 53740 163670 53770 163700
rect 53860 163670 53890 163700
rect 53980 163670 54010 163700
rect 54100 163670 54130 163700
rect 54220 163670 54250 163700
rect 54340 163670 54370 163700
rect 54460 163670 54490 163700
rect 54580 163670 54610 163700
rect 54700 163670 54730 163700
rect 54820 163670 54850 163700
rect 54940 163670 54970 163700
rect 55060 163670 55090 163700
rect 55180 163670 55210 163700
rect 55300 163670 55330 163700
rect 55420 163670 55450 163700
rect 55540 163670 55570 163700
rect 55660 163670 55690 163700
rect 55780 163670 55810 163700
rect 55900 163670 55930 163700
rect 56020 163670 56050 163700
rect 56140 163670 56170 163700
rect 56260 163670 56290 163700
rect 56380 163670 56410 163700
rect 56500 163670 56530 163700
rect 56620 163670 56650 163700
rect 56740 163670 56770 163700
rect 56860 163670 56890 163700
rect 56980 163670 57010 163700
rect 57100 163670 57130 163700
rect 57220 163670 57250 163700
rect 57340 163670 57370 163700
rect 57460 163670 57490 163700
rect 57580 163670 57610 163700
rect 57700 163670 57730 163700
rect 57820 163670 57850 163700
rect 57940 163670 57970 163700
rect 58060 163670 58090 163700
rect 58180 163670 58210 163700
rect 58300 163670 58330 163700
rect 58420 163670 58450 163700
rect 58540 163670 58570 163700
rect 58660 163670 58690 163700
rect 58780 163670 58810 163700
rect 58900 163670 58930 163700
rect 59020 163670 59050 163700
rect 59140 163670 59170 163700
rect 59260 163670 59290 163700
rect 59380 163670 59410 163700
rect 59500 163670 59530 163700
rect 59620 163670 59650 163700
rect 59740 163670 59770 163700
rect 48500 163640 48640 163650
rect 48710 163640 48790 163650
rect 49060 163640 49120 163670
rect 49180 163640 49240 163670
rect 49300 163640 49360 163670
rect 49420 163640 49480 163670
rect 49540 163640 49600 163670
rect 49660 163640 49720 163670
rect 49780 163640 49840 163670
rect 49900 163640 49960 163670
rect 50020 163640 50080 163670
rect 50140 163640 50200 163670
rect 50260 163640 50320 163670
rect 50380 163640 50440 163670
rect 50500 163640 50560 163670
rect 50620 163640 50680 163670
rect 50740 163640 50800 163670
rect 50860 163640 50920 163670
rect 50980 163640 51040 163670
rect 51100 163640 51160 163670
rect 51220 163640 51280 163670
rect 51340 163640 51400 163670
rect 51460 163640 51520 163670
rect 51580 163640 51640 163670
rect 51700 163640 51760 163670
rect 51820 163640 51880 163670
rect 51940 163640 52000 163670
rect 52060 163640 52120 163670
rect 52180 163640 52240 163670
rect 52300 163640 52360 163670
rect 52420 163640 52480 163670
rect 52540 163640 52600 163670
rect 52660 163640 52720 163670
rect 52780 163640 52840 163670
rect 52900 163640 52960 163670
rect 53020 163640 53080 163670
rect 53140 163640 53200 163670
rect 53260 163640 53320 163670
rect 53380 163640 53440 163670
rect 53500 163640 53560 163670
rect 53620 163640 53680 163670
rect 53740 163640 53800 163670
rect 53860 163640 53920 163670
rect 53980 163640 54040 163670
rect 54100 163640 54160 163670
rect 54220 163640 54280 163670
rect 54340 163640 54400 163670
rect 54460 163640 54520 163670
rect 54580 163640 54640 163670
rect 54700 163640 54760 163670
rect 54820 163640 54880 163670
rect 54940 163640 55000 163670
rect 55060 163640 55120 163670
rect 55180 163640 55240 163670
rect 55300 163640 55360 163670
rect 55420 163640 55480 163670
rect 55540 163640 55600 163670
rect 55660 163640 55720 163670
rect 55780 163640 55840 163670
rect 55900 163640 55960 163670
rect 56020 163640 56080 163670
rect 56140 163640 56200 163670
rect 56260 163640 56320 163670
rect 56380 163640 56440 163670
rect 56500 163640 56560 163670
rect 56620 163640 56680 163670
rect 56740 163640 56800 163670
rect 56860 163640 56920 163670
rect 56980 163640 57040 163670
rect 57100 163640 57160 163670
rect 57220 163640 57280 163670
rect 57340 163640 57400 163670
rect 57460 163640 57520 163670
rect 57580 163640 57640 163670
rect 57700 163640 57760 163670
rect 57820 163640 57880 163670
rect 57940 163640 58000 163670
rect 58060 163640 58120 163670
rect 58180 163640 58240 163670
rect 58300 163640 58360 163670
rect 58420 163640 58480 163670
rect 58540 163640 58600 163670
rect 58660 163640 58720 163670
rect 58780 163640 58840 163670
rect 58900 163640 58960 163670
rect 59020 163640 59080 163670
rect 59140 163640 59200 163670
rect 59260 163640 59320 163670
rect 59380 163640 59440 163670
rect 59500 163640 59560 163670
rect 59620 163640 59680 163670
rect 59740 163640 59800 163670
rect 60610 163669 60690 163679
rect 60930 163669 61010 163679
rect 61350 163669 61430 163679
rect 61670 163669 61750 163679
rect 62680 163670 62710 163700
rect 73245 163670 73270 163700
rect 60060 163640 60140 163650
rect 60210 163640 60290 163650
rect 60360 163640 60440 163650
rect 43060 163580 43140 163590
rect 43380 163580 43460 163590
rect 43140 163500 43150 163580
rect 43460 163500 43470 163580
rect 48500 163470 48605 163640
rect 48640 163560 48650 163640
rect 48790 163560 48800 163640
rect 49180 163550 49210 163580
rect 49300 163550 49330 163580
rect 49420 163550 49450 163580
rect 49540 163550 49570 163580
rect 49660 163550 49690 163580
rect 49780 163550 49810 163580
rect 49900 163550 49930 163580
rect 50020 163550 50050 163580
rect 50140 163550 50170 163580
rect 50260 163550 50290 163580
rect 50380 163550 50410 163580
rect 50500 163550 50530 163580
rect 50620 163550 50650 163580
rect 50740 163550 50770 163580
rect 50860 163550 50890 163580
rect 50980 163550 51010 163580
rect 51100 163550 51130 163580
rect 51220 163550 51250 163580
rect 51340 163550 51370 163580
rect 51460 163550 51490 163580
rect 51580 163550 51610 163580
rect 51700 163550 51730 163580
rect 51820 163550 51850 163580
rect 51940 163550 51970 163580
rect 52060 163550 52090 163580
rect 52180 163550 52210 163580
rect 52300 163550 52330 163580
rect 52420 163550 52450 163580
rect 52540 163550 52570 163580
rect 52660 163550 52690 163580
rect 52780 163550 52810 163580
rect 52900 163550 52930 163580
rect 53020 163550 53050 163580
rect 53140 163550 53170 163580
rect 53260 163550 53290 163580
rect 53380 163550 53410 163580
rect 53500 163550 53530 163580
rect 53620 163550 53650 163580
rect 53740 163550 53770 163580
rect 53860 163550 53890 163580
rect 53980 163550 54010 163580
rect 54100 163550 54130 163580
rect 54220 163550 54250 163580
rect 54340 163550 54370 163580
rect 54460 163550 54490 163580
rect 54580 163550 54610 163580
rect 54700 163550 54730 163580
rect 54820 163550 54850 163580
rect 54940 163550 54970 163580
rect 55060 163550 55090 163580
rect 55180 163550 55210 163580
rect 55300 163550 55330 163580
rect 55420 163550 55450 163580
rect 55540 163550 55570 163580
rect 55660 163550 55690 163580
rect 55780 163550 55810 163580
rect 55900 163550 55930 163580
rect 56020 163550 56050 163580
rect 56140 163550 56170 163580
rect 56260 163550 56290 163580
rect 56380 163550 56410 163580
rect 56500 163550 56530 163580
rect 56620 163550 56650 163580
rect 56740 163550 56770 163580
rect 56860 163550 56890 163580
rect 56980 163550 57010 163580
rect 57100 163550 57130 163580
rect 57220 163550 57250 163580
rect 57340 163550 57370 163580
rect 57460 163550 57490 163580
rect 57580 163550 57610 163580
rect 57700 163550 57730 163580
rect 57820 163550 57850 163580
rect 57940 163550 57970 163580
rect 58060 163550 58090 163580
rect 58180 163550 58210 163580
rect 58300 163550 58330 163580
rect 58420 163550 58450 163580
rect 58540 163550 58570 163580
rect 58660 163550 58690 163580
rect 58780 163550 58810 163580
rect 58900 163550 58930 163580
rect 59020 163550 59050 163580
rect 59140 163550 59170 163580
rect 59260 163550 59290 163580
rect 59380 163550 59410 163580
rect 59500 163550 59530 163580
rect 59620 163550 59650 163580
rect 59740 163550 59770 163580
rect 60140 163560 60150 163640
rect 60290 163560 60300 163640
rect 60440 163560 60450 163640
rect 60690 163589 60700 163669
rect 61010 163589 61020 163669
rect 61430 163589 61440 163669
rect 61750 163589 61760 163669
rect 62060 163640 62140 163650
rect 62210 163640 62290 163650
rect 62560 163640 62620 163670
rect 62680 163640 62740 163670
rect 73245 163640 73300 163670
rect 74110 163669 74190 163679
rect 74430 163669 74510 163679
rect 74850 163669 74930 163679
rect 75170 163669 75250 163679
rect 76180 163670 76210 163700
rect 86745 163670 86770 163700
rect 73560 163640 73640 163650
rect 73710 163640 73790 163650
rect 73860 163640 73940 163650
rect 62140 163560 62150 163640
rect 62290 163560 62300 163640
rect 62680 163550 62710 163580
rect 73245 163550 73270 163580
rect 73640 163560 73650 163640
rect 73790 163560 73800 163640
rect 73940 163560 73950 163640
rect 74190 163589 74200 163669
rect 74510 163589 74520 163669
rect 74930 163589 74940 163669
rect 75250 163589 75260 163669
rect 75560 163640 75640 163650
rect 75710 163640 75790 163650
rect 76060 163640 76120 163670
rect 76180 163640 76240 163670
rect 86745 163640 86800 163670
rect 87610 163669 87690 163679
rect 87930 163669 88010 163679
rect 88350 163669 88430 163679
rect 88670 163669 88750 163679
rect 89680 163670 89710 163700
rect 100245 163670 100270 163700
rect 87060 163640 87140 163650
rect 87210 163640 87290 163650
rect 87360 163640 87440 163650
rect 75640 163560 75650 163640
rect 75790 163560 75800 163640
rect 76180 163550 76210 163580
rect 86745 163550 86770 163580
rect 87140 163560 87150 163640
rect 87290 163560 87300 163640
rect 87440 163560 87450 163640
rect 87690 163589 87700 163669
rect 88010 163589 88020 163669
rect 88430 163589 88440 163669
rect 88750 163589 88760 163669
rect 89060 163640 89140 163650
rect 89210 163640 89290 163650
rect 89560 163640 89620 163670
rect 89680 163640 89740 163670
rect 100245 163640 100300 163670
rect 101110 163669 101190 163679
rect 101430 163669 101510 163679
rect 101850 163669 101930 163679
rect 102170 163669 102250 163679
rect 114610 163669 114690 163679
rect 114930 163669 115010 163679
rect 115350 163669 115430 163679
rect 115670 163669 115750 163679
rect 116680 163670 116710 163700
rect 127245 163670 127270 163700
rect 100560 163640 100640 163650
rect 100710 163640 100790 163650
rect 100860 163640 100940 163650
rect 89140 163560 89150 163640
rect 89290 163560 89300 163640
rect 89680 163550 89710 163580
rect 100245 163550 100270 163580
rect 100640 163560 100650 163640
rect 100790 163560 100800 163640
rect 100940 163560 100950 163640
rect 101190 163589 101200 163669
rect 101510 163589 101520 163669
rect 101930 163589 101940 163669
rect 102250 163589 102260 163669
rect 114690 163589 114700 163669
rect 115010 163589 115020 163669
rect 115430 163589 115440 163669
rect 115750 163589 115760 163669
rect 116060 163640 116140 163650
rect 116210 163640 116290 163650
rect 116560 163640 116620 163670
rect 116680 163640 116740 163670
rect 127245 163640 127300 163670
rect 128110 163669 128190 163679
rect 128430 163669 128510 163679
rect 128850 163669 128930 163679
rect 129170 163669 129250 163679
rect 130180 163670 130210 163700
rect 140740 163670 140770 163700
rect 141825 163670 141905 163680
rect 142145 163670 142200 163680
rect 145345 163670 145425 163680
rect 145665 163670 145745 163680
rect 145985 163670 146065 163680
rect 127560 163640 127640 163650
rect 127710 163640 127790 163650
rect 127860 163640 127940 163650
rect 116140 163560 116150 163640
rect 116290 163560 116300 163640
rect 116680 163550 116710 163580
rect 127245 163550 127270 163580
rect 127640 163560 127650 163640
rect 127790 163560 127800 163640
rect 127940 163560 127950 163640
rect 128190 163589 128200 163669
rect 128510 163589 128520 163669
rect 128930 163589 128940 163669
rect 129250 163589 129260 163669
rect 129560 163640 129640 163650
rect 129710 163640 129790 163650
rect 130060 163640 130120 163670
rect 130180 163640 130240 163670
rect 140740 163640 140800 163670
rect 141060 163640 141140 163650
rect 141210 163640 141290 163650
rect 141360 163640 141440 163650
rect 129640 163560 129650 163640
rect 129790 163560 129800 163640
rect 130180 163550 130210 163580
rect 140740 163550 140770 163580
rect 141140 163560 141150 163640
rect 141290 163560 141300 163640
rect 141440 163560 141450 163640
rect 141905 163590 141915 163670
rect 145425 163590 145435 163670
rect 145745 163590 145755 163670
rect 146065 163590 146075 163670
rect 146780 163660 146790 163740
rect 146540 163580 146620 163590
rect 146860 163580 146940 163590
rect 49060 163520 49120 163550
rect 49180 163520 49240 163550
rect 49300 163520 49360 163550
rect 49420 163520 49480 163550
rect 49540 163520 49600 163550
rect 49660 163520 49720 163550
rect 49780 163520 49840 163550
rect 49900 163520 49960 163550
rect 50020 163520 50080 163550
rect 50140 163520 50200 163550
rect 50260 163520 50320 163550
rect 50380 163520 50440 163550
rect 50500 163520 50560 163550
rect 50620 163520 50680 163550
rect 50740 163520 50800 163550
rect 50860 163520 50920 163550
rect 50980 163520 51040 163550
rect 51100 163520 51160 163550
rect 51220 163520 51280 163550
rect 51340 163520 51400 163550
rect 51460 163520 51520 163550
rect 51580 163520 51640 163550
rect 51700 163520 51760 163550
rect 51820 163520 51880 163550
rect 51940 163520 52000 163550
rect 52060 163520 52120 163550
rect 52180 163520 52240 163550
rect 52300 163520 52360 163550
rect 52420 163520 52480 163550
rect 52540 163520 52600 163550
rect 52660 163520 52720 163550
rect 52780 163520 52840 163550
rect 52900 163520 52960 163550
rect 53020 163520 53080 163550
rect 53140 163520 53200 163550
rect 53260 163520 53320 163550
rect 53380 163520 53440 163550
rect 53500 163520 53560 163550
rect 53620 163520 53680 163550
rect 53740 163520 53800 163550
rect 53860 163520 53920 163550
rect 53980 163520 54040 163550
rect 54100 163520 54160 163550
rect 54220 163520 54280 163550
rect 54340 163520 54400 163550
rect 54460 163520 54520 163550
rect 54580 163520 54640 163550
rect 54700 163520 54760 163550
rect 54820 163520 54880 163550
rect 54940 163520 55000 163550
rect 55060 163520 55120 163550
rect 55180 163520 55240 163550
rect 55300 163520 55360 163550
rect 55420 163520 55480 163550
rect 55540 163520 55600 163550
rect 55660 163520 55720 163550
rect 55780 163520 55840 163550
rect 55900 163520 55960 163550
rect 56020 163520 56080 163550
rect 56140 163520 56200 163550
rect 56260 163520 56320 163550
rect 56380 163520 56440 163550
rect 56500 163520 56560 163550
rect 56620 163520 56680 163550
rect 56740 163520 56800 163550
rect 56860 163520 56920 163550
rect 56980 163520 57040 163550
rect 57100 163520 57160 163550
rect 57220 163520 57280 163550
rect 57340 163520 57400 163550
rect 57460 163520 57520 163550
rect 57580 163520 57640 163550
rect 57700 163520 57760 163550
rect 57820 163520 57880 163550
rect 57940 163520 58000 163550
rect 58060 163520 58120 163550
rect 58180 163520 58240 163550
rect 58300 163520 58360 163550
rect 58420 163520 58480 163550
rect 58540 163520 58600 163550
rect 58660 163520 58720 163550
rect 58780 163520 58840 163550
rect 58900 163520 58960 163550
rect 59020 163520 59080 163550
rect 59140 163520 59200 163550
rect 59260 163520 59320 163550
rect 59380 163520 59440 163550
rect 59500 163520 59560 163550
rect 59620 163520 59680 163550
rect 59740 163520 59800 163550
rect 62560 163520 62620 163550
rect 62680 163520 62740 163550
rect 73245 163520 73300 163550
rect 76060 163520 76120 163550
rect 76180 163520 76240 163550
rect 86745 163520 86800 163550
rect 89560 163520 89620 163550
rect 89680 163520 89740 163550
rect 100245 163520 100300 163550
rect 116560 163520 116620 163550
rect 116680 163520 116740 163550
rect 127245 163520 127300 163550
rect 130060 163520 130120 163550
rect 130180 163520 130240 163550
rect 140740 163520 140800 163550
rect 146620 163500 146630 163580
rect 146940 163500 146950 163580
rect 48500 163460 48640 163470
rect 48710 163460 48790 163470
rect 60060 163460 60140 163470
rect 60210 163460 60290 163470
rect 60360 163460 60440 163470
rect 62060 163460 62140 163470
rect 62210 163460 62290 163470
rect 73560 163460 73640 163470
rect 73710 163460 73790 163470
rect 73860 163460 73940 163470
rect 75560 163460 75640 163470
rect 75710 163460 75790 163470
rect 87060 163460 87140 163470
rect 87210 163460 87290 163470
rect 87360 163460 87440 163470
rect 89060 163460 89140 163470
rect 89210 163460 89290 163470
rect 100560 163460 100640 163470
rect 100710 163460 100790 163470
rect 100860 163460 100940 163470
rect 116060 163460 116140 163470
rect 116210 163460 116290 163470
rect 127560 163460 127640 163470
rect 127710 163460 127790 163470
rect 127860 163460 127940 163470
rect 129560 163460 129640 163470
rect 129710 163460 129790 163470
rect 141060 163460 141140 163470
rect 141210 163460 141290 163470
rect 141360 163460 141440 163470
rect 48500 163300 48605 163460
rect 48640 163380 48650 163460
rect 48790 163380 48800 163460
rect 49180 163400 49210 163460
rect 49300 163400 49330 163460
rect 49420 163400 49450 163460
rect 49540 163400 49570 163460
rect 49660 163400 49690 163460
rect 49780 163400 49810 163460
rect 49900 163400 49930 163460
rect 50020 163400 50050 163460
rect 50140 163400 50170 163460
rect 50260 163400 50290 163460
rect 50380 163400 50410 163460
rect 50500 163400 50530 163460
rect 50620 163400 50650 163460
rect 50740 163400 50770 163460
rect 50860 163400 50890 163460
rect 50980 163400 51010 163460
rect 51100 163400 51130 163460
rect 51220 163400 51250 163460
rect 51340 163400 51370 163460
rect 51460 163400 51490 163460
rect 51580 163400 51610 163460
rect 51700 163400 51730 163460
rect 51820 163400 51850 163460
rect 51940 163400 51970 163460
rect 52060 163400 52090 163460
rect 52180 163400 52210 163460
rect 52300 163400 52330 163460
rect 52420 163400 52450 163460
rect 52540 163400 52570 163460
rect 52660 163400 52690 163460
rect 52780 163400 52810 163460
rect 52900 163400 52930 163460
rect 53020 163400 53050 163460
rect 53140 163400 53170 163460
rect 53260 163400 53290 163460
rect 53380 163400 53410 163460
rect 53500 163400 53530 163460
rect 53620 163400 53650 163460
rect 53740 163400 53770 163460
rect 53860 163400 53890 163460
rect 53980 163400 54010 163460
rect 54100 163400 54130 163460
rect 54220 163400 54250 163460
rect 54340 163400 54370 163460
rect 54460 163400 54490 163460
rect 54580 163400 54610 163460
rect 54700 163400 54730 163460
rect 54820 163400 54850 163460
rect 54940 163400 54970 163460
rect 55060 163400 55090 163460
rect 55180 163400 55210 163460
rect 55300 163400 55330 163460
rect 55420 163400 55450 163460
rect 55540 163400 55570 163460
rect 55660 163400 55690 163460
rect 55780 163400 55810 163460
rect 55900 163400 55930 163460
rect 56020 163400 56050 163460
rect 56140 163400 56170 163460
rect 56260 163400 56290 163460
rect 56380 163400 56410 163460
rect 56500 163400 56530 163460
rect 56620 163400 56650 163460
rect 56740 163400 56770 163460
rect 56860 163400 56890 163460
rect 56980 163400 57010 163460
rect 57100 163400 57130 163460
rect 57220 163400 57250 163460
rect 57340 163400 57370 163460
rect 57460 163400 57490 163460
rect 57580 163400 57610 163460
rect 57700 163400 57730 163460
rect 57820 163400 57850 163460
rect 57940 163400 57970 163460
rect 58060 163400 58090 163460
rect 58180 163400 58210 163460
rect 58300 163400 58330 163460
rect 58420 163400 58450 163460
rect 58540 163400 58570 163460
rect 58660 163400 58690 163460
rect 58780 163400 58810 163460
rect 58900 163400 58930 163460
rect 59020 163400 59050 163460
rect 59140 163400 59170 163460
rect 59260 163400 59290 163460
rect 59380 163400 59410 163460
rect 59500 163400 59530 163460
rect 59620 163400 59650 163460
rect 59740 163400 59770 163460
rect 60140 163380 60150 163460
rect 60290 163380 60300 163460
rect 60440 163380 60450 163460
rect 62140 163380 62150 163460
rect 62290 163380 62300 163460
rect 62680 163400 62710 163460
rect 73245 163400 73270 163460
rect 73640 163380 73650 163460
rect 73790 163380 73800 163460
rect 73940 163380 73950 163460
rect 75640 163380 75650 163460
rect 75790 163380 75800 163460
rect 76180 163400 76210 163460
rect 86745 163400 86770 163460
rect 87140 163380 87150 163460
rect 87290 163380 87300 163460
rect 87440 163380 87450 163460
rect 89140 163380 89150 163460
rect 89290 163380 89300 163460
rect 89680 163400 89710 163460
rect 100245 163400 100270 163460
rect 100640 163380 100650 163460
rect 100790 163380 100800 163460
rect 100940 163380 100950 163460
rect 116140 163380 116150 163460
rect 116290 163380 116300 163460
rect 116680 163400 116710 163460
rect 127245 163400 127270 163460
rect 127640 163380 127650 163460
rect 127790 163380 127800 163460
rect 127940 163380 127950 163460
rect 129640 163380 129650 163460
rect 129790 163380 129800 163460
rect 130180 163400 130210 163460
rect 140740 163400 140770 163460
rect 141140 163380 141150 163460
rect 141290 163380 141300 163460
rect 141440 163380 141450 163460
rect 62060 163299 62090 163300
rect 75560 163299 75590 163300
rect 89060 163299 89090 163300
rect 116060 163299 116090 163300
rect 129560 163299 129590 163300
rect 60085 162685 60165 162695
rect 60265 162685 60345 162695
rect 73585 162685 73665 162695
rect 73765 162685 73845 162695
rect 87085 162685 87165 162695
rect 87265 162685 87345 162695
rect 100585 162685 100665 162695
rect 100765 162685 100845 162695
rect 127585 162685 127665 162695
rect 127765 162685 127845 162695
rect 141085 162685 141165 162695
rect 141265 162685 141345 162695
rect 60165 162605 60175 162685
rect 60345 162605 60355 162685
rect 73665 162605 73675 162685
rect 73845 162605 73855 162685
rect 87165 162605 87175 162685
rect 87345 162605 87355 162685
rect 100665 162605 100675 162685
rect 100845 162605 100855 162685
rect 127665 162605 127675 162685
rect 127845 162605 127855 162685
rect 141165 162605 141175 162685
rect 141345 162605 141355 162685
rect 60085 162505 60165 162515
rect 60265 162505 60345 162515
rect 73585 162505 73665 162515
rect 73765 162505 73845 162515
rect 87085 162505 87165 162515
rect 87265 162505 87345 162515
rect 100585 162505 100665 162515
rect 100765 162505 100845 162515
rect 127585 162505 127665 162515
rect 127765 162505 127845 162515
rect 141085 162505 141165 162515
rect 141265 162505 141345 162515
rect 60165 162425 60175 162505
rect 60345 162425 60355 162505
rect 73665 162425 73675 162505
rect 73845 162425 73855 162505
rect 87165 162425 87175 162505
rect 87345 162425 87355 162505
rect 100665 162425 100675 162505
rect 100845 162425 100855 162505
rect 127665 162425 127675 162505
rect 127845 162425 127855 162505
rect 141165 162425 141175 162505
rect 141345 162425 141355 162505
rect 60085 162325 60165 162335
rect 60265 162325 60345 162335
rect 73585 162325 73665 162335
rect 73765 162325 73845 162335
rect 87085 162325 87165 162335
rect 87265 162325 87345 162335
rect 100585 162325 100665 162335
rect 100765 162325 100845 162335
rect 127585 162325 127665 162335
rect 127765 162325 127845 162335
rect 141085 162325 141165 162335
rect 141265 162325 141345 162335
rect 60165 162245 60175 162325
rect 60345 162245 60355 162325
rect 73665 162245 73675 162325
rect 73845 162245 73855 162325
rect 87165 162245 87175 162325
rect 87345 162245 87355 162325
rect 100665 162245 100675 162325
rect 100845 162245 100855 162325
rect 127665 162245 127675 162325
rect 127845 162245 127855 162325
rect 141165 162245 141175 162325
rect 141345 162245 141355 162325
rect 60085 162145 60165 162155
rect 60265 162145 60345 162155
rect 73585 162145 73665 162155
rect 73765 162145 73845 162155
rect 87085 162145 87165 162155
rect 87265 162145 87345 162155
rect 100585 162145 100665 162155
rect 100765 162145 100845 162155
rect 127585 162145 127665 162155
rect 127765 162145 127845 162155
rect 141085 162145 141165 162155
rect 141265 162145 141345 162155
rect 60165 162065 60175 162145
rect 60345 162065 60355 162145
rect 73665 162065 73675 162145
rect 73845 162065 73855 162145
rect 87165 162065 87175 162145
rect 87345 162065 87355 162145
rect 100665 162065 100675 162145
rect 100845 162065 100855 162145
rect 127665 162065 127675 162145
rect 127845 162065 127855 162145
rect 141165 162065 141175 162145
rect 141345 162065 141355 162145
rect 60085 161965 60165 161975
rect 60265 161965 60345 161975
rect 73585 161965 73665 161975
rect 73765 161965 73845 161975
rect 87085 161965 87165 161975
rect 87265 161965 87345 161975
rect 100585 161965 100665 161975
rect 100765 161965 100845 161975
rect 127585 161965 127665 161975
rect 127765 161965 127845 161975
rect 141085 161965 141165 161975
rect 141265 161965 141345 161975
rect 60165 161885 60175 161965
rect 60345 161885 60355 161965
rect 73665 161885 73675 161965
rect 73845 161885 73855 161965
rect 87165 161885 87175 161965
rect 87345 161885 87355 161965
rect 100665 161885 100675 161965
rect 100845 161885 100855 161965
rect 127665 161885 127675 161965
rect 127845 161885 127855 161965
rect 141165 161885 141175 161965
rect 141345 161885 141355 161965
rect 48685 161150 48765 161160
rect 62185 161150 62265 161160
rect 75685 161150 75765 161160
rect 89185 161150 89265 161160
rect 116185 161150 116265 161160
rect 129685 161150 129765 161160
rect 48765 161080 48775 161150
rect 62265 161080 62275 161150
rect 75765 161080 75775 161150
rect 89265 161080 89275 161150
rect 116265 161080 116275 161150
rect 129765 161080 129775 161150
rect 48685 161070 48775 161080
rect 62185 161070 62275 161080
rect 75685 161070 75775 161080
rect 89185 161070 89275 161080
rect 116185 161070 116275 161080
rect 129685 161070 129775 161080
rect 48685 160990 48765 161000
rect 62185 160990 62265 161000
rect 75685 160990 75765 161000
rect 89185 160990 89265 161000
rect 116185 160990 116265 161000
rect 129685 160990 129765 161000
rect 48765 160920 48775 160990
rect 62265 160920 62275 160990
rect 75765 160920 75775 160990
rect 89265 160920 89275 160990
rect 116265 160920 116275 160990
rect 129765 160920 129775 160990
rect 48685 160910 48775 160920
rect 62185 160910 62275 160920
rect 75685 160910 75775 160920
rect 89185 160910 89275 160920
rect 116185 160910 116275 160920
rect 129685 160910 129775 160920
rect 48685 160830 48765 160840
rect 62185 160830 62265 160840
rect 75685 160830 75765 160840
rect 89185 160830 89265 160840
rect 116185 160830 116265 160840
rect 129685 160830 129765 160840
rect 48765 160760 48775 160830
rect 62265 160760 62275 160830
rect 75765 160760 75775 160830
rect 89265 160760 89275 160830
rect 116265 160760 116275 160830
rect 129765 160760 129775 160830
rect 48685 160750 48775 160760
rect 62185 160750 62275 160760
rect 75685 160750 75775 160760
rect 89185 160750 89275 160760
rect 116185 160750 116275 160760
rect 129685 160750 129775 160760
rect 48685 160670 48765 160680
rect 62185 160670 62265 160680
rect 75685 160670 75765 160680
rect 89185 160670 89265 160680
rect 116185 160670 116265 160680
rect 129685 160670 129765 160680
rect 48765 160600 48775 160670
rect 62265 160600 62275 160670
rect 75765 160600 75775 160670
rect 89265 160600 89275 160670
rect 116265 160600 116275 160670
rect 129765 160600 129775 160670
rect 48685 160590 48775 160600
rect 62185 160590 62275 160600
rect 75685 160590 75775 160600
rect 89185 160590 89275 160600
rect 116185 160590 116275 160600
rect 129685 160590 129775 160600
rect 48685 160510 48765 160520
rect 62185 160510 62265 160520
rect 75685 160510 75765 160520
rect 89185 160510 89265 160520
rect 116185 160510 116265 160520
rect 129685 160510 129765 160520
rect 48765 160430 48775 160510
rect 62265 160430 62275 160510
rect 75765 160430 75775 160510
rect 89265 160430 89275 160510
rect 116265 160430 116275 160510
rect 129765 160430 129775 160510
rect 48500 159730 48605 159800
rect 48500 159720 48640 159730
rect 48710 159720 48790 159730
rect 60060 159720 60140 159730
rect 60210 159720 60290 159730
rect 60360 159720 60440 159730
rect 62060 159720 62140 159730
rect 62210 159720 62290 159730
rect 73560 159720 73640 159730
rect 73710 159720 73790 159730
rect 73860 159720 73940 159730
rect 75560 159720 75640 159730
rect 75710 159720 75790 159730
rect 87060 159720 87140 159730
rect 87210 159720 87290 159730
rect 87360 159720 87440 159730
rect 89060 159720 89140 159730
rect 89210 159720 89290 159730
rect 100560 159720 100640 159730
rect 100710 159720 100790 159730
rect 100860 159720 100940 159730
rect 116060 159720 116140 159730
rect 116210 159720 116290 159730
rect 127560 159720 127640 159730
rect 127710 159720 127790 159730
rect 127860 159720 127940 159730
rect 129560 159720 129640 159730
rect 129710 159720 129790 159730
rect 141060 159720 141140 159730
rect 141210 159720 141290 159730
rect 141360 159720 141440 159730
rect 43785 159640 43865 159650
rect 44105 159640 44185 159650
rect 44425 159640 44505 159650
rect 44745 159640 44825 159650
rect 45065 159640 45145 159650
rect 45385 159640 45465 159650
rect 45705 159640 45785 159650
rect 46025 159640 46105 159650
rect 46345 159640 46425 159650
rect 46665 159640 46745 159650
rect 46985 159640 47065 159650
rect 47305 159640 47385 159650
rect 47625 159640 47705 159650
rect 47945 159640 48025 159650
rect 48265 159640 48345 159650
rect 42950 159580 42980 159590
rect 43220 159580 43300 159590
rect 42980 159500 42990 159580
rect 43300 159500 43310 159580
rect 43865 159560 43875 159640
rect 44185 159560 44195 159640
rect 44505 159560 44515 159640
rect 44825 159560 44835 159640
rect 45145 159560 45155 159640
rect 45465 159560 45475 159640
rect 45785 159560 45795 159640
rect 46105 159560 46115 159640
rect 46425 159560 46435 159640
rect 46745 159560 46755 159640
rect 47065 159560 47075 159640
rect 47385 159560 47395 159640
rect 47705 159560 47715 159640
rect 48025 159560 48035 159640
rect 48345 159560 48355 159640
rect 48500 159550 48605 159720
rect 48640 159640 48650 159720
rect 48790 159640 48800 159720
rect 49180 159670 49210 159700
rect 49300 159670 49330 159700
rect 49420 159670 49450 159700
rect 49540 159670 49570 159700
rect 49660 159670 49690 159700
rect 49780 159670 49810 159700
rect 49900 159670 49930 159700
rect 50020 159670 50050 159700
rect 50140 159670 50170 159700
rect 50260 159670 50290 159700
rect 50380 159670 50410 159700
rect 50500 159670 50530 159700
rect 50620 159670 50650 159700
rect 50740 159670 50770 159700
rect 50860 159670 50890 159700
rect 50980 159670 51010 159700
rect 51100 159670 51130 159700
rect 51220 159670 51250 159700
rect 51340 159670 51370 159700
rect 51460 159670 51490 159700
rect 51580 159670 51610 159700
rect 51700 159670 51730 159700
rect 51820 159670 51850 159700
rect 51940 159670 51970 159700
rect 52060 159670 52090 159700
rect 52180 159670 52210 159700
rect 52300 159670 52330 159700
rect 52420 159670 52450 159700
rect 52540 159670 52570 159700
rect 52660 159670 52690 159700
rect 52780 159670 52810 159700
rect 52900 159670 52930 159700
rect 53020 159670 53050 159700
rect 53140 159670 53170 159700
rect 53260 159670 53290 159700
rect 53380 159670 53410 159700
rect 53500 159670 53530 159700
rect 53620 159670 53650 159700
rect 53740 159670 53770 159700
rect 53860 159670 53890 159700
rect 53980 159670 54010 159700
rect 54100 159670 54130 159700
rect 54220 159670 54250 159700
rect 54340 159670 54370 159700
rect 54460 159670 54490 159700
rect 54580 159670 54610 159700
rect 54700 159670 54730 159700
rect 54820 159670 54850 159700
rect 54940 159670 54970 159700
rect 55060 159670 55090 159700
rect 55180 159670 55210 159700
rect 55300 159670 55330 159700
rect 55420 159670 55450 159700
rect 55540 159670 55570 159700
rect 55660 159670 55690 159700
rect 55780 159670 55810 159700
rect 55900 159670 55930 159700
rect 56020 159670 56050 159700
rect 56140 159670 56170 159700
rect 56260 159670 56290 159700
rect 56380 159670 56410 159700
rect 56500 159670 56530 159700
rect 56620 159670 56650 159700
rect 56740 159670 56770 159700
rect 56860 159670 56890 159700
rect 56980 159670 57010 159700
rect 57100 159670 57130 159700
rect 57220 159670 57250 159700
rect 57340 159670 57370 159700
rect 57460 159670 57490 159700
rect 57580 159670 57610 159700
rect 57700 159670 57730 159700
rect 57820 159670 57850 159700
rect 57940 159670 57970 159700
rect 58060 159670 58090 159700
rect 58180 159670 58210 159700
rect 58300 159670 58330 159700
rect 58420 159670 58450 159700
rect 58540 159670 58570 159700
rect 58660 159670 58690 159700
rect 58780 159670 58810 159700
rect 58900 159670 58930 159700
rect 59020 159670 59050 159700
rect 59140 159670 59170 159700
rect 59260 159670 59290 159700
rect 59380 159670 59410 159700
rect 59500 159670 59530 159700
rect 59620 159670 59650 159700
rect 59740 159670 59770 159700
rect 59860 159670 59890 159700
rect 49060 159640 49120 159670
rect 49180 159640 49240 159670
rect 49300 159640 49360 159670
rect 49420 159640 49480 159670
rect 49540 159640 49600 159670
rect 49660 159640 49720 159670
rect 49780 159640 49840 159670
rect 49900 159640 49960 159670
rect 50020 159640 50080 159670
rect 50140 159640 50200 159670
rect 50260 159640 50320 159670
rect 50380 159640 50440 159670
rect 50500 159640 50560 159670
rect 50620 159640 50680 159670
rect 50740 159640 50800 159670
rect 50860 159640 50920 159670
rect 50980 159640 51040 159670
rect 51100 159640 51160 159670
rect 51220 159640 51280 159670
rect 51340 159640 51400 159670
rect 51460 159640 51520 159670
rect 51580 159640 51640 159670
rect 51700 159640 51760 159670
rect 51820 159640 51880 159670
rect 51940 159640 52000 159670
rect 52060 159640 52120 159670
rect 52180 159640 52240 159670
rect 52300 159640 52360 159670
rect 52420 159640 52480 159670
rect 52540 159640 52600 159670
rect 52660 159640 52720 159670
rect 52780 159640 52840 159670
rect 52900 159640 52960 159670
rect 53020 159640 53080 159670
rect 53140 159640 53200 159670
rect 53260 159640 53320 159670
rect 53380 159640 53440 159670
rect 53500 159640 53560 159670
rect 53620 159640 53680 159670
rect 53740 159640 53800 159670
rect 53860 159640 53920 159670
rect 53980 159640 54040 159670
rect 54100 159640 54160 159670
rect 54220 159640 54280 159670
rect 54340 159640 54400 159670
rect 54460 159640 54520 159670
rect 54580 159640 54640 159670
rect 54700 159640 54760 159670
rect 54820 159640 54880 159670
rect 54940 159640 55000 159670
rect 55060 159640 55120 159670
rect 55180 159640 55240 159670
rect 55300 159640 55360 159670
rect 55420 159640 55480 159670
rect 55540 159640 55600 159670
rect 55660 159640 55720 159670
rect 55780 159640 55840 159670
rect 55900 159640 55960 159670
rect 56020 159640 56080 159670
rect 56140 159640 56200 159670
rect 56260 159640 56320 159670
rect 56380 159640 56440 159670
rect 56500 159640 56560 159670
rect 56620 159640 56680 159670
rect 56740 159640 56800 159670
rect 56860 159640 56920 159670
rect 56980 159640 57040 159670
rect 57100 159640 57160 159670
rect 57220 159640 57280 159670
rect 57340 159640 57400 159670
rect 57460 159640 57520 159670
rect 57580 159640 57640 159670
rect 57700 159640 57760 159670
rect 57820 159640 57880 159670
rect 57940 159640 58000 159670
rect 58060 159640 58120 159670
rect 58180 159640 58240 159670
rect 58300 159640 58360 159670
rect 58420 159640 58480 159670
rect 58540 159640 58600 159670
rect 58660 159640 58720 159670
rect 58780 159640 58840 159670
rect 58900 159640 58960 159670
rect 59020 159640 59080 159670
rect 59140 159640 59200 159670
rect 59260 159640 59320 159670
rect 59380 159640 59440 159670
rect 59500 159640 59560 159670
rect 59620 159640 59680 159670
rect 59740 159640 59800 159670
rect 59860 159640 59920 159670
rect 60140 159640 60150 159720
rect 60290 159640 60300 159720
rect 60440 159640 60450 159720
rect 60580 159639 60660 159649
rect 60900 159639 60980 159649
rect 61320 159639 61400 159649
rect 61640 159639 61720 159649
rect 62140 159640 62150 159720
rect 62290 159640 62300 159720
rect 62680 159670 62710 159700
rect 73245 159670 73270 159700
rect 73360 159670 73390 159700
rect 62560 159640 62620 159670
rect 62680 159640 62740 159670
rect 73245 159640 73300 159670
rect 73360 159640 73420 159670
rect 73640 159640 73650 159720
rect 73790 159640 73800 159720
rect 73940 159640 73950 159720
rect 74080 159639 74160 159649
rect 74400 159639 74480 159649
rect 74820 159639 74900 159649
rect 75140 159639 75220 159649
rect 75640 159640 75650 159720
rect 75790 159640 75800 159720
rect 76180 159670 76210 159700
rect 86745 159670 86770 159700
rect 86860 159670 86890 159700
rect 76060 159640 76120 159670
rect 76180 159640 76240 159670
rect 86745 159640 86800 159670
rect 86860 159640 86920 159670
rect 87140 159640 87150 159720
rect 87290 159640 87300 159720
rect 87440 159640 87450 159720
rect 87580 159639 87660 159649
rect 87900 159639 87980 159649
rect 88320 159639 88400 159649
rect 88640 159639 88720 159649
rect 89140 159640 89150 159720
rect 89290 159640 89300 159720
rect 89680 159670 89710 159700
rect 100245 159670 100270 159700
rect 100360 159670 100390 159700
rect 89560 159640 89620 159670
rect 89680 159640 89740 159670
rect 100245 159640 100300 159670
rect 100360 159640 100420 159670
rect 100640 159640 100650 159720
rect 100790 159640 100800 159720
rect 100940 159640 100950 159720
rect 101080 159639 101160 159649
rect 101400 159639 101480 159649
rect 101820 159639 101900 159649
rect 102140 159639 102220 159649
rect 114580 159639 114660 159649
rect 114900 159639 114980 159649
rect 115320 159639 115400 159649
rect 115640 159639 115720 159649
rect 116140 159640 116150 159720
rect 116290 159640 116300 159720
rect 116680 159670 116710 159700
rect 127245 159670 127270 159700
rect 127360 159670 127390 159700
rect 116560 159640 116620 159670
rect 116680 159640 116740 159670
rect 127245 159640 127300 159670
rect 127360 159640 127420 159670
rect 127640 159640 127650 159720
rect 127790 159640 127800 159720
rect 127940 159640 127950 159720
rect 128080 159639 128160 159649
rect 128400 159639 128480 159649
rect 128820 159639 128900 159649
rect 129140 159639 129220 159649
rect 129640 159640 129650 159720
rect 129790 159640 129800 159720
rect 130180 159670 130210 159700
rect 140740 159670 140770 159700
rect 140860 159670 140890 159700
rect 130060 159640 130120 159670
rect 130180 159640 130240 159670
rect 140740 159640 140800 159670
rect 140860 159640 140920 159670
rect 141140 159640 141150 159720
rect 141290 159640 141300 159720
rect 141440 159640 141450 159720
rect 141545 159640 141625 159650
rect 141865 159640 141945 159650
rect 142185 159640 142200 159650
rect 145385 159640 145465 159650
rect 145705 159640 145785 159650
rect 146025 159640 146105 159650
rect 49180 159550 49210 159580
rect 49300 159550 49330 159580
rect 49420 159550 49450 159580
rect 49540 159550 49570 159580
rect 49660 159550 49690 159580
rect 49780 159550 49810 159580
rect 49900 159550 49930 159580
rect 50020 159550 50050 159580
rect 50140 159550 50170 159580
rect 50260 159550 50290 159580
rect 50380 159550 50410 159580
rect 50500 159550 50530 159580
rect 50620 159550 50650 159580
rect 50740 159550 50770 159580
rect 50860 159550 50890 159580
rect 50980 159550 51010 159580
rect 51100 159550 51130 159580
rect 51220 159550 51250 159580
rect 51340 159550 51370 159580
rect 51460 159550 51490 159580
rect 51580 159550 51610 159580
rect 51700 159550 51730 159580
rect 51820 159550 51850 159580
rect 51940 159550 51970 159580
rect 52060 159550 52090 159580
rect 52180 159550 52210 159580
rect 52300 159550 52330 159580
rect 52420 159550 52450 159580
rect 52540 159550 52570 159580
rect 52660 159550 52690 159580
rect 52780 159550 52810 159580
rect 52900 159550 52930 159580
rect 53020 159550 53050 159580
rect 53140 159550 53170 159580
rect 53260 159550 53290 159580
rect 53380 159550 53410 159580
rect 53500 159550 53530 159580
rect 53620 159550 53650 159580
rect 53740 159550 53770 159580
rect 53860 159550 53890 159580
rect 53980 159550 54010 159580
rect 54100 159550 54130 159580
rect 54220 159550 54250 159580
rect 54340 159550 54370 159580
rect 54460 159550 54490 159580
rect 54580 159550 54610 159580
rect 54700 159550 54730 159580
rect 54820 159550 54850 159580
rect 54940 159550 54970 159580
rect 55060 159550 55090 159580
rect 55180 159550 55210 159580
rect 55300 159550 55330 159580
rect 55420 159550 55450 159580
rect 55540 159550 55570 159580
rect 55660 159550 55690 159580
rect 55780 159550 55810 159580
rect 55900 159550 55930 159580
rect 56020 159550 56050 159580
rect 56140 159550 56170 159580
rect 56260 159550 56290 159580
rect 56380 159550 56410 159580
rect 56500 159550 56530 159580
rect 56620 159550 56650 159580
rect 56740 159550 56770 159580
rect 56860 159550 56890 159580
rect 56980 159550 57010 159580
rect 57100 159550 57130 159580
rect 57220 159550 57250 159580
rect 57340 159550 57370 159580
rect 57460 159550 57490 159580
rect 57580 159550 57610 159580
rect 57700 159550 57730 159580
rect 57820 159550 57850 159580
rect 57940 159550 57970 159580
rect 58060 159550 58090 159580
rect 58180 159550 58210 159580
rect 58300 159550 58330 159580
rect 58420 159550 58450 159580
rect 58540 159550 58570 159580
rect 58660 159550 58690 159580
rect 58780 159550 58810 159580
rect 58900 159550 58930 159580
rect 59020 159550 59050 159580
rect 59140 159550 59170 159580
rect 59260 159550 59290 159580
rect 59380 159550 59410 159580
rect 59500 159550 59530 159580
rect 59620 159550 59650 159580
rect 59740 159550 59770 159580
rect 59860 159550 59890 159580
rect 60660 159559 60670 159639
rect 60980 159559 60990 159639
rect 61400 159559 61410 159639
rect 61720 159559 61730 159639
rect 62680 159550 62710 159580
rect 73245 159550 73270 159580
rect 73360 159550 73390 159580
rect 74160 159559 74170 159639
rect 74480 159559 74490 159639
rect 74900 159559 74910 159639
rect 75220 159559 75230 159639
rect 76180 159550 76210 159580
rect 86745 159550 86770 159580
rect 86860 159550 86890 159580
rect 87660 159559 87670 159639
rect 87980 159559 87990 159639
rect 88400 159559 88410 159639
rect 88720 159559 88730 159639
rect 89680 159550 89710 159580
rect 100245 159550 100270 159580
rect 100360 159550 100390 159580
rect 101160 159559 101170 159639
rect 101480 159559 101490 159639
rect 101900 159559 101910 159639
rect 102220 159559 102230 159639
rect 114660 159559 114670 159639
rect 114980 159559 114990 159639
rect 115400 159559 115410 159639
rect 115720 159559 115730 159639
rect 116680 159550 116710 159580
rect 127245 159550 127270 159580
rect 127360 159550 127390 159580
rect 128160 159559 128170 159639
rect 128480 159559 128490 159639
rect 128900 159559 128910 159639
rect 129220 159559 129230 159639
rect 130180 159550 130210 159580
rect 140740 159550 140770 159580
rect 140860 159550 140890 159580
rect 141625 159560 141635 159640
rect 141945 159560 141955 159640
rect 145465 159560 145475 159640
rect 145785 159560 145795 159640
rect 146105 159560 146115 159640
rect 146700 159580 146780 159590
rect 48500 159540 48640 159550
rect 48710 159540 48790 159550
rect 43945 159480 44025 159490
rect 44265 159480 44345 159490
rect 44585 159480 44665 159490
rect 44905 159480 44985 159490
rect 45225 159480 45305 159490
rect 45545 159480 45625 159490
rect 45865 159480 45945 159490
rect 46185 159480 46265 159490
rect 46505 159480 46585 159490
rect 46825 159480 46905 159490
rect 47145 159480 47225 159490
rect 47465 159480 47545 159490
rect 47785 159480 47865 159490
rect 48105 159480 48185 159490
rect 43060 159420 43140 159430
rect 43380 159420 43460 159430
rect 43140 159340 43150 159420
rect 43460 159340 43470 159420
rect 44025 159400 44035 159480
rect 44345 159400 44355 159480
rect 44665 159400 44675 159480
rect 44985 159400 44995 159480
rect 45305 159400 45315 159480
rect 45625 159400 45635 159480
rect 45945 159400 45955 159480
rect 46265 159400 46275 159480
rect 46585 159400 46595 159480
rect 46905 159400 46915 159480
rect 47225 159400 47235 159480
rect 47545 159400 47555 159480
rect 47865 159400 47875 159480
rect 48185 159400 48195 159480
rect 48500 159370 48605 159540
rect 48640 159460 48650 159540
rect 48790 159460 48800 159540
rect 49060 159520 49120 159550
rect 49180 159520 49240 159550
rect 49300 159520 49360 159550
rect 49420 159520 49480 159550
rect 49540 159520 49600 159550
rect 49660 159520 49720 159550
rect 49780 159520 49840 159550
rect 49900 159520 49960 159550
rect 50020 159520 50080 159550
rect 50140 159520 50200 159550
rect 50260 159520 50320 159550
rect 50380 159520 50440 159550
rect 50500 159520 50560 159550
rect 50620 159520 50680 159550
rect 50740 159520 50800 159550
rect 50860 159520 50920 159550
rect 50980 159520 51040 159550
rect 51100 159520 51160 159550
rect 51220 159520 51280 159550
rect 51340 159520 51400 159550
rect 51460 159520 51520 159550
rect 51580 159520 51640 159550
rect 51700 159520 51760 159550
rect 51820 159520 51880 159550
rect 51940 159520 52000 159550
rect 52060 159520 52120 159550
rect 52180 159520 52240 159550
rect 52300 159520 52360 159550
rect 52420 159520 52480 159550
rect 52540 159520 52600 159550
rect 52660 159520 52720 159550
rect 52780 159520 52840 159550
rect 52900 159520 52960 159550
rect 53020 159520 53080 159550
rect 53140 159520 53200 159550
rect 53260 159520 53320 159550
rect 53380 159520 53440 159550
rect 53500 159520 53560 159550
rect 53620 159520 53680 159550
rect 53740 159520 53800 159550
rect 53860 159520 53920 159550
rect 53980 159520 54040 159550
rect 54100 159520 54160 159550
rect 54220 159520 54280 159550
rect 54340 159520 54400 159550
rect 54460 159520 54520 159550
rect 54580 159520 54640 159550
rect 54700 159520 54760 159550
rect 54820 159520 54880 159550
rect 54940 159520 55000 159550
rect 55060 159520 55120 159550
rect 55180 159520 55240 159550
rect 55300 159520 55360 159550
rect 55420 159520 55480 159550
rect 55540 159520 55600 159550
rect 55660 159520 55720 159550
rect 55780 159520 55840 159550
rect 55900 159520 55960 159550
rect 56020 159520 56080 159550
rect 56140 159520 56200 159550
rect 56260 159520 56320 159550
rect 56380 159520 56440 159550
rect 56500 159520 56560 159550
rect 56620 159520 56680 159550
rect 56740 159520 56800 159550
rect 56860 159520 56920 159550
rect 56980 159520 57040 159550
rect 57100 159520 57160 159550
rect 57220 159520 57280 159550
rect 57340 159520 57400 159550
rect 57460 159520 57520 159550
rect 57580 159520 57640 159550
rect 57700 159520 57760 159550
rect 57820 159520 57880 159550
rect 57940 159520 58000 159550
rect 58060 159520 58120 159550
rect 58180 159520 58240 159550
rect 58300 159520 58360 159550
rect 58420 159520 58480 159550
rect 58540 159520 58600 159550
rect 58660 159520 58720 159550
rect 58780 159520 58840 159550
rect 58900 159520 58960 159550
rect 59020 159520 59080 159550
rect 59140 159520 59200 159550
rect 59260 159520 59320 159550
rect 59380 159520 59440 159550
rect 59500 159520 59560 159550
rect 59620 159520 59680 159550
rect 59740 159520 59800 159550
rect 59860 159520 59920 159550
rect 60060 159540 60140 159550
rect 60210 159540 60290 159550
rect 60360 159540 60440 159550
rect 62060 159540 62140 159550
rect 62210 159540 62290 159550
rect 60140 159460 60150 159540
rect 60290 159460 60300 159540
rect 60440 159460 60450 159540
rect 60740 159479 60820 159489
rect 61060 159479 61140 159489
rect 61480 159479 61560 159489
rect 61800 159479 61880 159489
rect 49180 159400 49210 159460
rect 49300 159400 49330 159460
rect 49420 159400 49450 159460
rect 49540 159400 49570 159460
rect 49660 159400 49690 159460
rect 49780 159400 49810 159460
rect 49900 159400 49930 159460
rect 50020 159400 50050 159460
rect 50140 159400 50170 159460
rect 50260 159400 50290 159460
rect 50380 159400 50410 159460
rect 50500 159400 50530 159460
rect 50620 159400 50650 159460
rect 50740 159400 50770 159460
rect 50860 159400 50890 159460
rect 50980 159400 51010 159460
rect 51100 159400 51130 159460
rect 51220 159400 51250 159460
rect 51340 159400 51370 159460
rect 51460 159400 51490 159460
rect 51580 159400 51610 159460
rect 51700 159400 51730 159460
rect 51820 159400 51850 159460
rect 51940 159400 51970 159460
rect 52060 159400 52090 159460
rect 52180 159400 52210 159460
rect 52300 159400 52330 159460
rect 52420 159400 52450 159460
rect 52540 159400 52570 159460
rect 52660 159400 52690 159460
rect 52780 159400 52810 159460
rect 52900 159400 52930 159460
rect 53020 159400 53050 159460
rect 53140 159400 53170 159460
rect 53260 159400 53290 159460
rect 53380 159400 53410 159460
rect 53500 159400 53530 159460
rect 53620 159400 53650 159460
rect 53740 159400 53770 159460
rect 53860 159400 53890 159460
rect 53980 159400 54010 159460
rect 54100 159400 54130 159460
rect 54220 159400 54250 159460
rect 54340 159400 54370 159460
rect 54460 159400 54490 159460
rect 54580 159400 54610 159460
rect 54700 159400 54730 159460
rect 54820 159400 54850 159460
rect 54940 159400 54970 159460
rect 55060 159400 55090 159460
rect 55180 159400 55210 159460
rect 55300 159400 55330 159460
rect 55420 159400 55450 159460
rect 55540 159400 55570 159460
rect 55660 159400 55690 159460
rect 55780 159400 55810 159460
rect 55900 159400 55930 159460
rect 56020 159400 56050 159460
rect 56140 159400 56170 159460
rect 56260 159400 56290 159460
rect 56380 159400 56410 159460
rect 56500 159400 56530 159460
rect 56620 159400 56650 159460
rect 56740 159400 56770 159460
rect 56860 159400 56890 159460
rect 56980 159400 57010 159460
rect 57100 159400 57130 159460
rect 57220 159400 57250 159460
rect 57340 159400 57370 159460
rect 57460 159400 57490 159460
rect 57580 159400 57610 159460
rect 57700 159400 57730 159460
rect 57820 159400 57850 159460
rect 57940 159400 57970 159460
rect 58060 159400 58090 159460
rect 58180 159400 58210 159460
rect 58300 159400 58330 159460
rect 58420 159400 58450 159460
rect 58540 159400 58570 159460
rect 58660 159400 58690 159460
rect 58780 159400 58810 159460
rect 58900 159400 58930 159460
rect 59020 159400 59050 159460
rect 59140 159400 59170 159460
rect 59260 159400 59290 159460
rect 59380 159400 59410 159460
rect 59500 159400 59530 159460
rect 59620 159400 59650 159460
rect 59740 159400 59770 159460
rect 59860 159400 59890 159460
rect 60820 159399 60830 159479
rect 61140 159399 61150 159479
rect 61560 159399 61570 159479
rect 61880 159399 61890 159479
rect 62140 159460 62150 159540
rect 62290 159460 62300 159540
rect 62560 159520 62620 159550
rect 62680 159520 62740 159550
rect 73245 159520 73300 159550
rect 73360 159520 73420 159550
rect 73560 159540 73640 159550
rect 73710 159540 73790 159550
rect 73860 159540 73940 159550
rect 75560 159540 75640 159550
rect 75710 159540 75790 159550
rect 73640 159460 73650 159540
rect 73790 159460 73800 159540
rect 73940 159460 73950 159540
rect 74240 159479 74320 159489
rect 74560 159479 74640 159489
rect 74980 159479 75060 159489
rect 75300 159479 75380 159489
rect 62680 159400 62710 159460
rect 73245 159400 73270 159460
rect 73360 159400 73390 159460
rect 74320 159399 74330 159479
rect 74640 159399 74650 159479
rect 75060 159399 75070 159479
rect 75380 159399 75390 159479
rect 75640 159460 75650 159540
rect 75790 159460 75800 159540
rect 76060 159520 76120 159550
rect 76180 159520 76240 159550
rect 86745 159520 86800 159550
rect 86860 159520 86920 159550
rect 87060 159540 87140 159550
rect 87210 159540 87290 159550
rect 87360 159540 87440 159550
rect 89060 159540 89140 159550
rect 89210 159540 89290 159550
rect 87140 159460 87150 159540
rect 87290 159460 87300 159540
rect 87440 159460 87450 159540
rect 87740 159479 87820 159489
rect 88060 159479 88140 159489
rect 88480 159479 88560 159489
rect 88800 159479 88880 159489
rect 76180 159400 76210 159460
rect 86745 159400 86770 159460
rect 86860 159400 86890 159460
rect 87820 159399 87830 159479
rect 88140 159399 88150 159479
rect 88560 159399 88570 159479
rect 88880 159399 88890 159479
rect 89140 159460 89150 159540
rect 89290 159460 89300 159540
rect 89560 159520 89620 159550
rect 89680 159520 89740 159550
rect 100245 159520 100300 159550
rect 100360 159520 100420 159550
rect 100560 159540 100640 159550
rect 100710 159540 100790 159550
rect 100860 159540 100940 159550
rect 116060 159540 116140 159550
rect 116210 159540 116290 159550
rect 100640 159460 100650 159540
rect 100790 159460 100800 159540
rect 100940 159460 100950 159540
rect 101240 159479 101320 159489
rect 101560 159479 101640 159489
rect 101980 159479 102060 159489
rect 102300 159479 102380 159489
rect 114740 159479 114820 159489
rect 115060 159479 115140 159489
rect 115480 159479 115560 159489
rect 115800 159479 115880 159489
rect 89680 159400 89710 159460
rect 100245 159400 100270 159460
rect 100360 159400 100390 159460
rect 101320 159399 101330 159479
rect 101640 159399 101650 159479
rect 102060 159399 102070 159479
rect 102380 159399 102390 159479
rect 114820 159399 114830 159479
rect 115140 159399 115150 159479
rect 115560 159399 115570 159479
rect 115880 159399 115890 159479
rect 116140 159460 116150 159540
rect 116290 159460 116300 159540
rect 116560 159520 116620 159550
rect 116680 159520 116740 159550
rect 127245 159520 127300 159550
rect 127360 159520 127420 159550
rect 127560 159540 127640 159550
rect 127710 159540 127790 159550
rect 127860 159540 127940 159550
rect 129560 159540 129640 159550
rect 129710 159540 129790 159550
rect 127640 159460 127650 159540
rect 127790 159460 127800 159540
rect 127940 159460 127950 159540
rect 128240 159479 128320 159489
rect 128560 159479 128640 159489
rect 128980 159479 129060 159489
rect 129300 159479 129380 159489
rect 116680 159400 116710 159460
rect 127245 159400 127270 159460
rect 127360 159400 127390 159460
rect 128320 159399 128330 159479
rect 128640 159399 128650 159479
rect 129060 159399 129070 159479
rect 129380 159399 129390 159479
rect 129640 159460 129650 159540
rect 129790 159460 129800 159540
rect 130060 159520 130120 159550
rect 130180 159520 130240 159550
rect 140740 159520 140800 159550
rect 140860 159520 140920 159550
rect 141060 159540 141140 159550
rect 141210 159540 141290 159550
rect 141360 159540 141440 159550
rect 141140 159460 141150 159540
rect 141290 159460 141300 159540
rect 141440 159460 141450 159540
rect 146780 159500 146790 159580
rect 141705 159480 141785 159490
rect 142025 159480 142105 159490
rect 145225 159480 145305 159490
rect 145545 159480 145625 159490
rect 145865 159480 145945 159490
rect 130180 159400 130210 159460
rect 140740 159400 140770 159460
rect 140860 159400 140890 159460
rect 141785 159400 141795 159480
rect 142105 159400 142115 159480
rect 145305 159400 145315 159480
rect 145625 159400 145635 159480
rect 145945 159400 145955 159480
rect 146540 159420 146620 159430
rect 146860 159420 146940 159430
rect 48500 159360 48640 159370
rect 48710 159360 48790 159370
rect 60060 159360 60140 159370
rect 60210 159360 60290 159370
rect 60360 159360 60440 159370
rect 62060 159360 62140 159370
rect 62210 159360 62290 159370
rect 73560 159360 73640 159370
rect 73710 159360 73790 159370
rect 73860 159360 73940 159370
rect 75560 159360 75640 159370
rect 75710 159360 75790 159370
rect 87060 159360 87140 159370
rect 87210 159360 87290 159370
rect 87360 159360 87440 159370
rect 89060 159360 89140 159370
rect 89210 159360 89290 159370
rect 100560 159360 100640 159370
rect 100710 159360 100790 159370
rect 100860 159360 100940 159370
rect 116060 159360 116140 159370
rect 116210 159360 116290 159370
rect 127560 159360 127640 159370
rect 127710 159360 127790 159370
rect 127860 159360 127940 159370
rect 129560 159360 129640 159370
rect 129710 159360 129790 159370
rect 141060 159360 141140 159370
rect 141210 159360 141290 159370
rect 141360 159360 141440 159370
rect 43785 159320 43865 159330
rect 44105 159320 44185 159330
rect 44425 159320 44505 159330
rect 44745 159320 44825 159330
rect 45065 159320 45145 159330
rect 45385 159320 45465 159330
rect 45705 159320 45785 159330
rect 46025 159320 46105 159330
rect 46345 159320 46425 159330
rect 46665 159320 46745 159330
rect 46985 159320 47065 159330
rect 47305 159320 47385 159330
rect 47625 159320 47705 159330
rect 47945 159320 48025 159330
rect 48265 159320 48345 159330
rect 42950 159260 42980 159270
rect 43220 159260 43300 159270
rect 42980 159180 42990 159260
rect 43300 159180 43310 159260
rect 43865 159240 43875 159320
rect 44185 159240 44195 159320
rect 44505 159240 44515 159320
rect 44825 159240 44835 159320
rect 45145 159240 45155 159320
rect 45465 159240 45475 159320
rect 45785 159240 45795 159320
rect 46105 159240 46115 159320
rect 46425 159240 46435 159320
rect 46745 159240 46755 159320
rect 47065 159240 47075 159320
rect 47385 159240 47395 159320
rect 47705 159240 47715 159320
rect 48025 159240 48035 159320
rect 48345 159240 48355 159320
rect 48500 159190 48605 159360
rect 48640 159280 48650 159360
rect 48790 159280 48800 159360
rect 60140 159280 60150 159360
rect 60290 159280 60300 159360
rect 60440 159280 60450 159360
rect 60580 159319 60660 159329
rect 60900 159319 60980 159329
rect 61320 159319 61400 159329
rect 61640 159319 61720 159329
rect 60660 159239 60670 159319
rect 60980 159239 60990 159319
rect 61400 159239 61410 159319
rect 61720 159239 61730 159319
rect 62140 159280 62150 159360
rect 62290 159280 62300 159360
rect 73640 159280 73650 159360
rect 73790 159280 73800 159360
rect 73940 159280 73950 159360
rect 74080 159319 74160 159329
rect 74400 159319 74480 159329
rect 74820 159319 74900 159329
rect 75140 159319 75220 159329
rect 74160 159239 74170 159319
rect 74480 159239 74490 159319
rect 74900 159239 74910 159319
rect 75220 159239 75230 159319
rect 75640 159280 75650 159360
rect 75790 159280 75800 159360
rect 87140 159280 87150 159360
rect 87290 159280 87300 159360
rect 87440 159280 87450 159360
rect 87580 159319 87660 159329
rect 87900 159319 87980 159329
rect 88320 159319 88400 159329
rect 88640 159319 88720 159329
rect 87660 159239 87670 159319
rect 87980 159239 87990 159319
rect 88400 159239 88410 159319
rect 88720 159239 88730 159319
rect 89140 159280 89150 159360
rect 89290 159280 89300 159360
rect 100640 159280 100650 159360
rect 100790 159280 100800 159360
rect 100940 159280 100950 159360
rect 101080 159319 101160 159329
rect 101400 159319 101480 159329
rect 101820 159319 101900 159329
rect 102140 159319 102220 159329
rect 114580 159319 114660 159329
rect 114900 159319 114980 159329
rect 115320 159319 115400 159329
rect 115640 159319 115720 159329
rect 101160 159239 101170 159319
rect 101480 159239 101490 159319
rect 101900 159239 101910 159319
rect 102220 159239 102230 159319
rect 114660 159239 114670 159319
rect 114980 159239 114990 159319
rect 115400 159239 115410 159319
rect 115720 159239 115730 159319
rect 116140 159280 116150 159360
rect 116290 159280 116300 159360
rect 127640 159280 127650 159360
rect 127790 159280 127800 159360
rect 127940 159280 127950 159360
rect 128080 159319 128160 159329
rect 128400 159319 128480 159329
rect 128820 159319 128900 159329
rect 129140 159319 129220 159329
rect 128160 159239 128170 159319
rect 128480 159239 128490 159319
rect 128900 159239 128910 159319
rect 129220 159239 129230 159319
rect 129640 159280 129650 159360
rect 129790 159280 129800 159360
rect 141140 159280 141150 159360
rect 141290 159280 141300 159360
rect 141440 159280 141450 159360
rect 146620 159340 146630 159420
rect 146940 159340 146950 159420
rect 141545 159320 141625 159330
rect 141865 159320 141945 159330
rect 142185 159320 142200 159330
rect 145385 159320 145465 159330
rect 145705 159320 145785 159330
rect 146025 159320 146105 159330
rect 141625 159240 141635 159320
rect 141945 159240 141955 159320
rect 145465 159240 145475 159320
rect 145785 159240 145795 159320
rect 146105 159240 146115 159320
rect 146700 159260 146780 159270
rect 48500 159180 48640 159190
rect 48710 159180 48790 159190
rect 60060 159180 60140 159190
rect 60210 159180 60290 159190
rect 60360 159180 60440 159190
rect 62060 159180 62140 159190
rect 62210 159180 62290 159190
rect 73560 159180 73640 159190
rect 73710 159180 73790 159190
rect 73860 159180 73940 159190
rect 75560 159180 75640 159190
rect 75710 159180 75790 159190
rect 87060 159180 87140 159190
rect 87210 159180 87290 159190
rect 87360 159180 87440 159190
rect 89060 159180 89140 159190
rect 89210 159180 89290 159190
rect 100560 159180 100640 159190
rect 100710 159180 100790 159190
rect 100860 159180 100940 159190
rect 116060 159180 116140 159190
rect 116210 159180 116290 159190
rect 127560 159180 127640 159190
rect 127710 159180 127790 159190
rect 127860 159180 127940 159190
rect 129560 159180 129640 159190
rect 129710 159180 129790 159190
rect 141060 159180 141140 159190
rect 141210 159180 141290 159190
rect 141360 159180 141440 159190
rect 146780 159180 146790 159260
rect 43945 159160 44025 159170
rect 44265 159160 44345 159170
rect 44585 159160 44665 159170
rect 44905 159160 44985 159170
rect 45225 159160 45305 159170
rect 45545 159160 45625 159170
rect 45865 159160 45945 159170
rect 46185 159160 46265 159170
rect 46505 159160 46585 159170
rect 46825 159160 46905 159170
rect 47145 159160 47225 159170
rect 47465 159160 47545 159170
rect 47785 159160 47865 159170
rect 48105 159160 48185 159170
rect 43060 159100 43140 159110
rect 43380 159100 43460 159110
rect 43140 159020 43150 159100
rect 43460 159020 43470 159100
rect 44025 159080 44035 159160
rect 44345 159080 44355 159160
rect 44665 159080 44675 159160
rect 44985 159080 44995 159160
rect 45305 159080 45315 159160
rect 45625 159080 45635 159160
rect 45945 159080 45955 159160
rect 46265 159080 46275 159160
rect 46585 159080 46595 159160
rect 46905 159080 46915 159160
rect 47225 159080 47235 159160
rect 47545 159080 47555 159160
rect 47865 159080 47875 159160
rect 48185 159080 48195 159160
rect 48500 159010 48605 159180
rect 48640 159100 48650 159180
rect 48790 159100 48800 159180
rect 60140 159100 60150 159180
rect 60290 159100 60300 159180
rect 60440 159100 60450 159180
rect 60740 159159 60820 159169
rect 61060 159159 61140 159169
rect 61480 159159 61560 159169
rect 61800 159159 61880 159169
rect 60820 159079 60830 159159
rect 61140 159079 61150 159159
rect 61560 159079 61570 159159
rect 61880 159079 61890 159159
rect 62140 159100 62150 159180
rect 62290 159100 62300 159180
rect 73640 159100 73650 159180
rect 73790 159100 73800 159180
rect 73940 159100 73950 159180
rect 74240 159159 74320 159169
rect 74560 159159 74640 159169
rect 74980 159159 75060 159169
rect 75300 159159 75380 159169
rect 74320 159079 74330 159159
rect 74640 159079 74650 159159
rect 75060 159079 75070 159159
rect 75380 159079 75390 159159
rect 75640 159100 75650 159180
rect 75790 159100 75800 159180
rect 87140 159100 87150 159180
rect 87290 159100 87300 159180
rect 87440 159100 87450 159180
rect 87740 159159 87820 159169
rect 88060 159159 88140 159169
rect 88480 159159 88560 159169
rect 88800 159159 88880 159169
rect 87820 159079 87830 159159
rect 88140 159079 88150 159159
rect 88560 159079 88570 159159
rect 88880 159079 88890 159159
rect 89140 159100 89150 159180
rect 89290 159100 89300 159180
rect 100640 159100 100650 159180
rect 100790 159100 100800 159180
rect 100940 159100 100950 159180
rect 101240 159159 101320 159169
rect 101560 159159 101640 159169
rect 101980 159159 102060 159169
rect 102300 159159 102380 159169
rect 114740 159159 114820 159169
rect 115060 159159 115140 159169
rect 115480 159159 115560 159169
rect 115800 159159 115880 159169
rect 101320 159079 101330 159159
rect 101640 159079 101650 159159
rect 102060 159079 102070 159159
rect 102380 159079 102390 159159
rect 114820 159079 114830 159159
rect 115140 159079 115150 159159
rect 115560 159079 115570 159159
rect 115880 159079 115890 159159
rect 116140 159100 116150 159180
rect 116290 159100 116300 159180
rect 127640 159100 127650 159180
rect 127790 159100 127800 159180
rect 127940 159100 127950 159180
rect 128240 159159 128320 159169
rect 128560 159159 128640 159169
rect 128980 159159 129060 159169
rect 129300 159159 129380 159169
rect 128320 159079 128330 159159
rect 128640 159079 128650 159159
rect 129060 159079 129070 159159
rect 129380 159079 129390 159159
rect 129640 159100 129650 159180
rect 129790 159100 129800 159180
rect 141140 159100 141150 159180
rect 141290 159100 141300 159180
rect 141440 159100 141450 159180
rect 141705 159160 141785 159170
rect 142025 159160 142105 159170
rect 145225 159160 145305 159170
rect 145545 159160 145625 159170
rect 145865 159160 145945 159170
rect 141785 159080 141795 159160
rect 142105 159080 142115 159160
rect 145305 159080 145315 159160
rect 145625 159080 145635 159160
rect 145945 159080 145955 159160
rect 146540 159100 146620 159110
rect 146860 159100 146940 159110
rect 146620 159020 146630 159100
rect 146940 159020 146950 159100
rect 43785 159000 43865 159010
rect 44105 159000 44185 159010
rect 44425 159000 44505 159010
rect 44745 159000 44825 159010
rect 45065 159000 45145 159010
rect 45385 159000 45465 159010
rect 45705 159000 45785 159010
rect 46025 159000 46105 159010
rect 46345 159000 46425 159010
rect 46665 159000 46745 159010
rect 46985 159000 47065 159010
rect 47305 159000 47385 159010
rect 47625 159000 47705 159010
rect 47945 159000 48025 159010
rect 48265 159000 48345 159010
rect 48500 159000 48640 159010
rect 48710 159000 48790 159010
rect 60060 159000 60140 159010
rect 60210 159000 60290 159010
rect 60360 159000 60440 159010
rect 42950 158940 42980 158950
rect 43220 158940 43300 158950
rect 42980 158860 42990 158940
rect 43300 158860 43310 158940
rect 43865 158920 43875 159000
rect 44185 158920 44195 159000
rect 44505 158920 44515 159000
rect 44825 158920 44835 159000
rect 45145 158920 45155 159000
rect 45465 158920 45475 159000
rect 45785 158920 45795 159000
rect 46105 158920 46115 159000
rect 46425 158920 46435 159000
rect 46745 158920 46755 159000
rect 47065 158920 47075 159000
rect 47385 158920 47395 159000
rect 47705 158920 47715 159000
rect 48025 158920 48035 159000
rect 48345 158920 48355 159000
rect 43945 158840 44025 158850
rect 44265 158840 44345 158850
rect 44585 158840 44665 158850
rect 44905 158840 44985 158850
rect 45225 158840 45305 158850
rect 45545 158840 45625 158850
rect 45865 158840 45945 158850
rect 46185 158840 46265 158850
rect 46505 158840 46585 158850
rect 46825 158840 46905 158850
rect 47145 158840 47225 158850
rect 47465 158840 47545 158850
rect 47785 158840 47865 158850
rect 48105 158840 48185 158850
rect 43060 158780 43140 158790
rect 43380 158780 43460 158790
rect 43140 158700 43150 158780
rect 43460 158700 43470 158780
rect 44025 158760 44035 158840
rect 44345 158760 44355 158840
rect 44665 158760 44675 158840
rect 44985 158760 44995 158840
rect 45305 158760 45315 158840
rect 45625 158760 45635 158840
rect 45945 158760 45955 158840
rect 46265 158760 46275 158840
rect 46585 158760 46595 158840
rect 46905 158760 46915 158840
rect 47225 158760 47235 158840
rect 47545 158760 47555 158840
rect 47865 158760 47875 158840
rect 48185 158760 48195 158840
rect 48500 158830 48605 159000
rect 48640 158920 48650 159000
rect 48790 158920 48800 159000
rect 49240 158900 59760 158990
rect 60140 158920 60150 159000
rect 60290 158920 60300 159000
rect 60440 158920 60450 159000
rect 60580 158999 60660 159009
rect 60900 158999 60980 159009
rect 61320 158999 61400 159009
rect 61640 158999 61720 159009
rect 62060 159000 62140 159010
rect 62210 159000 62290 159010
rect 73560 159000 73640 159010
rect 73710 159000 73790 159010
rect 73860 159000 73940 159010
rect 60660 158919 60670 158999
rect 60980 158919 60990 158999
rect 61400 158919 61410 158999
rect 61720 158919 61730 158999
rect 62140 158920 62150 159000
rect 62290 158920 62300 159000
rect 62740 158900 62755 158990
rect 49560 158830 49590 158900
rect 48500 158820 48640 158830
rect 48710 158820 48790 158830
rect 49270 158820 49350 158830
rect 49420 158820 49500 158830
rect 49560 158820 49650 158830
rect 49660 158820 49690 158900
rect 43785 158680 43865 158690
rect 44105 158680 44185 158690
rect 44425 158680 44505 158690
rect 44745 158680 44825 158690
rect 45065 158680 45145 158690
rect 45385 158680 45465 158690
rect 45705 158680 45785 158690
rect 46025 158680 46105 158690
rect 46345 158680 46425 158690
rect 46665 158680 46745 158690
rect 46985 158680 47065 158690
rect 47305 158680 47385 158690
rect 47625 158680 47705 158690
rect 47945 158680 48025 158690
rect 48265 158680 48345 158690
rect 42950 158620 42980 158630
rect 43220 158620 43300 158630
rect 42980 158540 42990 158620
rect 43300 158540 43310 158620
rect 43865 158600 43875 158680
rect 44185 158600 44195 158680
rect 44505 158600 44515 158680
rect 44825 158600 44835 158680
rect 45145 158600 45155 158680
rect 45465 158600 45475 158680
rect 45785 158600 45795 158680
rect 46105 158600 46115 158680
rect 46425 158600 46435 158680
rect 46745 158600 46755 158680
rect 47065 158600 47075 158680
rect 47385 158600 47395 158680
rect 47705 158600 47715 158680
rect 48025 158600 48035 158680
rect 48345 158600 48355 158680
rect 48500 158650 48605 158820
rect 48640 158740 48650 158820
rect 48790 158740 48800 158820
rect 49350 158740 49360 158820
rect 49500 158740 49510 158820
rect 49560 158650 49590 158820
rect 49650 158740 49690 158820
rect 48500 158640 48640 158650
rect 48710 158640 48790 158650
rect 49270 158640 49350 158650
rect 49420 158640 49500 158650
rect 49560 158640 49650 158650
rect 49660 158640 49690 158740
rect 43945 158520 44025 158530
rect 44265 158520 44345 158530
rect 44585 158520 44665 158530
rect 44905 158520 44985 158530
rect 45225 158520 45305 158530
rect 45545 158520 45625 158530
rect 45865 158520 45945 158530
rect 46185 158520 46265 158530
rect 46505 158520 46585 158530
rect 46825 158520 46905 158530
rect 47145 158520 47225 158530
rect 47465 158520 47545 158530
rect 47785 158520 47865 158530
rect 48105 158520 48185 158530
rect 43060 158460 43140 158470
rect 43380 158460 43460 158470
rect 43140 158380 43150 158460
rect 43460 158380 43470 158460
rect 44025 158440 44035 158520
rect 44345 158440 44355 158520
rect 44665 158440 44675 158520
rect 44985 158440 44995 158520
rect 45305 158440 45315 158520
rect 45625 158440 45635 158520
rect 45945 158440 45955 158520
rect 46265 158440 46275 158520
rect 46585 158440 46595 158520
rect 46905 158440 46915 158520
rect 47225 158440 47235 158520
rect 47545 158440 47555 158520
rect 47865 158440 47875 158520
rect 48185 158440 48195 158520
rect 48500 158470 48605 158640
rect 48640 158560 48650 158640
rect 48790 158560 48800 158640
rect 49350 158560 49360 158640
rect 49500 158560 49510 158640
rect 49560 158470 49590 158640
rect 49650 158560 49690 158640
rect 48500 158460 48640 158470
rect 48710 158460 48790 158470
rect 49270 158460 49350 158470
rect 49420 158460 49500 158470
rect 49560 158460 49650 158470
rect 49660 158460 49690 158560
rect 43785 158360 43865 158370
rect 44105 158360 44185 158370
rect 44425 158360 44505 158370
rect 44745 158360 44825 158370
rect 45065 158360 45145 158370
rect 45385 158360 45465 158370
rect 45705 158360 45785 158370
rect 46025 158360 46105 158370
rect 46345 158360 46425 158370
rect 46665 158360 46745 158370
rect 46985 158360 47065 158370
rect 47305 158360 47385 158370
rect 47625 158360 47705 158370
rect 47945 158360 48025 158370
rect 48265 158360 48345 158370
rect 42950 158300 42980 158310
rect 43220 158300 43300 158310
rect 42980 158220 42990 158300
rect 43300 158220 43310 158300
rect 43865 158280 43875 158360
rect 44185 158280 44195 158360
rect 44505 158280 44515 158360
rect 44825 158280 44835 158360
rect 45145 158280 45155 158360
rect 45465 158280 45475 158360
rect 45785 158280 45795 158360
rect 46105 158280 46115 158360
rect 46425 158280 46435 158360
rect 46745 158280 46755 158360
rect 47065 158280 47075 158360
rect 47385 158280 47395 158360
rect 47705 158280 47715 158360
rect 48025 158280 48035 158360
rect 48345 158280 48355 158360
rect 48500 158290 48605 158460
rect 48640 158380 48650 158460
rect 48790 158380 48800 158460
rect 49350 158380 49360 158460
rect 49500 158380 49510 158460
rect 49560 158290 49590 158460
rect 49650 158380 49690 158460
rect 48500 158280 48640 158290
rect 48710 158280 48790 158290
rect 49270 158280 49350 158290
rect 49420 158280 49500 158290
rect 49560 158280 49650 158290
rect 49660 158280 49690 158380
rect 43945 158200 44025 158210
rect 44265 158200 44345 158210
rect 44585 158200 44665 158210
rect 44905 158200 44985 158210
rect 45225 158200 45305 158210
rect 45545 158200 45625 158210
rect 45865 158200 45945 158210
rect 46185 158200 46265 158210
rect 46505 158200 46585 158210
rect 46825 158200 46905 158210
rect 47145 158200 47225 158210
rect 47465 158200 47545 158210
rect 47785 158200 47865 158210
rect 48105 158200 48185 158210
rect 43060 158140 43140 158150
rect 43380 158140 43460 158150
rect 43140 158060 43150 158140
rect 43460 158060 43470 158140
rect 44025 158120 44035 158200
rect 44345 158120 44355 158200
rect 44665 158120 44675 158200
rect 44985 158120 44995 158200
rect 45305 158120 45315 158200
rect 45625 158120 45635 158200
rect 45945 158120 45955 158200
rect 46265 158120 46275 158200
rect 46585 158120 46595 158200
rect 46905 158120 46915 158200
rect 47225 158120 47235 158200
rect 47545 158120 47555 158200
rect 47865 158120 47875 158200
rect 48185 158120 48195 158200
rect 48500 158110 48605 158280
rect 48640 158200 48650 158280
rect 48790 158200 48800 158280
rect 49350 158200 49360 158280
rect 49500 158200 49510 158280
rect 49560 158110 49590 158280
rect 49650 158200 49690 158280
rect 48500 158100 48640 158110
rect 48710 158100 48790 158110
rect 49270 158100 49350 158110
rect 49420 158100 49500 158110
rect 49560 158100 49650 158110
rect 49660 158100 49690 158200
rect 43785 158040 43865 158050
rect 44105 158040 44185 158050
rect 44425 158040 44505 158050
rect 44745 158040 44825 158050
rect 45065 158040 45145 158050
rect 45385 158040 45465 158050
rect 45705 158040 45785 158050
rect 46025 158040 46105 158050
rect 46345 158040 46425 158050
rect 46665 158040 46745 158050
rect 46985 158040 47065 158050
rect 47305 158040 47385 158050
rect 47625 158040 47705 158050
rect 47945 158040 48025 158050
rect 48265 158040 48345 158050
rect 42950 157980 42980 157990
rect 43220 157980 43300 157990
rect 42980 157900 42990 157980
rect 43300 157900 43310 157980
rect 43865 157960 43875 158040
rect 44185 157960 44195 158040
rect 44505 157960 44515 158040
rect 44825 157960 44835 158040
rect 45145 157960 45155 158040
rect 45465 157960 45475 158040
rect 45785 157960 45795 158040
rect 46105 157960 46115 158040
rect 46425 157960 46435 158040
rect 46745 157960 46755 158040
rect 47065 157960 47075 158040
rect 47385 157960 47395 158040
rect 47705 157960 47715 158040
rect 48025 157960 48035 158040
rect 48345 157960 48355 158040
rect 48500 157930 48605 158100
rect 48640 158020 48650 158100
rect 48790 158020 48800 158100
rect 49350 158020 49360 158100
rect 49500 158020 49510 158100
rect 49560 157930 49590 158100
rect 49650 158020 49690 158100
rect 48500 157920 48640 157930
rect 48710 157920 48790 157930
rect 49270 157920 49350 157930
rect 49420 157920 49500 157930
rect 49560 157920 49650 157930
rect 49660 157920 49690 158020
rect 43945 157880 44025 157890
rect 44265 157880 44345 157890
rect 44585 157880 44665 157890
rect 44905 157880 44985 157890
rect 45225 157880 45305 157890
rect 45545 157880 45625 157890
rect 45865 157880 45945 157890
rect 46185 157880 46265 157890
rect 46505 157880 46585 157890
rect 46825 157880 46905 157890
rect 47145 157880 47225 157890
rect 47465 157880 47545 157890
rect 47785 157880 47865 157890
rect 48105 157880 48185 157890
rect 43060 157820 43140 157830
rect 43380 157820 43460 157830
rect 43140 157740 43150 157820
rect 43460 157740 43470 157820
rect 44025 157800 44035 157880
rect 44345 157800 44355 157880
rect 44665 157800 44675 157880
rect 44985 157800 44995 157880
rect 45305 157800 45315 157880
rect 45625 157800 45635 157880
rect 45945 157800 45955 157880
rect 46265 157800 46275 157880
rect 46585 157800 46595 157880
rect 46905 157800 46915 157880
rect 47225 157800 47235 157880
rect 47545 157800 47555 157880
rect 47865 157800 47875 157880
rect 48185 157800 48195 157880
rect 48500 157750 48605 157920
rect 48640 157840 48650 157920
rect 48790 157840 48800 157920
rect 49350 157840 49360 157920
rect 49500 157840 49510 157920
rect 49560 157750 49590 157920
rect 49650 157840 49690 157920
rect 48500 157740 48640 157750
rect 48710 157740 48790 157750
rect 49270 157740 49350 157750
rect 49420 157740 49500 157750
rect 49560 157740 49650 157750
rect 49660 157740 49690 157840
rect 43785 157720 43865 157730
rect 44105 157720 44185 157730
rect 44425 157720 44505 157730
rect 44745 157720 44825 157730
rect 45065 157720 45145 157730
rect 45385 157720 45465 157730
rect 45705 157720 45785 157730
rect 46025 157720 46105 157730
rect 46345 157720 46425 157730
rect 46665 157720 46745 157730
rect 46985 157720 47065 157730
rect 47305 157720 47385 157730
rect 47625 157720 47705 157730
rect 47945 157720 48025 157730
rect 48265 157720 48345 157730
rect 42950 157660 42980 157670
rect 43220 157660 43300 157670
rect 42980 157580 42990 157660
rect 43300 157580 43310 157660
rect 43865 157640 43875 157720
rect 44185 157640 44195 157720
rect 44505 157640 44515 157720
rect 44825 157640 44835 157720
rect 45145 157640 45155 157720
rect 45465 157640 45475 157720
rect 45785 157640 45795 157720
rect 46105 157640 46115 157720
rect 46425 157640 46435 157720
rect 46745 157640 46755 157720
rect 47065 157640 47075 157720
rect 47385 157640 47395 157720
rect 47705 157640 47715 157720
rect 48025 157640 48035 157720
rect 48345 157640 48355 157720
rect 48500 157570 48605 157740
rect 48640 157660 48650 157740
rect 48790 157660 48800 157740
rect 49350 157660 49360 157740
rect 49500 157660 49510 157740
rect 49560 157570 49590 157740
rect 49650 157660 49690 157740
rect 43945 157560 44025 157570
rect 44265 157560 44345 157570
rect 44585 157560 44665 157570
rect 44905 157560 44985 157570
rect 45225 157560 45305 157570
rect 45545 157560 45625 157570
rect 45865 157560 45945 157570
rect 46185 157560 46265 157570
rect 46505 157560 46585 157570
rect 46825 157560 46905 157570
rect 47145 157560 47225 157570
rect 47465 157560 47545 157570
rect 47785 157560 47865 157570
rect 48105 157560 48185 157570
rect 48500 157560 48640 157570
rect 48710 157560 48790 157570
rect 49270 157560 49350 157570
rect 49420 157560 49500 157570
rect 49560 157560 49650 157570
rect 49660 157560 49690 157660
rect 43060 157500 43140 157510
rect 43380 157500 43460 157510
rect 43140 157420 43150 157500
rect 43460 157420 43470 157500
rect 44025 157480 44035 157560
rect 44345 157480 44355 157560
rect 44665 157480 44675 157560
rect 44985 157480 44995 157560
rect 45305 157480 45315 157560
rect 45625 157480 45635 157560
rect 45945 157480 45955 157560
rect 46265 157480 46275 157560
rect 46585 157480 46595 157560
rect 46905 157480 46915 157560
rect 47225 157480 47235 157560
rect 47545 157480 47555 157560
rect 47865 157480 47875 157560
rect 48185 157480 48195 157560
rect 43785 157400 43865 157410
rect 44105 157400 44185 157410
rect 44425 157400 44505 157410
rect 44745 157400 44825 157410
rect 45065 157400 45145 157410
rect 45385 157400 45465 157410
rect 45705 157400 45785 157410
rect 46025 157400 46105 157410
rect 46345 157400 46425 157410
rect 46665 157400 46745 157410
rect 46985 157400 47065 157410
rect 47305 157400 47385 157410
rect 47625 157400 47705 157410
rect 47945 157400 48025 157410
rect 48265 157400 48345 157410
rect 42950 157340 42980 157350
rect 43220 157340 43300 157350
rect 42980 157260 42990 157340
rect 43300 157260 43310 157340
rect 43865 157320 43875 157400
rect 44185 157320 44195 157400
rect 44505 157320 44515 157400
rect 44825 157320 44835 157400
rect 45145 157320 45155 157400
rect 45465 157320 45475 157400
rect 45785 157320 45795 157400
rect 46105 157320 46115 157400
rect 46425 157320 46435 157400
rect 46745 157320 46755 157400
rect 47065 157320 47075 157400
rect 47385 157320 47395 157400
rect 47705 157320 47715 157400
rect 48025 157320 48035 157400
rect 48345 157320 48355 157400
rect 48500 157390 48605 157560
rect 48640 157480 48650 157560
rect 48790 157480 48800 157560
rect 49350 157480 49360 157560
rect 49500 157480 49510 157560
rect 49560 157390 49590 157560
rect 49650 157480 49690 157560
rect 48500 157380 48640 157390
rect 48710 157380 48790 157390
rect 49270 157380 49350 157390
rect 49420 157380 49500 157390
rect 49560 157380 49650 157390
rect 49660 157380 49690 157480
rect 43945 157240 44025 157250
rect 44265 157240 44345 157250
rect 44585 157240 44665 157250
rect 44905 157240 44985 157250
rect 45225 157240 45305 157250
rect 45545 157240 45625 157250
rect 45865 157240 45945 157250
rect 46185 157240 46265 157250
rect 46505 157240 46585 157250
rect 46825 157240 46905 157250
rect 47145 157240 47225 157250
rect 47465 157240 47545 157250
rect 47785 157240 47865 157250
rect 48105 157240 48185 157250
rect 43060 157180 43140 157190
rect 43380 157180 43460 157190
rect 43140 157100 43150 157180
rect 43460 157100 43470 157180
rect 44025 157160 44035 157240
rect 44345 157160 44355 157240
rect 44665 157160 44675 157240
rect 44985 157160 44995 157240
rect 45305 157160 45315 157240
rect 45625 157160 45635 157240
rect 45945 157160 45955 157240
rect 46265 157160 46275 157240
rect 46585 157160 46595 157240
rect 46905 157160 46915 157240
rect 47225 157160 47235 157240
rect 47545 157160 47555 157240
rect 47865 157160 47875 157240
rect 48185 157160 48195 157240
rect 48500 157210 48605 157380
rect 48640 157300 48650 157380
rect 48790 157300 48800 157380
rect 49350 157300 49360 157380
rect 49500 157300 49510 157380
rect 49560 157210 49590 157380
rect 49650 157300 49690 157380
rect 48500 157200 48640 157210
rect 48710 157200 48790 157210
rect 49270 157200 49350 157210
rect 49420 157200 49500 157210
rect 49560 157200 49650 157210
rect 49660 157200 49690 157300
rect 43785 157080 43865 157090
rect 44105 157080 44185 157090
rect 44425 157080 44505 157090
rect 44745 157080 44825 157090
rect 45065 157080 45145 157090
rect 45385 157080 45465 157090
rect 45705 157080 45785 157090
rect 46025 157080 46105 157090
rect 46345 157080 46425 157090
rect 46665 157080 46745 157090
rect 46985 157080 47065 157090
rect 47305 157080 47385 157090
rect 47625 157080 47705 157090
rect 47945 157080 48025 157090
rect 48265 157080 48345 157090
rect 42950 157020 42980 157030
rect 43220 157020 43300 157030
rect 42980 156940 42990 157020
rect 43300 156940 43310 157020
rect 43865 157000 43875 157080
rect 44185 157000 44195 157080
rect 44505 157000 44515 157080
rect 44825 157000 44835 157080
rect 45145 157000 45155 157080
rect 45465 157000 45475 157080
rect 45785 157000 45795 157080
rect 46105 157000 46115 157080
rect 46425 157000 46435 157080
rect 46745 157000 46755 157080
rect 47065 157000 47075 157080
rect 47385 157000 47395 157080
rect 47705 157000 47715 157080
rect 48025 157000 48035 157080
rect 48345 157000 48355 157080
rect 48500 157030 48605 157200
rect 48640 157120 48650 157200
rect 48790 157120 48800 157200
rect 49350 157120 49360 157200
rect 49500 157120 49510 157200
rect 49560 157030 49590 157200
rect 49650 157120 49690 157200
rect 48500 157020 48640 157030
rect 48710 157020 48790 157030
rect 49270 157020 49350 157030
rect 49420 157020 49500 157030
rect 49560 157020 49650 157030
rect 49660 157020 49690 157120
rect 43945 156920 44025 156930
rect 44265 156920 44345 156930
rect 44585 156920 44665 156930
rect 44905 156920 44985 156930
rect 45225 156920 45305 156930
rect 45545 156920 45625 156930
rect 45865 156920 45945 156930
rect 46185 156920 46265 156930
rect 46505 156920 46585 156930
rect 46825 156920 46905 156930
rect 47145 156920 47225 156930
rect 47465 156920 47545 156930
rect 47785 156920 47865 156930
rect 48105 156920 48185 156930
rect 43060 156860 43140 156870
rect 43380 156860 43460 156870
rect 43140 156780 43150 156860
rect 43460 156780 43470 156860
rect 44025 156840 44035 156920
rect 44345 156840 44355 156920
rect 44665 156840 44675 156920
rect 44985 156840 44995 156920
rect 45305 156840 45315 156920
rect 45625 156840 45635 156920
rect 45945 156840 45955 156920
rect 46265 156840 46275 156920
rect 46585 156840 46595 156920
rect 46905 156840 46915 156920
rect 47225 156840 47235 156920
rect 47545 156840 47555 156920
rect 47865 156840 47875 156920
rect 48185 156840 48195 156920
rect 48500 156850 48605 157020
rect 48640 156940 48650 157020
rect 48790 156940 48800 157020
rect 49350 156940 49360 157020
rect 49500 156940 49510 157020
rect 49560 156850 49590 157020
rect 49650 156940 49690 157020
rect 48500 156840 48640 156850
rect 48710 156840 48790 156850
rect 49270 156840 49350 156850
rect 49420 156840 49500 156850
rect 49560 156840 49650 156850
rect 49660 156840 49690 156940
rect 43785 156760 43865 156770
rect 44105 156760 44185 156770
rect 44425 156760 44505 156770
rect 44745 156760 44825 156770
rect 45065 156760 45145 156770
rect 45385 156760 45465 156770
rect 45705 156760 45785 156770
rect 46025 156760 46105 156770
rect 46345 156760 46425 156770
rect 46665 156760 46745 156770
rect 46985 156760 47065 156770
rect 47305 156760 47385 156770
rect 47625 156760 47705 156770
rect 47945 156760 48025 156770
rect 48265 156760 48345 156770
rect 42950 156700 42980 156710
rect 43220 156700 43300 156710
rect 42980 156620 42990 156700
rect 43300 156620 43310 156700
rect 43865 156680 43875 156760
rect 44185 156680 44195 156760
rect 44505 156680 44515 156760
rect 44825 156680 44835 156760
rect 45145 156680 45155 156760
rect 45465 156680 45475 156760
rect 45785 156680 45795 156760
rect 46105 156680 46115 156760
rect 46425 156680 46435 156760
rect 46745 156680 46755 156760
rect 47065 156680 47075 156760
rect 47385 156680 47395 156760
rect 47705 156680 47715 156760
rect 48025 156680 48035 156760
rect 48345 156680 48355 156760
rect 48500 156670 48605 156840
rect 48640 156760 48650 156840
rect 48790 156760 48800 156840
rect 49350 156760 49360 156840
rect 49500 156760 49510 156840
rect 49560 156670 49590 156840
rect 49650 156760 49690 156840
rect 48500 156660 48640 156670
rect 48710 156660 48790 156670
rect 49270 156660 49350 156670
rect 49420 156660 49500 156670
rect 49560 156660 49650 156670
rect 49660 156660 49690 156760
rect 43945 156600 44025 156610
rect 44265 156600 44345 156610
rect 44585 156600 44665 156610
rect 44905 156600 44985 156610
rect 45225 156600 45305 156610
rect 45545 156600 45625 156610
rect 45865 156600 45945 156610
rect 46185 156600 46265 156610
rect 46505 156600 46585 156610
rect 46825 156600 46905 156610
rect 47145 156600 47225 156610
rect 47465 156600 47545 156610
rect 47785 156600 47865 156610
rect 48105 156600 48185 156610
rect 43060 156540 43140 156550
rect 43380 156540 43460 156550
rect 43140 156460 43150 156540
rect 43460 156460 43470 156540
rect 44025 156520 44035 156600
rect 44345 156520 44355 156600
rect 44665 156520 44675 156600
rect 44985 156520 44995 156600
rect 45305 156520 45315 156600
rect 45625 156520 45635 156600
rect 45945 156520 45955 156600
rect 46265 156520 46275 156600
rect 46585 156520 46595 156600
rect 46905 156520 46915 156600
rect 47225 156520 47235 156600
rect 47545 156520 47555 156600
rect 47865 156520 47875 156600
rect 48185 156520 48195 156600
rect 48500 156490 48605 156660
rect 48640 156580 48650 156660
rect 48790 156580 48800 156660
rect 49350 156580 49360 156660
rect 49500 156580 49510 156660
rect 49560 156490 49590 156660
rect 49650 156580 49690 156660
rect 48500 156480 48640 156490
rect 48710 156480 48790 156490
rect 49270 156480 49350 156490
rect 49420 156480 49500 156490
rect 49560 156480 49650 156490
rect 49660 156480 49690 156580
rect 43785 156440 43865 156450
rect 44105 156440 44185 156450
rect 44425 156440 44505 156450
rect 44745 156440 44825 156450
rect 45065 156440 45145 156450
rect 45385 156440 45465 156450
rect 45705 156440 45785 156450
rect 46025 156440 46105 156450
rect 46345 156440 46425 156450
rect 46665 156440 46745 156450
rect 46985 156440 47065 156450
rect 47305 156440 47385 156450
rect 47625 156440 47705 156450
rect 47945 156440 48025 156450
rect 48265 156440 48345 156450
rect 42950 156380 42980 156390
rect 43220 156380 43300 156390
rect 42980 156300 42990 156380
rect 43300 156300 43310 156380
rect 43865 156360 43875 156440
rect 44185 156360 44195 156440
rect 44505 156360 44515 156440
rect 44825 156360 44835 156440
rect 45145 156360 45155 156440
rect 45465 156360 45475 156440
rect 45785 156360 45795 156440
rect 46105 156360 46115 156440
rect 46425 156360 46435 156440
rect 46745 156360 46755 156440
rect 47065 156360 47075 156440
rect 47385 156360 47395 156440
rect 47705 156360 47715 156440
rect 48025 156360 48035 156440
rect 48345 156360 48355 156440
rect 48500 156310 48605 156480
rect 48640 156400 48650 156480
rect 48790 156400 48800 156480
rect 49350 156400 49360 156480
rect 49500 156400 49510 156480
rect 49560 156310 49590 156480
rect 49650 156400 49690 156480
rect 48500 156300 48640 156310
rect 48710 156300 48790 156310
rect 49270 156300 49350 156310
rect 49420 156300 49500 156310
rect 49560 156300 49650 156310
rect 49660 156300 49690 156400
rect 43945 156280 44025 156290
rect 44265 156280 44345 156290
rect 44585 156280 44665 156290
rect 44905 156280 44985 156290
rect 45225 156280 45305 156290
rect 45545 156280 45625 156290
rect 45865 156280 45945 156290
rect 46185 156280 46265 156290
rect 46505 156280 46585 156290
rect 46825 156280 46905 156290
rect 47145 156280 47225 156290
rect 47465 156280 47545 156290
rect 47785 156280 47865 156290
rect 48105 156280 48185 156290
rect 43060 156220 43140 156230
rect 43380 156220 43460 156230
rect 43140 156140 43150 156220
rect 43460 156140 43470 156220
rect 44025 156200 44035 156280
rect 44345 156200 44355 156280
rect 44665 156200 44675 156280
rect 44985 156200 44995 156280
rect 45305 156200 45315 156280
rect 45625 156200 45635 156280
rect 45945 156200 45955 156280
rect 46265 156200 46275 156280
rect 46585 156200 46595 156280
rect 46905 156200 46915 156280
rect 47225 156200 47235 156280
rect 47545 156200 47555 156280
rect 47865 156200 47875 156280
rect 48185 156200 48195 156280
rect 48500 156130 48605 156300
rect 48640 156220 48650 156300
rect 48790 156220 48800 156300
rect 49350 156220 49360 156300
rect 49500 156220 49510 156300
rect 49560 156130 49590 156300
rect 49650 156220 49690 156300
rect 43785 156120 43865 156130
rect 44105 156120 44185 156130
rect 44425 156120 44505 156130
rect 44745 156120 44825 156130
rect 45065 156120 45145 156130
rect 45385 156120 45465 156130
rect 45705 156120 45785 156130
rect 46025 156120 46105 156130
rect 46345 156120 46425 156130
rect 46665 156120 46745 156130
rect 46985 156120 47065 156130
rect 47305 156120 47385 156130
rect 47625 156120 47705 156130
rect 47945 156120 48025 156130
rect 48265 156120 48345 156130
rect 48500 156120 48640 156130
rect 48710 156120 48790 156130
rect 49270 156120 49350 156130
rect 49420 156120 49500 156130
rect 49560 156120 49650 156130
rect 49660 156120 49690 156220
rect 42950 156060 42980 156070
rect 43220 156060 43300 156070
rect 36260 155980 36270 156000
rect 36580 155980 36590 156000
rect 36900 155980 36910 156000
rect 37220 155980 37230 156000
rect 37540 155980 37550 156000
rect 37860 155980 37870 156000
rect 38180 155980 38190 156000
rect 38500 155980 38510 156000
rect 38820 155980 38830 156000
rect 39140 155980 39150 156000
rect 39460 155980 39470 156000
rect 39780 155980 39790 156000
rect 40100 155980 40110 156000
rect 40420 155980 40430 156000
rect 40740 155980 40750 156000
rect 41060 155980 41070 156000
rect 41380 155980 41390 156000
rect 41700 155980 41710 156000
rect 42020 155980 42030 156000
rect 42340 155980 42350 156000
rect 42660 155980 42670 156000
rect 42980 155980 42990 156060
rect 43300 155980 43310 156060
rect 43865 156040 43875 156120
rect 44185 156040 44195 156120
rect 44505 156040 44515 156120
rect 44825 156040 44835 156120
rect 45145 156040 45155 156120
rect 45465 156040 45475 156120
rect 45785 156040 45795 156120
rect 46105 156040 46115 156120
rect 46425 156040 46435 156120
rect 46745 156040 46755 156120
rect 47065 156040 47075 156120
rect 47385 156040 47395 156120
rect 47705 156040 47715 156120
rect 48025 156040 48035 156120
rect 48345 156040 48355 156120
rect 43945 155960 44025 155970
rect 44265 155960 44345 155970
rect 44585 155960 44665 155970
rect 44905 155960 44985 155970
rect 45225 155960 45305 155970
rect 45545 155960 45625 155970
rect 45865 155960 45945 155970
rect 46185 155960 46265 155970
rect 46505 155960 46585 155970
rect 46825 155960 46905 155970
rect 47145 155960 47225 155970
rect 47465 155960 47545 155970
rect 47785 155960 47865 155970
rect 48105 155960 48185 155970
rect 36020 155900 36100 155910
rect 36340 155900 36420 155910
rect 36660 155900 36740 155910
rect 36980 155900 37060 155910
rect 37300 155900 37380 155910
rect 37620 155900 37700 155910
rect 37940 155900 38020 155910
rect 38260 155900 38340 155910
rect 38580 155900 38660 155910
rect 38900 155900 38980 155910
rect 39220 155900 39300 155910
rect 39540 155900 39620 155910
rect 39860 155900 39940 155910
rect 40180 155900 40260 155910
rect 40500 155900 40580 155910
rect 40820 155900 40900 155910
rect 41140 155900 41220 155910
rect 41460 155900 41540 155910
rect 41780 155900 41860 155910
rect 42100 155900 42180 155910
rect 42420 155900 42500 155910
rect 42740 155900 42820 155910
rect 43060 155900 43140 155910
rect 43380 155900 43460 155910
rect 36100 155820 36110 155900
rect 36420 155820 36430 155900
rect 36740 155820 36750 155900
rect 37060 155820 37070 155900
rect 37380 155820 37390 155900
rect 37700 155820 37710 155900
rect 38020 155820 38030 155900
rect 38340 155820 38350 155900
rect 38660 155820 38670 155900
rect 38980 155820 38990 155900
rect 39300 155820 39310 155900
rect 39620 155820 39630 155900
rect 39940 155820 39950 155900
rect 40260 155820 40270 155900
rect 40580 155820 40590 155900
rect 40900 155820 40910 155900
rect 41220 155820 41230 155900
rect 41540 155820 41550 155900
rect 41860 155820 41870 155900
rect 42180 155820 42190 155900
rect 42500 155820 42510 155900
rect 42820 155820 42830 155900
rect 43140 155820 43150 155900
rect 43460 155820 43470 155900
rect 44025 155880 44035 155960
rect 44345 155880 44355 155960
rect 44665 155880 44675 155960
rect 44985 155880 44995 155960
rect 45305 155880 45315 155960
rect 45625 155880 45635 155960
rect 45945 155880 45955 155960
rect 46265 155880 46275 155960
rect 46585 155880 46595 155960
rect 46905 155880 46915 155960
rect 47225 155880 47235 155960
rect 47545 155880 47555 155960
rect 47865 155880 47875 155960
rect 48185 155880 48195 155960
rect 48500 155950 48605 156120
rect 48640 156040 48650 156120
rect 48790 156040 48800 156120
rect 49350 156040 49360 156120
rect 49500 156040 49510 156120
rect 49560 155950 49590 156120
rect 49650 156040 49690 156120
rect 48500 155940 48640 155950
rect 48710 155940 48790 155950
rect 49270 155940 49350 155950
rect 49420 155940 49500 155950
rect 49560 155940 49650 155950
rect 49660 155940 49690 156040
rect 43785 155800 43865 155810
rect 44105 155800 44185 155810
rect 44425 155800 44505 155810
rect 44745 155800 44825 155810
rect 45065 155800 45145 155810
rect 45385 155800 45465 155810
rect 45705 155800 45785 155810
rect 46025 155800 46105 155810
rect 46345 155800 46425 155810
rect 46665 155800 46745 155810
rect 46985 155800 47065 155810
rect 47305 155800 47385 155810
rect 47625 155800 47705 155810
rect 47945 155800 48025 155810
rect 48265 155800 48345 155810
rect 36180 155740 36260 155750
rect 36500 155740 36580 155750
rect 36820 155740 36900 155750
rect 37140 155740 37220 155750
rect 37460 155740 37540 155750
rect 37780 155740 37860 155750
rect 38100 155740 38180 155750
rect 38420 155740 38500 155750
rect 38740 155740 38820 155750
rect 39060 155740 39140 155750
rect 39380 155740 39460 155750
rect 39700 155740 39780 155750
rect 40020 155740 40100 155750
rect 40340 155740 40420 155750
rect 40660 155740 40740 155750
rect 40980 155740 41060 155750
rect 41300 155740 41380 155750
rect 41620 155740 41700 155750
rect 41940 155740 42020 155750
rect 42260 155740 42340 155750
rect 42580 155740 42660 155750
rect 42900 155740 42980 155750
rect 43220 155740 43300 155750
rect 36260 155660 36270 155740
rect 36580 155660 36590 155740
rect 36900 155660 36910 155740
rect 37220 155660 37230 155740
rect 37540 155660 37550 155740
rect 37860 155660 37870 155740
rect 38180 155660 38190 155740
rect 38500 155660 38510 155740
rect 38820 155660 38830 155740
rect 39140 155660 39150 155740
rect 39460 155660 39470 155740
rect 39780 155660 39790 155740
rect 40100 155660 40110 155740
rect 40420 155660 40430 155740
rect 40740 155660 40750 155740
rect 41060 155660 41070 155740
rect 41380 155660 41390 155740
rect 41700 155660 41710 155740
rect 42020 155660 42030 155740
rect 42340 155660 42350 155740
rect 42660 155660 42670 155740
rect 42980 155660 42990 155740
rect 43300 155660 43310 155740
rect 43865 155720 43875 155800
rect 44185 155720 44195 155800
rect 44505 155720 44515 155800
rect 44825 155720 44835 155800
rect 45145 155720 45155 155800
rect 45465 155720 45475 155800
rect 45785 155720 45795 155800
rect 46105 155720 46115 155800
rect 46425 155720 46435 155800
rect 46745 155720 46755 155800
rect 47065 155720 47075 155800
rect 47385 155720 47395 155800
rect 47705 155720 47715 155800
rect 48025 155720 48035 155800
rect 48345 155720 48355 155800
rect 48500 155770 48605 155940
rect 48640 155860 48650 155940
rect 48790 155860 48800 155940
rect 49350 155860 49360 155940
rect 49500 155860 49510 155940
rect 49560 155770 49590 155940
rect 49650 155860 49690 155940
rect 48500 155760 48640 155770
rect 48710 155760 48790 155770
rect 49270 155760 49350 155770
rect 49420 155760 49500 155770
rect 49560 155760 49650 155770
rect 49660 155760 49690 155860
rect 43945 155640 44025 155650
rect 44265 155640 44345 155650
rect 44585 155640 44665 155650
rect 44905 155640 44985 155650
rect 45225 155640 45305 155650
rect 45545 155640 45625 155650
rect 45865 155640 45945 155650
rect 46185 155640 46265 155650
rect 46505 155640 46585 155650
rect 46825 155640 46905 155650
rect 47145 155640 47225 155650
rect 47465 155640 47545 155650
rect 47785 155640 47865 155650
rect 48105 155640 48185 155650
rect 36020 155580 36100 155590
rect 36340 155580 36420 155590
rect 36660 155580 36740 155590
rect 36980 155580 37060 155590
rect 37300 155580 37380 155590
rect 37620 155580 37700 155590
rect 37940 155580 38020 155590
rect 38260 155580 38340 155590
rect 38580 155580 38660 155590
rect 38900 155580 38980 155590
rect 39220 155580 39300 155590
rect 39540 155580 39620 155590
rect 39860 155580 39940 155590
rect 40180 155580 40260 155590
rect 40500 155580 40580 155590
rect 40820 155580 40900 155590
rect 41140 155580 41220 155590
rect 41460 155580 41540 155590
rect 41780 155580 41860 155590
rect 42100 155580 42180 155590
rect 42420 155580 42500 155590
rect 42740 155580 42820 155590
rect 43060 155580 43140 155590
rect 43380 155580 43460 155590
rect 36100 155500 36110 155580
rect 36420 155500 36430 155580
rect 36740 155500 36750 155580
rect 37060 155500 37070 155580
rect 37380 155500 37390 155580
rect 37700 155500 37710 155580
rect 38020 155500 38030 155580
rect 38340 155500 38350 155580
rect 38660 155500 38670 155580
rect 38980 155500 38990 155580
rect 39300 155500 39310 155580
rect 39620 155500 39630 155580
rect 39940 155500 39950 155580
rect 40260 155500 40270 155580
rect 40580 155500 40590 155580
rect 40900 155500 40910 155580
rect 41220 155500 41230 155580
rect 41540 155500 41550 155580
rect 41860 155500 41870 155580
rect 42180 155500 42190 155580
rect 42500 155500 42510 155580
rect 42820 155500 42830 155580
rect 43140 155500 43150 155580
rect 43460 155500 43470 155580
rect 44025 155560 44035 155640
rect 44345 155560 44355 155640
rect 44665 155560 44675 155640
rect 44985 155560 44995 155640
rect 45305 155560 45315 155640
rect 45625 155560 45635 155640
rect 45945 155560 45955 155640
rect 46265 155560 46275 155640
rect 46585 155560 46595 155640
rect 46905 155560 46915 155640
rect 47225 155560 47235 155640
rect 47545 155560 47555 155640
rect 47865 155560 47875 155640
rect 48185 155560 48195 155640
rect 48500 155590 48605 155760
rect 48640 155680 48650 155760
rect 48790 155680 48800 155760
rect 49350 155680 49360 155760
rect 49500 155680 49510 155760
rect 49560 155590 49590 155760
rect 49650 155680 49690 155760
rect 48500 155580 48640 155590
rect 48710 155580 48790 155590
rect 49270 155580 49350 155590
rect 49420 155580 49500 155590
rect 49560 155580 49650 155590
rect 49660 155580 49690 155680
rect 43785 155480 43865 155490
rect 44105 155480 44185 155490
rect 44425 155480 44505 155490
rect 44745 155480 44825 155490
rect 45065 155480 45145 155490
rect 45385 155480 45465 155490
rect 45705 155480 45785 155490
rect 46025 155480 46105 155490
rect 46345 155480 46425 155490
rect 46665 155480 46745 155490
rect 46985 155480 47065 155490
rect 47305 155480 47385 155490
rect 47625 155480 47705 155490
rect 47945 155480 48025 155490
rect 48265 155480 48345 155490
rect 36180 155420 36260 155430
rect 36500 155420 36580 155430
rect 36820 155420 36900 155430
rect 37140 155420 37220 155430
rect 37460 155420 37540 155430
rect 37780 155420 37860 155430
rect 38100 155420 38180 155430
rect 38420 155420 38500 155430
rect 38740 155420 38820 155430
rect 39060 155420 39140 155430
rect 39380 155420 39460 155430
rect 39700 155420 39780 155430
rect 40020 155420 40100 155430
rect 40340 155420 40420 155430
rect 40660 155420 40740 155430
rect 40980 155420 41060 155430
rect 41300 155420 41380 155430
rect 41620 155420 41700 155430
rect 41940 155420 42020 155430
rect 42260 155420 42340 155430
rect 42580 155420 42660 155430
rect 42900 155420 42980 155430
rect 43220 155420 43300 155430
rect 36260 155340 36270 155420
rect 36580 155340 36590 155420
rect 36900 155340 36910 155420
rect 37220 155340 37230 155420
rect 37540 155340 37550 155420
rect 37860 155340 37870 155420
rect 38180 155340 38190 155420
rect 38500 155340 38510 155420
rect 38820 155340 38830 155420
rect 39140 155340 39150 155420
rect 39460 155340 39470 155420
rect 39780 155340 39790 155420
rect 40100 155340 40110 155420
rect 40420 155340 40430 155420
rect 40740 155340 40750 155420
rect 41060 155340 41070 155420
rect 41380 155340 41390 155420
rect 41700 155340 41710 155420
rect 42020 155340 42030 155420
rect 42340 155340 42350 155420
rect 42660 155340 42670 155420
rect 42980 155340 42990 155420
rect 43300 155340 43310 155420
rect 43865 155400 43875 155480
rect 44185 155400 44195 155480
rect 44505 155400 44515 155480
rect 44825 155400 44835 155480
rect 45145 155400 45155 155480
rect 45465 155400 45475 155480
rect 45785 155400 45795 155480
rect 46105 155400 46115 155480
rect 46425 155400 46435 155480
rect 46745 155400 46755 155480
rect 47065 155400 47075 155480
rect 47385 155400 47395 155480
rect 47705 155400 47715 155480
rect 48025 155400 48035 155480
rect 48345 155400 48355 155480
rect 48500 155410 48605 155580
rect 48640 155500 48650 155580
rect 48790 155500 48800 155580
rect 49350 155500 49360 155580
rect 49500 155500 49510 155580
rect 49560 155410 49590 155580
rect 49650 155500 49690 155580
rect 48500 155400 48640 155410
rect 48710 155400 48790 155410
rect 49270 155400 49350 155410
rect 49420 155400 49500 155410
rect 49560 155400 49650 155410
rect 49660 155400 49690 155500
rect 43945 155320 44025 155330
rect 44265 155320 44345 155330
rect 44585 155320 44665 155330
rect 44905 155320 44985 155330
rect 45225 155320 45305 155330
rect 45545 155320 45625 155330
rect 45865 155320 45945 155330
rect 46185 155320 46265 155330
rect 46505 155320 46585 155330
rect 46825 155320 46905 155330
rect 47145 155320 47225 155330
rect 47465 155320 47545 155330
rect 47785 155320 47865 155330
rect 48105 155320 48185 155330
rect 36020 155260 36100 155270
rect 36340 155260 36420 155270
rect 36660 155260 36740 155270
rect 36980 155260 37060 155270
rect 37300 155260 37380 155270
rect 37620 155260 37700 155270
rect 37940 155260 38020 155270
rect 38260 155260 38340 155270
rect 38580 155260 38660 155270
rect 38900 155260 38980 155270
rect 39220 155260 39300 155270
rect 39540 155260 39620 155270
rect 39860 155260 39940 155270
rect 40180 155260 40260 155270
rect 40500 155260 40580 155270
rect 40820 155260 40900 155270
rect 41140 155260 41220 155270
rect 41460 155260 41540 155270
rect 41780 155260 41860 155270
rect 42100 155260 42180 155270
rect 42420 155260 42500 155270
rect 42740 155260 42820 155270
rect 43060 155260 43140 155270
rect 43380 155260 43460 155270
rect 36100 155180 36110 155260
rect 36420 155180 36430 155260
rect 36740 155180 36750 155260
rect 37060 155180 37070 155260
rect 37380 155180 37390 155260
rect 37700 155180 37710 155260
rect 38020 155180 38030 155260
rect 38340 155180 38350 155260
rect 38660 155180 38670 155260
rect 38980 155180 38990 155260
rect 39300 155180 39310 155260
rect 39620 155180 39630 155260
rect 39940 155180 39950 155260
rect 40260 155180 40270 155260
rect 40580 155180 40590 155260
rect 40900 155180 40910 155260
rect 41220 155180 41230 155260
rect 41540 155180 41550 155260
rect 41860 155180 41870 155260
rect 42180 155180 42190 155260
rect 42500 155180 42510 155260
rect 42820 155180 42830 155260
rect 43140 155180 43150 155260
rect 43460 155180 43470 155260
rect 44025 155240 44035 155320
rect 44345 155240 44355 155320
rect 44665 155240 44675 155320
rect 44985 155240 44995 155320
rect 45305 155240 45315 155320
rect 45625 155240 45635 155320
rect 45945 155240 45955 155320
rect 46265 155240 46275 155320
rect 46585 155240 46595 155320
rect 46905 155240 46915 155320
rect 47225 155240 47235 155320
rect 47545 155240 47555 155320
rect 47865 155240 47875 155320
rect 48185 155240 48195 155320
rect 48500 155230 48605 155400
rect 48640 155320 48650 155400
rect 48790 155320 48800 155400
rect 49350 155320 49360 155400
rect 49500 155320 49510 155400
rect 49560 155230 49590 155400
rect 49650 155320 49690 155400
rect 48500 155220 48640 155230
rect 48710 155220 48790 155230
rect 49270 155220 49350 155230
rect 49420 155220 49500 155230
rect 49560 155220 49650 155230
rect 49660 155220 49690 155320
rect 43785 155160 43865 155170
rect 44105 155160 44185 155170
rect 44425 155160 44505 155170
rect 44745 155160 44825 155170
rect 45065 155160 45145 155170
rect 45385 155160 45465 155170
rect 45705 155160 45785 155170
rect 46025 155160 46105 155170
rect 46345 155160 46425 155170
rect 46665 155160 46745 155170
rect 46985 155160 47065 155170
rect 47305 155160 47385 155170
rect 47625 155160 47705 155170
rect 47945 155160 48025 155170
rect 48265 155160 48345 155170
rect 36180 155100 36260 155110
rect 36500 155100 36580 155110
rect 36820 155100 36900 155110
rect 37140 155100 37220 155110
rect 37460 155100 37540 155110
rect 37780 155100 37860 155110
rect 38100 155100 38180 155110
rect 38420 155100 38500 155110
rect 38740 155100 38820 155110
rect 39060 155100 39140 155110
rect 39380 155100 39460 155110
rect 39700 155100 39780 155110
rect 40020 155100 40100 155110
rect 40340 155100 40420 155110
rect 40660 155100 40740 155110
rect 40980 155100 41060 155110
rect 41300 155100 41380 155110
rect 41620 155100 41700 155110
rect 41940 155100 42020 155110
rect 42260 155100 42340 155110
rect 42580 155100 42660 155110
rect 42900 155100 42980 155110
rect 43220 155100 43300 155110
rect 36260 155020 36270 155100
rect 36580 155020 36590 155100
rect 36900 155020 36910 155100
rect 37220 155020 37230 155100
rect 37540 155020 37550 155100
rect 37860 155020 37870 155100
rect 38180 155020 38190 155100
rect 38500 155020 38510 155100
rect 38820 155020 38830 155100
rect 39140 155020 39150 155100
rect 39460 155020 39470 155100
rect 39780 155020 39790 155100
rect 40100 155020 40110 155100
rect 40420 155020 40430 155100
rect 40740 155020 40750 155100
rect 41060 155020 41070 155100
rect 41380 155020 41390 155100
rect 41700 155020 41710 155100
rect 42020 155020 42030 155100
rect 42340 155020 42350 155100
rect 42660 155020 42670 155100
rect 42980 155020 42990 155100
rect 43300 155020 43310 155100
rect 43865 155080 43875 155160
rect 44185 155080 44195 155160
rect 44505 155080 44515 155160
rect 44825 155080 44835 155160
rect 45145 155080 45155 155160
rect 45465 155080 45475 155160
rect 45785 155080 45795 155160
rect 46105 155080 46115 155160
rect 46425 155080 46435 155160
rect 46745 155080 46755 155160
rect 47065 155080 47075 155160
rect 47385 155080 47395 155160
rect 47705 155080 47715 155160
rect 48025 155080 48035 155160
rect 48345 155080 48355 155160
rect 48500 155050 48605 155220
rect 48640 155140 48650 155220
rect 48790 155140 48800 155220
rect 49350 155140 49360 155220
rect 49500 155140 49510 155220
rect 49560 155050 49590 155220
rect 49650 155140 49690 155220
rect 48500 155040 48640 155050
rect 48710 155040 48790 155050
rect 49270 155040 49350 155050
rect 49420 155040 49500 155050
rect 49560 155040 49650 155050
rect 49660 155040 49690 155140
rect 43945 155000 44025 155010
rect 44265 155000 44345 155010
rect 44585 155000 44665 155010
rect 44905 155000 44985 155010
rect 45225 155000 45305 155010
rect 45545 155000 45625 155010
rect 45865 155000 45945 155010
rect 46185 155000 46265 155010
rect 46505 155000 46585 155010
rect 46825 155000 46905 155010
rect 47145 155000 47225 155010
rect 47465 155000 47545 155010
rect 47785 155000 47865 155010
rect 48105 155000 48185 155010
rect 36020 154940 36100 154950
rect 36340 154940 36420 154950
rect 36660 154940 36740 154950
rect 36980 154940 37060 154950
rect 37300 154940 37380 154950
rect 37620 154940 37700 154950
rect 37940 154940 38020 154950
rect 38260 154940 38340 154950
rect 38580 154940 38660 154950
rect 38900 154940 38980 154950
rect 39220 154940 39300 154950
rect 39540 154940 39620 154950
rect 39860 154940 39940 154950
rect 40180 154940 40260 154950
rect 40500 154940 40580 154950
rect 40820 154940 40900 154950
rect 41140 154940 41220 154950
rect 41460 154940 41540 154950
rect 41780 154940 41860 154950
rect 42100 154940 42180 154950
rect 42420 154940 42500 154950
rect 42740 154940 42820 154950
rect 43060 154940 43140 154950
rect 43380 154940 43460 154950
rect 36100 154860 36110 154940
rect 36420 154860 36430 154940
rect 36740 154860 36750 154940
rect 37060 154860 37070 154940
rect 37380 154860 37390 154940
rect 37700 154860 37710 154940
rect 38020 154860 38030 154940
rect 38340 154860 38350 154940
rect 38660 154860 38670 154940
rect 38980 154860 38990 154940
rect 39300 154860 39310 154940
rect 39620 154860 39630 154940
rect 39940 154860 39950 154940
rect 40260 154860 40270 154940
rect 40580 154860 40590 154940
rect 40900 154860 40910 154940
rect 41220 154860 41230 154940
rect 41540 154860 41550 154940
rect 41860 154860 41870 154940
rect 42180 154860 42190 154940
rect 42500 154860 42510 154940
rect 42820 154860 42830 154940
rect 43140 154860 43150 154940
rect 43460 154860 43470 154940
rect 44025 154920 44035 155000
rect 44345 154920 44355 155000
rect 44665 154920 44675 155000
rect 44985 154920 44995 155000
rect 45305 154920 45315 155000
rect 45625 154920 45635 155000
rect 45945 154920 45955 155000
rect 46265 154920 46275 155000
rect 46585 154920 46595 155000
rect 46905 154920 46915 155000
rect 47225 154920 47235 155000
rect 47545 154920 47555 155000
rect 47865 154920 47875 155000
rect 48185 154920 48195 155000
rect 48500 154870 48605 155040
rect 48640 154960 48650 155040
rect 48790 154960 48800 155040
rect 49350 154960 49360 155040
rect 49500 154960 49510 155040
rect 49560 154870 49590 155040
rect 49650 154960 49690 155040
rect 48500 154860 48640 154870
rect 48710 154860 48790 154870
rect 49270 154860 49350 154870
rect 49420 154860 49500 154870
rect 49560 154860 49650 154870
rect 49660 154860 49690 154960
rect 43785 154840 43865 154850
rect 44105 154840 44185 154850
rect 44425 154840 44505 154850
rect 44745 154840 44825 154850
rect 45065 154840 45145 154850
rect 45385 154840 45465 154850
rect 45705 154840 45785 154850
rect 46025 154840 46105 154850
rect 46345 154840 46425 154850
rect 46665 154840 46745 154850
rect 46985 154840 47065 154850
rect 47305 154840 47385 154850
rect 47625 154840 47705 154850
rect 47945 154840 48025 154850
rect 48265 154840 48345 154850
rect 36180 154780 36260 154790
rect 36500 154780 36580 154790
rect 36820 154780 36900 154790
rect 37140 154780 37220 154790
rect 37460 154780 37540 154790
rect 37780 154780 37860 154790
rect 38100 154780 38180 154790
rect 38420 154780 38500 154790
rect 38740 154780 38820 154790
rect 39060 154780 39140 154790
rect 39380 154780 39460 154790
rect 39700 154780 39780 154790
rect 40020 154780 40100 154790
rect 40340 154780 40420 154790
rect 40660 154780 40740 154790
rect 40980 154780 41060 154790
rect 41300 154780 41380 154790
rect 41620 154780 41700 154790
rect 41940 154780 42020 154790
rect 42260 154780 42340 154790
rect 42580 154780 42660 154790
rect 42900 154780 42980 154790
rect 43220 154780 43300 154790
rect 36260 154700 36270 154780
rect 36580 154700 36590 154780
rect 36900 154700 36910 154780
rect 37220 154700 37230 154780
rect 37540 154700 37550 154780
rect 37860 154700 37870 154780
rect 38180 154700 38190 154780
rect 38500 154700 38510 154780
rect 38820 154700 38830 154780
rect 39140 154700 39150 154780
rect 39460 154700 39470 154780
rect 39780 154700 39790 154780
rect 40100 154700 40110 154780
rect 40420 154700 40430 154780
rect 40740 154700 40750 154780
rect 41060 154700 41070 154780
rect 41380 154700 41390 154780
rect 41700 154700 41710 154780
rect 42020 154700 42030 154780
rect 42340 154700 42350 154780
rect 42660 154700 42670 154780
rect 42980 154700 42990 154780
rect 43300 154700 43310 154780
rect 43865 154760 43875 154840
rect 44185 154760 44195 154840
rect 44505 154760 44515 154840
rect 44825 154760 44835 154840
rect 45145 154760 45155 154840
rect 45465 154760 45475 154840
rect 45785 154760 45795 154840
rect 46105 154760 46115 154840
rect 46425 154760 46435 154840
rect 46745 154760 46755 154840
rect 47065 154760 47075 154840
rect 47385 154760 47395 154840
rect 47705 154760 47715 154840
rect 48025 154760 48035 154840
rect 48345 154760 48355 154840
rect 48500 154690 48605 154860
rect 48640 154780 48650 154860
rect 48790 154780 48800 154860
rect 49350 154780 49360 154860
rect 49500 154780 49510 154860
rect 49560 154690 49590 154860
rect 49650 154780 49690 154860
rect 43945 154680 44025 154690
rect 44265 154680 44345 154690
rect 44585 154680 44665 154690
rect 44905 154680 44985 154690
rect 45225 154680 45305 154690
rect 45545 154680 45625 154690
rect 45865 154680 45945 154690
rect 46185 154680 46265 154690
rect 46505 154680 46585 154690
rect 46825 154680 46905 154690
rect 47145 154680 47225 154690
rect 47465 154680 47545 154690
rect 47785 154680 47865 154690
rect 48105 154680 48185 154690
rect 48500 154680 48640 154690
rect 48710 154680 48790 154690
rect 49270 154680 49350 154690
rect 49420 154680 49500 154690
rect 49560 154680 49650 154690
rect 49660 154680 49690 154780
rect 36020 154620 36100 154630
rect 36340 154620 36420 154630
rect 36660 154620 36740 154630
rect 36980 154620 37060 154630
rect 37300 154620 37380 154630
rect 37620 154620 37700 154630
rect 37940 154620 38020 154630
rect 38260 154620 38340 154630
rect 38580 154620 38660 154630
rect 38900 154620 38980 154630
rect 39220 154620 39300 154630
rect 39540 154620 39620 154630
rect 39860 154620 39940 154630
rect 40180 154620 40260 154630
rect 40500 154620 40580 154630
rect 40820 154620 40900 154630
rect 41140 154620 41220 154630
rect 41460 154620 41540 154630
rect 41780 154620 41860 154630
rect 42100 154620 42180 154630
rect 42420 154620 42500 154630
rect 42740 154620 42820 154630
rect 43060 154620 43140 154630
rect 43380 154620 43460 154630
rect 36100 154540 36110 154620
rect 36420 154540 36430 154620
rect 36740 154540 36750 154620
rect 37060 154540 37070 154620
rect 37380 154540 37390 154620
rect 37700 154540 37710 154620
rect 38020 154540 38030 154620
rect 38340 154540 38350 154620
rect 38660 154540 38670 154620
rect 38980 154540 38990 154620
rect 39300 154540 39310 154620
rect 39620 154540 39630 154620
rect 39940 154540 39950 154620
rect 40260 154540 40270 154620
rect 40580 154540 40590 154620
rect 40900 154540 40910 154620
rect 41220 154540 41230 154620
rect 41540 154540 41550 154620
rect 41860 154540 41870 154620
rect 42180 154540 42190 154620
rect 42500 154540 42510 154620
rect 42820 154540 42830 154620
rect 43140 154540 43150 154620
rect 43460 154540 43470 154620
rect 44025 154600 44035 154680
rect 44345 154600 44355 154680
rect 44665 154600 44675 154680
rect 44985 154600 44995 154680
rect 45305 154600 45315 154680
rect 45625 154600 45635 154680
rect 45945 154600 45955 154680
rect 46265 154600 46275 154680
rect 46585 154600 46595 154680
rect 46905 154600 46915 154680
rect 47225 154600 47235 154680
rect 47545 154600 47555 154680
rect 47865 154600 47875 154680
rect 48185 154600 48195 154680
rect 43785 154520 43865 154530
rect 44105 154520 44185 154530
rect 44425 154520 44505 154530
rect 44745 154520 44825 154530
rect 45065 154520 45145 154530
rect 45385 154520 45465 154530
rect 45705 154520 45785 154530
rect 46025 154520 46105 154530
rect 46345 154520 46425 154530
rect 46665 154520 46745 154530
rect 46985 154520 47065 154530
rect 47305 154520 47385 154530
rect 47625 154520 47705 154530
rect 47945 154520 48025 154530
rect 48265 154520 48345 154530
rect 36180 154460 36260 154470
rect 36500 154460 36580 154470
rect 36820 154460 36900 154470
rect 37140 154460 37220 154470
rect 37460 154460 37540 154470
rect 37780 154460 37860 154470
rect 38100 154460 38180 154470
rect 38420 154460 38500 154470
rect 38740 154460 38820 154470
rect 39060 154460 39140 154470
rect 39380 154460 39460 154470
rect 39700 154460 39780 154470
rect 40020 154460 40100 154470
rect 40340 154460 40420 154470
rect 40660 154460 40740 154470
rect 40980 154460 41060 154470
rect 41300 154460 41380 154470
rect 41620 154460 41700 154470
rect 41940 154460 42020 154470
rect 42260 154460 42340 154470
rect 42580 154460 42660 154470
rect 42900 154460 42980 154470
rect 43220 154460 43300 154470
rect 36260 154380 36270 154460
rect 36580 154380 36590 154460
rect 36900 154380 36910 154460
rect 37220 154380 37230 154460
rect 37540 154380 37550 154460
rect 37860 154380 37870 154460
rect 38180 154380 38190 154460
rect 38500 154380 38510 154460
rect 38820 154380 38830 154460
rect 39140 154380 39150 154460
rect 39460 154380 39470 154460
rect 39780 154380 39790 154460
rect 40100 154380 40110 154460
rect 40420 154380 40430 154460
rect 40740 154380 40750 154460
rect 41060 154380 41070 154460
rect 41380 154380 41390 154460
rect 41700 154380 41710 154460
rect 42020 154380 42030 154460
rect 42340 154380 42350 154460
rect 42660 154380 42670 154460
rect 42980 154380 42990 154460
rect 43300 154380 43310 154460
rect 43865 154440 43875 154520
rect 44185 154440 44195 154520
rect 44505 154440 44515 154520
rect 44825 154440 44835 154520
rect 45145 154440 45155 154520
rect 45465 154440 45475 154520
rect 45785 154440 45795 154520
rect 46105 154440 46115 154520
rect 46425 154440 46435 154520
rect 46745 154440 46755 154520
rect 47065 154440 47075 154520
rect 47385 154440 47395 154520
rect 47705 154440 47715 154520
rect 48025 154440 48035 154520
rect 48345 154440 48355 154520
rect 48500 154510 48605 154680
rect 48640 154600 48650 154680
rect 48790 154600 48800 154680
rect 49350 154600 49360 154680
rect 49500 154600 49510 154680
rect 49560 154510 49590 154680
rect 49650 154600 49690 154680
rect 48500 154500 48640 154510
rect 48710 154500 48790 154510
rect 49270 154500 49350 154510
rect 49420 154500 49500 154510
rect 49560 154500 49650 154510
rect 49660 154500 49690 154600
rect 43945 154360 44025 154370
rect 44265 154360 44345 154370
rect 44585 154360 44665 154370
rect 44905 154360 44985 154370
rect 45225 154360 45305 154370
rect 45545 154360 45625 154370
rect 45865 154360 45945 154370
rect 46185 154360 46265 154370
rect 46505 154360 46585 154370
rect 46825 154360 46905 154370
rect 47145 154360 47225 154370
rect 47465 154360 47545 154370
rect 47785 154360 47865 154370
rect 48105 154360 48185 154370
rect 36020 154300 36100 154310
rect 36340 154300 36420 154310
rect 36660 154300 36740 154310
rect 36980 154300 37060 154310
rect 37300 154300 37380 154310
rect 37620 154300 37700 154310
rect 37940 154300 38020 154310
rect 38260 154300 38340 154310
rect 38580 154300 38660 154310
rect 38900 154300 38980 154310
rect 39220 154300 39300 154310
rect 39540 154300 39620 154310
rect 39860 154300 39940 154310
rect 40180 154300 40260 154310
rect 40500 154300 40580 154310
rect 40820 154300 40900 154310
rect 41140 154300 41220 154310
rect 41460 154300 41540 154310
rect 41780 154300 41860 154310
rect 42100 154300 42180 154310
rect 42420 154300 42500 154310
rect 42740 154300 42820 154310
rect 43060 154300 43140 154310
rect 43380 154300 43460 154310
rect 36100 154220 36110 154300
rect 36420 154220 36430 154300
rect 36740 154220 36750 154300
rect 37060 154220 37070 154300
rect 37380 154220 37390 154300
rect 37700 154220 37710 154300
rect 38020 154220 38030 154300
rect 38340 154220 38350 154300
rect 38660 154220 38670 154300
rect 38980 154220 38990 154300
rect 39300 154220 39310 154300
rect 39620 154220 39630 154300
rect 39940 154220 39950 154300
rect 40260 154220 40270 154300
rect 40580 154220 40590 154300
rect 40900 154220 40910 154300
rect 41220 154220 41230 154300
rect 41540 154220 41550 154300
rect 41860 154220 41870 154300
rect 42180 154220 42190 154300
rect 42500 154220 42510 154300
rect 42820 154220 42830 154300
rect 43140 154220 43150 154300
rect 43460 154220 43470 154300
rect 44025 154280 44035 154360
rect 44345 154280 44355 154360
rect 44665 154280 44675 154360
rect 44985 154280 44995 154360
rect 45305 154280 45315 154360
rect 45625 154280 45635 154360
rect 45945 154280 45955 154360
rect 46265 154280 46275 154360
rect 46585 154280 46595 154360
rect 46905 154280 46915 154360
rect 47225 154280 47235 154360
rect 47545 154280 47555 154360
rect 47865 154280 47875 154360
rect 48185 154280 48195 154360
rect 48500 154330 48605 154500
rect 48640 154420 48650 154500
rect 48790 154420 48800 154500
rect 49350 154420 49360 154500
rect 49500 154420 49510 154500
rect 49560 154330 49590 154500
rect 49650 154420 49690 154500
rect 48500 154320 48640 154330
rect 48710 154320 48790 154330
rect 49270 154320 49350 154330
rect 49420 154320 49500 154330
rect 49560 154320 49650 154330
rect 49660 154320 49690 154420
rect 43785 154200 43865 154210
rect 44105 154200 44185 154210
rect 44425 154200 44505 154210
rect 44745 154200 44825 154210
rect 45065 154200 45145 154210
rect 45385 154200 45465 154210
rect 45705 154200 45785 154210
rect 46025 154200 46105 154210
rect 46345 154200 46425 154210
rect 46665 154200 46745 154210
rect 46985 154200 47065 154210
rect 47305 154200 47385 154210
rect 47625 154200 47705 154210
rect 47945 154200 48025 154210
rect 48265 154200 48345 154210
rect 36180 154140 36260 154150
rect 36500 154140 36580 154150
rect 36820 154140 36900 154150
rect 37140 154140 37220 154150
rect 37460 154140 37540 154150
rect 37780 154140 37860 154150
rect 38100 154140 38180 154150
rect 38420 154140 38500 154150
rect 38740 154140 38820 154150
rect 39060 154140 39140 154150
rect 39380 154140 39460 154150
rect 39700 154140 39780 154150
rect 40020 154140 40100 154150
rect 40340 154140 40420 154150
rect 40660 154140 40740 154150
rect 40980 154140 41060 154150
rect 41300 154140 41380 154150
rect 41620 154140 41700 154150
rect 41940 154140 42020 154150
rect 42260 154140 42340 154150
rect 42580 154140 42660 154150
rect 42900 154140 42980 154150
rect 43220 154140 43300 154150
rect 36260 154060 36270 154140
rect 36580 154060 36590 154140
rect 36900 154060 36910 154140
rect 37220 154060 37230 154140
rect 37540 154060 37550 154140
rect 37860 154060 37870 154140
rect 38180 154060 38190 154140
rect 38500 154060 38510 154140
rect 38820 154060 38830 154140
rect 39140 154060 39150 154140
rect 39460 154060 39470 154140
rect 39780 154060 39790 154140
rect 40100 154060 40110 154140
rect 40420 154060 40430 154140
rect 40740 154060 40750 154140
rect 41060 154060 41070 154140
rect 41380 154060 41390 154140
rect 41700 154060 41710 154140
rect 42020 154060 42030 154140
rect 42340 154060 42350 154140
rect 42660 154060 42670 154140
rect 42980 154060 42990 154140
rect 43300 154060 43310 154140
rect 43865 154120 43875 154200
rect 44185 154120 44195 154200
rect 44505 154120 44515 154200
rect 44825 154120 44835 154200
rect 45145 154120 45155 154200
rect 45465 154120 45475 154200
rect 45785 154120 45795 154200
rect 46105 154120 46115 154200
rect 46425 154120 46435 154200
rect 46745 154120 46755 154200
rect 47065 154120 47075 154200
rect 47385 154120 47395 154200
rect 47705 154120 47715 154200
rect 48025 154120 48035 154200
rect 48345 154120 48355 154200
rect 48500 154150 48605 154320
rect 48640 154240 48650 154320
rect 48790 154240 48800 154320
rect 49350 154240 49360 154320
rect 49500 154240 49510 154320
rect 49560 154150 49590 154320
rect 49650 154240 49690 154320
rect 48500 154140 48640 154150
rect 48710 154140 48790 154150
rect 49270 154140 49350 154150
rect 49420 154140 49500 154150
rect 49560 154140 49650 154150
rect 49660 154140 49690 154240
rect 43945 154040 44025 154050
rect 44265 154040 44345 154050
rect 44585 154040 44665 154050
rect 44905 154040 44985 154050
rect 45225 154040 45305 154050
rect 45545 154040 45625 154050
rect 45865 154040 45945 154050
rect 46185 154040 46265 154050
rect 46505 154040 46585 154050
rect 46825 154040 46905 154050
rect 47145 154040 47225 154050
rect 47465 154040 47545 154050
rect 47785 154040 47865 154050
rect 48105 154040 48185 154050
rect 36020 153980 36100 153990
rect 36340 153980 36420 153990
rect 36660 153980 36740 153990
rect 36980 153980 37060 153990
rect 37300 153980 37380 153990
rect 37620 153980 37700 153990
rect 37940 153980 38020 153990
rect 38260 153980 38340 153990
rect 38580 153980 38660 153990
rect 38900 153980 38980 153990
rect 39220 153980 39300 153990
rect 39540 153980 39620 153990
rect 39860 153980 39940 153990
rect 40180 153980 40260 153990
rect 40500 153980 40580 153990
rect 40820 153980 40900 153990
rect 41140 153980 41220 153990
rect 41460 153980 41540 153990
rect 41780 153980 41860 153990
rect 42100 153980 42180 153990
rect 42420 153980 42500 153990
rect 42740 153980 42820 153990
rect 43060 153980 43140 153990
rect 43380 153980 43460 153990
rect 36100 153900 36110 153980
rect 36420 153900 36430 153980
rect 36740 153900 36750 153980
rect 37060 153900 37070 153980
rect 37380 153900 37390 153980
rect 37700 153900 37710 153980
rect 38020 153900 38030 153980
rect 38340 153900 38350 153980
rect 38660 153900 38670 153980
rect 38980 153900 38990 153980
rect 39300 153900 39310 153980
rect 39620 153900 39630 153980
rect 39940 153900 39950 153980
rect 40260 153900 40270 153980
rect 40580 153900 40590 153980
rect 40900 153900 40910 153980
rect 41220 153900 41230 153980
rect 41540 153900 41550 153980
rect 41860 153900 41870 153980
rect 42180 153900 42190 153980
rect 42500 153900 42510 153980
rect 42820 153900 42830 153980
rect 43140 153900 43150 153980
rect 43460 153900 43470 153980
rect 44025 153960 44035 154040
rect 44345 153960 44355 154040
rect 44665 153960 44675 154040
rect 44985 153960 44995 154040
rect 45305 153960 45315 154040
rect 45625 153960 45635 154040
rect 45945 153960 45955 154040
rect 46265 153960 46275 154040
rect 46585 153960 46595 154040
rect 46905 153960 46915 154040
rect 47225 153960 47235 154040
rect 47545 153960 47555 154040
rect 47865 153960 47875 154040
rect 48185 153960 48195 154040
rect 48500 153970 48605 154140
rect 48640 154060 48650 154140
rect 48790 154060 48800 154140
rect 49350 154060 49360 154140
rect 49500 154060 49510 154140
rect 49560 153970 49590 154140
rect 49650 154060 49690 154140
rect 48500 153960 48640 153970
rect 48710 153960 48790 153970
rect 49270 153960 49350 153970
rect 49420 153960 49500 153970
rect 49560 153960 49650 153970
rect 49660 153960 49690 154060
rect 43785 153880 43865 153890
rect 44105 153880 44185 153890
rect 44425 153880 44505 153890
rect 44745 153880 44825 153890
rect 45065 153880 45145 153890
rect 45385 153880 45465 153890
rect 45705 153880 45785 153890
rect 46025 153880 46105 153890
rect 46345 153880 46425 153890
rect 46665 153880 46745 153890
rect 46985 153880 47065 153890
rect 47305 153880 47385 153890
rect 47625 153880 47705 153890
rect 47945 153880 48025 153890
rect 48265 153880 48345 153890
rect 36180 153820 36260 153830
rect 36500 153820 36580 153830
rect 36820 153820 36900 153830
rect 37140 153820 37220 153830
rect 37460 153820 37540 153830
rect 37780 153820 37860 153830
rect 38100 153820 38180 153830
rect 38420 153820 38500 153830
rect 38740 153820 38820 153830
rect 39060 153820 39140 153830
rect 39380 153820 39460 153830
rect 39700 153820 39780 153830
rect 40020 153820 40100 153830
rect 40340 153820 40420 153830
rect 40660 153820 40740 153830
rect 40980 153820 41060 153830
rect 41300 153820 41380 153830
rect 41620 153820 41700 153830
rect 41940 153820 42020 153830
rect 42260 153820 42340 153830
rect 42580 153820 42660 153830
rect 42900 153820 42980 153830
rect 43220 153820 43300 153830
rect 36260 153740 36270 153820
rect 36580 153740 36590 153820
rect 36900 153740 36910 153820
rect 37220 153740 37230 153820
rect 37540 153740 37550 153820
rect 37860 153740 37870 153820
rect 38180 153740 38190 153820
rect 38500 153740 38510 153820
rect 38820 153740 38830 153820
rect 39140 153740 39150 153820
rect 39460 153740 39470 153820
rect 39780 153740 39790 153820
rect 40100 153740 40110 153820
rect 40420 153740 40430 153820
rect 40740 153740 40750 153820
rect 41060 153740 41070 153820
rect 41380 153740 41390 153820
rect 41700 153740 41710 153820
rect 42020 153740 42030 153820
rect 42340 153740 42350 153820
rect 42660 153740 42670 153820
rect 42980 153740 42990 153820
rect 43300 153740 43310 153820
rect 43865 153800 43875 153880
rect 44185 153800 44195 153880
rect 44505 153800 44515 153880
rect 44825 153800 44835 153880
rect 45145 153800 45155 153880
rect 45465 153800 45475 153880
rect 45785 153800 45795 153880
rect 46105 153800 46115 153880
rect 46425 153800 46435 153880
rect 46745 153800 46755 153880
rect 47065 153800 47075 153880
rect 47385 153800 47395 153880
rect 47705 153800 47715 153880
rect 48025 153800 48035 153880
rect 48345 153800 48355 153880
rect 48500 153790 48605 153960
rect 48640 153880 48650 153960
rect 48790 153880 48800 153960
rect 49350 153880 49360 153960
rect 49500 153880 49510 153960
rect 49560 153790 49590 153960
rect 49650 153880 49690 153960
rect 48500 153780 48640 153790
rect 48710 153780 48790 153790
rect 49270 153780 49350 153790
rect 49420 153780 49500 153790
rect 49560 153780 49650 153790
rect 49660 153780 49690 153880
rect 43945 153720 44025 153730
rect 44265 153720 44345 153730
rect 44585 153720 44665 153730
rect 44905 153720 44985 153730
rect 45225 153720 45305 153730
rect 45545 153720 45625 153730
rect 45865 153720 45945 153730
rect 46185 153720 46265 153730
rect 46505 153720 46585 153730
rect 46825 153720 46905 153730
rect 47145 153720 47225 153730
rect 47465 153720 47545 153730
rect 47785 153720 47865 153730
rect 48105 153720 48185 153730
rect 36020 153660 36100 153670
rect 36340 153660 36420 153670
rect 36660 153660 36740 153670
rect 36980 153660 37060 153670
rect 37300 153660 37380 153670
rect 37620 153660 37700 153670
rect 37940 153660 38020 153670
rect 38260 153660 38340 153670
rect 38580 153660 38660 153670
rect 38900 153660 38980 153670
rect 39220 153660 39300 153670
rect 39540 153660 39620 153670
rect 39860 153660 39940 153670
rect 40180 153660 40260 153670
rect 40500 153660 40580 153670
rect 40820 153660 40900 153670
rect 41140 153660 41220 153670
rect 41460 153660 41540 153670
rect 41780 153660 41860 153670
rect 42100 153660 42180 153670
rect 42420 153660 42500 153670
rect 42740 153660 42820 153670
rect 43060 153660 43140 153670
rect 43380 153660 43460 153670
rect 36100 153580 36110 153660
rect 36420 153580 36430 153660
rect 36740 153580 36750 153660
rect 37060 153580 37070 153660
rect 37380 153580 37390 153660
rect 37700 153580 37710 153660
rect 38020 153580 38030 153660
rect 38340 153580 38350 153660
rect 38660 153580 38670 153660
rect 38980 153580 38990 153660
rect 39300 153580 39310 153660
rect 39620 153580 39630 153660
rect 39940 153580 39950 153660
rect 40260 153580 40270 153660
rect 40580 153580 40590 153660
rect 40900 153580 40910 153660
rect 41220 153580 41230 153660
rect 41540 153580 41550 153660
rect 41860 153580 41870 153660
rect 42180 153580 42190 153660
rect 42500 153580 42510 153660
rect 42820 153580 42830 153660
rect 43140 153580 43150 153660
rect 43460 153580 43470 153660
rect 44025 153640 44035 153720
rect 44345 153640 44355 153720
rect 44665 153640 44675 153720
rect 44985 153640 44995 153720
rect 45305 153640 45315 153720
rect 45625 153640 45635 153720
rect 45945 153640 45955 153720
rect 46265 153640 46275 153720
rect 46585 153640 46595 153720
rect 46905 153640 46915 153720
rect 47225 153640 47235 153720
rect 47545 153640 47555 153720
rect 47865 153640 47875 153720
rect 48185 153640 48195 153720
rect 48500 153610 48605 153780
rect 48640 153700 48650 153780
rect 48790 153700 48800 153780
rect 49350 153700 49360 153780
rect 49500 153700 49510 153780
rect 49560 153610 49590 153780
rect 49650 153700 49690 153780
rect 48500 153600 48640 153610
rect 48710 153600 48790 153610
rect 49270 153600 49350 153610
rect 49420 153600 49500 153610
rect 49560 153600 49650 153610
rect 49660 153600 49690 153700
rect 43785 153560 43865 153570
rect 44105 153560 44185 153570
rect 44425 153560 44505 153570
rect 44745 153560 44825 153570
rect 45065 153560 45145 153570
rect 45385 153560 45465 153570
rect 45705 153560 45785 153570
rect 46025 153560 46105 153570
rect 46345 153560 46425 153570
rect 46665 153560 46745 153570
rect 46985 153560 47065 153570
rect 47305 153560 47385 153570
rect 47625 153560 47705 153570
rect 47945 153560 48025 153570
rect 48265 153560 48345 153570
rect 36180 153500 36260 153510
rect 36500 153500 36580 153510
rect 36820 153500 36900 153510
rect 37140 153500 37220 153510
rect 37460 153500 37540 153510
rect 37780 153500 37860 153510
rect 38100 153500 38180 153510
rect 38420 153500 38500 153510
rect 38740 153500 38820 153510
rect 39060 153500 39140 153510
rect 39380 153500 39460 153510
rect 39700 153500 39780 153510
rect 40020 153500 40100 153510
rect 40340 153500 40420 153510
rect 40660 153500 40740 153510
rect 40980 153500 41060 153510
rect 41300 153500 41380 153510
rect 41620 153500 41700 153510
rect 41940 153500 42020 153510
rect 42260 153500 42340 153510
rect 42580 153500 42660 153510
rect 42900 153500 42980 153510
rect 43220 153500 43300 153510
rect 36260 153420 36270 153500
rect 36580 153420 36590 153500
rect 36900 153420 36910 153500
rect 37220 153420 37230 153500
rect 37540 153420 37550 153500
rect 37860 153420 37870 153500
rect 38180 153420 38190 153500
rect 38500 153420 38510 153500
rect 38820 153420 38830 153500
rect 39140 153420 39150 153500
rect 39460 153420 39470 153500
rect 39780 153420 39790 153500
rect 40100 153420 40110 153500
rect 40420 153420 40430 153500
rect 40740 153420 40750 153500
rect 41060 153420 41070 153500
rect 41380 153420 41390 153500
rect 41700 153420 41710 153500
rect 42020 153420 42030 153500
rect 42340 153420 42350 153500
rect 42660 153420 42670 153500
rect 42980 153420 42990 153500
rect 43300 153420 43310 153500
rect 43865 153480 43875 153560
rect 44185 153480 44195 153560
rect 44505 153480 44515 153560
rect 44825 153480 44835 153560
rect 45145 153480 45155 153560
rect 45465 153480 45475 153560
rect 45785 153480 45795 153560
rect 46105 153480 46115 153560
rect 46425 153480 46435 153560
rect 46745 153480 46755 153560
rect 47065 153480 47075 153560
rect 47385 153480 47395 153560
rect 47705 153480 47715 153560
rect 48025 153480 48035 153560
rect 48345 153480 48355 153560
rect 48500 153430 48605 153600
rect 48640 153520 48650 153600
rect 48790 153520 48800 153600
rect 49350 153520 49360 153600
rect 49500 153520 49510 153600
rect 49560 153430 49590 153600
rect 49650 153520 49690 153600
rect 48500 153420 48640 153430
rect 48710 153420 48790 153430
rect 49270 153420 49350 153430
rect 49420 153420 49500 153430
rect 49560 153420 49650 153430
rect 49660 153420 49690 153520
rect 43945 153400 44025 153410
rect 44265 153400 44345 153410
rect 44585 153400 44665 153410
rect 44905 153400 44985 153410
rect 45225 153400 45305 153410
rect 45545 153400 45625 153410
rect 45865 153400 45945 153410
rect 46185 153400 46265 153410
rect 46505 153400 46585 153410
rect 46825 153400 46905 153410
rect 47145 153400 47225 153410
rect 47465 153400 47545 153410
rect 47785 153400 47865 153410
rect 48105 153400 48185 153410
rect 36020 153340 36100 153350
rect 36340 153340 36420 153350
rect 36660 153340 36740 153350
rect 36980 153340 37060 153350
rect 37300 153340 37380 153350
rect 37620 153340 37700 153350
rect 37940 153340 38020 153350
rect 38260 153340 38340 153350
rect 38580 153340 38660 153350
rect 38900 153340 38980 153350
rect 39220 153340 39300 153350
rect 39540 153340 39620 153350
rect 39860 153340 39940 153350
rect 40180 153340 40260 153350
rect 40500 153340 40580 153350
rect 40820 153340 40900 153350
rect 41140 153340 41220 153350
rect 41460 153340 41540 153350
rect 41780 153340 41860 153350
rect 42100 153340 42180 153350
rect 42420 153340 42500 153350
rect 42740 153340 42820 153350
rect 43060 153340 43140 153350
rect 43380 153340 43460 153350
rect 36100 153260 36110 153340
rect 36420 153260 36430 153340
rect 36740 153260 36750 153340
rect 37060 153260 37070 153340
rect 37380 153260 37390 153340
rect 37700 153260 37710 153340
rect 38020 153260 38030 153340
rect 38340 153260 38350 153340
rect 38660 153260 38670 153340
rect 38980 153260 38990 153340
rect 39300 153260 39310 153340
rect 39620 153260 39630 153340
rect 39940 153260 39950 153340
rect 40260 153260 40270 153340
rect 40580 153260 40590 153340
rect 40900 153260 40910 153340
rect 41220 153260 41230 153340
rect 41540 153260 41550 153340
rect 41860 153260 41870 153340
rect 42180 153260 42190 153340
rect 42500 153260 42510 153340
rect 42820 153260 42830 153340
rect 43140 153260 43150 153340
rect 43460 153260 43470 153340
rect 44025 153320 44035 153400
rect 44345 153320 44355 153400
rect 44665 153320 44675 153400
rect 44985 153320 44995 153400
rect 45305 153320 45315 153400
rect 45625 153320 45635 153400
rect 45945 153320 45955 153400
rect 46265 153320 46275 153400
rect 46585 153320 46595 153400
rect 46905 153320 46915 153400
rect 47225 153320 47235 153400
rect 47545 153320 47555 153400
rect 47865 153320 47875 153400
rect 48185 153320 48195 153400
rect 48500 153250 48605 153420
rect 48640 153340 48650 153420
rect 48790 153340 48800 153420
rect 49350 153340 49360 153420
rect 49500 153340 49510 153420
rect 49560 153250 49590 153420
rect 49650 153340 49690 153420
rect 43785 153240 43865 153250
rect 44105 153240 44185 153250
rect 44425 153240 44505 153250
rect 44745 153240 44825 153250
rect 45065 153240 45145 153250
rect 45385 153240 45465 153250
rect 45705 153240 45785 153250
rect 46025 153240 46105 153250
rect 46345 153240 46425 153250
rect 46665 153240 46745 153250
rect 46985 153240 47065 153250
rect 47305 153240 47385 153250
rect 47625 153240 47705 153250
rect 47945 153240 48025 153250
rect 48265 153240 48345 153250
rect 48500 153240 48640 153250
rect 48710 153240 48790 153250
rect 49270 153240 49350 153250
rect 49420 153240 49500 153250
rect 49560 153240 49650 153250
rect 49660 153240 49690 153340
rect 36180 153180 36260 153190
rect 36500 153180 36580 153190
rect 36820 153180 36900 153190
rect 37140 153180 37220 153190
rect 37460 153180 37540 153190
rect 37780 153180 37860 153190
rect 38100 153180 38180 153190
rect 38420 153180 38500 153190
rect 38740 153180 38820 153190
rect 39060 153180 39140 153190
rect 39380 153180 39460 153190
rect 39700 153180 39780 153190
rect 40020 153180 40100 153190
rect 40340 153180 40420 153190
rect 40660 153180 40740 153190
rect 40980 153180 41060 153190
rect 41300 153180 41380 153190
rect 41620 153180 41700 153190
rect 41940 153180 42020 153190
rect 42260 153180 42340 153190
rect 42580 153180 42660 153190
rect 42900 153180 42980 153190
rect 43220 153180 43300 153190
rect 36260 153100 36270 153180
rect 36580 153100 36590 153180
rect 36900 153100 36910 153180
rect 37220 153100 37230 153180
rect 37540 153100 37550 153180
rect 37860 153100 37870 153180
rect 38180 153100 38190 153180
rect 38500 153100 38510 153180
rect 38820 153100 38830 153180
rect 39140 153100 39150 153180
rect 39460 153100 39470 153180
rect 39780 153100 39790 153180
rect 40100 153100 40110 153180
rect 40420 153100 40430 153180
rect 40740 153100 40750 153180
rect 41060 153100 41070 153180
rect 41380 153100 41390 153180
rect 41700 153100 41710 153180
rect 42020 153100 42030 153180
rect 42340 153100 42350 153180
rect 42660 153100 42670 153180
rect 42980 153100 42990 153180
rect 43300 153100 43310 153180
rect 43865 153160 43875 153240
rect 44185 153160 44195 153240
rect 44505 153160 44515 153240
rect 44825 153160 44835 153240
rect 45145 153160 45155 153240
rect 45465 153160 45475 153240
rect 45785 153160 45795 153240
rect 46105 153160 46115 153240
rect 46425 153160 46435 153240
rect 46745 153160 46755 153240
rect 47065 153160 47075 153240
rect 47385 153160 47395 153240
rect 47705 153160 47715 153240
rect 48025 153160 48035 153240
rect 48345 153160 48355 153240
rect 43945 153080 44025 153090
rect 44265 153080 44345 153090
rect 44585 153080 44665 153090
rect 44905 153080 44985 153090
rect 45225 153080 45305 153090
rect 45545 153080 45625 153090
rect 45865 153080 45945 153090
rect 46185 153080 46265 153090
rect 46505 153080 46585 153090
rect 46825 153080 46905 153090
rect 47145 153080 47225 153090
rect 47465 153080 47545 153090
rect 47785 153080 47865 153090
rect 48105 153080 48185 153090
rect 36020 153020 36100 153030
rect 36340 153020 36420 153030
rect 36660 153020 36740 153030
rect 36980 153020 37060 153030
rect 37300 153020 37380 153030
rect 37620 153020 37700 153030
rect 37940 153020 38020 153030
rect 38260 153020 38340 153030
rect 38580 153020 38660 153030
rect 38900 153020 38980 153030
rect 39220 153020 39300 153030
rect 39540 153020 39620 153030
rect 39860 153020 39940 153030
rect 40180 153020 40260 153030
rect 40500 153020 40580 153030
rect 40820 153020 40900 153030
rect 41140 153020 41220 153030
rect 41460 153020 41540 153030
rect 41780 153020 41860 153030
rect 42100 153020 42180 153030
rect 42420 153020 42500 153030
rect 42740 153020 42820 153030
rect 43060 153020 43140 153030
rect 43380 153020 43460 153030
rect 36100 152940 36110 153020
rect 36420 152940 36430 153020
rect 36740 152940 36750 153020
rect 37060 152940 37070 153020
rect 37380 152940 37390 153020
rect 37700 152940 37710 153020
rect 38020 152940 38030 153020
rect 38340 152940 38350 153020
rect 38660 152940 38670 153020
rect 38980 152940 38990 153020
rect 39300 152940 39310 153020
rect 39620 152940 39630 153020
rect 39940 152940 39950 153020
rect 40260 152940 40270 153020
rect 40580 152940 40590 153020
rect 40900 152940 40910 153020
rect 41220 152940 41230 153020
rect 41540 152940 41550 153020
rect 41860 152940 41870 153020
rect 42180 152940 42190 153020
rect 42500 152940 42510 153020
rect 42820 152940 42830 153020
rect 43140 152940 43150 153020
rect 43460 152940 43470 153020
rect 44025 153000 44035 153080
rect 44345 153000 44355 153080
rect 44665 153000 44675 153080
rect 44985 153000 44995 153080
rect 45305 153000 45315 153080
rect 45625 153000 45635 153080
rect 45945 153000 45955 153080
rect 46265 153000 46275 153080
rect 46585 153000 46595 153080
rect 46905 153000 46915 153080
rect 47225 153000 47235 153080
rect 47545 153000 47555 153080
rect 47865 153000 47875 153080
rect 48185 153000 48195 153080
rect 48500 153070 48605 153240
rect 48640 153160 48650 153240
rect 48790 153160 48800 153240
rect 49350 153160 49360 153240
rect 49500 153160 49510 153240
rect 49560 153070 49590 153240
rect 49650 153160 49690 153240
rect 48500 153060 48640 153070
rect 48710 153060 48790 153070
rect 49270 153060 49350 153070
rect 49420 153060 49500 153070
rect 49560 153060 49650 153070
rect 49660 153060 49690 153160
rect 43785 152920 43865 152930
rect 44105 152920 44185 152930
rect 44425 152920 44505 152930
rect 44745 152920 44825 152930
rect 45065 152920 45145 152930
rect 45385 152920 45465 152930
rect 45705 152920 45785 152930
rect 46025 152920 46105 152930
rect 46345 152920 46425 152930
rect 46665 152920 46745 152930
rect 46985 152920 47065 152930
rect 47305 152920 47385 152930
rect 47625 152920 47705 152930
rect 47945 152920 48025 152930
rect 48265 152920 48345 152930
rect 36180 152860 36260 152870
rect 36500 152860 36580 152870
rect 36820 152860 36900 152870
rect 37140 152860 37220 152870
rect 37460 152860 37540 152870
rect 37780 152860 37860 152870
rect 38100 152860 38180 152870
rect 38420 152860 38500 152870
rect 38740 152860 38820 152870
rect 39060 152860 39140 152870
rect 39380 152860 39460 152870
rect 39700 152860 39780 152870
rect 40020 152860 40100 152870
rect 40340 152860 40420 152870
rect 40660 152860 40740 152870
rect 40980 152860 41060 152870
rect 41300 152860 41380 152870
rect 41620 152860 41700 152870
rect 41940 152860 42020 152870
rect 42260 152860 42340 152870
rect 42580 152860 42660 152870
rect 42900 152860 42980 152870
rect 43220 152860 43300 152870
rect 36260 152780 36270 152860
rect 36580 152780 36590 152860
rect 36900 152780 36910 152860
rect 37220 152780 37230 152860
rect 37540 152780 37550 152860
rect 37860 152780 37870 152860
rect 38180 152780 38190 152860
rect 38500 152780 38510 152860
rect 38820 152780 38830 152860
rect 39140 152780 39150 152860
rect 39460 152780 39470 152860
rect 39780 152780 39790 152860
rect 40100 152780 40110 152860
rect 40420 152780 40430 152860
rect 40740 152780 40750 152860
rect 41060 152780 41070 152860
rect 41380 152780 41390 152860
rect 41700 152780 41710 152860
rect 42020 152780 42030 152860
rect 42340 152780 42350 152860
rect 42660 152780 42670 152860
rect 42980 152780 42990 152860
rect 43300 152780 43310 152860
rect 43865 152840 43875 152920
rect 44185 152840 44195 152920
rect 44505 152840 44515 152920
rect 44825 152840 44835 152920
rect 45145 152840 45155 152920
rect 45465 152840 45475 152920
rect 45785 152840 45795 152920
rect 46105 152840 46115 152920
rect 46425 152840 46435 152920
rect 46745 152840 46755 152920
rect 47065 152840 47075 152920
rect 47385 152840 47395 152920
rect 47705 152840 47715 152920
rect 48025 152840 48035 152920
rect 48345 152840 48355 152920
rect 48500 152890 48605 153060
rect 48640 152980 48650 153060
rect 48790 152980 48800 153060
rect 49350 152980 49360 153060
rect 49500 152980 49510 153060
rect 49560 152900 49590 153060
rect 49650 152980 49690 153060
rect 49660 152900 49690 152980
rect 49790 152900 49800 158900
rect 49890 158820 49970 158830
rect 50210 158820 50290 158830
rect 49970 158740 49980 158820
rect 50290 158740 50300 158820
rect 49890 158640 49970 158650
rect 50210 158640 50290 158650
rect 49970 158560 49980 158640
rect 50290 158560 50300 158640
rect 49890 158460 49970 158470
rect 50210 158460 50290 158470
rect 49970 158380 49980 158460
rect 50290 158380 50300 158460
rect 49890 158280 49970 158290
rect 50210 158280 50290 158290
rect 49970 158200 49980 158280
rect 50290 158200 50300 158280
rect 49890 158100 49970 158110
rect 50210 158100 50290 158110
rect 49970 158020 49980 158100
rect 50290 158020 50300 158100
rect 49890 157920 49970 157930
rect 50210 157920 50290 157930
rect 49970 157840 49980 157920
rect 50290 157840 50300 157920
rect 49890 157740 49970 157750
rect 50210 157740 50290 157750
rect 49970 157660 49980 157740
rect 50290 157660 50300 157740
rect 49890 157560 49970 157570
rect 50210 157560 50290 157570
rect 49970 157480 49980 157560
rect 50290 157480 50300 157560
rect 49890 157380 49970 157390
rect 50210 157380 50290 157390
rect 49970 157300 49980 157380
rect 50290 157300 50300 157380
rect 49890 157200 49970 157210
rect 50210 157200 50290 157210
rect 49970 157120 49980 157200
rect 50290 157120 50300 157200
rect 49890 157020 49970 157030
rect 50210 157020 50290 157030
rect 49970 156940 49980 157020
rect 50290 156940 50300 157020
rect 49890 156840 49970 156850
rect 50210 156840 50290 156850
rect 49970 156760 49980 156840
rect 50290 156760 50300 156840
rect 49890 156660 49970 156670
rect 50210 156660 50290 156670
rect 49970 156580 49980 156660
rect 50290 156580 50300 156660
rect 49890 156480 49970 156490
rect 50210 156480 50290 156490
rect 49970 156400 49980 156480
rect 50290 156400 50300 156480
rect 49890 156300 49970 156310
rect 50210 156300 50290 156310
rect 49970 156220 49980 156300
rect 50290 156220 50300 156300
rect 49890 156120 49970 156130
rect 50210 156120 50290 156130
rect 49970 156040 49980 156120
rect 50290 156040 50300 156120
rect 49890 155940 49970 155950
rect 50210 155940 50290 155950
rect 49970 155860 49980 155940
rect 50290 155860 50300 155940
rect 49890 155760 49970 155770
rect 50210 155760 50290 155770
rect 49970 155680 49980 155760
rect 50290 155680 50300 155760
rect 49890 155580 49970 155590
rect 50210 155580 50290 155590
rect 49970 155500 49980 155580
rect 50290 155500 50300 155580
rect 49890 155400 49970 155410
rect 50210 155400 50290 155410
rect 49970 155320 49980 155400
rect 50290 155320 50300 155400
rect 49890 155220 49970 155230
rect 50210 155220 50290 155230
rect 49970 155140 49980 155220
rect 50290 155140 50300 155220
rect 49890 155040 49970 155050
rect 50210 155040 50290 155050
rect 49970 154960 49980 155040
rect 50290 154960 50300 155040
rect 49890 154860 49970 154870
rect 50210 154860 50290 154870
rect 49970 154780 49980 154860
rect 50290 154780 50300 154860
rect 49890 154680 49970 154690
rect 50210 154680 50290 154690
rect 49970 154600 49980 154680
rect 50290 154600 50300 154680
rect 49890 154500 49970 154510
rect 50210 154500 50290 154510
rect 49970 154420 49980 154500
rect 50290 154420 50300 154500
rect 49890 154320 49970 154330
rect 50210 154320 50290 154330
rect 49970 154240 49980 154320
rect 50290 154240 50300 154320
rect 49890 154140 49970 154150
rect 50210 154140 50290 154150
rect 49970 154060 49980 154140
rect 50290 154060 50300 154140
rect 49890 153960 49970 153970
rect 50210 153960 50290 153970
rect 49970 153880 49980 153960
rect 50290 153880 50300 153960
rect 49890 153780 49970 153790
rect 50210 153780 50290 153790
rect 49970 153700 49980 153780
rect 50290 153700 50300 153780
rect 49890 153600 49970 153610
rect 50210 153600 50290 153610
rect 49970 153520 49980 153600
rect 50290 153520 50300 153600
rect 49890 153420 49970 153430
rect 50210 153420 50290 153430
rect 49970 153340 49980 153420
rect 50290 153340 50300 153420
rect 49890 153240 49970 153250
rect 50210 153240 50290 153250
rect 49970 153160 49980 153240
rect 50290 153160 50300 153240
rect 49890 153060 49970 153070
rect 50210 153060 50290 153070
rect 49970 152980 49980 153060
rect 50290 152980 50300 153060
rect 50470 152900 50480 158900
rect 50490 152900 50520 158900
rect 50590 158830 50620 158900
rect 50820 158830 50850 158900
rect 50530 158820 50620 158830
rect 50680 158820 50760 158830
rect 50820 158820 50910 158830
rect 50920 158820 50950 158900
rect 50590 158650 50620 158820
rect 50760 158740 50770 158820
rect 50820 158650 50850 158820
rect 50910 158740 50950 158820
rect 50530 158640 50620 158650
rect 50680 158640 50760 158650
rect 50820 158640 50910 158650
rect 50920 158640 50950 158740
rect 50590 158470 50620 158640
rect 50760 158560 50770 158640
rect 50820 158470 50850 158640
rect 50910 158560 50950 158640
rect 50530 158460 50620 158470
rect 50680 158460 50760 158470
rect 50820 158460 50910 158470
rect 50920 158460 50950 158560
rect 50590 158290 50620 158460
rect 50760 158380 50770 158460
rect 50820 158290 50850 158460
rect 50910 158380 50950 158460
rect 50530 158280 50620 158290
rect 50680 158280 50760 158290
rect 50820 158280 50910 158290
rect 50920 158280 50950 158380
rect 50590 158110 50620 158280
rect 50760 158200 50770 158280
rect 50820 158110 50850 158280
rect 50910 158200 50950 158280
rect 50530 158100 50620 158110
rect 50680 158100 50760 158110
rect 50820 158100 50910 158110
rect 50920 158100 50950 158200
rect 50590 157930 50620 158100
rect 50760 158020 50770 158100
rect 50820 157930 50850 158100
rect 50910 158020 50950 158100
rect 50530 157920 50620 157930
rect 50680 157920 50760 157930
rect 50820 157920 50910 157930
rect 50920 157920 50950 158020
rect 50590 157750 50620 157920
rect 50760 157840 50770 157920
rect 50820 157750 50850 157920
rect 50910 157840 50950 157920
rect 50530 157740 50620 157750
rect 50680 157740 50760 157750
rect 50820 157740 50910 157750
rect 50920 157740 50950 157840
rect 50590 157570 50620 157740
rect 50760 157660 50770 157740
rect 50820 157570 50850 157740
rect 50910 157660 50950 157740
rect 50530 157560 50620 157570
rect 50680 157560 50760 157570
rect 50820 157560 50910 157570
rect 50920 157560 50950 157660
rect 50590 157390 50620 157560
rect 50760 157480 50770 157560
rect 50820 157390 50850 157560
rect 50910 157480 50950 157560
rect 50530 157380 50620 157390
rect 50680 157380 50760 157390
rect 50820 157380 50910 157390
rect 50920 157380 50950 157480
rect 50590 157210 50620 157380
rect 50760 157300 50770 157380
rect 50820 157210 50850 157380
rect 50910 157300 50950 157380
rect 50530 157200 50620 157210
rect 50680 157200 50760 157210
rect 50820 157200 50910 157210
rect 50920 157200 50950 157300
rect 50590 157030 50620 157200
rect 50760 157120 50770 157200
rect 50820 157030 50850 157200
rect 50910 157120 50950 157200
rect 50530 157020 50620 157030
rect 50680 157020 50760 157030
rect 50820 157020 50910 157030
rect 50920 157020 50950 157120
rect 50590 156850 50620 157020
rect 50760 156940 50770 157020
rect 50820 156850 50850 157020
rect 50910 156940 50950 157020
rect 50530 156840 50620 156850
rect 50680 156840 50760 156850
rect 50820 156840 50910 156850
rect 50920 156840 50950 156940
rect 50590 156670 50620 156840
rect 50760 156760 50770 156840
rect 50820 156670 50850 156840
rect 50910 156760 50950 156840
rect 50530 156660 50620 156670
rect 50680 156660 50760 156670
rect 50820 156660 50910 156670
rect 50920 156660 50950 156760
rect 50590 156490 50620 156660
rect 50760 156580 50770 156660
rect 50820 156490 50850 156660
rect 50910 156580 50950 156660
rect 50530 156480 50620 156490
rect 50680 156480 50760 156490
rect 50820 156480 50910 156490
rect 50920 156480 50950 156580
rect 50590 156310 50620 156480
rect 50760 156400 50770 156480
rect 50820 156310 50850 156480
rect 50910 156400 50950 156480
rect 50530 156300 50620 156310
rect 50680 156300 50760 156310
rect 50820 156300 50910 156310
rect 50920 156300 50950 156400
rect 50590 156130 50620 156300
rect 50760 156220 50770 156300
rect 50820 156130 50850 156300
rect 50910 156220 50950 156300
rect 50530 156120 50620 156130
rect 50680 156120 50760 156130
rect 50820 156120 50910 156130
rect 50920 156120 50950 156220
rect 50590 155950 50620 156120
rect 50760 156040 50770 156120
rect 50820 155950 50850 156120
rect 50910 156040 50950 156120
rect 50530 155940 50620 155950
rect 50680 155940 50760 155950
rect 50820 155940 50910 155950
rect 50920 155940 50950 156040
rect 50590 155770 50620 155940
rect 50760 155860 50770 155940
rect 50820 155770 50850 155940
rect 50910 155860 50950 155940
rect 50530 155760 50620 155770
rect 50680 155760 50760 155770
rect 50820 155760 50910 155770
rect 50920 155760 50950 155860
rect 50590 155590 50620 155760
rect 50760 155680 50770 155760
rect 50820 155590 50850 155760
rect 50910 155680 50950 155760
rect 50530 155580 50620 155590
rect 50680 155580 50760 155590
rect 50820 155580 50910 155590
rect 50920 155580 50950 155680
rect 50590 155410 50620 155580
rect 50760 155500 50770 155580
rect 50820 155410 50850 155580
rect 50910 155500 50950 155580
rect 50530 155400 50620 155410
rect 50680 155400 50760 155410
rect 50820 155400 50910 155410
rect 50920 155400 50950 155500
rect 50590 155230 50620 155400
rect 50760 155320 50770 155400
rect 50820 155230 50850 155400
rect 50910 155320 50950 155400
rect 50530 155220 50620 155230
rect 50680 155220 50760 155230
rect 50820 155220 50910 155230
rect 50920 155220 50950 155320
rect 50590 155050 50620 155220
rect 50760 155140 50770 155220
rect 50820 155050 50850 155220
rect 50910 155140 50950 155220
rect 50530 155040 50620 155050
rect 50680 155040 50760 155050
rect 50820 155040 50910 155050
rect 50920 155040 50950 155140
rect 50590 154870 50620 155040
rect 50760 154960 50770 155040
rect 50820 154870 50850 155040
rect 50910 154960 50950 155040
rect 50530 154860 50620 154870
rect 50680 154860 50760 154870
rect 50820 154860 50910 154870
rect 50920 154860 50950 154960
rect 50590 154690 50620 154860
rect 50760 154780 50770 154860
rect 50820 154690 50850 154860
rect 50910 154780 50950 154860
rect 50530 154680 50620 154690
rect 50680 154680 50760 154690
rect 50820 154680 50910 154690
rect 50920 154680 50950 154780
rect 50590 154510 50620 154680
rect 50760 154600 50770 154680
rect 50820 154510 50850 154680
rect 50910 154600 50950 154680
rect 50530 154500 50620 154510
rect 50680 154500 50760 154510
rect 50820 154500 50910 154510
rect 50920 154500 50950 154600
rect 50590 154330 50620 154500
rect 50760 154420 50770 154500
rect 50820 154330 50850 154500
rect 50910 154420 50950 154500
rect 50530 154320 50620 154330
rect 50680 154320 50760 154330
rect 50820 154320 50910 154330
rect 50920 154320 50950 154420
rect 50590 154150 50620 154320
rect 50760 154240 50770 154320
rect 50820 154150 50850 154320
rect 50910 154240 50950 154320
rect 50530 154140 50620 154150
rect 50680 154140 50760 154150
rect 50820 154140 50910 154150
rect 50920 154140 50950 154240
rect 50590 153970 50620 154140
rect 50760 154060 50770 154140
rect 50820 153970 50850 154140
rect 50910 154060 50950 154140
rect 50530 153960 50620 153970
rect 50680 153960 50760 153970
rect 50820 153960 50910 153970
rect 50920 153960 50950 154060
rect 50590 153790 50620 153960
rect 50760 153880 50770 153960
rect 50820 153790 50850 153960
rect 50910 153880 50950 153960
rect 50530 153780 50620 153790
rect 50680 153780 50760 153790
rect 50820 153780 50910 153790
rect 50920 153780 50950 153880
rect 50590 153610 50620 153780
rect 50760 153700 50770 153780
rect 50820 153610 50850 153780
rect 50910 153700 50950 153780
rect 50530 153600 50620 153610
rect 50680 153600 50760 153610
rect 50820 153600 50910 153610
rect 50920 153600 50950 153700
rect 50590 153430 50620 153600
rect 50760 153520 50770 153600
rect 50820 153430 50850 153600
rect 50910 153520 50950 153600
rect 50530 153420 50620 153430
rect 50680 153420 50760 153430
rect 50820 153420 50910 153430
rect 50920 153420 50950 153520
rect 50590 153250 50620 153420
rect 50760 153340 50770 153420
rect 50820 153250 50850 153420
rect 50910 153340 50950 153420
rect 50530 153240 50620 153250
rect 50680 153240 50760 153250
rect 50820 153240 50910 153250
rect 50920 153240 50950 153340
rect 50590 153070 50620 153240
rect 50760 153160 50770 153240
rect 50820 153070 50850 153240
rect 50910 153160 50950 153240
rect 50530 153060 50620 153070
rect 50680 153060 50760 153070
rect 50820 153060 50910 153070
rect 50920 153060 50950 153160
rect 50590 152900 50620 153060
rect 50760 152980 50770 153060
rect 50820 152900 50850 153060
rect 50910 152980 50950 153060
rect 50920 152900 50950 152980
rect 51050 152900 51060 158900
rect 51150 158820 51230 158830
rect 51470 158820 51550 158830
rect 51230 158740 51240 158820
rect 51550 158740 51560 158820
rect 51150 158640 51230 158650
rect 51470 158640 51550 158650
rect 51230 158560 51240 158640
rect 51550 158560 51560 158640
rect 51150 158460 51230 158470
rect 51470 158460 51550 158470
rect 51230 158380 51240 158460
rect 51550 158380 51560 158460
rect 51150 158280 51230 158290
rect 51470 158280 51550 158290
rect 51230 158200 51240 158280
rect 51550 158200 51560 158280
rect 51150 158100 51230 158110
rect 51470 158100 51550 158110
rect 51230 158020 51240 158100
rect 51550 158020 51560 158100
rect 51150 157920 51230 157930
rect 51470 157920 51550 157930
rect 51230 157840 51240 157920
rect 51550 157840 51560 157920
rect 51150 157740 51230 157750
rect 51470 157740 51550 157750
rect 51230 157660 51240 157740
rect 51550 157660 51560 157740
rect 51150 157560 51230 157570
rect 51470 157560 51550 157570
rect 51230 157480 51240 157560
rect 51550 157480 51560 157560
rect 51150 157380 51230 157390
rect 51470 157380 51550 157390
rect 51230 157300 51240 157380
rect 51550 157300 51560 157380
rect 51150 157200 51230 157210
rect 51470 157200 51550 157210
rect 51230 157120 51240 157200
rect 51550 157120 51560 157200
rect 51150 157020 51230 157030
rect 51470 157020 51550 157030
rect 51230 156940 51240 157020
rect 51550 156940 51560 157020
rect 51150 156840 51230 156850
rect 51470 156840 51550 156850
rect 51230 156760 51240 156840
rect 51550 156760 51560 156840
rect 51150 156660 51230 156670
rect 51470 156660 51550 156670
rect 51230 156580 51240 156660
rect 51550 156580 51560 156660
rect 51150 156480 51230 156490
rect 51470 156480 51550 156490
rect 51230 156400 51240 156480
rect 51550 156400 51560 156480
rect 51150 156300 51230 156310
rect 51470 156300 51550 156310
rect 51230 156220 51240 156300
rect 51550 156220 51560 156300
rect 51150 156120 51230 156130
rect 51470 156120 51550 156130
rect 51230 156040 51240 156120
rect 51550 156040 51560 156120
rect 51150 155940 51230 155950
rect 51470 155940 51550 155950
rect 51230 155860 51240 155940
rect 51550 155860 51560 155940
rect 51150 155760 51230 155770
rect 51470 155760 51550 155770
rect 51230 155680 51240 155760
rect 51550 155680 51560 155760
rect 51150 155580 51230 155590
rect 51470 155580 51550 155590
rect 51230 155500 51240 155580
rect 51550 155500 51560 155580
rect 51150 155400 51230 155410
rect 51470 155400 51550 155410
rect 51230 155320 51240 155400
rect 51550 155320 51560 155400
rect 51150 155220 51230 155230
rect 51470 155220 51550 155230
rect 51230 155140 51240 155220
rect 51550 155140 51560 155220
rect 51150 155040 51230 155050
rect 51470 155040 51550 155050
rect 51230 154960 51240 155040
rect 51550 154960 51560 155040
rect 51150 154860 51230 154870
rect 51470 154860 51550 154870
rect 51230 154780 51240 154860
rect 51550 154780 51560 154860
rect 51150 154680 51230 154690
rect 51470 154680 51550 154690
rect 51230 154600 51240 154680
rect 51550 154600 51560 154680
rect 51150 154500 51230 154510
rect 51470 154500 51550 154510
rect 51230 154420 51240 154500
rect 51550 154420 51560 154500
rect 51150 154320 51230 154330
rect 51470 154320 51550 154330
rect 51230 154240 51240 154320
rect 51550 154240 51560 154320
rect 51150 154140 51230 154150
rect 51470 154140 51550 154150
rect 51230 154060 51240 154140
rect 51550 154060 51560 154140
rect 51150 153960 51230 153970
rect 51470 153960 51550 153970
rect 51230 153880 51240 153960
rect 51550 153880 51560 153960
rect 51150 153780 51230 153790
rect 51470 153780 51550 153790
rect 51230 153700 51240 153780
rect 51550 153700 51560 153780
rect 51150 153600 51230 153610
rect 51470 153600 51550 153610
rect 51230 153520 51240 153600
rect 51550 153520 51560 153600
rect 51150 153420 51230 153430
rect 51470 153420 51550 153430
rect 51230 153340 51240 153420
rect 51550 153340 51560 153420
rect 51150 153240 51230 153250
rect 51470 153240 51550 153250
rect 51230 153160 51240 153240
rect 51550 153160 51560 153240
rect 51150 153060 51230 153070
rect 51470 153060 51550 153070
rect 51230 152980 51240 153060
rect 51550 152980 51560 153060
rect 51730 152900 51740 158900
rect 51750 152900 51780 158900
rect 51850 158830 51880 158900
rect 52080 158830 52110 158900
rect 51790 158820 51880 158830
rect 51940 158820 52020 158830
rect 52080 158820 52170 158830
rect 52180 158820 52210 158900
rect 51850 158650 51880 158820
rect 52020 158740 52030 158820
rect 52080 158650 52110 158820
rect 52170 158740 52210 158820
rect 51790 158640 51880 158650
rect 51940 158640 52020 158650
rect 52080 158640 52170 158650
rect 52180 158640 52210 158740
rect 51850 158470 51880 158640
rect 52020 158560 52030 158640
rect 52080 158470 52110 158640
rect 52170 158560 52210 158640
rect 51790 158460 51880 158470
rect 51940 158460 52020 158470
rect 52080 158460 52170 158470
rect 52180 158460 52210 158560
rect 51850 158290 51880 158460
rect 52020 158380 52030 158460
rect 52080 158290 52110 158460
rect 52170 158380 52210 158460
rect 51790 158280 51880 158290
rect 51940 158280 52020 158290
rect 52080 158280 52170 158290
rect 52180 158280 52210 158380
rect 51850 158110 51880 158280
rect 52020 158200 52030 158280
rect 52080 158110 52110 158280
rect 52170 158200 52210 158280
rect 51790 158100 51880 158110
rect 51940 158100 52020 158110
rect 52080 158100 52170 158110
rect 52180 158100 52210 158200
rect 51850 157930 51880 158100
rect 52020 158020 52030 158100
rect 52080 157930 52110 158100
rect 52170 158020 52210 158100
rect 51790 157920 51880 157930
rect 51940 157920 52020 157930
rect 52080 157920 52170 157930
rect 52180 157920 52210 158020
rect 51850 157750 51880 157920
rect 52020 157840 52030 157920
rect 52080 157750 52110 157920
rect 52170 157840 52210 157920
rect 51790 157740 51880 157750
rect 51940 157740 52020 157750
rect 52080 157740 52170 157750
rect 52180 157740 52210 157840
rect 51850 157570 51880 157740
rect 52020 157660 52030 157740
rect 52080 157570 52110 157740
rect 52170 157660 52210 157740
rect 51790 157560 51880 157570
rect 51940 157560 52020 157570
rect 52080 157560 52170 157570
rect 52180 157560 52210 157660
rect 51850 157390 51880 157560
rect 52020 157480 52030 157560
rect 52080 157390 52110 157560
rect 52170 157480 52210 157560
rect 51790 157380 51880 157390
rect 51940 157380 52020 157390
rect 52080 157380 52170 157390
rect 52180 157380 52210 157480
rect 51850 157210 51880 157380
rect 52020 157300 52030 157380
rect 52080 157210 52110 157380
rect 52170 157300 52210 157380
rect 51790 157200 51880 157210
rect 51940 157200 52020 157210
rect 52080 157200 52170 157210
rect 52180 157200 52210 157300
rect 51850 157030 51880 157200
rect 52020 157120 52030 157200
rect 52080 157030 52110 157200
rect 52170 157120 52210 157200
rect 51790 157020 51880 157030
rect 51940 157020 52020 157030
rect 52080 157020 52170 157030
rect 52180 157020 52210 157120
rect 51850 156850 51880 157020
rect 52020 156940 52030 157020
rect 52080 156850 52110 157020
rect 52170 156940 52210 157020
rect 51790 156840 51880 156850
rect 51940 156840 52020 156850
rect 52080 156840 52170 156850
rect 52180 156840 52210 156940
rect 51850 156670 51880 156840
rect 52020 156760 52030 156840
rect 52080 156670 52110 156840
rect 52170 156760 52210 156840
rect 51790 156660 51880 156670
rect 51940 156660 52020 156670
rect 52080 156660 52170 156670
rect 52180 156660 52210 156760
rect 51850 156490 51880 156660
rect 52020 156580 52030 156660
rect 52080 156490 52110 156660
rect 52170 156580 52210 156660
rect 51790 156480 51880 156490
rect 51940 156480 52020 156490
rect 52080 156480 52170 156490
rect 52180 156480 52210 156580
rect 51850 156310 51880 156480
rect 52020 156400 52030 156480
rect 52080 156310 52110 156480
rect 52170 156400 52210 156480
rect 51790 156300 51880 156310
rect 51940 156300 52020 156310
rect 52080 156300 52170 156310
rect 52180 156300 52210 156400
rect 51850 156130 51880 156300
rect 52020 156220 52030 156300
rect 52080 156130 52110 156300
rect 52170 156220 52210 156300
rect 51790 156120 51880 156130
rect 51940 156120 52020 156130
rect 52080 156120 52170 156130
rect 52180 156120 52210 156220
rect 51850 155950 51880 156120
rect 52020 156040 52030 156120
rect 52080 155950 52110 156120
rect 52170 156040 52210 156120
rect 51790 155940 51880 155950
rect 51940 155940 52020 155950
rect 52080 155940 52170 155950
rect 52180 155940 52210 156040
rect 51850 155770 51880 155940
rect 52020 155860 52030 155940
rect 52080 155770 52110 155940
rect 52170 155860 52210 155940
rect 51790 155760 51880 155770
rect 51940 155760 52020 155770
rect 52080 155760 52170 155770
rect 52180 155760 52210 155860
rect 51850 155590 51880 155760
rect 52020 155680 52030 155760
rect 52080 155590 52110 155760
rect 52170 155680 52210 155760
rect 51790 155580 51880 155590
rect 51940 155580 52020 155590
rect 52080 155580 52170 155590
rect 52180 155580 52210 155680
rect 51850 155410 51880 155580
rect 52020 155500 52030 155580
rect 52080 155410 52110 155580
rect 52170 155500 52210 155580
rect 51790 155400 51880 155410
rect 51940 155400 52020 155410
rect 52080 155400 52170 155410
rect 52180 155400 52210 155500
rect 51850 155230 51880 155400
rect 52020 155320 52030 155400
rect 52080 155230 52110 155400
rect 52170 155320 52210 155400
rect 51790 155220 51880 155230
rect 51940 155220 52020 155230
rect 52080 155220 52170 155230
rect 52180 155220 52210 155320
rect 51850 155050 51880 155220
rect 52020 155140 52030 155220
rect 52080 155050 52110 155220
rect 52170 155140 52210 155220
rect 51790 155040 51880 155050
rect 51940 155040 52020 155050
rect 52080 155040 52170 155050
rect 52180 155040 52210 155140
rect 51850 154870 51880 155040
rect 52020 154960 52030 155040
rect 52080 154870 52110 155040
rect 52170 154960 52210 155040
rect 51790 154860 51880 154870
rect 51940 154860 52020 154870
rect 52080 154860 52170 154870
rect 52180 154860 52210 154960
rect 51850 154690 51880 154860
rect 52020 154780 52030 154860
rect 52080 154690 52110 154860
rect 52170 154780 52210 154860
rect 51790 154680 51880 154690
rect 51940 154680 52020 154690
rect 52080 154680 52170 154690
rect 52180 154680 52210 154780
rect 51850 154510 51880 154680
rect 52020 154600 52030 154680
rect 52080 154510 52110 154680
rect 52170 154600 52210 154680
rect 51790 154500 51880 154510
rect 51940 154500 52020 154510
rect 52080 154500 52170 154510
rect 52180 154500 52210 154600
rect 51850 154330 51880 154500
rect 52020 154420 52030 154500
rect 52080 154330 52110 154500
rect 52170 154420 52210 154500
rect 51790 154320 51880 154330
rect 51940 154320 52020 154330
rect 52080 154320 52170 154330
rect 52180 154320 52210 154420
rect 51850 154150 51880 154320
rect 52020 154240 52030 154320
rect 52080 154150 52110 154320
rect 52170 154240 52210 154320
rect 51790 154140 51880 154150
rect 51940 154140 52020 154150
rect 52080 154140 52170 154150
rect 52180 154140 52210 154240
rect 51850 153970 51880 154140
rect 52020 154060 52030 154140
rect 52080 153970 52110 154140
rect 52170 154060 52210 154140
rect 51790 153960 51880 153970
rect 51940 153960 52020 153970
rect 52080 153960 52170 153970
rect 52180 153960 52210 154060
rect 51850 153790 51880 153960
rect 52020 153880 52030 153960
rect 52080 153790 52110 153960
rect 52170 153880 52210 153960
rect 51790 153780 51880 153790
rect 51940 153780 52020 153790
rect 52080 153780 52170 153790
rect 52180 153780 52210 153880
rect 51850 153610 51880 153780
rect 52020 153700 52030 153780
rect 52080 153610 52110 153780
rect 52170 153700 52210 153780
rect 51790 153600 51880 153610
rect 51940 153600 52020 153610
rect 52080 153600 52170 153610
rect 52180 153600 52210 153700
rect 51850 153430 51880 153600
rect 52020 153520 52030 153600
rect 52080 153430 52110 153600
rect 52170 153520 52210 153600
rect 51790 153420 51880 153430
rect 51940 153420 52020 153430
rect 52080 153420 52170 153430
rect 52180 153420 52210 153520
rect 51850 153250 51880 153420
rect 52020 153340 52030 153420
rect 52080 153250 52110 153420
rect 52170 153340 52210 153420
rect 51790 153240 51880 153250
rect 51940 153240 52020 153250
rect 52080 153240 52170 153250
rect 52180 153240 52210 153340
rect 51850 153070 51880 153240
rect 52020 153160 52030 153240
rect 52080 153070 52110 153240
rect 52170 153160 52210 153240
rect 51790 153060 51880 153070
rect 51940 153060 52020 153070
rect 52080 153060 52170 153070
rect 52180 153060 52210 153160
rect 51850 152900 51880 153060
rect 52020 152980 52030 153060
rect 52080 152900 52110 153060
rect 52170 152980 52210 153060
rect 52180 152900 52210 152980
rect 52310 152900 52320 158900
rect 52410 158820 52490 158830
rect 52730 158820 52810 158830
rect 52490 158740 52500 158820
rect 52810 158740 52820 158820
rect 52410 158640 52490 158650
rect 52730 158640 52810 158650
rect 52490 158560 52500 158640
rect 52810 158560 52820 158640
rect 52410 158460 52490 158470
rect 52730 158460 52810 158470
rect 52490 158380 52500 158460
rect 52810 158380 52820 158460
rect 52410 158280 52490 158290
rect 52730 158280 52810 158290
rect 52490 158200 52500 158280
rect 52810 158200 52820 158280
rect 52410 158100 52490 158110
rect 52730 158100 52810 158110
rect 52490 158020 52500 158100
rect 52810 158020 52820 158100
rect 52410 157920 52490 157930
rect 52730 157920 52810 157930
rect 52490 157840 52500 157920
rect 52810 157840 52820 157920
rect 52410 157740 52490 157750
rect 52730 157740 52810 157750
rect 52490 157660 52500 157740
rect 52810 157660 52820 157740
rect 52410 157560 52490 157570
rect 52730 157560 52810 157570
rect 52490 157480 52500 157560
rect 52810 157480 52820 157560
rect 52410 157380 52490 157390
rect 52730 157380 52810 157390
rect 52490 157300 52500 157380
rect 52810 157300 52820 157380
rect 52410 157200 52490 157210
rect 52730 157200 52810 157210
rect 52490 157120 52500 157200
rect 52810 157120 52820 157200
rect 52410 157020 52490 157030
rect 52730 157020 52810 157030
rect 52490 156940 52500 157020
rect 52810 156940 52820 157020
rect 52410 156840 52490 156850
rect 52730 156840 52810 156850
rect 52490 156760 52500 156840
rect 52810 156760 52820 156840
rect 52410 156660 52490 156670
rect 52730 156660 52810 156670
rect 52490 156580 52500 156660
rect 52810 156580 52820 156660
rect 52410 156480 52490 156490
rect 52730 156480 52810 156490
rect 52490 156400 52500 156480
rect 52810 156400 52820 156480
rect 52410 156300 52490 156310
rect 52730 156300 52810 156310
rect 52490 156220 52500 156300
rect 52810 156220 52820 156300
rect 52410 156120 52490 156130
rect 52730 156120 52810 156130
rect 52490 156040 52500 156120
rect 52810 156040 52820 156120
rect 52410 155940 52490 155950
rect 52730 155940 52810 155950
rect 52490 155860 52500 155940
rect 52810 155860 52820 155940
rect 52410 155760 52490 155770
rect 52730 155760 52810 155770
rect 52490 155680 52500 155760
rect 52810 155680 52820 155760
rect 52410 155580 52490 155590
rect 52730 155580 52810 155590
rect 52490 155500 52500 155580
rect 52810 155500 52820 155580
rect 52410 155400 52490 155410
rect 52730 155400 52810 155410
rect 52490 155320 52500 155400
rect 52810 155320 52820 155400
rect 52410 155220 52490 155230
rect 52730 155220 52810 155230
rect 52490 155140 52500 155220
rect 52810 155140 52820 155220
rect 52410 155040 52490 155050
rect 52730 155040 52810 155050
rect 52490 154960 52500 155040
rect 52810 154960 52820 155040
rect 52410 154860 52490 154870
rect 52730 154860 52810 154870
rect 52490 154780 52500 154860
rect 52810 154780 52820 154860
rect 52410 154680 52490 154690
rect 52730 154680 52810 154690
rect 52490 154600 52500 154680
rect 52810 154600 52820 154680
rect 52410 154500 52490 154510
rect 52730 154500 52810 154510
rect 52490 154420 52500 154500
rect 52810 154420 52820 154500
rect 52410 154320 52490 154330
rect 52730 154320 52810 154330
rect 52490 154240 52500 154320
rect 52810 154240 52820 154320
rect 52410 154140 52490 154150
rect 52730 154140 52810 154150
rect 52490 154060 52500 154140
rect 52810 154060 52820 154140
rect 52410 153960 52490 153970
rect 52730 153960 52810 153970
rect 52490 153880 52500 153960
rect 52810 153880 52820 153960
rect 52410 153780 52490 153790
rect 52730 153780 52810 153790
rect 52490 153700 52500 153780
rect 52810 153700 52820 153780
rect 52410 153600 52490 153610
rect 52730 153600 52810 153610
rect 52490 153520 52500 153600
rect 52810 153520 52820 153600
rect 52410 153420 52490 153430
rect 52730 153420 52810 153430
rect 52490 153340 52500 153420
rect 52810 153340 52820 153420
rect 52410 153240 52490 153250
rect 52730 153240 52810 153250
rect 52490 153160 52500 153240
rect 52810 153160 52820 153240
rect 52410 153060 52490 153070
rect 52730 153060 52810 153070
rect 52490 152980 52500 153060
rect 52810 152980 52820 153060
rect 52990 152900 53000 158900
rect 53010 152900 53040 158900
rect 53110 158830 53140 158900
rect 53340 158830 53370 158900
rect 53050 158820 53140 158830
rect 53200 158820 53280 158830
rect 53340 158820 53430 158830
rect 53440 158820 53470 158900
rect 53110 158650 53140 158820
rect 53280 158740 53290 158820
rect 53340 158650 53370 158820
rect 53430 158740 53470 158820
rect 53050 158640 53140 158650
rect 53200 158640 53280 158650
rect 53340 158640 53430 158650
rect 53440 158640 53470 158740
rect 53110 158470 53140 158640
rect 53280 158560 53290 158640
rect 53340 158470 53370 158640
rect 53430 158560 53470 158640
rect 53050 158460 53140 158470
rect 53200 158460 53280 158470
rect 53340 158460 53430 158470
rect 53440 158460 53470 158560
rect 53110 158290 53140 158460
rect 53280 158380 53290 158460
rect 53340 158290 53370 158460
rect 53430 158380 53470 158460
rect 53050 158280 53140 158290
rect 53200 158280 53280 158290
rect 53340 158280 53430 158290
rect 53440 158280 53470 158380
rect 53110 158110 53140 158280
rect 53280 158200 53290 158280
rect 53340 158110 53370 158280
rect 53430 158200 53470 158280
rect 53050 158100 53140 158110
rect 53200 158100 53280 158110
rect 53340 158100 53430 158110
rect 53440 158100 53470 158200
rect 53110 157930 53140 158100
rect 53280 158020 53290 158100
rect 53340 157930 53370 158100
rect 53430 158020 53470 158100
rect 53050 157920 53140 157930
rect 53200 157920 53280 157930
rect 53340 157920 53430 157930
rect 53440 157920 53470 158020
rect 53110 157750 53140 157920
rect 53280 157840 53290 157920
rect 53340 157750 53370 157920
rect 53430 157840 53470 157920
rect 53050 157740 53140 157750
rect 53200 157740 53280 157750
rect 53340 157740 53430 157750
rect 53440 157740 53470 157840
rect 53110 157570 53140 157740
rect 53280 157660 53290 157740
rect 53340 157570 53370 157740
rect 53430 157660 53470 157740
rect 53050 157560 53140 157570
rect 53200 157560 53280 157570
rect 53340 157560 53430 157570
rect 53440 157560 53470 157660
rect 53110 157390 53140 157560
rect 53280 157480 53290 157560
rect 53340 157390 53370 157560
rect 53430 157480 53470 157560
rect 53050 157380 53140 157390
rect 53200 157380 53280 157390
rect 53340 157380 53430 157390
rect 53440 157380 53470 157480
rect 53110 157210 53140 157380
rect 53280 157300 53290 157380
rect 53340 157210 53370 157380
rect 53430 157300 53470 157380
rect 53050 157200 53140 157210
rect 53200 157200 53280 157210
rect 53340 157200 53430 157210
rect 53440 157200 53470 157300
rect 53110 157030 53140 157200
rect 53280 157120 53290 157200
rect 53340 157030 53370 157200
rect 53430 157120 53470 157200
rect 53050 157020 53140 157030
rect 53200 157020 53280 157030
rect 53340 157020 53430 157030
rect 53440 157020 53470 157120
rect 53110 156850 53140 157020
rect 53280 156940 53290 157020
rect 53340 156850 53370 157020
rect 53430 156940 53470 157020
rect 53050 156840 53140 156850
rect 53200 156840 53280 156850
rect 53340 156840 53430 156850
rect 53440 156840 53470 156940
rect 53110 156670 53140 156840
rect 53280 156760 53290 156840
rect 53340 156670 53370 156840
rect 53430 156760 53470 156840
rect 53050 156660 53140 156670
rect 53200 156660 53280 156670
rect 53340 156660 53430 156670
rect 53440 156660 53470 156760
rect 53110 156490 53140 156660
rect 53280 156580 53290 156660
rect 53340 156490 53370 156660
rect 53430 156580 53470 156660
rect 53050 156480 53140 156490
rect 53200 156480 53280 156490
rect 53340 156480 53430 156490
rect 53440 156480 53470 156580
rect 53110 156310 53140 156480
rect 53280 156400 53290 156480
rect 53340 156310 53370 156480
rect 53430 156400 53470 156480
rect 53050 156300 53140 156310
rect 53200 156300 53280 156310
rect 53340 156300 53430 156310
rect 53440 156300 53470 156400
rect 53110 156130 53140 156300
rect 53280 156220 53290 156300
rect 53340 156130 53370 156300
rect 53430 156220 53470 156300
rect 53050 156120 53140 156130
rect 53200 156120 53280 156130
rect 53340 156120 53430 156130
rect 53440 156120 53470 156220
rect 53110 155950 53140 156120
rect 53280 156040 53290 156120
rect 53340 155950 53370 156120
rect 53430 156040 53470 156120
rect 53050 155940 53140 155950
rect 53200 155940 53280 155950
rect 53340 155940 53430 155950
rect 53440 155940 53470 156040
rect 53110 155770 53140 155940
rect 53280 155860 53290 155940
rect 53340 155770 53370 155940
rect 53430 155860 53470 155940
rect 53050 155760 53140 155770
rect 53200 155760 53280 155770
rect 53340 155760 53430 155770
rect 53440 155760 53470 155860
rect 53110 155590 53140 155760
rect 53280 155680 53290 155760
rect 53340 155590 53370 155760
rect 53430 155680 53470 155760
rect 53050 155580 53140 155590
rect 53200 155580 53280 155590
rect 53340 155580 53430 155590
rect 53440 155580 53470 155680
rect 53110 155410 53140 155580
rect 53280 155500 53290 155580
rect 53340 155410 53370 155580
rect 53430 155500 53470 155580
rect 53050 155400 53140 155410
rect 53200 155400 53280 155410
rect 53340 155400 53430 155410
rect 53440 155400 53470 155500
rect 53110 155230 53140 155400
rect 53280 155320 53290 155400
rect 53340 155230 53370 155400
rect 53430 155320 53470 155400
rect 53050 155220 53140 155230
rect 53200 155220 53280 155230
rect 53340 155220 53430 155230
rect 53440 155220 53470 155320
rect 53110 155050 53140 155220
rect 53280 155140 53290 155220
rect 53340 155050 53370 155220
rect 53430 155140 53470 155220
rect 53050 155040 53140 155050
rect 53200 155040 53280 155050
rect 53340 155040 53430 155050
rect 53440 155040 53470 155140
rect 53110 154870 53140 155040
rect 53280 154960 53290 155040
rect 53340 154870 53370 155040
rect 53430 154960 53470 155040
rect 53050 154860 53140 154870
rect 53200 154860 53280 154870
rect 53340 154860 53430 154870
rect 53440 154860 53470 154960
rect 53110 154690 53140 154860
rect 53280 154780 53290 154860
rect 53340 154690 53370 154860
rect 53430 154780 53470 154860
rect 53050 154680 53140 154690
rect 53200 154680 53280 154690
rect 53340 154680 53430 154690
rect 53440 154680 53470 154780
rect 53110 154510 53140 154680
rect 53280 154600 53290 154680
rect 53340 154510 53370 154680
rect 53430 154600 53470 154680
rect 53050 154500 53140 154510
rect 53200 154500 53280 154510
rect 53340 154500 53430 154510
rect 53440 154500 53470 154600
rect 53110 154330 53140 154500
rect 53280 154420 53290 154500
rect 53340 154330 53370 154500
rect 53430 154420 53470 154500
rect 53050 154320 53140 154330
rect 53200 154320 53280 154330
rect 53340 154320 53430 154330
rect 53440 154320 53470 154420
rect 53110 154150 53140 154320
rect 53280 154240 53290 154320
rect 53340 154150 53370 154320
rect 53430 154240 53470 154320
rect 53050 154140 53140 154150
rect 53200 154140 53280 154150
rect 53340 154140 53430 154150
rect 53440 154140 53470 154240
rect 53110 153970 53140 154140
rect 53280 154060 53290 154140
rect 53340 153970 53370 154140
rect 53430 154060 53470 154140
rect 53050 153960 53140 153970
rect 53200 153960 53280 153970
rect 53340 153960 53430 153970
rect 53440 153960 53470 154060
rect 53110 153790 53140 153960
rect 53280 153880 53290 153960
rect 53340 153790 53370 153960
rect 53430 153880 53470 153960
rect 53050 153780 53140 153790
rect 53200 153780 53280 153790
rect 53340 153780 53430 153790
rect 53440 153780 53470 153880
rect 53110 153610 53140 153780
rect 53280 153700 53290 153780
rect 53340 153610 53370 153780
rect 53430 153700 53470 153780
rect 53050 153600 53140 153610
rect 53200 153600 53280 153610
rect 53340 153600 53430 153610
rect 53440 153600 53470 153700
rect 53110 153430 53140 153600
rect 53280 153520 53290 153600
rect 53340 153430 53370 153600
rect 53430 153520 53470 153600
rect 53050 153420 53140 153430
rect 53200 153420 53280 153430
rect 53340 153420 53430 153430
rect 53440 153420 53470 153520
rect 53110 153250 53140 153420
rect 53280 153340 53290 153420
rect 53340 153250 53370 153420
rect 53430 153340 53470 153420
rect 53050 153240 53140 153250
rect 53200 153240 53280 153250
rect 53340 153240 53430 153250
rect 53440 153240 53470 153340
rect 53110 153070 53140 153240
rect 53280 153160 53290 153240
rect 53340 153070 53370 153240
rect 53430 153160 53470 153240
rect 53050 153060 53140 153070
rect 53200 153060 53280 153070
rect 53340 153060 53430 153070
rect 53440 153060 53470 153160
rect 53110 152900 53140 153060
rect 53280 152980 53290 153060
rect 53340 152900 53370 153060
rect 53430 152980 53470 153060
rect 53440 152900 53470 152980
rect 53570 152900 53580 158900
rect 53670 158820 53750 158830
rect 53990 158820 54070 158830
rect 53750 158740 53760 158820
rect 54070 158740 54080 158820
rect 53670 158640 53750 158650
rect 53990 158640 54070 158650
rect 53750 158560 53760 158640
rect 54070 158560 54080 158640
rect 53670 158460 53750 158470
rect 53990 158460 54070 158470
rect 53750 158380 53760 158460
rect 54070 158380 54080 158460
rect 53670 158280 53750 158290
rect 53990 158280 54070 158290
rect 53750 158200 53760 158280
rect 54070 158200 54080 158280
rect 53670 158100 53750 158110
rect 53990 158100 54070 158110
rect 53750 158020 53760 158100
rect 54070 158020 54080 158100
rect 53670 157920 53750 157930
rect 53990 157920 54070 157930
rect 53750 157840 53760 157920
rect 54070 157840 54080 157920
rect 53670 157740 53750 157750
rect 53990 157740 54070 157750
rect 53750 157660 53760 157740
rect 54070 157660 54080 157740
rect 53670 157560 53750 157570
rect 53990 157560 54070 157570
rect 53750 157480 53760 157560
rect 54070 157480 54080 157560
rect 53670 157380 53750 157390
rect 53990 157380 54070 157390
rect 53750 157300 53760 157380
rect 54070 157300 54080 157380
rect 53670 157200 53750 157210
rect 53990 157200 54070 157210
rect 53750 157120 53760 157200
rect 54070 157120 54080 157200
rect 53670 157020 53750 157030
rect 53990 157020 54070 157030
rect 53750 156940 53760 157020
rect 54070 156940 54080 157020
rect 53670 156840 53750 156850
rect 53990 156840 54070 156850
rect 53750 156760 53760 156840
rect 54070 156760 54080 156840
rect 53670 156660 53750 156670
rect 53990 156660 54070 156670
rect 53750 156580 53760 156660
rect 54070 156580 54080 156660
rect 53670 156480 53750 156490
rect 53990 156480 54070 156490
rect 53750 156400 53760 156480
rect 54070 156400 54080 156480
rect 53670 156300 53750 156310
rect 53990 156300 54070 156310
rect 53750 156220 53760 156300
rect 54070 156220 54080 156300
rect 53670 156120 53750 156130
rect 53990 156120 54070 156130
rect 53750 156040 53760 156120
rect 54070 156040 54080 156120
rect 53670 155940 53750 155950
rect 53990 155940 54070 155950
rect 53750 155860 53760 155940
rect 54070 155860 54080 155940
rect 53670 155760 53750 155770
rect 53990 155760 54070 155770
rect 53750 155680 53760 155760
rect 54070 155680 54080 155760
rect 53670 155580 53750 155590
rect 53990 155580 54070 155590
rect 53750 155500 53760 155580
rect 54070 155500 54080 155580
rect 53670 155400 53750 155410
rect 53990 155400 54070 155410
rect 53750 155320 53760 155400
rect 54070 155320 54080 155400
rect 53670 155220 53750 155230
rect 53990 155220 54070 155230
rect 53750 155140 53760 155220
rect 54070 155140 54080 155220
rect 53670 155040 53750 155050
rect 53990 155040 54070 155050
rect 53750 154960 53760 155040
rect 54070 154960 54080 155040
rect 53670 154860 53750 154870
rect 53990 154860 54070 154870
rect 53750 154780 53760 154860
rect 54070 154780 54080 154860
rect 53670 154680 53750 154690
rect 53990 154680 54070 154690
rect 53750 154600 53760 154680
rect 54070 154600 54080 154680
rect 53670 154500 53750 154510
rect 53990 154500 54070 154510
rect 53750 154420 53760 154500
rect 54070 154420 54080 154500
rect 53670 154320 53750 154330
rect 53990 154320 54070 154330
rect 53750 154240 53760 154320
rect 54070 154240 54080 154320
rect 53670 154140 53750 154150
rect 53990 154140 54070 154150
rect 53750 154060 53760 154140
rect 54070 154060 54080 154140
rect 53670 153960 53750 153970
rect 53990 153960 54070 153970
rect 53750 153880 53760 153960
rect 54070 153880 54080 153960
rect 53670 153780 53750 153790
rect 53990 153780 54070 153790
rect 53750 153700 53760 153780
rect 54070 153700 54080 153780
rect 53670 153600 53750 153610
rect 53990 153600 54070 153610
rect 53750 153520 53760 153600
rect 54070 153520 54080 153600
rect 53670 153420 53750 153430
rect 53990 153420 54070 153430
rect 53750 153340 53760 153420
rect 54070 153340 54080 153420
rect 53670 153240 53750 153250
rect 53990 153240 54070 153250
rect 53750 153160 53760 153240
rect 54070 153160 54080 153240
rect 53670 153060 53750 153070
rect 53990 153060 54070 153070
rect 53750 152980 53760 153060
rect 54070 152980 54080 153060
rect 54250 152900 54260 158900
rect 54270 152900 54300 158900
rect 54370 158830 54400 158900
rect 54600 158830 54630 158900
rect 54310 158820 54400 158830
rect 54460 158820 54540 158830
rect 54600 158820 54690 158830
rect 54700 158820 54730 158900
rect 54370 158650 54400 158820
rect 54540 158740 54550 158820
rect 54600 158650 54630 158820
rect 54690 158740 54730 158820
rect 54310 158640 54400 158650
rect 54460 158640 54540 158650
rect 54600 158640 54690 158650
rect 54700 158640 54730 158740
rect 54370 158470 54400 158640
rect 54540 158560 54550 158640
rect 54600 158470 54630 158640
rect 54690 158560 54730 158640
rect 54310 158460 54400 158470
rect 54460 158460 54540 158470
rect 54600 158460 54690 158470
rect 54700 158460 54730 158560
rect 54370 158290 54400 158460
rect 54540 158380 54550 158460
rect 54600 158290 54630 158460
rect 54690 158380 54730 158460
rect 54310 158280 54400 158290
rect 54460 158280 54540 158290
rect 54600 158280 54690 158290
rect 54700 158280 54730 158380
rect 54370 158110 54400 158280
rect 54540 158200 54550 158280
rect 54600 158110 54630 158280
rect 54690 158200 54730 158280
rect 54310 158100 54400 158110
rect 54460 158100 54540 158110
rect 54600 158100 54690 158110
rect 54700 158100 54730 158200
rect 54370 157930 54400 158100
rect 54540 158020 54550 158100
rect 54600 157930 54630 158100
rect 54690 158020 54730 158100
rect 54310 157920 54400 157930
rect 54460 157920 54540 157930
rect 54600 157920 54690 157930
rect 54700 157920 54730 158020
rect 54370 157750 54400 157920
rect 54540 157840 54550 157920
rect 54600 157750 54630 157920
rect 54690 157840 54730 157920
rect 54310 157740 54400 157750
rect 54460 157740 54540 157750
rect 54600 157740 54690 157750
rect 54700 157740 54730 157840
rect 54370 157570 54400 157740
rect 54540 157660 54550 157740
rect 54600 157570 54630 157740
rect 54690 157660 54730 157740
rect 54310 157560 54400 157570
rect 54460 157560 54540 157570
rect 54600 157560 54690 157570
rect 54700 157560 54730 157660
rect 54370 157390 54400 157560
rect 54540 157480 54550 157560
rect 54600 157390 54630 157560
rect 54690 157480 54730 157560
rect 54310 157380 54400 157390
rect 54460 157380 54540 157390
rect 54600 157380 54690 157390
rect 54700 157380 54730 157480
rect 54370 157210 54400 157380
rect 54540 157300 54550 157380
rect 54600 157210 54630 157380
rect 54690 157300 54730 157380
rect 54310 157200 54400 157210
rect 54460 157200 54540 157210
rect 54600 157200 54690 157210
rect 54700 157200 54730 157300
rect 54370 157030 54400 157200
rect 54540 157120 54550 157200
rect 54600 157030 54630 157200
rect 54690 157120 54730 157200
rect 54310 157020 54400 157030
rect 54460 157020 54540 157030
rect 54600 157020 54690 157030
rect 54700 157020 54730 157120
rect 54370 156850 54400 157020
rect 54540 156940 54550 157020
rect 54600 156850 54630 157020
rect 54690 156940 54730 157020
rect 54310 156840 54400 156850
rect 54460 156840 54540 156850
rect 54600 156840 54690 156850
rect 54700 156840 54730 156940
rect 54370 156670 54400 156840
rect 54540 156760 54550 156840
rect 54600 156670 54630 156840
rect 54690 156760 54730 156840
rect 54310 156660 54400 156670
rect 54460 156660 54540 156670
rect 54600 156660 54690 156670
rect 54700 156660 54730 156760
rect 54370 156490 54400 156660
rect 54540 156580 54550 156660
rect 54600 156490 54630 156660
rect 54690 156580 54730 156660
rect 54310 156480 54400 156490
rect 54460 156480 54540 156490
rect 54600 156480 54690 156490
rect 54700 156480 54730 156580
rect 54370 156310 54400 156480
rect 54540 156400 54550 156480
rect 54600 156310 54630 156480
rect 54690 156400 54730 156480
rect 54310 156300 54400 156310
rect 54460 156300 54540 156310
rect 54600 156300 54690 156310
rect 54700 156300 54730 156400
rect 54370 156130 54400 156300
rect 54540 156220 54550 156300
rect 54600 156130 54630 156300
rect 54690 156220 54730 156300
rect 54310 156120 54400 156130
rect 54460 156120 54540 156130
rect 54600 156120 54690 156130
rect 54700 156120 54730 156220
rect 54370 155950 54400 156120
rect 54540 156040 54550 156120
rect 54600 155950 54630 156120
rect 54690 156040 54730 156120
rect 54310 155940 54400 155950
rect 54460 155940 54540 155950
rect 54600 155940 54690 155950
rect 54700 155940 54730 156040
rect 54370 155770 54400 155940
rect 54540 155860 54550 155940
rect 54600 155770 54630 155940
rect 54690 155860 54730 155940
rect 54310 155760 54400 155770
rect 54460 155760 54540 155770
rect 54600 155760 54690 155770
rect 54700 155760 54730 155860
rect 54370 155590 54400 155760
rect 54540 155680 54550 155760
rect 54600 155590 54630 155760
rect 54690 155680 54730 155760
rect 54310 155580 54400 155590
rect 54460 155580 54540 155590
rect 54600 155580 54690 155590
rect 54700 155580 54730 155680
rect 54370 155410 54400 155580
rect 54540 155500 54550 155580
rect 54600 155410 54630 155580
rect 54690 155500 54730 155580
rect 54310 155400 54400 155410
rect 54460 155400 54540 155410
rect 54600 155400 54690 155410
rect 54700 155400 54730 155500
rect 54370 155230 54400 155400
rect 54540 155320 54550 155400
rect 54600 155230 54630 155400
rect 54690 155320 54730 155400
rect 54310 155220 54400 155230
rect 54460 155220 54540 155230
rect 54600 155220 54690 155230
rect 54700 155220 54730 155320
rect 54370 155050 54400 155220
rect 54540 155140 54550 155220
rect 54600 155050 54630 155220
rect 54690 155140 54730 155220
rect 54310 155040 54400 155050
rect 54460 155040 54540 155050
rect 54600 155040 54690 155050
rect 54700 155040 54730 155140
rect 54370 154870 54400 155040
rect 54540 154960 54550 155040
rect 54600 154870 54630 155040
rect 54690 154960 54730 155040
rect 54310 154860 54400 154870
rect 54460 154860 54540 154870
rect 54600 154860 54690 154870
rect 54700 154860 54730 154960
rect 54370 154690 54400 154860
rect 54540 154780 54550 154860
rect 54600 154690 54630 154860
rect 54690 154780 54730 154860
rect 54310 154680 54400 154690
rect 54460 154680 54540 154690
rect 54600 154680 54690 154690
rect 54700 154680 54730 154780
rect 54370 154510 54400 154680
rect 54540 154600 54550 154680
rect 54600 154510 54630 154680
rect 54690 154600 54730 154680
rect 54310 154500 54400 154510
rect 54460 154500 54540 154510
rect 54600 154500 54690 154510
rect 54700 154500 54730 154600
rect 54370 154330 54400 154500
rect 54540 154420 54550 154500
rect 54600 154330 54630 154500
rect 54690 154420 54730 154500
rect 54310 154320 54400 154330
rect 54460 154320 54540 154330
rect 54600 154320 54690 154330
rect 54700 154320 54730 154420
rect 54370 154150 54400 154320
rect 54540 154240 54550 154320
rect 54600 154150 54630 154320
rect 54690 154240 54730 154320
rect 54310 154140 54400 154150
rect 54460 154140 54540 154150
rect 54600 154140 54690 154150
rect 54700 154140 54730 154240
rect 54370 153970 54400 154140
rect 54540 154060 54550 154140
rect 54600 153970 54630 154140
rect 54690 154060 54730 154140
rect 54310 153960 54400 153970
rect 54460 153960 54540 153970
rect 54600 153960 54690 153970
rect 54700 153960 54730 154060
rect 54370 153790 54400 153960
rect 54540 153880 54550 153960
rect 54600 153790 54630 153960
rect 54690 153880 54730 153960
rect 54310 153780 54400 153790
rect 54460 153780 54540 153790
rect 54600 153780 54690 153790
rect 54700 153780 54730 153880
rect 54370 153610 54400 153780
rect 54540 153700 54550 153780
rect 54600 153610 54630 153780
rect 54690 153700 54730 153780
rect 54310 153600 54400 153610
rect 54460 153600 54540 153610
rect 54600 153600 54690 153610
rect 54700 153600 54730 153700
rect 54370 153430 54400 153600
rect 54540 153520 54550 153600
rect 54600 153430 54630 153600
rect 54690 153520 54730 153600
rect 54310 153420 54400 153430
rect 54460 153420 54540 153430
rect 54600 153420 54690 153430
rect 54700 153420 54730 153520
rect 54370 153250 54400 153420
rect 54540 153340 54550 153420
rect 54600 153250 54630 153420
rect 54690 153340 54730 153420
rect 54310 153240 54400 153250
rect 54460 153240 54540 153250
rect 54600 153240 54690 153250
rect 54700 153240 54730 153340
rect 54370 153070 54400 153240
rect 54540 153160 54550 153240
rect 54600 153070 54630 153240
rect 54690 153160 54730 153240
rect 54310 153060 54400 153070
rect 54460 153060 54540 153070
rect 54600 153060 54690 153070
rect 54700 153060 54730 153160
rect 54370 152900 54400 153060
rect 54540 152980 54550 153060
rect 54600 152900 54630 153060
rect 54690 152980 54730 153060
rect 54700 152900 54730 152980
rect 54830 152900 54840 158900
rect 54930 158820 55010 158830
rect 55250 158820 55330 158830
rect 55010 158740 55020 158820
rect 55330 158740 55340 158820
rect 54930 158640 55010 158650
rect 55250 158640 55330 158650
rect 55010 158560 55020 158640
rect 55330 158560 55340 158640
rect 54930 158460 55010 158470
rect 55250 158460 55330 158470
rect 55010 158380 55020 158460
rect 55330 158380 55340 158460
rect 54930 158280 55010 158290
rect 55250 158280 55330 158290
rect 55010 158200 55020 158280
rect 55330 158200 55340 158280
rect 54930 158100 55010 158110
rect 55250 158100 55330 158110
rect 55010 158020 55020 158100
rect 55330 158020 55340 158100
rect 54930 157920 55010 157930
rect 55250 157920 55330 157930
rect 55010 157840 55020 157920
rect 55330 157840 55340 157920
rect 54930 157740 55010 157750
rect 55250 157740 55330 157750
rect 55010 157660 55020 157740
rect 55330 157660 55340 157740
rect 54930 157560 55010 157570
rect 55250 157560 55330 157570
rect 55010 157480 55020 157560
rect 55330 157480 55340 157560
rect 54930 157380 55010 157390
rect 55250 157380 55330 157390
rect 55010 157300 55020 157380
rect 55330 157300 55340 157380
rect 54930 157200 55010 157210
rect 55250 157200 55330 157210
rect 55010 157120 55020 157200
rect 55330 157120 55340 157200
rect 54930 157020 55010 157030
rect 55250 157020 55330 157030
rect 55010 156940 55020 157020
rect 55330 156940 55340 157020
rect 54930 156840 55010 156850
rect 55250 156840 55330 156850
rect 55010 156760 55020 156840
rect 55330 156760 55340 156840
rect 54930 156660 55010 156670
rect 55250 156660 55330 156670
rect 55010 156580 55020 156660
rect 55330 156580 55340 156660
rect 54930 156480 55010 156490
rect 55250 156480 55330 156490
rect 55010 156400 55020 156480
rect 55330 156400 55340 156480
rect 54930 156300 55010 156310
rect 55250 156300 55330 156310
rect 55010 156220 55020 156300
rect 55330 156220 55340 156300
rect 54930 156120 55010 156130
rect 55250 156120 55330 156130
rect 55010 156040 55020 156120
rect 55330 156040 55340 156120
rect 54930 155940 55010 155950
rect 55250 155940 55330 155950
rect 55010 155860 55020 155940
rect 55330 155860 55340 155940
rect 54930 155760 55010 155770
rect 55250 155760 55330 155770
rect 55010 155680 55020 155760
rect 55330 155680 55340 155760
rect 54930 155580 55010 155590
rect 55250 155580 55330 155590
rect 55010 155500 55020 155580
rect 55330 155500 55340 155580
rect 54930 155400 55010 155410
rect 55250 155400 55330 155410
rect 55010 155320 55020 155400
rect 55330 155320 55340 155400
rect 54930 155220 55010 155230
rect 55250 155220 55330 155230
rect 55010 155140 55020 155220
rect 55330 155140 55340 155220
rect 54930 155040 55010 155050
rect 55250 155040 55330 155050
rect 55010 154960 55020 155040
rect 55330 154960 55340 155040
rect 54930 154860 55010 154870
rect 55250 154860 55330 154870
rect 55010 154780 55020 154860
rect 55330 154780 55340 154860
rect 54930 154680 55010 154690
rect 55250 154680 55330 154690
rect 55010 154600 55020 154680
rect 55330 154600 55340 154680
rect 54930 154500 55010 154510
rect 55250 154500 55330 154510
rect 55010 154420 55020 154500
rect 55330 154420 55340 154500
rect 54930 154320 55010 154330
rect 55250 154320 55330 154330
rect 55010 154240 55020 154320
rect 55330 154240 55340 154320
rect 54930 154140 55010 154150
rect 55250 154140 55330 154150
rect 55010 154060 55020 154140
rect 55330 154060 55340 154140
rect 54930 153960 55010 153970
rect 55250 153960 55330 153970
rect 55010 153880 55020 153960
rect 55330 153880 55340 153960
rect 54930 153780 55010 153790
rect 55250 153780 55330 153790
rect 55010 153700 55020 153780
rect 55330 153700 55340 153780
rect 54930 153600 55010 153610
rect 55250 153600 55330 153610
rect 55010 153520 55020 153600
rect 55330 153520 55340 153600
rect 54930 153420 55010 153430
rect 55250 153420 55330 153430
rect 55010 153340 55020 153420
rect 55330 153340 55340 153420
rect 54930 153240 55010 153250
rect 55250 153240 55330 153250
rect 55010 153160 55020 153240
rect 55330 153160 55340 153240
rect 54930 153060 55010 153070
rect 55250 153060 55330 153070
rect 55010 152980 55020 153060
rect 55330 152980 55340 153060
rect 55510 152900 55520 158900
rect 55530 152900 55560 158900
rect 55630 158830 55660 158900
rect 55860 158830 55890 158900
rect 55570 158820 55660 158830
rect 55720 158820 55800 158830
rect 55860 158820 55950 158830
rect 55960 158820 55990 158900
rect 55630 158650 55660 158820
rect 55800 158740 55810 158820
rect 55860 158650 55890 158820
rect 55950 158740 55990 158820
rect 55570 158640 55660 158650
rect 55720 158640 55800 158650
rect 55860 158640 55950 158650
rect 55960 158640 55990 158740
rect 55630 158470 55660 158640
rect 55800 158560 55810 158640
rect 55860 158470 55890 158640
rect 55950 158560 55990 158640
rect 55570 158460 55660 158470
rect 55720 158460 55800 158470
rect 55860 158460 55950 158470
rect 55960 158460 55990 158560
rect 55630 158290 55660 158460
rect 55800 158380 55810 158460
rect 55860 158290 55890 158460
rect 55950 158380 55990 158460
rect 55570 158280 55660 158290
rect 55720 158280 55800 158290
rect 55860 158280 55950 158290
rect 55960 158280 55990 158380
rect 55630 158110 55660 158280
rect 55800 158200 55810 158280
rect 55860 158110 55890 158280
rect 55950 158200 55990 158280
rect 55570 158100 55660 158110
rect 55720 158100 55800 158110
rect 55860 158100 55950 158110
rect 55960 158100 55990 158200
rect 55630 157930 55660 158100
rect 55800 158020 55810 158100
rect 55860 157930 55890 158100
rect 55950 158020 55990 158100
rect 55570 157920 55660 157930
rect 55720 157920 55800 157930
rect 55860 157920 55950 157930
rect 55960 157920 55990 158020
rect 55630 157750 55660 157920
rect 55800 157840 55810 157920
rect 55860 157750 55890 157920
rect 55950 157840 55990 157920
rect 55570 157740 55660 157750
rect 55720 157740 55800 157750
rect 55860 157740 55950 157750
rect 55960 157740 55990 157840
rect 55630 157570 55660 157740
rect 55800 157660 55810 157740
rect 55860 157570 55890 157740
rect 55950 157660 55990 157740
rect 55570 157560 55660 157570
rect 55720 157560 55800 157570
rect 55860 157560 55950 157570
rect 55960 157560 55990 157660
rect 55630 157390 55660 157560
rect 55800 157480 55810 157560
rect 55860 157390 55890 157560
rect 55950 157480 55990 157560
rect 55570 157380 55660 157390
rect 55720 157380 55800 157390
rect 55860 157380 55950 157390
rect 55960 157380 55990 157480
rect 55630 157210 55660 157380
rect 55800 157300 55810 157380
rect 55860 157210 55890 157380
rect 55950 157300 55990 157380
rect 55570 157200 55660 157210
rect 55720 157200 55800 157210
rect 55860 157200 55950 157210
rect 55960 157200 55990 157300
rect 55630 157030 55660 157200
rect 55800 157120 55810 157200
rect 55860 157030 55890 157200
rect 55950 157120 55990 157200
rect 55570 157020 55660 157030
rect 55720 157020 55800 157030
rect 55860 157020 55950 157030
rect 55960 157020 55990 157120
rect 55630 156850 55660 157020
rect 55800 156940 55810 157020
rect 55860 156850 55890 157020
rect 55950 156940 55990 157020
rect 55570 156840 55660 156850
rect 55720 156840 55800 156850
rect 55860 156840 55950 156850
rect 55960 156840 55990 156940
rect 55630 156670 55660 156840
rect 55800 156760 55810 156840
rect 55860 156670 55890 156840
rect 55950 156760 55990 156840
rect 55570 156660 55660 156670
rect 55720 156660 55800 156670
rect 55860 156660 55950 156670
rect 55960 156660 55990 156760
rect 55630 156490 55660 156660
rect 55800 156580 55810 156660
rect 55860 156490 55890 156660
rect 55950 156580 55990 156660
rect 55570 156480 55660 156490
rect 55720 156480 55800 156490
rect 55860 156480 55950 156490
rect 55960 156480 55990 156580
rect 55630 156310 55660 156480
rect 55800 156400 55810 156480
rect 55860 156310 55890 156480
rect 55950 156400 55990 156480
rect 55570 156300 55660 156310
rect 55720 156300 55800 156310
rect 55860 156300 55950 156310
rect 55960 156300 55990 156400
rect 55630 156130 55660 156300
rect 55800 156220 55810 156300
rect 55860 156130 55890 156300
rect 55950 156220 55990 156300
rect 55570 156120 55660 156130
rect 55720 156120 55800 156130
rect 55860 156120 55950 156130
rect 55960 156120 55990 156220
rect 55630 155950 55660 156120
rect 55800 156040 55810 156120
rect 55860 155950 55890 156120
rect 55950 156040 55990 156120
rect 55570 155940 55660 155950
rect 55720 155940 55800 155950
rect 55860 155940 55950 155950
rect 55960 155940 55990 156040
rect 55630 155770 55660 155940
rect 55800 155860 55810 155940
rect 55860 155770 55890 155940
rect 55950 155860 55990 155940
rect 55570 155760 55660 155770
rect 55720 155760 55800 155770
rect 55860 155760 55950 155770
rect 55960 155760 55990 155860
rect 55630 155590 55660 155760
rect 55800 155680 55810 155760
rect 55860 155590 55890 155760
rect 55950 155680 55990 155760
rect 55570 155580 55660 155590
rect 55720 155580 55800 155590
rect 55860 155580 55950 155590
rect 55960 155580 55990 155680
rect 55630 155410 55660 155580
rect 55800 155500 55810 155580
rect 55860 155410 55890 155580
rect 55950 155500 55990 155580
rect 55570 155400 55660 155410
rect 55720 155400 55800 155410
rect 55860 155400 55950 155410
rect 55960 155400 55990 155500
rect 55630 155230 55660 155400
rect 55800 155320 55810 155400
rect 55860 155230 55890 155400
rect 55950 155320 55990 155400
rect 55570 155220 55660 155230
rect 55720 155220 55800 155230
rect 55860 155220 55950 155230
rect 55960 155220 55990 155320
rect 55630 155050 55660 155220
rect 55800 155140 55810 155220
rect 55860 155050 55890 155220
rect 55950 155140 55990 155220
rect 55570 155040 55660 155050
rect 55720 155040 55800 155050
rect 55860 155040 55950 155050
rect 55960 155040 55990 155140
rect 55630 154870 55660 155040
rect 55800 154960 55810 155040
rect 55860 154870 55890 155040
rect 55950 154960 55990 155040
rect 55570 154860 55660 154870
rect 55720 154860 55800 154870
rect 55860 154860 55950 154870
rect 55960 154860 55990 154960
rect 55630 154690 55660 154860
rect 55800 154780 55810 154860
rect 55860 154690 55890 154860
rect 55950 154780 55990 154860
rect 55570 154680 55660 154690
rect 55720 154680 55800 154690
rect 55860 154680 55950 154690
rect 55960 154680 55990 154780
rect 55630 154510 55660 154680
rect 55800 154600 55810 154680
rect 55860 154510 55890 154680
rect 55950 154600 55990 154680
rect 55570 154500 55660 154510
rect 55720 154500 55800 154510
rect 55860 154500 55950 154510
rect 55960 154500 55990 154600
rect 55630 154330 55660 154500
rect 55800 154420 55810 154500
rect 55860 154330 55890 154500
rect 55950 154420 55990 154500
rect 55570 154320 55660 154330
rect 55720 154320 55800 154330
rect 55860 154320 55950 154330
rect 55960 154320 55990 154420
rect 55630 154150 55660 154320
rect 55800 154240 55810 154320
rect 55860 154150 55890 154320
rect 55950 154240 55990 154320
rect 55570 154140 55660 154150
rect 55720 154140 55800 154150
rect 55860 154140 55950 154150
rect 55960 154140 55990 154240
rect 55630 153970 55660 154140
rect 55800 154060 55810 154140
rect 55860 153970 55890 154140
rect 55950 154060 55990 154140
rect 55570 153960 55660 153970
rect 55720 153960 55800 153970
rect 55860 153960 55950 153970
rect 55960 153960 55990 154060
rect 55630 153790 55660 153960
rect 55800 153880 55810 153960
rect 55860 153790 55890 153960
rect 55950 153880 55990 153960
rect 55570 153780 55660 153790
rect 55720 153780 55800 153790
rect 55860 153780 55950 153790
rect 55960 153780 55990 153880
rect 55630 153610 55660 153780
rect 55800 153700 55810 153780
rect 55860 153610 55890 153780
rect 55950 153700 55990 153780
rect 55570 153600 55660 153610
rect 55720 153600 55800 153610
rect 55860 153600 55950 153610
rect 55960 153600 55990 153700
rect 55630 153430 55660 153600
rect 55800 153520 55810 153600
rect 55860 153430 55890 153600
rect 55950 153520 55990 153600
rect 55570 153420 55660 153430
rect 55720 153420 55800 153430
rect 55860 153420 55950 153430
rect 55960 153420 55990 153520
rect 55630 153250 55660 153420
rect 55800 153340 55810 153420
rect 55860 153250 55890 153420
rect 55950 153340 55990 153420
rect 55570 153240 55660 153250
rect 55720 153240 55800 153250
rect 55860 153240 55950 153250
rect 55960 153240 55990 153340
rect 55630 153070 55660 153240
rect 55800 153160 55810 153240
rect 55860 153070 55890 153240
rect 55950 153160 55990 153240
rect 55570 153060 55660 153070
rect 55720 153060 55800 153070
rect 55860 153060 55950 153070
rect 55960 153060 55990 153160
rect 55630 152900 55660 153060
rect 55800 152980 55810 153060
rect 55860 152900 55890 153060
rect 55950 152980 55990 153060
rect 55960 152900 55990 152980
rect 56090 152900 56100 158900
rect 56190 158820 56270 158830
rect 56510 158820 56590 158830
rect 56270 158740 56280 158820
rect 56590 158740 56600 158820
rect 56190 158640 56270 158650
rect 56510 158640 56590 158650
rect 56270 158560 56280 158640
rect 56590 158560 56600 158640
rect 56190 158460 56270 158470
rect 56510 158460 56590 158470
rect 56270 158380 56280 158460
rect 56590 158380 56600 158460
rect 56190 158280 56270 158290
rect 56510 158280 56590 158290
rect 56270 158200 56280 158280
rect 56590 158200 56600 158280
rect 56190 158100 56270 158110
rect 56510 158100 56590 158110
rect 56270 158020 56280 158100
rect 56590 158020 56600 158100
rect 56190 157920 56270 157930
rect 56510 157920 56590 157930
rect 56270 157840 56280 157920
rect 56590 157840 56600 157920
rect 56190 157740 56270 157750
rect 56510 157740 56590 157750
rect 56270 157660 56280 157740
rect 56590 157660 56600 157740
rect 56190 157560 56270 157570
rect 56510 157560 56590 157570
rect 56270 157480 56280 157560
rect 56590 157480 56600 157560
rect 56190 157380 56270 157390
rect 56510 157380 56590 157390
rect 56270 157300 56280 157380
rect 56590 157300 56600 157380
rect 56190 157200 56270 157210
rect 56510 157200 56590 157210
rect 56270 157120 56280 157200
rect 56590 157120 56600 157200
rect 56190 157020 56270 157030
rect 56510 157020 56590 157030
rect 56270 156940 56280 157020
rect 56590 156940 56600 157020
rect 56190 156840 56270 156850
rect 56510 156840 56590 156850
rect 56270 156760 56280 156840
rect 56590 156760 56600 156840
rect 56190 156660 56270 156670
rect 56510 156660 56590 156670
rect 56270 156580 56280 156660
rect 56590 156580 56600 156660
rect 56190 156480 56270 156490
rect 56510 156480 56590 156490
rect 56270 156400 56280 156480
rect 56590 156400 56600 156480
rect 56190 156300 56270 156310
rect 56510 156300 56590 156310
rect 56270 156220 56280 156300
rect 56590 156220 56600 156300
rect 56190 156120 56270 156130
rect 56510 156120 56590 156130
rect 56270 156040 56280 156120
rect 56590 156040 56600 156120
rect 56190 155940 56270 155950
rect 56510 155940 56590 155950
rect 56270 155860 56280 155940
rect 56590 155860 56600 155940
rect 56190 155760 56270 155770
rect 56510 155760 56590 155770
rect 56270 155680 56280 155760
rect 56590 155680 56600 155760
rect 56190 155580 56270 155590
rect 56510 155580 56590 155590
rect 56270 155500 56280 155580
rect 56590 155500 56600 155580
rect 56190 155400 56270 155410
rect 56510 155400 56590 155410
rect 56270 155320 56280 155400
rect 56590 155320 56600 155400
rect 56190 155220 56270 155230
rect 56510 155220 56590 155230
rect 56270 155140 56280 155220
rect 56590 155140 56600 155220
rect 56190 155040 56270 155050
rect 56510 155040 56590 155050
rect 56270 154960 56280 155040
rect 56590 154960 56600 155040
rect 56190 154860 56270 154870
rect 56510 154860 56590 154870
rect 56270 154780 56280 154860
rect 56590 154780 56600 154860
rect 56190 154680 56270 154690
rect 56510 154680 56590 154690
rect 56270 154600 56280 154680
rect 56590 154600 56600 154680
rect 56190 154500 56270 154510
rect 56510 154500 56590 154510
rect 56270 154420 56280 154500
rect 56590 154420 56600 154500
rect 56190 154320 56270 154330
rect 56510 154320 56590 154330
rect 56270 154240 56280 154320
rect 56590 154240 56600 154320
rect 56190 154140 56270 154150
rect 56510 154140 56590 154150
rect 56270 154060 56280 154140
rect 56590 154060 56600 154140
rect 56190 153960 56270 153970
rect 56510 153960 56590 153970
rect 56270 153880 56280 153960
rect 56590 153880 56600 153960
rect 56190 153780 56270 153790
rect 56510 153780 56590 153790
rect 56270 153700 56280 153780
rect 56590 153700 56600 153780
rect 56190 153600 56270 153610
rect 56510 153600 56590 153610
rect 56270 153520 56280 153600
rect 56590 153520 56600 153600
rect 56190 153420 56270 153430
rect 56510 153420 56590 153430
rect 56270 153340 56280 153420
rect 56590 153340 56600 153420
rect 56190 153240 56270 153250
rect 56510 153240 56590 153250
rect 56270 153160 56280 153240
rect 56590 153160 56600 153240
rect 56190 153060 56270 153070
rect 56510 153060 56590 153070
rect 56270 152980 56280 153060
rect 56590 152980 56600 153060
rect 56770 152900 56780 158900
rect 56790 152900 56820 158900
rect 56890 158830 56920 158900
rect 57120 158830 57150 158900
rect 56830 158820 56920 158830
rect 56980 158820 57060 158830
rect 57120 158820 57210 158830
rect 57220 158820 57250 158900
rect 56890 158650 56920 158820
rect 57060 158740 57070 158820
rect 57120 158650 57150 158820
rect 57210 158740 57250 158820
rect 56830 158640 56920 158650
rect 56980 158640 57060 158650
rect 57120 158640 57210 158650
rect 57220 158640 57250 158740
rect 56890 158470 56920 158640
rect 57060 158560 57070 158640
rect 57120 158470 57150 158640
rect 57210 158560 57250 158640
rect 56830 158460 56920 158470
rect 56980 158460 57060 158470
rect 57120 158460 57210 158470
rect 57220 158460 57250 158560
rect 56890 158290 56920 158460
rect 57060 158380 57070 158460
rect 57120 158290 57150 158460
rect 57210 158380 57250 158460
rect 56830 158280 56920 158290
rect 56980 158280 57060 158290
rect 57120 158280 57210 158290
rect 57220 158280 57250 158380
rect 56890 158110 56920 158280
rect 57060 158200 57070 158280
rect 57120 158110 57150 158280
rect 57210 158200 57250 158280
rect 56830 158100 56920 158110
rect 56980 158100 57060 158110
rect 57120 158100 57210 158110
rect 57220 158100 57250 158200
rect 56890 157930 56920 158100
rect 57060 158020 57070 158100
rect 57120 157930 57150 158100
rect 57210 158020 57250 158100
rect 56830 157920 56920 157930
rect 56980 157920 57060 157930
rect 57120 157920 57210 157930
rect 57220 157920 57250 158020
rect 56890 157750 56920 157920
rect 57060 157840 57070 157920
rect 57120 157750 57150 157920
rect 57210 157840 57250 157920
rect 56830 157740 56920 157750
rect 56980 157740 57060 157750
rect 57120 157740 57210 157750
rect 57220 157740 57250 157840
rect 56890 157570 56920 157740
rect 57060 157660 57070 157740
rect 57120 157570 57150 157740
rect 57210 157660 57250 157740
rect 56830 157560 56920 157570
rect 56980 157560 57060 157570
rect 57120 157560 57210 157570
rect 57220 157560 57250 157660
rect 56890 157390 56920 157560
rect 57060 157480 57070 157560
rect 57120 157390 57150 157560
rect 57210 157480 57250 157560
rect 56830 157380 56920 157390
rect 56980 157380 57060 157390
rect 57120 157380 57210 157390
rect 57220 157380 57250 157480
rect 56890 157210 56920 157380
rect 57060 157300 57070 157380
rect 57120 157210 57150 157380
rect 57210 157300 57250 157380
rect 56830 157200 56920 157210
rect 56980 157200 57060 157210
rect 57120 157200 57210 157210
rect 57220 157200 57250 157300
rect 56890 157030 56920 157200
rect 57060 157120 57070 157200
rect 57120 157030 57150 157200
rect 57210 157120 57250 157200
rect 56830 157020 56920 157030
rect 56980 157020 57060 157030
rect 57120 157020 57210 157030
rect 57220 157020 57250 157120
rect 56890 156850 56920 157020
rect 57060 156940 57070 157020
rect 57120 156850 57150 157020
rect 57210 156940 57250 157020
rect 56830 156840 56920 156850
rect 56980 156840 57060 156850
rect 57120 156840 57210 156850
rect 57220 156840 57250 156940
rect 56890 156670 56920 156840
rect 57060 156760 57070 156840
rect 57120 156670 57150 156840
rect 57210 156760 57250 156840
rect 56830 156660 56920 156670
rect 56980 156660 57060 156670
rect 57120 156660 57210 156670
rect 57220 156660 57250 156760
rect 56890 156490 56920 156660
rect 57060 156580 57070 156660
rect 57120 156490 57150 156660
rect 57210 156580 57250 156660
rect 56830 156480 56920 156490
rect 56980 156480 57060 156490
rect 57120 156480 57210 156490
rect 57220 156480 57250 156580
rect 56890 156310 56920 156480
rect 57060 156400 57070 156480
rect 57120 156310 57150 156480
rect 57210 156400 57250 156480
rect 56830 156300 56920 156310
rect 56980 156300 57060 156310
rect 57120 156300 57210 156310
rect 57220 156300 57250 156400
rect 56890 156130 56920 156300
rect 57060 156220 57070 156300
rect 57120 156130 57150 156300
rect 57210 156220 57250 156300
rect 56830 156120 56920 156130
rect 56980 156120 57060 156130
rect 57120 156120 57210 156130
rect 57220 156120 57250 156220
rect 56890 155950 56920 156120
rect 57060 156040 57070 156120
rect 57120 155950 57150 156120
rect 57210 156040 57250 156120
rect 56830 155940 56920 155950
rect 56980 155940 57060 155950
rect 57120 155940 57210 155950
rect 57220 155940 57250 156040
rect 56890 155770 56920 155940
rect 57060 155860 57070 155940
rect 57120 155770 57150 155940
rect 57210 155860 57250 155940
rect 56830 155760 56920 155770
rect 56980 155760 57060 155770
rect 57120 155760 57210 155770
rect 57220 155760 57250 155860
rect 56890 155590 56920 155760
rect 57060 155680 57070 155760
rect 57120 155590 57150 155760
rect 57210 155680 57250 155760
rect 56830 155580 56920 155590
rect 56980 155580 57060 155590
rect 57120 155580 57210 155590
rect 57220 155580 57250 155680
rect 56890 155410 56920 155580
rect 57060 155500 57070 155580
rect 57120 155410 57150 155580
rect 57210 155500 57250 155580
rect 56830 155400 56920 155410
rect 56980 155400 57060 155410
rect 57120 155400 57210 155410
rect 57220 155400 57250 155500
rect 56890 155230 56920 155400
rect 57060 155320 57070 155400
rect 57120 155230 57150 155400
rect 57210 155320 57250 155400
rect 56830 155220 56920 155230
rect 56980 155220 57060 155230
rect 57120 155220 57210 155230
rect 57220 155220 57250 155320
rect 56890 155050 56920 155220
rect 57060 155140 57070 155220
rect 57120 155050 57150 155220
rect 57210 155140 57250 155220
rect 56830 155040 56920 155050
rect 56980 155040 57060 155050
rect 57120 155040 57210 155050
rect 57220 155040 57250 155140
rect 56890 154870 56920 155040
rect 57060 154960 57070 155040
rect 57120 154870 57150 155040
rect 57210 154960 57250 155040
rect 56830 154860 56920 154870
rect 56980 154860 57060 154870
rect 57120 154860 57210 154870
rect 57220 154860 57250 154960
rect 56890 154690 56920 154860
rect 57060 154780 57070 154860
rect 57120 154690 57150 154860
rect 57210 154780 57250 154860
rect 56830 154680 56920 154690
rect 56980 154680 57060 154690
rect 57120 154680 57210 154690
rect 57220 154680 57250 154780
rect 56890 154510 56920 154680
rect 57060 154600 57070 154680
rect 57120 154510 57150 154680
rect 57210 154600 57250 154680
rect 56830 154500 56920 154510
rect 56980 154500 57060 154510
rect 57120 154500 57210 154510
rect 57220 154500 57250 154600
rect 56890 154330 56920 154500
rect 57060 154420 57070 154500
rect 57120 154330 57150 154500
rect 57210 154420 57250 154500
rect 56830 154320 56920 154330
rect 56980 154320 57060 154330
rect 57120 154320 57210 154330
rect 57220 154320 57250 154420
rect 56890 154150 56920 154320
rect 57060 154240 57070 154320
rect 57120 154150 57150 154320
rect 57210 154240 57250 154320
rect 56830 154140 56920 154150
rect 56980 154140 57060 154150
rect 57120 154140 57210 154150
rect 57220 154140 57250 154240
rect 56890 153970 56920 154140
rect 57060 154060 57070 154140
rect 57120 153970 57150 154140
rect 57210 154060 57250 154140
rect 56830 153960 56920 153970
rect 56980 153960 57060 153970
rect 57120 153960 57210 153970
rect 57220 153960 57250 154060
rect 56890 153790 56920 153960
rect 57060 153880 57070 153960
rect 57120 153790 57150 153960
rect 57210 153880 57250 153960
rect 56830 153780 56920 153790
rect 56980 153780 57060 153790
rect 57120 153780 57210 153790
rect 57220 153780 57250 153880
rect 56890 153610 56920 153780
rect 57060 153700 57070 153780
rect 57120 153610 57150 153780
rect 57210 153700 57250 153780
rect 56830 153600 56920 153610
rect 56980 153600 57060 153610
rect 57120 153600 57210 153610
rect 57220 153600 57250 153700
rect 56890 153430 56920 153600
rect 57060 153520 57070 153600
rect 57120 153430 57150 153600
rect 57210 153520 57250 153600
rect 56830 153420 56920 153430
rect 56980 153420 57060 153430
rect 57120 153420 57210 153430
rect 57220 153420 57250 153520
rect 56890 153250 56920 153420
rect 57060 153340 57070 153420
rect 57120 153250 57150 153420
rect 57210 153340 57250 153420
rect 56830 153240 56920 153250
rect 56980 153240 57060 153250
rect 57120 153240 57210 153250
rect 57220 153240 57250 153340
rect 56890 153070 56920 153240
rect 57060 153160 57070 153240
rect 57120 153070 57150 153240
rect 57210 153160 57250 153240
rect 56830 153060 56920 153070
rect 56980 153060 57060 153070
rect 57120 153060 57210 153070
rect 57220 153060 57250 153160
rect 56890 152900 56920 153060
rect 57060 152980 57070 153060
rect 57120 152900 57150 153060
rect 57210 152980 57250 153060
rect 57220 152900 57250 152980
rect 57350 152900 57360 158900
rect 57450 158820 57530 158830
rect 57770 158820 57850 158830
rect 57530 158740 57540 158820
rect 57850 158740 57860 158820
rect 57450 158640 57530 158650
rect 57770 158640 57850 158650
rect 57530 158560 57540 158640
rect 57850 158560 57860 158640
rect 57450 158460 57530 158470
rect 57770 158460 57850 158470
rect 57530 158380 57540 158460
rect 57850 158380 57860 158460
rect 57450 158280 57530 158290
rect 57770 158280 57850 158290
rect 57530 158200 57540 158280
rect 57850 158200 57860 158280
rect 57450 158100 57530 158110
rect 57770 158100 57850 158110
rect 57530 158020 57540 158100
rect 57850 158020 57860 158100
rect 57450 157920 57530 157930
rect 57770 157920 57850 157930
rect 57530 157840 57540 157920
rect 57850 157840 57860 157920
rect 57450 157740 57530 157750
rect 57770 157740 57850 157750
rect 57530 157660 57540 157740
rect 57850 157660 57860 157740
rect 57450 157560 57530 157570
rect 57770 157560 57850 157570
rect 57530 157480 57540 157560
rect 57850 157480 57860 157560
rect 57450 157380 57530 157390
rect 57770 157380 57850 157390
rect 57530 157300 57540 157380
rect 57850 157300 57860 157380
rect 57450 157200 57530 157210
rect 57770 157200 57850 157210
rect 57530 157120 57540 157200
rect 57850 157120 57860 157200
rect 57450 157020 57530 157030
rect 57770 157020 57850 157030
rect 57530 156940 57540 157020
rect 57850 156940 57860 157020
rect 57450 156840 57530 156850
rect 57770 156840 57850 156850
rect 57530 156760 57540 156840
rect 57850 156760 57860 156840
rect 57450 156660 57530 156670
rect 57770 156660 57850 156670
rect 57530 156580 57540 156660
rect 57850 156580 57860 156660
rect 57450 156480 57530 156490
rect 57770 156480 57850 156490
rect 57530 156400 57540 156480
rect 57850 156400 57860 156480
rect 57450 156300 57530 156310
rect 57770 156300 57850 156310
rect 57530 156220 57540 156300
rect 57850 156220 57860 156300
rect 57450 156120 57530 156130
rect 57770 156120 57850 156130
rect 57530 156040 57540 156120
rect 57850 156040 57860 156120
rect 57450 155940 57530 155950
rect 57770 155940 57850 155950
rect 57530 155860 57540 155940
rect 57850 155860 57860 155940
rect 57450 155760 57530 155770
rect 57770 155760 57850 155770
rect 57530 155680 57540 155760
rect 57850 155680 57860 155760
rect 57450 155580 57530 155590
rect 57770 155580 57850 155590
rect 57530 155500 57540 155580
rect 57850 155500 57860 155580
rect 57450 155400 57530 155410
rect 57770 155400 57850 155410
rect 57530 155320 57540 155400
rect 57850 155320 57860 155400
rect 57450 155220 57530 155230
rect 57770 155220 57850 155230
rect 57530 155140 57540 155220
rect 57850 155140 57860 155220
rect 57450 155040 57530 155050
rect 57770 155040 57850 155050
rect 57530 154960 57540 155040
rect 57850 154960 57860 155040
rect 57450 154860 57530 154870
rect 57770 154860 57850 154870
rect 57530 154780 57540 154860
rect 57850 154780 57860 154860
rect 57450 154680 57530 154690
rect 57770 154680 57850 154690
rect 57530 154600 57540 154680
rect 57850 154600 57860 154680
rect 57450 154500 57530 154510
rect 57770 154500 57850 154510
rect 57530 154420 57540 154500
rect 57850 154420 57860 154500
rect 57450 154320 57530 154330
rect 57770 154320 57850 154330
rect 57530 154240 57540 154320
rect 57850 154240 57860 154320
rect 57450 154140 57530 154150
rect 57770 154140 57850 154150
rect 57530 154060 57540 154140
rect 57850 154060 57860 154140
rect 57450 153960 57530 153970
rect 57770 153960 57850 153970
rect 57530 153880 57540 153960
rect 57850 153880 57860 153960
rect 57450 153780 57530 153790
rect 57770 153780 57850 153790
rect 57530 153700 57540 153780
rect 57850 153700 57860 153780
rect 57450 153600 57530 153610
rect 57770 153600 57850 153610
rect 57530 153520 57540 153600
rect 57850 153520 57860 153600
rect 57450 153420 57530 153430
rect 57770 153420 57850 153430
rect 57530 153340 57540 153420
rect 57850 153340 57860 153420
rect 57450 153240 57530 153250
rect 57770 153240 57850 153250
rect 57530 153160 57540 153240
rect 57850 153160 57860 153240
rect 57450 153060 57530 153070
rect 57770 153060 57850 153070
rect 57530 152980 57540 153060
rect 57850 152980 57860 153060
rect 58030 152900 58040 158900
rect 58050 152900 58080 158900
rect 58150 158830 58180 158900
rect 58380 158830 58410 158900
rect 58090 158820 58180 158830
rect 58240 158820 58320 158830
rect 58380 158820 58470 158830
rect 58480 158820 58510 158900
rect 58150 158650 58180 158820
rect 58320 158740 58330 158820
rect 58380 158650 58410 158820
rect 58470 158740 58510 158820
rect 58090 158640 58180 158650
rect 58240 158640 58320 158650
rect 58380 158640 58470 158650
rect 58480 158640 58510 158740
rect 58150 158470 58180 158640
rect 58320 158560 58330 158640
rect 58380 158470 58410 158640
rect 58470 158560 58510 158640
rect 58090 158460 58180 158470
rect 58240 158460 58320 158470
rect 58380 158460 58470 158470
rect 58480 158460 58510 158560
rect 58150 158290 58180 158460
rect 58320 158380 58330 158460
rect 58380 158290 58410 158460
rect 58470 158380 58510 158460
rect 58090 158280 58180 158290
rect 58240 158280 58320 158290
rect 58380 158280 58470 158290
rect 58480 158280 58510 158380
rect 58150 158110 58180 158280
rect 58320 158200 58330 158280
rect 58380 158110 58410 158280
rect 58470 158200 58510 158280
rect 58090 158100 58180 158110
rect 58240 158100 58320 158110
rect 58380 158100 58470 158110
rect 58480 158100 58510 158200
rect 58150 157930 58180 158100
rect 58320 158020 58330 158100
rect 58380 157930 58410 158100
rect 58470 158020 58510 158100
rect 58090 157920 58180 157930
rect 58240 157920 58320 157930
rect 58380 157920 58470 157930
rect 58480 157920 58510 158020
rect 58150 157750 58180 157920
rect 58320 157840 58330 157920
rect 58380 157750 58410 157920
rect 58470 157840 58510 157920
rect 58090 157740 58180 157750
rect 58240 157740 58320 157750
rect 58380 157740 58470 157750
rect 58480 157740 58510 157840
rect 58150 157570 58180 157740
rect 58320 157660 58330 157740
rect 58380 157570 58410 157740
rect 58470 157660 58510 157740
rect 58090 157560 58180 157570
rect 58240 157560 58320 157570
rect 58380 157560 58470 157570
rect 58480 157560 58510 157660
rect 58150 157390 58180 157560
rect 58320 157480 58330 157560
rect 58380 157390 58410 157560
rect 58470 157480 58510 157560
rect 58090 157380 58180 157390
rect 58240 157380 58320 157390
rect 58380 157380 58470 157390
rect 58480 157380 58510 157480
rect 58150 157210 58180 157380
rect 58320 157300 58330 157380
rect 58380 157210 58410 157380
rect 58470 157300 58510 157380
rect 58090 157200 58180 157210
rect 58240 157200 58320 157210
rect 58380 157200 58470 157210
rect 58480 157200 58510 157300
rect 58150 157030 58180 157200
rect 58320 157120 58330 157200
rect 58380 157030 58410 157200
rect 58470 157120 58510 157200
rect 58090 157020 58180 157030
rect 58240 157020 58320 157030
rect 58380 157020 58470 157030
rect 58480 157020 58510 157120
rect 58150 156850 58180 157020
rect 58320 156940 58330 157020
rect 58380 156850 58410 157020
rect 58470 156940 58510 157020
rect 58090 156840 58180 156850
rect 58240 156840 58320 156850
rect 58380 156840 58470 156850
rect 58480 156840 58510 156940
rect 58150 156670 58180 156840
rect 58320 156760 58330 156840
rect 58380 156670 58410 156840
rect 58470 156760 58510 156840
rect 58090 156660 58180 156670
rect 58240 156660 58320 156670
rect 58380 156660 58470 156670
rect 58480 156660 58510 156760
rect 58150 156490 58180 156660
rect 58320 156580 58330 156660
rect 58380 156490 58410 156660
rect 58470 156580 58510 156660
rect 58090 156480 58180 156490
rect 58240 156480 58320 156490
rect 58380 156480 58470 156490
rect 58480 156480 58510 156580
rect 58150 156310 58180 156480
rect 58320 156400 58330 156480
rect 58380 156310 58410 156480
rect 58470 156400 58510 156480
rect 58090 156300 58180 156310
rect 58240 156300 58320 156310
rect 58380 156300 58470 156310
rect 58480 156300 58510 156400
rect 58150 156130 58180 156300
rect 58320 156220 58330 156300
rect 58380 156130 58410 156300
rect 58470 156220 58510 156300
rect 58090 156120 58180 156130
rect 58240 156120 58320 156130
rect 58380 156120 58470 156130
rect 58480 156120 58510 156220
rect 58150 155950 58180 156120
rect 58320 156040 58330 156120
rect 58380 155950 58410 156120
rect 58470 156040 58510 156120
rect 58090 155940 58180 155950
rect 58240 155940 58320 155950
rect 58380 155940 58470 155950
rect 58480 155940 58510 156040
rect 58150 155770 58180 155940
rect 58320 155860 58330 155940
rect 58380 155770 58410 155940
rect 58470 155860 58510 155940
rect 58090 155760 58180 155770
rect 58240 155760 58320 155770
rect 58380 155760 58470 155770
rect 58480 155760 58510 155860
rect 58150 155590 58180 155760
rect 58320 155680 58330 155760
rect 58380 155590 58410 155760
rect 58470 155680 58510 155760
rect 58090 155580 58180 155590
rect 58240 155580 58320 155590
rect 58380 155580 58470 155590
rect 58480 155580 58510 155680
rect 58150 155410 58180 155580
rect 58320 155500 58330 155580
rect 58380 155410 58410 155580
rect 58470 155500 58510 155580
rect 58090 155400 58180 155410
rect 58240 155400 58320 155410
rect 58380 155400 58470 155410
rect 58480 155400 58510 155500
rect 58150 155230 58180 155400
rect 58320 155320 58330 155400
rect 58380 155230 58410 155400
rect 58470 155320 58510 155400
rect 58090 155220 58180 155230
rect 58240 155220 58320 155230
rect 58380 155220 58470 155230
rect 58480 155220 58510 155320
rect 58150 155050 58180 155220
rect 58320 155140 58330 155220
rect 58380 155050 58410 155220
rect 58470 155140 58510 155220
rect 58090 155040 58180 155050
rect 58240 155040 58320 155050
rect 58380 155040 58470 155050
rect 58480 155040 58510 155140
rect 58150 154870 58180 155040
rect 58320 154960 58330 155040
rect 58380 154870 58410 155040
rect 58470 154960 58510 155040
rect 58090 154860 58180 154870
rect 58240 154860 58320 154870
rect 58380 154860 58470 154870
rect 58480 154860 58510 154960
rect 58150 154690 58180 154860
rect 58320 154780 58330 154860
rect 58380 154690 58410 154860
rect 58470 154780 58510 154860
rect 58090 154680 58180 154690
rect 58240 154680 58320 154690
rect 58380 154680 58470 154690
rect 58480 154680 58510 154780
rect 58150 154510 58180 154680
rect 58320 154600 58330 154680
rect 58380 154510 58410 154680
rect 58470 154600 58510 154680
rect 58090 154500 58180 154510
rect 58240 154500 58320 154510
rect 58380 154500 58470 154510
rect 58480 154500 58510 154600
rect 58150 154330 58180 154500
rect 58320 154420 58330 154500
rect 58380 154330 58410 154500
rect 58470 154420 58510 154500
rect 58090 154320 58180 154330
rect 58240 154320 58320 154330
rect 58380 154320 58470 154330
rect 58480 154320 58510 154420
rect 58150 154150 58180 154320
rect 58320 154240 58330 154320
rect 58380 154150 58410 154320
rect 58470 154240 58510 154320
rect 58090 154140 58180 154150
rect 58240 154140 58320 154150
rect 58380 154140 58470 154150
rect 58480 154140 58510 154240
rect 58150 153970 58180 154140
rect 58320 154060 58330 154140
rect 58380 153970 58410 154140
rect 58470 154060 58510 154140
rect 58090 153960 58180 153970
rect 58240 153960 58320 153970
rect 58380 153960 58470 153970
rect 58480 153960 58510 154060
rect 58150 153790 58180 153960
rect 58320 153880 58330 153960
rect 58380 153790 58410 153960
rect 58470 153880 58510 153960
rect 58090 153780 58180 153790
rect 58240 153780 58320 153790
rect 58380 153780 58470 153790
rect 58480 153780 58510 153880
rect 58150 153610 58180 153780
rect 58320 153700 58330 153780
rect 58380 153610 58410 153780
rect 58470 153700 58510 153780
rect 58090 153600 58180 153610
rect 58240 153600 58320 153610
rect 58380 153600 58470 153610
rect 58480 153600 58510 153700
rect 58150 153430 58180 153600
rect 58320 153520 58330 153600
rect 58380 153430 58410 153600
rect 58470 153520 58510 153600
rect 58090 153420 58180 153430
rect 58240 153420 58320 153430
rect 58380 153420 58470 153430
rect 58480 153420 58510 153520
rect 58150 153250 58180 153420
rect 58320 153340 58330 153420
rect 58380 153250 58410 153420
rect 58470 153340 58510 153420
rect 58090 153240 58180 153250
rect 58240 153240 58320 153250
rect 58380 153240 58470 153250
rect 58480 153240 58510 153340
rect 58150 153070 58180 153240
rect 58320 153160 58330 153240
rect 58380 153070 58410 153240
rect 58470 153160 58510 153240
rect 58090 153060 58180 153070
rect 58240 153060 58320 153070
rect 58380 153060 58470 153070
rect 58480 153060 58510 153160
rect 58150 152900 58180 153060
rect 58320 152980 58330 153060
rect 58380 152900 58410 153060
rect 58470 152980 58510 153060
rect 58480 152900 58510 152980
rect 58610 152900 58620 158900
rect 58710 158820 58790 158830
rect 59030 158820 59110 158830
rect 58790 158740 58800 158820
rect 59110 158740 59120 158820
rect 58710 158640 58790 158650
rect 59030 158640 59110 158650
rect 58790 158560 58800 158640
rect 59110 158560 59120 158640
rect 58710 158460 58790 158470
rect 59030 158460 59110 158470
rect 58790 158380 58800 158460
rect 59110 158380 59120 158460
rect 58710 158280 58790 158290
rect 59030 158280 59110 158290
rect 58790 158200 58800 158280
rect 59110 158200 59120 158280
rect 58710 158100 58790 158110
rect 59030 158100 59110 158110
rect 58790 158020 58800 158100
rect 59110 158020 59120 158100
rect 58710 157920 58790 157930
rect 59030 157920 59110 157930
rect 58790 157840 58800 157920
rect 59110 157840 59120 157920
rect 58710 157740 58790 157750
rect 59030 157740 59110 157750
rect 58790 157660 58800 157740
rect 59110 157660 59120 157740
rect 58710 157560 58790 157570
rect 59030 157560 59110 157570
rect 58790 157480 58800 157560
rect 59110 157480 59120 157560
rect 58710 157380 58790 157390
rect 59030 157380 59110 157390
rect 58790 157300 58800 157380
rect 59110 157300 59120 157380
rect 58710 157200 58790 157210
rect 59030 157200 59110 157210
rect 58790 157120 58800 157200
rect 59110 157120 59120 157200
rect 58710 157020 58790 157030
rect 59030 157020 59110 157030
rect 58790 156940 58800 157020
rect 59110 156940 59120 157020
rect 58710 156840 58790 156850
rect 59030 156840 59110 156850
rect 58790 156760 58800 156840
rect 59110 156760 59120 156840
rect 58710 156660 58790 156670
rect 59030 156660 59110 156670
rect 58790 156580 58800 156660
rect 59110 156580 59120 156660
rect 58710 156480 58790 156490
rect 59030 156480 59110 156490
rect 58790 156400 58800 156480
rect 59110 156400 59120 156480
rect 58710 156300 58790 156310
rect 59030 156300 59110 156310
rect 58790 156220 58800 156300
rect 59110 156220 59120 156300
rect 58710 156120 58790 156130
rect 59030 156120 59110 156130
rect 58790 156040 58800 156120
rect 59110 156040 59120 156120
rect 58710 155940 58790 155950
rect 59030 155940 59110 155950
rect 58790 155860 58800 155940
rect 59110 155860 59120 155940
rect 58710 155760 58790 155770
rect 59030 155760 59110 155770
rect 58790 155680 58800 155760
rect 59110 155680 59120 155760
rect 58710 155580 58790 155590
rect 59030 155580 59110 155590
rect 58790 155500 58800 155580
rect 59110 155500 59120 155580
rect 58710 155400 58790 155410
rect 59030 155400 59110 155410
rect 58790 155320 58800 155400
rect 59110 155320 59120 155400
rect 58710 155220 58790 155230
rect 59030 155220 59110 155230
rect 58790 155140 58800 155220
rect 59110 155140 59120 155220
rect 58710 155040 58790 155050
rect 59030 155040 59110 155050
rect 58790 154960 58800 155040
rect 59110 154960 59120 155040
rect 58710 154860 58790 154870
rect 59030 154860 59110 154870
rect 58790 154780 58800 154860
rect 59110 154780 59120 154860
rect 58710 154680 58790 154690
rect 59030 154680 59110 154690
rect 58790 154600 58800 154680
rect 59110 154600 59120 154680
rect 58710 154500 58790 154510
rect 59030 154500 59110 154510
rect 58790 154420 58800 154500
rect 59110 154420 59120 154500
rect 58710 154320 58790 154330
rect 59030 154320 59110 154330
rect 58790 154240 58800 154320
rect 59110 154240 59120 154320
rect 58710 154140 58790 154150
rect 59030 154140 59110 154150
rect 58790 154060 58800 154140
rect 59110 154060 59120 154140
rect 58710 153960 58790 153970
rect 59030 153960 59110 153970
rect 58790 153880 58800 153960
rect 59110 153880 59120 153960
rect 58710 153780 58790 153790
rect 59030 153780 59110 153790
rect 58790 153700 58800 153780
rect 59110 153700 59120 153780
rect 58710 153600 58790 153610
rect 59030 153600 59110 153610
rect 58790 153520 58800 153600
rect 59110 153520 59120 153600
rect 58710 153420 58790 153430
rect 59030 153420 59110 153430
rect 58790 153340 58800 153420
rect 59110 153340 59120 153420
rect 58710 153240 58790 153250
rect 59030 153240 59110 153250
rect 58790 153160 58800 153240
rect 59110 153160 59120 153240
rect 58710 153060 58790 153070
rect 59030 153060 59110 153070
rect 58790 152980 58800 153060
rect 59110 152980 59120 153060
rect 59290 152900 59300 158900
rect 59310 152900 59340 158900
rect 59410 158830 59440 158900
rect 59670 158830 59760 158900
rect 60740 158839 60820 158849
rect 61060 158839 61140 158849
rect 61480 158839 61560 158849
rect 61800 158839 61880 158849
rect 59350 158820 59440 158830
rect 59500 158820 59580 158830
rect 59650 158820 59760 158830
rect 60060 158820 60140 158830
rect 60210 158820 60290 158830
rect 60360 158820 60440 158830
rect 59410 158650 59440 158820
rect 59580 158740 59590 158820
rect 59670 158650 59760 158820
rect 60140 158740 60150 158820
rect 60290 158740 60300 158820
rect 60440 158740 60450 158820
rect 60820 158759 60830 158839
rect 61140 158759 61150 158839
rect 61560 158759 61570 158839
rect 61880 158759 61890 158839
rect 62060 158820 62140 158830
rect 62210 158820 62290 158830
rect 62140 158740 62150 158820
rect 62290 158740 62300 158820
rect 60580 158679 60660 158689
rect 60900 158679 60980 158689
rect 61320 158679 61400 158689
rect 61640 158679 61720 158689
rect 59350 158640 59440 158650
rect 59500 158640 59580 158650
rect 59650 158640 59760 158650
rect 60060 158640 60140 158650
rect 60210 158640 60290 158650
rect 60360 158640 60440 158650
rect 59410 158470 59440 158640
rect 59580 158560 59590 158640
rect 59670 158470 59760 158640
rect 60140 158560 60150 158640
rect 60290 158560 60300 158640
rect 60440 158560 60450 158640
rect 60660 158599 60670 158679
rect 60980 158599 60990 158679
rect 61400 158599 61410 158679
rect 61720 158599 61730 158679
rect 62060 158640 62140 158650
rect 62210 158640 62290 158650
rect 62140 158560 62150 158640
rect 62290 158560 62300 158640
rect 60740 158519 60820 158529
rect 61060 158519 61140 158529
rect 61480 158519 61560 158529
rect 61800 158519 61880 158529
rect 59350 158460 59440 158470
rect 59500 158460 59580 158470
rect 59650 158460 59760 158470
rect 60060 158460 60140 158470
rect 60210 158460 60290 158470
rect 60360 158460 60440 158470
rect 59410 158290 59440 158460
rect 59580 158380 59590 158460
rect 59670 158290 59760 158460
rect 60140 158380 60150 158460
rect 60290 158380 60300 158460
rect 60440 158380 60450 158460
rect 60820 158439 60830 158519
rect 61140 158439 61150 158519
rect 61560 158439 61570 158519
rect 61880 158439 61890 158519
rect 62060 158460 62140 158470
rect 62210 158460 62290 158470
rect 62140 158380 62150 158460
rect 62290 158380 62300 158460
rect 60580 158359 60660 158369
rect 60900 158359 60980 158369
rect 61320 158359 61400 158369
rect 61640 158359 61720 158369
rect 59350 158280 59440 158290
rect 59500 158280 59580 158290
rect 59650 158280 59760 158290
rect 60060 158280 60140 158290
rect 60210 158280 60290 158290
rect 60360 158280 60440 158290
rect 59410 158110 59440 158280
rect 59580 158200 59590 158280
rect 59670 158110 59760 158280
rect 60140 158200 60150 158280
rect 60290 158200 60300 158280
rect 60440 158200 60450 158280
rect 60660 158279 60670 158359
rect 60980 158279 60990 158359
rect 61400 158279 61410 158359
rect 61720 158279 61730 158359
rect 62060 158280 62140 158290
rect 62210 158280 62290 158290
rect 60740 158199 60820 158209
rect 61060 158199 61140 158209
rect 61480 158199 61560 158209
rect 61800 158199 61880 158209
rect 62140 158200 62150 158280
rect 62290 158200 62300 158280
rect 60820 158119 60830 158199
rect 61140 158119 61150 158199
rect 61560 158119 61570 158199
rect 61880 158119 61890 158199
rect 59350 158100 59440 158110
rect 59500 158100 59580 158110
rect 59650 158100 59760 158110
rect 60060 158100 60140 158110
rect 60210 158100 60290 158110
rect 60360 158100 60440 158110
rect 62060 158100 62140 158110
rect 62210 158100 62290 158110
rect 59410 157930 59440 158100
rect 59580 158020 59590 158100
rect 59670 157930 59760 158100
rect 60140 158020 60150 158100
rect 60290 158020 60300 158100
rect 60440 158020 60450 158100
rect 60580 158039 60660 158049
rect 60900 158039 60980 158049
rect 61320 158039 61400 158049
rect 61640 158039 61720 158049
rect 60660 157959 60670 158039
rect 60980 157959 60990 158039
rect 61400 157959 61410 158039
rect 61720 157959 61730 158039
rect 62140 158020 62150 158100
rect 62290 158020 62300 158100
rect 59350 157920 59440 157930
rect 59500 157920 59580 157930
rect 59650 157920 59760 157930
rect 60060 157920 60140 157930
rect 60210 157920 60290 157930
rect 60360 157920 60440 157930
rect 62060 157920 62140 157930
rect 62210 157920 62290 157930
rect 59410 157750 59440 157920
rect 59580 157840 59590 157920
rect 59670 157750 59760 157920
rect 60140 157840 60150 157920
rect 60290 157840 60300 157920
rect 60440 157840 60450 157920
rect 60740 157879 60820 157889
rect 61060 157879 61140 157889
rect 61480 157879 61560 157889
rect 61800 157879 61880 157889
rect 60820 157799 60830 157879
rect 61140 157799 61150 157879
rect 61560 157799 61570 157879
rect 61880 157799 61890 157879
rect 62140 157840 62150 157920
rect 62290 157840 62300 157920
rect 59350 157740 59440 157750
rect 59500 157740 59580 157750
rect 59650 157740 59760 157750
rect 60060 157740 60140 157750
rect 60210 157740 60290 157750
rect 60360 157740 60440 157750
rect 62060 157740 62140 157750
rect 62210 157740 62290 157750
rect 59410 157570 59440 157740
rect 59580 157660 59590 157740
rect 59670 157570 59760 157740
rect 60140 157660 60150 157740
rect 60290 157660 60300 157740
rect 60440 157660 60450 157740
rect 60580 157719 60660 157729
rect 60900 157719 60980 157729
rect 61320 157719 61400 157729
rect 61640 157719 61720 157729
rect 60660 157639 60670 157719
rect 60980 157639 60990 157719
rect 61400 157639 61410 157719
rect 61720 157639 61730 157719
rect 62140 157660 62150 157740
rect 62290 157660 62300 157740
rect 59350 157560 59440 157570
rect 59500 157560 59580 157570
rect 59650 157560 59760 157570
rect 60060 157560 60140 157570
rect 60210 157560 60290 157570
rect 60360 157560 60440 157570
rect 59410 157390 59440 157560
rect 59580 157480 59590 157560
rect 59670 157390 59760 157560
rect 60140 157480 60150 157560
rect 60290 157480 60300 157560
rect 60440 157480 60450 157560
rect 60740 157559 60820 157569
rect 61060 157559 61140 157569
rect 61480 157559 61560 157569
rect 61800 157559 61880 157569
rect 62060 157560 62140 157570
rect 62210 157560 62290 157570
rect 60820 157479 60830 157559
rect 61140 157479 61150 157559
rect 61560 157479 61570 157559
rect 61880 157479 61890 157559
rect 62140 157480 62150 157560
rect 62290 157480 62300 157560
rect 60580 157399 60660 157409
rect 60900 157399 60980 157409
rect 61320 157399 61400 157409
rect 61640 157399 61720 157409
rect 59350 157380 59440 157390
rect 59500 157380 59580 157390
rect 59650 157380 59760 157390
rect 60060 157380 60140 157390
rect 60210 157380 60290 157390
rect 60360 157380 60440 157390
rect 59410 157210 59440 157380
rect 59580 157300 59590 157380
rect 59670 157210 59760 157380
rect 60140 157300 60150 157380
rect 60290 157300 60300 157380
rect 60440 157300 60450 157380
rect 60660 157319 60670 157399
rect 60980 157319 60990 157399
rect 61400 157319 61410 157399
rect 61720 157319 61730 157399
rect 62060 157380 62140 157390
rect 62210 157380 62290 157390
rect 62140 157300 62150 157380
rect 62290 157300 62300 157380
rect 60740 157239 60820 157249
rect 61060 157239 61140 157249
rect 61480 157239 61560 157249
rect 61800 157239 61880 157249
rect 59350 157200 59440 157210
rect 59500 157200 59580 157210
rect 59650 157200 59760 157210
rect 60060 157200 60140 157210
rect 60210 157200 60290 157210
rect 60360 157200 60440 157210
rect 59410 157030 59440 157200
rect 59580 157120 59590 157200
rect 59670 157030 59760 157200
rect 60140 157120 60150 157200
rect 60290 157120 60300 157200
rect 60440 157120 60450 157200
rect 60820 157159 60830 157239
rect 61140 157159 61150 157239
rect 61560 157159 61570 157239
rect 61880 157159 61890 157239
rect 62060 157200 62140 157210
rect 62210 157200 62290 157210
rect 62140 157120 62150 157200
rect 62290 157120 62300 157200
rect 60580 157079 60660 157089
rect 60900 157079 60980 157089
rect 61320 157079 61400 157089
rect 61640 157079 61720 157089
rect 59350 157020 59440 157030
rect 59500 157020 59580 157030
rect 59650 157020 59760 157030
rect 60060 157020 60140 157030
rect 60210 157020 60290 157030
rect 60360 157020 60440 157030
rect 59410 156850 59440 157020
rect 59580 156940 59590 157020
rect 59670 156850 59760 157020
rect 60140 156940 60150 157020
rect 60290 156940 60300 157020
rect 60440 156940 60450 157020
rect 60660 156999 60670 157079
rect 60980 156999 60990 157079
rect 61400 156999 61410 157079
rect 61720 156999 61730 157079
rect 62060 157020 62140 157030
rect 62210 157020 62290 157030
rect 62140 156940 62150 157020
rect 62290 156940 62300 157020
rect 60740 156919 60820 156929
rect 61060 156919 61140 156929
rect 61480 156919 61560 156929
rect 61800 156919 61880 156929
rect 59350 156840 59440 156850
rect 59500 156840 59580 156850
rect 59650 156840 59760 156850
rect 60060 156840 60140 156850
rect 60210 156840 60290 156850
rect 60360 156840 60440 156850
rect 59410 156670 59440 156840
rect 59580 156760 59590 156840
rect 59670 156670 59760 156840
rect 60140 156760 60150 156840
rect 60290 156760 60300 156840
rect 60440 156760 60450 156840
rect 60820 156839 60830 156919
rect 61140 156839 61150 156919
rect 61560 156839 61570 156919
rect 61880 156839 61890 156919
rect 62060 156840 62140 156850
rect 62210 156840 62290 156850
rect 60580 156759 60660 156769
rect 60900 156759 60980 156769
rect 61320 156759 61400 156769
rect 61640 156759 61720 156769
rect 62140 156760 62150 156840
rect 62290 156760 62300 156840
rect 60660 156679 60670 156759
rect 60980 156679 60990 156759
rect 61400 156679 61410 156759
rect 61720 156679 61730 156759
rect 59350 156660 59440 156670
rect 59500 156660 59580 156670
rect 59650 156660 59760 156670
rect 60060 156660 60140 156670
rect 60210 156660 60290 156670
rect 60360 156660 60440 156670
rect 62060 156660 62140 156670
rect 62210 156660 62290 156670
rect 59410 156490 59440 156660
rect 59580 156580 59590 156660
rect 59670 156490 59760 156660
rect 60140 156580 60150 156660
rect 60290 156580 60300 156660
rect 60440 156580 60450 156660
rect 60740 156599 60820 156609
rect 61060 156599 61140 156609
rect 61480 156599 61560 156609
rect 61800 156599 61880 156609
rect 60820 156519 60830 156599
rect 61140 156519 61150 156599
rect 61560 156519 61570 156599
rect 61880 156519 61890 156599
rect 62140 156580 62150 156660
rect 62290 156580 62300 156660
rect 59350 156480 59440 156490
rect 59500 156480 59580 156490
rect 59650 156480 59760 156490
rect 60060 156480 60140 156490
rect 60210 156480 60290 156490
rect 60360 156480 60440 156490
rect 62060 156480 62140 156490
rect 62210 156480 62290 156490
rect 59410 156310 59440 156480
rect 59580 156400 59590 156480
rect 59670 156310 59760 156480
rect 60140 156400 60150 156480
rect 60290 156400 60300 156480
rect 60440 156400 60450 156480
rect 60580 156439 60660 156449
rect 60900 156439 60980 156449
rect 61320 156439 61400 156449
rect 61640 156439 61720 156449
rect 60660 156359 60670 156439
rect 60980 156359 60990 156439
rect 61400 156359 61410 156439
rect 61720 156359 61730 156439
rect 62140 156400 62150 156480
rect 62290 156400 62300 156480
rect 59350 156300 59440 156310
rect 59500 156300 59580 156310
rect 59650 156300 59760 156310
rect 60060 156300 60140 156310
rect 60210 156300 60290 156310
rect 60360 156300 60440 156310
rect 62060 156300 62140 156310
rect 62210 156300 62290 156310
rect 59410 156130 59440 156300
rect 59580 156220 59590 156300
rect 59670 156130 59760 156300
rect 60140 156220 60150 156300
rect 60290 156220 60300 156300
rect 60440 156220 60450 156300
rect 60740 156279 60820 156289
rect 61060 156279 61140 156289
rect 61480 156279 61560 156289
rect 61800 156279 61880 156289
rect 60820 156199 60830 156279
rect 61140 156199 61150 156279
rect 61560 156199 61570 156279
rect 61880 156199 61890 156279
rect 62140 156220 62150 156300
rect 62290 156220 62300 156300
rect 59350 156120 59440 156130
rect 59500 156120 59580 156130
rect 59650 156120 59760 156130
rect 60060 156120 60140 156130
rect 60210 156120 60290 156130
rect 60360 156120 60440 156130
rect 59410 155950 59440 156120
rect 59580 156040 59590 156120
rect 59670 155950 59760 156120
rect 60140 156040 60150 156120
rect 60290 156040 60300 156120
rect 60440 156040 60450 156120
rect 60580 156119 60660 156129
rect 60900 156119 60980 156129
rect 61320 156119 61400 156129
rect 61640 156119 61720 156129
rect 62060 156120 62140 156130
rect 62210 156120 62290 156130
rect 60660 156039 60670 156119
rect 60980 156039 60990 156119
rect 61400 156039 61410 156119
rect 61720 156039 61730 156119
rect 62140 156040 62150 156120
rect 62290 156040 62300 156120
rect 60740 155959 60820 155969
rect 61060 155959 61140 155969
rect 61480 155959 61560 155969
rect 61800 155959 61880 155969
rect 59350 155940 59440 155950
rect 59500 155940 59580 155950
rect 59650 155940 59760 155950
rect 60060 155940 60140 155950
rect 60210 155940 60290 155950
rect 60360 155940 60440 155950
rect 59410 155770 59440 155940
rect 59580 155860 59590 155940
rect 59670 155770 59760 155940
rect 60140 155860 60150 155940
rect 60290 155860 60300 155940
rect 60440 155860 60450 155940
rect 60820 155879 60830 155959
rect 61140 155879 61150 155959
rect 61560 155879 61570 155959
rect 61880 155879 61890 155959
rect 62060 155940 62140 155950
rect 62210 155940 62290 155950
rect 62140 155860 62150 155940
rect 62290 155860 62300 155940
rect 60580 155799 60660 155809
rect 60900 155799 60980 155809
rect 61320 155799 61400 155809
rect 61640 155799 61720 155809
rect 59350 155760 59440 155770
rect 59500 155760 59580 155770
rect 59650 155760 59760 155770
rect 60060 155760 60140 155770
rect 60210 155760 60290 155770
rect 60360 155760 60440 155770
rect 59410 155590 59440 155760
rect 59580 155680 59590 155760
rect 59670 155590 59760 155760
rect 60140 155680 60150 155760
rect 60290 155680 60300 155760
rect 60440 155680 60450 155760
rect 60660 155719 60670 155799
rect 60980 155719 60990 155799
rect 61400 155719 61410 155799
rect 61720 155719 61730 155799
rect 62060 155760 62140 155770
rect 62210 155760 62290 155770
rect 62140 155680 62150 155760
rect 62290 155680 62300 155760
rect 60740 155639 60820 155649
rect 61060 155639 61140 155649
rect 61480 155639 61560 155649
rect 61800 155639 61880 155649
rect 59350 155580 59440 155590
rect 59500 155580 59580 155590
rect 59650 155580 59760 155590
rect 60060 155580 60140 155590
rect 60210 155580 60290 155590
rect 60360 155580 60440 155590
rect 59410 155410 59440 155580
rect 59580 155500 59590 155580
rect 59670 155410 59760 155580
rect 60140 155500 60150 155580
rect 60290 155500 60300 155580
rect 60440 155500 60450 155580
rect 60820 155559 60830 155639
rect 61140 155559 61150 155639
rect 61560 155559 61570 155639
rect 61880 155559 61890 155639
rect 62060 155580 62140 155590
rect 62210 155580 62290 155590
rect 62140 155500 62150 155580
rect 62290 155500 62300 155580
rect 60580 155479 60660 155489
rect 60900 155479 60980 155489
rect 61320 155479 61400 155489
rect 61640 155479 61720 155489
rect 59350 155400 59440 155410
rect 59500 155400 59580 155410
rect 59650 155400 59760 155410
rect 60060 155400 60140 155410
rect 60210 155400 60290 155410
rect 60360 155400 60440 155410
rect 59410 155230 59440 155400
rect 59580 155320 59590 155400
rect 59670 155230 59760 155400
rect 60140 155320 60150 155400
rect 60290 155320 60300 155400
rect 60440 155320 60450 155400
rect 60660 155399 60670 155479
rect 60980 155399 60990 155479
rect 61400 155399 61410 155479
rect 61720 155399 61730 155479
rect 62060 155400 62140 155410
rect 62210 155400 62290 155410
rect 60740 155319 60820 155329
rect 61060 155319 61140 155329
rect 61480 155319 61560 155329
rect 61800 155319 61880 155329
rect 62140 155320 62150 155400
rect 62290 155320 62300 155400
rect 60820 155239 60830 155319
rect 61140 155239 61150 155319
rect 61560 155239 61570 155319
rect 61880 155239 61890 155319
rect 59350 155220 59440 155230
rect 59500 155220 59580 155230
rect 59650 155220 59760 155230
rect 60060 155220 60140 155230
rect 60210 155220 60290 155230
rect 60360 155220 60440 155230
rect 62060 155220 62140 155230
rect 62210 155220 62290 155230
rect 59410 155050 59440 155220
rect 59580 155140 59590 155220
rect 59670 155050 59760 155220
rect 60140 155140 60150 155220
rect 60290 155140 60300 155220
rect 60440 155140 60450 155220
rect 60580 155159 60660 155169
rect 60900 155159 60980 155169
rect 61320 155159 61400 155169
rect 61640 155159 61720 155169
rect 60660 155079 60670 155159
rect 60980 155079 60990 155159
rect 61400 155079 61410 155159
rect 61720 155079 61730 155159
rect 62140 155140 62150 155220
rect 62290 155140 62300 155220
rect 59350 155040 59440 155050
rect 59500 155040 59580 155050
rect 59650 155040 59760 155050
rect 60060 155040 60140 155050
rect 60210 155040 60290 155050
rect 60360 155040 60440 155050
rect 62060 155040 62140 155050
rect 62210 155040 62290 155050
rect 59410 154870 59440 155040
rect 59580 154960 59590 155040
rect 59670 154870 59760 155040
rect 60140 154960 60150 155040
rect 60290 154960 60300 155040
rect 60440 154960 60450 155040
rect 60740 154999 60820 155009
rect 61060 154999 61140 155009
rect 61480 154999 61560 155009
rect 61800 154999 61880 155009
rect 60820 154919 60830 154999
rect 61140 154919 61150 154999
rect 61560 154919 61570 154999
rect 61880 154919 61890 154999
rect 62140 154960 62150 155040
rect 62290 154960 62300 155040
rect 59350 154860 59440 154870
rect 59500 154860 59580 154870
rect 59650 154860 59760 154870
rect 60060 154860 60140 154870
rect 60210 154860 60290 154870
rect 60360 154860 60440 154870
rect 62060 154860 62140 154870
rect 62210 154860 62290 154870
rect 59410 154690 59440 154860
rect 59580 154780 59590 154860
rect 59670 154690 59760 154860
rect 60140 154780 60150 154860
rect 60290 154780 60300 154860
rect 60440 154780 60450 154860
rect 60580 154839 60660 154849
rect 60900 154839 60980 154849
rect 61320 154839 61400 154849
rect 61640 154839 61720 154849
rect 60660 154759 60670 154839
rect 60980 154759 60990 154839
rect 61400 154759 61410 154839
rect 61720 154759 61730 154839
rect 62140 154780 62150 154860
rect 62290 154780 62300 154860
rect 59350 154680 59440 154690
rect 59500 154680 59580 154690
rect 59650 154680 59760 154690
rect 60060 154680 60140 154690
rect 60210 154680 60290 154690
rect 60360 154680 60440 154690
rect 59410 154510 59440 154680
rect 59580 154600 59590 154680
rect 59670 154510 59760 154680
rect 60140 154600 60150 154680
rect 60290 154600 60300 154680
rect 60440 154600 60450 154680
rect 60740 154679 60820 154689
rect 61060 154679 61140 154689
rect 61480 154679 61560 154689
rect 61800 154679 61880 154689
rect 62060 154680 62140 154690
rect 62210 154680 62290 154690
rect 60820 154599 60830 154679
rect 61140 154599 61150 154679
rect 61560 154599 61570 154679
rect 61880 154599 61890 154679
rect 62140 154600 62150 154680
rect 62290 154600 62300 154680
rect 60580 154519 60660 154529
rect 60900 154519 60980 154529
rect 61320 154519 61400 154529
rect 61640 154519 61720 154529
rect 59350 154500 59440 154510
rect 59500 154500 59580 154510
rect 59650 154500 59760 154510
rect 60060 154500 60140 154510
rect 60210 154500 60290 154510
rect 60360 154500 60440 154510
rect 59410 154330 59440 154500
rect 59580 154420 59590 154500
rect 59670 154330 59760 154500
rect 60140 154420 60150 154500
rect 60290 154420 60300 154500
rect 60440 154420 60450 154500
rect 60660 154439 60670 154519
rect 60980 154439 60990 154519
rect 61400 154439 61410 154519
rect 61720 154439 61730 154519
rect 62060 154500 62140 154510
rect 62210 154500 62290 154510
rect 62140 154420 62150 154500
rect 62290 154420 62300 154500
rect 60740 154359 60820 154369
rect 61060 154359 61140 154369
rect 61480 154359 61560 154369
rect 61800 154359 61880 154369
rect 59350 154320 59440 154330
rect 59500 154320 59580 154330
rect 59650 154320 59760 154330
rect 60060 154320 60140 154330
rect 60210 154320 60290 154330
rect 60360 154320 60440 154330
rect 59410 154150 59440 154320
rect 59580 154240 59590 154320
rect 59670 154150 59760 154320
rect 60140 154240 60150 154320
rect 60290 154240 60300 154320
rect 60440 154240 60450 154320
rect 60820 154279 60830 154359
rect 61140 154279 61150 154359
rect 61560 154279 61570 154359
rect 61880 154279 61890 154359
rect 62060 154320 62140 154330
rect 62210 154320 62290 154330
rect 62140 154240 62150 154320
rect 62290 154240 62300 154320
rect 60580 154199 60660 154209
rect 60900 154199 60980 154209
rect 61320 154199 61400 154209
rect 61640 154199 61720 154209
rect 59350 154140 59440 154150
rect 59500 154140 59580 154150
rect 59650 154140 59760 154150
rect 60060 154140 60140 154150
rect 60210 154140 60290 154150
rect 60360 154140 60440 154150
rect 59410 153970 59440 154140
rect 59580 154060 59590 154140
rect 59670 153970 59760 154140
rect 60140 154060 60150 154140
rect 60290 154060 60300 154140
rect 60440 154060 60450 154140
rect 60660 154119 60670 154199
rect 60980 154119 60990 154199
rect 61400 154119 61410 154199
rect 61720 154119 61730 154199
rect 62060 154140 62140 154150
rect 62210 154140 62290 154150
rect 62140 154060 62150 154140
rect 62290 154060 62300 154140
rect 60740 154039 60820 154049
rect 61060 154039 61140 154049
rect 61480 154039 61560 154049
rect 61800 154039 61880 154049
rect 59350 153960 59440 153970
rect 59500 153960 59580 153970
rect 59650 153960 59760 153970
rect 60060 153960 60140 153970
rect 60210 153960 60290 153970
rect 60360 153960 60440 153970
rect 59410 153790 59440 153960
rect 59580 153880 59590 153960
rect 59670 153790 59760 153960
rect 60140 153880 60150 153960
rect 60290 153880 60300 153960
rect 60440 153880 60450 153960
rect 60820 153959 60830 154039
rect 61140 153959 61150 154039
rect 61560 153959 61570 154039
rect 61880 153959 61890 154039
rect 62060 153960 62140 153970
rect 62210 153960 62290 153970
rect 60580 153879 60660 153889
rect 60900 153879 60980 153889
rect 61320 153879 61400 153889
rect 61640 153879 61720 153889
rect 62140 153880 62150 153960
rect 62290 153880 62300 153960
rect 60660 153799 60670 153879
rect 60980 153799 60990 153879
rect 61400 153799 61410 153879
rect 61720 153799 61730 153879
rect 59350 153780 59440 153790
rect 59500 153780 59580 153790
rect 59650 153780 59760 153790
rect 60060 153780 60140 153790
rect 60210 153780 60290 153790
rect 60360 153780 60440 153790
rect 62060 153780 62140 153790
rect 62210 153780 62290 153790
rect 59410 153610 59440 153780
rect 59580 153700 59590 153780
rect 59670 153610 59760 153780
rect 60140 153700 60150 153780
rect 60290 153700 60300 153780
rect 60440 153700 60450 153780
rect 60740 153719 60820 153729
rect 61060 153719 61140 153729
rect 61480 153719 61560 153729
rect 61800 153719 61880 153729
rect 60820 153639 60830 153719
rect 61140 153639 61150 153719
rect 61560 153639 61570 153719
rect 61880 153639 61890 153719
rect 62140 153700 62150 153780
rect 62290 153700 62300 153780
rect 59350 153600 59440 153610
rect 59500 153600 59580 153610
rect 59650 153600 59760 153610
rect 60060 153600 60140 153610
rect 60210 153600 60290 153610
rect 60360 153600 60440 153610
rect 62060 153600 62140 153610
rect 62210 153600 62290 153610
rect 59410 153430 59440 153600
rect 59580 153520 59590 153600
rect 59670 153430 59760 153600
rect 60140 153520 60150 153600
rect 60290 153520 60300 153600
rect 60440 153520 60450 153600
rect 60580 153559 60660 153569
rect 60900 153559 60980 153569
rect 61320 153559 61400 153569
rect 61640 153559 61720 153569
rect 60660 153479 60670 153559
rect 60980 153479 60990 153559
rect 61400 153479 61410 153559
rect 61720 153479 61730 153559
rect 62140 153520 62150 153600
rect 62290 153520 62300 153600
rect 59350 153420 59440 153430
rect 59500 153420 59580 153430
rect 59650 153420 59760 153430
rect 60060 153420 60140 153430
rect 60210 153420 60290 153430
rect 60360 153420 60440 153430
rect 62060 153420 62140 153430
rect 62210 153420 62290 153430
rect 59410 153250 59440 153420
rect 59580 153340 59590 153420
rect 59670 153250 59760 153420
rect 60140 153340 60150 153420
rect 60290 153340 60300 153420
rect 60440 153340 60450 153420
rect 60740 153399 60820 153409
rect 61060 153399 61140 153409
rect 61480 153399 61560 153409
rect 61800 153399 61880 153409
rect 60820 153319 60830 153399
rect 61140 153319 61150 153399
rect 61560 153319 61570 153399
rect 61880 153319 61890 153399
rect 62140 153340 62150 153420
rect 62290 153340 62300 153420
rect 59350 153240 59440 153250
rect 59500 153240 59580 153250
rect 59650 153240 59760 153250
rect 60060 153240 60140 153250
rect 60210 153240 60290 153250
rect 60360 153240 60440 153250
rect 59410 153070 59440 153240
rect 59580 153160 59590 153240
rect 59670 153070 59760 153240
rect 60140 153160 60150 153240
rect 60290 153160 60300 153240
rect 60440 153160 60450 153240
rect 60580 153239 60660 153249
rect 60900 153239 60980 153249
rect 61320 153239 61400 153249
rect 61640 153239 61720 153249
rect 62060 153240 62140 153250
rect 62210 153240 62290 153250
rect 60660 153159 60670 153239
rect 60980 153159 60990 153239
rect 61400 153159 61410 153239
rect 61720 153159 61730 153239
rect 62140 153160 62150 153240
rect 62290 153160 62300 153240
rect 60740 153079 60820 153089
rect 61060 153079 61140 153089
rect 61480 153079 61560 153089
rect 61800 153079 61880 153089
rect 59350 153060 59440 153070
rect 59500 153060 59580 153070
rect 59650 153060 59760 153070
rect 60060 153060 60140 153070
rect 60210 153060 60290 153070
rect 60360 153060 60440 153070
rect 59410 152900 59440 153060
rect 59580 152980 59590 153060
rect 59670 152900 59760 153060
rect 60140 152980 60150 153060
rect 60290 152980 60300 153060
rect 60440 152980 60450 153060
rect 60820 152999 60830 153079
rect 61140 152999 61150 153079
rect 61560 152999 61570 153079
rect 61880 152999 61890 153079
rect 62060 153060 62140 153070
rect 62210 153060 62290 153070
rect 62140 152980 62150 153060
rect 62290 152980 62300 153060
rect 60580 152919 60660 152929
rect 60900 152919 60980 152929
rect 61320 152919 61400 152929
rect 61640 152919 61720 152929
rect 48500 152880 48640 152890
rect 48710 152880 48790 152890
rect 60060 152880 60140 152890
rect 60210 152880 60290 152890
rect 60360 152880 60440 152890
rect 43945 152760 44025 152770
rect 44265 152760 44345 152770
rect 44585 152760 44665 152770
rect 44905 152760 44985 152770
rect 45225 152760 45305 152770
rect 45545 152760 45625 152770
rect 45865 152760 45945 152770
rect 46185 152760 46265 152770
rect 46505 152760 46585 152770
rect 46825 152760 46905 152770
rect 47145 152760 47225 152770
rect 47465 152760 47545 152770
rect 47785 152760 47865 152770
rect 48105 152760 48185 152770
rect 36020 152700 36100 152710
rect 36340 152700 36420 152710
rect 36660 152700 36740 152710
rect 36980 152700 37060 152710
rect 37300 152700 37380 152710
rect 37620 152700 37700 152710
rect 37940 152700 38020 152710
rect 38260 152700 38340 152710
rect 38580 152700 38660 152710
rect 38900 152700 38980 152710
rect 39220 152700 39300 152710
rect 39540 152700 39620 152710
rect 39860 152700 39940 152710
rect 40180 152700 40260 152710
rect 40500 152700 40580 152710
rect 40820 152700 40900 152710
rect 41140 152700 41220 152710
rect 41460 152700 41540 152710
rect 41780 152700 41860 152710
rect 42100 152700 42180 152710
rect 42420 152700 42500 152710
rect 42740 152700 42820 152710
rect 43060 152700 43140 152710
rect 43380 152700 43460 152710
rect 36100 152620 36110 152700
rect 36420 152620 36430 152700
rect 36740 152620 36750 152700
rect 37060 152620 37070 152700
rect 37380 152620 37390 152700
rect 37700 152620 37710 152700
rect 38020 152620 38030 152700
rect 38340 152620 38350 152700
rect 38660 152620 38670 152700
rect 38980 152620 38990 152700
rect 39300 152620 39310 152700
rect 39620 152620 39630 152700
rect 39940 152620 39950 152700
rect 40260 152620 40270 152700
rect 40580 152620 40590 152700
rect 40900 152620 40910 152700
rect 41220 152620 41230 152700
rect 41540 152620 41550 152700
rect 41860 152620 41870 152700
rect 42180 152620 42190 152700
rect 42500 152620 42510 152700
rect 42820 152620 42830 152700
rect 43140 152620 43150 152700
rect 43460 152620 43470 152700
rect 44025 152680 44035 152760
rect 44345 152680 44355 152760
rect 44665 152680 44675 152760
rect 44985 152680 44995 152760
rect 45305 152680 45315 152760
rect 45625 152680 45635 152760
rect 45945 152680 45955 152760
rect 46265 152680 46275 152760
rect 46585 152680 46595 152760
rect 46905 152680 46915 152760
rect 47225 152680 47235 152760
rect 47545 152680 47555 152760
rect 47865 152680 47875 152760
rect 48185 152680 48195 152760
rect 48500 152710 48605 152880
rect 48640 152800 48650 152880
rect 48790 152800 48800 152880
rect 60140 152800 60150 152880
rect 60290 152800 60300 152880
rect 60440 152800 60450 152880
rect 60660 152839 60670 152919
rect 60980 152839 60990 152919
rect 61400 152839 61410 152919
rect 61720 152839 61730 152919
rect 73245 152900 73260 158990
rect 73640 158920 73650 159000
rect 73790 158920 73800 159000
rect 73940 158920 73950 159000
rect 74080 158999 74160 159009
rect 74400 158999 74480 159009
rect 74820 158999 74900 159009
rect 75140 158999 75220 159009
rect 75560 159000 75640 159010
rect 75710 159000 75790 159010
rect 87060 159000 87140 159010
rect 87210 159000 87290 159010
rect 87360 159000 87440 159010
rect 74160 158919 74170 158999
rect 74480 158919 74490 158999
rect 74900 158919 74910 158999
rect 75220 158919 75230 158999
rect 75640 158920 75650 159000
rect 75790 158920 75800 159000
rect 76240 158900 76255 158990
rect 74240 158839 74320 158849
rect 74560 158839 74640 158849
rect 74980 158839 75060 158849
rect 75300 158839 75380 158849
rect 73560 158820 73640 158830
rect 73710 158820 73790 158830
rect 73860 158820 73940 158830
rect 73640 158740 73650 158820
rect 73790 158740 73800 158820
rect 73940 158740 73950 158820
rect 74320 158759 74330 158839
rect 74640 158759 74650 158839
rect 75060 158759 75070 158839
rect 75380 158759 75390 158839
rect 75560 158820 75640 158830
rect 75710 158820 75790 158830
rect 75640 158740 75650 158820
rect 75790 158740 75800 158820
rect 74080 158679 74160 158689
rect 74400 158679 74480 158689
rect 74820 158679 74900 158689
rect 75140 158679 75220 158689
rect 73560 158640 73640 158650
rect 73710 158640 73790 158650
rect 73860 158640 73940 158650
rect 73640 158560 73650 158640
rect 73790 158560 73800 158640
rect 73940 158560 73950 158640
rect 74160 158599 74170 158679
rect 74480 158599 74490 158679
rect 74900 158599 74910 158679
rect 75220 158599 75230 158679
rect 75560 158640 75640 158650
rect 75710 158640 75790 158650
rect 75640 158560 75650 158640
rect 75790 158560 75800 158640
rect 74240 158519 74320 158529
rect 74560 158519 74640 158529
rect 74980 158519 75060 158529
rect 75300 158519 75380 158529
rect 73560 158460 73640 158470
rect 73710 158460 73790 158470
rect 73860 158460 73940 158470
rect 73640 158380 73650 158460
rect 73790 158380 73800 158460
rect 73940 158380 73950 158460
rect 74320 158439 74330 158519
rect 74640 158439 74650 158519
rect 75060 158439 75070 158519
rect 75380 158439 75390 158519
rect 75560 158460 75640 158470
rect 75710 158460 75790 158470
rect 75640 158380 75650 158460
rect 75790 158380 75800 158460
rect 74080 158359 74160 158369
rect 74400 158359 74480 158369
rect 74820 158359 74900 158369
rect 75140 158359 75220 158369
rect 73560 158280 73640 158290
rect 73710 158280 73790 158290
rect 73860 158280 73940 158290
rect 73640 158200 73650 158280
rect 73790 158200 73800 158280
rect 73940 158200 73950 158280
rect 74160 158279 74170 158359
rect 74480 158279 74490 158359
rect 74900 158279 74910 158359
rect 75220 158279 75230 158359
rect 75560 158280 75640 158290
rect 75710 158280 75790 158290
rect 74240 158199 74320 158209
rect 74560 158199 74640 158209
rect 74980 158199 75060 158209
rect 75300 158199 75380 158209
rect 75640 158200 75650 158280
rect 75790 158200 75800 158280
rect 74320 158119 74330 158199
rect 74640 158119 74650 158199
rect 75060 158119 75070 158199
rect 75380 158119 75390 158199
rect 73560 158100 73640 158110
rect 73710 158100 73790 158110
rect 73860 158100 73940 158110
rect 75560 158100 75640 158110
rect 75710 158100 75790 158110
rect 73640 158020 73650 158100
rect 73790 158020 73800 158100
rect 73940 158020 73950 158100
rect 74080 158039 74160 158049
rect 74400 158039 74480 158049
rect 74820 158039 74900 158049
rect 75140 158039 75220 158049
rect 74160 157959 74170 158039
rect 74480 157959 74490 158039
rect 74900 157959 74910 158039
rect 75220 157959 75230 158039
rect 75640 158020 75650 158100
rect 75790 158020 75800 158100
rect 73560 157920 73640 157930
rect 73710 157920 73790 157930
rect 73860 157920 73940 157930
rect 75560 157920 75640 157930
rect 75710 157920 75790 157930
rect 73640 157840 73650 157920
rect 73790 157840 73800 157920
rect 73940 157840 73950 157920
rect 74240 157879 74320 157889
rect 74560 157879 74640 157889
rect 74980 157879 75060 157889
rect 75300 157879 75380 157889
rect 74320 157799 74330 157879
rect 74640 157799 74650 157879
rect 75060 157799 75070 157879
rect 75380 157799 75390 157879
rect 75640 157840 75650 157920
rect 75790 157840 75800 157920
rect 73560 157740 73640 157750
rect 73710 157740 73790 157750
rect 73860 157740 73940 157750
rect 75560 157740 75640 157750
rect 75710 157740 75790 157750
rect 73640 157660 73650 157740
rect 73790 157660 73800 157740
rect 73940 157660 73950 157740
rect 74080 157719 74160 157729
rect 74400 157719 74480 157729
rect 74820 157719 74900 157729
rect 75140 157719 75220 157729
rect 74160 157639 74170 157719
rect 74480 157639 74490 157719
rect 74900 157639 74910 157719
rect 75220 157639 75230 157719
rect 75640 157660 75650 157740
rect 75790 157660 75800 157740
rect 73560 157560 73640 157570
rect 73710 157560 73790 157570
rect 73860 157560 73940 157570
rect 73640 157480 73650 157560
rect 73790 157480 73800 157560
rect 73940 157480 73950 157560
rect 74240 157559 74320 157569
rect 74560 157559 74640 157569
rect 74980 157559 75060 157569
rect 75300 157559 75380 157569
rect 75560 157560 75640 157570
rect 75710 157560 75790 157570
rect 74320 157479 74330 157559
rect 74640 157479 74650 157559
rect 75060 157479 75070 157559
rect 75380 157479 75390 157559
rect 75640 157480 75650 157560
rect 75790 157480 75800 157560
rect 74080 157399 74160 157409
rect 74400 157399 74480 157409
rect 74820 157399 74900 157409
rect 75140 157399 75220 157409
rect 73560 157380 73640 157390
rect 73710 157380 73790 157390
rect 73860 157380 73940 157390
rect 73640 157300 73650 157380
rect 73790 157300 73800 157380
rect 73940 157300 73950 157380
rect 74160 157319 74170 157399
rect 74480 157319 74490 157399
rect 74900 157319 74910 157399
rect 75220 157319 75230 157399
rect 75560 157380 75640 157390
rect 75710 157380 75790 157390
rect 75640 157300 75650 157380
rect 75790 157300 75800 157380
rect 74240 157239 74320 157249
rect 74560 157239 74640 157249
rect 74980 157239 75060 157249
rect 75300 157239 75380 157249
rect 73560 157200 73640 157210
rect 73710 157200 73790 157210
rect 73860 157200 73940 157210
rect 73640 157120 73650 157200
rect 73790 157120 73800 157200
rect 73940 157120 73950 157200
rect 74320 157159 74330 157239
rect 74640 157159 74650 157239
rect 75060 157159 75070 157239
rect 75380 157159 75390 157239
rect 75560 157200 75640 157210
rect 75710 157200 75790 157210
rect 75640 157120 75650 157200
rect 75790 157120 75800 157200
rect 74080 157079 74160 157089
rect 74400 157079 74480 157089
rect 74820 157079 74900 157089
rect 75140 157079 75220 157089
rect 73560 157020 73640 157030
rect 73710 157020 73790 157030
rect 73860 157020 73940 157030
rect 73640 156940 73650 157020
rect 73790 156940 73800 157020
rect 73940 156940 73950 157020
rect 74160 156999 74170 157079
rect 74480 156999 74490 157079
rect 74900 156999 74910 157079
rect 75220 156999 75230 157079
rect 75560 157020 75640 157030
rect 75710 157020 75790 157030
rect 75640 156940 75650 157020
rect 75790 156940 75800 157020
rect 74240 156919 74320 156929
rect 74560 156919 74640 156929
rect 74980 156919 75060 156929
rect 75300 156919 75380 156929
rect 73560 156840 73640 156850
rect 73710 156840 73790 156850
rect 73860 156840 73940 156850
rect 73640 156760 73650 156840
rect 73790 156760 73800 156840
rect 73940 156760 73950 156840
rect 74320 156839 74330 156919
rect 74640 156839 74650 156919
rect 75060 156839 75070 156919
rect 75380 156839 75390 156919
rect 75560 156840 75640 156850
rect 75710 156840 75790 156850
rect 74080 156759 74160 156769
rect 74400 156759 74480 156769
rect 74820 156759 74900 156769
rect 75140 156759 75220 156769
rect 75640 156760 75650 156840
rect 75790 156760 75800 156840
rect 74160 156679 74170 156759
rect 74480 156679 74490 156759
rect 74900 156679 74910 156759
rect 75220 156679 75230 156759
rect 73560 156660 73640 156670
rect 73710 156660 73790 156670
rect 73860 156660 73940 156670
rect 75560 156660 75640 156670
rect 75710 156660 75790 156670
rect 73640 156580 73650 156660
rect 73790 156580 73800 156660
rect 73940 156580 73950 156660
rect 74240 156599 74320 156609
rect 74560 156599 74640 156609
rect 74980 156599 75060 156609
rect 75300 156599 75380 156609
rect 74320 156519 74330 156599
rect 74640 156519 74650 156599
rect 75060 156519 75070 156599
rect 75380 156519 75390 156599
rect 75640 156580 75650 156660
rect 75790 156580 75800 156660
rect 73560 156480 73640 156490
rect 73710 156480 73790 156490
rect 73860 156480 73940 156490
rect 75560 156480 75640 156490
rect 75710 156480 75790 156490
rect 73640 156400 73650 156480
rect 73790 156400 73800 156480
rect 73940 156400 73950 156480
rect 74080 156439 74160 156449
rect 74400 156439 74480 156449
rect 74820 156439 74900 156449
rect 75140 156439 75220 156449
rect 74160 156359 74170 156439
rect 74480 156359 74490 156439
rect 74900 156359 74910 156439
rect 75220 156359 75230 156439
rect 75640 156400 75650 156480
rect 75790 156400 75800 156480
rect 73560 156300 73640 156310
rect 73710 156300 73790 156310
rect 73860 156300 73940 156310
rect 75560 156300 75640 156310
rect 75710 156300 75790 156310
rect 73640 156220 73650 156300
rect 73790 156220 73800 156300
rect 73940 156220 73950 156300
rect 74240 156279 74320 156289
rect 74560 156279 74640 156289
rect 74980 156279 75060 156289
rect 75300 156279 75380 156289
rect 74320 156199 74330 156279
rect 74640 156199 74650 156279
rect 75060 156199 75070 156279
rect 75380 156199 75390 156279
rect 75640 156220 75650 156300
rect 75790 156220 75800 156300
rect 73560 156120 73640 156130
rect 73710 156120 73790 156130
rect 73860 156120 73940 156130
rect 73640 156040 73650 156120
rect 73790 156040 73800 156120
rect 73940 156040 73950 156120
rect 74080 156119 74160 156129
rect 74400 156119 74480 156129
rect 74820 156119 74900 156129
rect 75140 156119 75220 156129
rect 75560 156120 75640 156130
rect 75710 156120 75790 156130
rect 74160 156039 74170 156119
rect 74480 156039 74490 156119
rect 74900 156039 74910 156119
rect 75220 156039 75230 156119
rect 75640 156040 75650 156120
rect 75790 156040 75800 156120
rect 74240 155959 74320 155969
rect 74560 155959 74640 155969
rect 74980 155959 75060 155969
rect 75300 155959 75380 155969
rect 73560 155940 73640 155950
rect 73710 155940 73790 155950
rect 73860 155940 73940 155950
rect 73640 155860 73650 155940
rect 73790 155860 73800 155940
rect 73940 155860 73950 155940
rect 74320 155879 74330 155959
rect 74640 155879 74650 155959
rect 75060 155879 75070 155959
rect 75380 155879 75390 155959
rect 75560 155940 75640 155950
rect 75710 155940 75790 155950
rect 75640 155860 75650 155940
rect 75790 155860 75800 155940
rect 74080 155799 74160 155809
rect 74400 155799 74480 155809
rect 74820 155799 74900 155809
rect 75140 155799 75220 155809
rect 73560 155760 73640 155770
rect 73710 155760 73790 155770
rect 73860 155760 73940 155770
rect 73640 155680 73650 155760
rect 73790 155680 73800 155760
rect 73940 155680 73950 155760
rect 74160 155719 74170 155799
rect 74480 155719 74490 155799
rect 74900 155719 74910 155799
rect 75220 155719 75230 155799
rect 75560 155760 75640 155770
rect 75710 155760 75790 155770
rect 75640 155680 75650 155760
rect 75790 155680 75800 155760
rect 74240 155639 74320 155649
rect 74560 155639 74640 155649
rect 74980 155639 75060 155649
rect 75300 155639 75380 155649
rect 73560 155580 73640 155590
rect 73710 155580 73790 155590
rect 73860 155580 73940 155590
rect 73640 155500 73650 155580
rect 73790 155500 73800 155580
rect 73940 155500 73950 155580
rect 74320 155559 74330 155639
rect 74640 155559 74650 155639
rect 75060 155559 75070 155639
rect 75380 155559 75390 155639
rect 75560 155580 75640 155590
rect 75710 155580 75790 155590
rect 75640 155500 75650 155580
rect 75790 155500 75800 155580
rect 74080 155479 74160 155489
rect 74400 155479 74480 155489
rect 74820 155479 74900 155489
rect 75140 155479 75220 155489
rect 73560 155400 73640 155410
rect 73710 155400 73790 155410
rect 73860 155400 73940 155410
rect 73640 155320 73650 155400
rect 73790 155320 73800 155400
rect 73940 155320 73950 155400
rect 74160 155399 74170 155479
rect 74480 155399 74490 155479
rect 74900 155399 74910 155479
rect 75220 155399 75230 155479
rect 75560 155400 75640 155410
rect 75710 155400 75790 155410
rect 74240 155319 74320 155329
rect 74560 155319 74640 155329
rect 74980 155319 75060 155329
rect 75300 155319 75380 155329
rect 75640 155320 75650 155400
rect 75790 155320 75800 155400
rect 74320 155239 74330 155319
rect 74640 155239 74650 155319
rect 75060 155239 75070 155319
rect 75380 155239 75390 155319
rect 73560 155220 73640 155230
rect 73710 155220 73790 155230
rect 73860 155220 73940 155230
rect 75560 155220 75640 155230
rect 75710 155220 75790 155230
rect 73640 155140 73650 155220
rect 73790 155140 73800 155220
rect 73940 155140 73950 155220
rect 74080 155159 74160 155169
rect 74400 155159 74480 155169
rect 74820 155159 74900 155169
rect 75140 155159 75220 155169
rect 74160 155079 74170 155159
rect 74480 155079 74490 155159
rect 74900 155079 74910 155159
rect 75220 155079 75230 155159
rect 75640 155140 75650 155220
rect 75790 155140 75800 155220
rect 73560 155040 73640 155050
rect 73710 155040 73790 155050
rect 73860 155040 73940 155050
rect 75560 155040 75640 155050
rect 75710 155040 75790 155050
rect 73640 154960 73650 155040
rect 73790 154960 73800 155040
rect 73940 154960 73950 155040
rect 74240 154999 74320 155009
rect 74560 154999 74640 155009
rect 74980 154999 75060 155009
rect 75300 154999 75380 155009
rect 74320 154919 74330 154999
rect 74640 154919 74650 154999
rect 75060 154919 75070 154999
rect 75380 154919 75390 154999
rect 75640 154960 75650 155040
rect 75790 154960 75800 155040
rect 73560 154860 73640 154870
rect 73710 154860 73790 154870
rect 73860 154860 73940 154870
rect 75560 154860 75640 154870
rect 75710 154860 75790 154870
rect 73640 154780 73650 154860
rect 73790 154780 73800 154860
rect 73940 154780 73950 154860
rect 74080 154839 74160 154849
rect 74400 154839 74480 154849
rect 74820 154839 74900 154849
rect 75140 154839 75220 154849
rect 74160 154759 74170 154839
rect 74480 154759 74490 154839
rect 74900 154759 74910 154839
rect 75220 154759 75230 154839
rect 75640 154780 75650 154860
rect 75790 154780 75800 154860
rect 73560 154680 73640 154690
rect 73710 154680 73790 154690
rect 73860 154680 73940 154690
rect 73640 154600 73650 154680
rect 73790 154600 73800 154680
rect 73940 154600 73950 154680
rect 74240 154679 74320 154689
rect 74560 154679 74640 154689
rect 74980 154679 75060 154689
rect 75300 154679 75380 154689
rect 75560 154680 75640 154690
rect 75710 154680 75790 154690
rect 74320 154599 74330 154679
rect 74640 154599 74650 154679
rect 75060 154599 75070 154679
rect 75380 154599 75390 154679
rect 75640 154600 75650 154680
rect 75790 154600 75800 154680
rect 74080 154519 74160 154529
rect 74400 154519 74480 154529
rect 74820 154519 74900 154529
rect 75140 154519 75220 154529
rect 73560 154500 73640 154510
rect 73710 154500 73790 154510
rect 73860 154500 73940 154510
rect 73640 154420 73650 154500
rect 73790 154420 73800 154500
rect 73940 154420 73950 154500
rect 74160 154439 74170 154519
rect 74480 154439 74490 154519
rect 74900 154439 74910 154519
rect 75220 154439 75230 154519
rect 75560 154500 75640 154510
rect 75710 154500 75790 154510
rect 75640 154420 75650 154500
rect 75790 154420 75800 154500
rect 74240 154359 74320 154369
rect 74560 154359 74640 154369
rect 74980 154359 75060 154369
rect 75300 154359 75380 154369
rect 73560 154320 73640 154330
rect 73710 154320 73790 154330
rect 73860 154320 73940 154330
rect 73640 154240 73650 154320
rect 73790 154240 73800 154320
rect 73940 154240 73950 154320
rect 74320 154279 74330 154359
rect 74640 154279 74650 154359
rect 75060 154279 75070 154359
rect 75380 154279 75390 154359
rect 75560 154320 75640 154330
rect 75710 154320 75790 154330
rect 75640 154240 75650 154320
rect 75790 154240 75800 154320
rect 74080 154199 74160 154209
rect 74400 154199 74480 154209
rect 74820 154199 74900 154209
rect 75140 154199 75220 154209
rect 73560 154140 73640 154150
rect 73710 154140 73790 154150
rect 73860 154140 73940 154150
rect 73640 154060 73650 154140
rect 73790 154060 73800 154140
rect 73940 154060 73950 154140
rect 74160 154119 74170 154199
rect 74480 154119 74490 154199
rect 74900 154119 74910 154199
rect 75220 154119 75230 154199
rect 75560 154140 75640 154150
rect 75710 154140 75790 154150
rect 75640 154060 75650 154140
rect 75790 154060 75800 154140
rect 74240 154039 74320 154049
rect 74560 154039 74640 154049
rect 74980 154039 75060 154049
rect 75300 154039 75380 154049
rect 73560 153960 73640 153970
rect 73710 153960 73790 153970
rect 73860 153960 73940 153970
rect 73640 153880 73650 153960
rect 73790 153880 73800 153960
rect 73940 153880 73950 153960
rect 74320 153959 74330 154039
rect 74640 153959 74650 154039
rect 75060 153959 75070 154039
rect 75380 153959 75390 154039
rect 75560 153960 75640 153970
rect 75710 153960 75790 153970
rect 74080 153879 74160 153889
rect 74400 153879 74480 153889
rect 74820 153879 74900 153889
rect 75140 153879 75220 153889
rect 75640 153880 75650 153960
rect 75790 153880 75800 153960
rect 74160 153799 74170 153879
rect 74480 153799 74490 153879
rect 74900 153799 74910 153879
rect 75220 153799 75230 153879
rect 73560 153780 73640 153790
rect 73710 153780 73790 153790
rect 73860 153780 73940 153790
rect 75560 153780 75640 153790
rect 75710 153780 75790 153790
rect 73640 153700 73650 153780
rect 73790 153700 73800 153780
rect 73940 153700 73950 153780
rect 74240 153719 74320 153729
rect 74560 153719 74640 153729
rect 74980 153719 75060 153729
rect 75300 153719 75380 153729
rect 74320 153639 74330 153719
rect 74640 153639 74650 153719
rect 75060 153639 75070 153719
rect 75380 153639 75390 153719
rect 75640 153700 75650 153780
rect 75790 153700 75800 153780
rect 73560 153600 73640 153610
rect 73710 153600 73790 153610
rect 73860 153600 73940 153610
rect 75560 153600 75640 153610
rect 75710 153600 75790 153610
rect 73640 153520 73650 153600
rect 73790 153520 73800 153600
rect 73940 153520 73950 153600
rect 74080 153559 74160 153569
rect 74400 153559 74480 153569
rect 74820 153559 74900 153569
rect 75140 153559 75220 153569
rect 74160 153479 74170 153559
rect 74480 153479 74490 153559
rect 74900 153479 74910 153559
rect 75220 153479 75230 153559
rect 75640 153520 75650 153600
rect 75790 153520 75800 153600
rect 73560 153420 73640 153430
rect 73710 153420 73790 153430
rect 73860 153420 73940 153430
rect 75560 153420 75640 153430
rect 75710 153420 75790 153430
rect 73640 153340 73650 153420
rect 73790 153340 73800 153420
rect 73940 153340 73950 153420
rect 74240 153399 74320 153409
rect 74560 153399 74640 153409
rect 74980 153399 75060 153409
rect 75300 153399 75380 153409
rect 74320 153319 74330 153399
rect 74640 153319 74650 153399
rect 75060 153319 75070 153399
rect 75380 153319 75390 153399
rect 75640 153340 75650 153420
rect 75790 153340 75800 153420
rect 73560 153240 73640 153250
rect 73710 153240 73790 153250
rect 73860 153240 73940 153250
rect 73640 153160 73650 153240
rect 73790 153160 73800 153240
rect 73940 153160 73950 153240
rect 74080 153239 74160 153249
rect 74400 153239 74480 153249
rect 74820 153239 74900 153249
rect 75140 153239 75220 153249
rect 75560 153240 75640 153250
rect 75710 153240 75790 153250
rect 74160 153159 74170 153239
rect 74480 153159 74490 153239
rect 74900 153159 74910 153239
rect 75220 153159 75230 153239
rect 75640 153160 75650 153240
rect 75790 153160 75800 153240
rect 74240 153079 74320 153089
rect 74560 153079 74640 153089
rect 74980 153079 75060 153089
rect 75300 153079 75380 153089
rect 73560 153060 73640 153070
rect 73710 153060 73790 153070
rect 73860 153060 73940 153070
rect 73640 152980 73650 153060
rect 73790 152980 73800 153060
rect 73940 152980 73950 153060
rect 74320 152999 74330 153079
rect 74640 152999 74650 153079
rect 75060 152999 75070 153079
rect 75380 152999 75390 153079
rect 75560 153060 75640 153070
rect 75710 153060 75790 153070
rect 75640 152980 75650 153060
rect 75790 152980 75800 153060
rect 74080 152919 74160 152929
rect 74400 152919 74480 152929
rect 74820 152919 74900 152929
rect 75140 152919 75220 152929
rect 62060 152880 62140 152890
rect 62210 152880 62290 152890
rect 73560 152880 73640 152890
rect 73710 152880 73790 152890
rect 73860 152880 73940 152890
rect 62140 152800 62150 152880
rect 62290 152800 62300 152880
rect 73640 152800 73650 152880
rect 73790 152800 73800 152880
rect 73940 152800 73950 152880
rect 74160 152839 74170 152919
rect 74480 152839 74490 152919
rect 74900 152839 74910 152919
rect 75220 152839 75230 152919
rect 86745 152900 86760 158990
rect 87140 158920 87150 159000
rect 87290 158920 87300 159000
rect 87440 158920 87450 159000
rect 87580 158999 87660 159009
rect 87900 158999 87980 159009
rect 88320 158999 88400 159009
rect 88640 158999 88720 159009
rect 89060 159000 89140 159010
rect 89210 159000 89290 159010
rect 100560 159000 100640 159010
rect 100710 159000 100790 159010
rect 100860 159000 100940 159010
rect 87660 158919 87670 158999
rect 87980 158919 87990 158999
rect 88400 158919 88410 158999
rect 88720 158919 88730 158999
rect 89140 158920 89150 159000
rect 89290 158920 89300 159000
rect 89740 158900 89755 158990
rect 87740 158839 87820 158849
rect 88060 158839 88140 158849
rect 88480 158839 88560 158849
rect 88800 158839 88880 158849
rect 87060 158820 87140 158830
rect 87210 158820 87290 158830
rect 87360 158820 87440 158830
rect 87140 158740 87150 158820
rect 87290 158740 87300 158820
rect 87440 158740 87450 158820
rect 87820 158759 87830 158839
rect 88140 158759 88150 158839
rect 88560 158759 88570 158839
rect 88880 158759 88890 158839
rect 89060 158820 89140 158830
rect 89210 158820 89290 158830
rect 89140 158740 89150 158820
rect 89290 158740 89300 158820
rect 87580 158679 87660 158689
rect 87900 158679 87980 158689
rect 88320 158679 88400 158689
rect 88640 158679 88720 158689
rect 87060 158640 87140 158650
rect 87210 158640 87290 158650
rect 87360 158640 87440 158650
rect 87140 158560 87150 158640
rect 87290 158560 87300 158640
rect 87440 158560 87450 158640
rect 87660 158599 87670 158679
rect 87980 158599 87990 158679
rect 88400 158599 88410 158679
rect 88720 158599 88730 158679
rect 89060 158640 89140 158650
rect 89210 158640 89290 158650
rect 89140 158560 89150 158640
rect 89290 158560 89300 158640
rect 87740 158519 87820 158529
rect 88060 158519 88140 158529
rect 88480 158519 88560 158529
rect 88800 158519 88880 158529
rect 87060 158460 87140 158470
rect 87210 158460 87290 158470
rect 87360 158460 87440 158470
rect 87140 158380 87150 158460
rect 87290 158380 87300 158460
rect 87440 158380 87450 158460
rect 87820 158439 87830 158519
rect 88140 158439 88150 158519
rect 88560 158439 88570 158519
rect 88880 158439 88890 158519
rect 89060 158460 89140 158470
rect 89210 158460 89290 158470
rect 89140 158380 89150 158460
rect 89290 158380 89300 158460
rect 87580 158359 87660 158369
rect 87900 158359 87980 158369
rect 88320 158359 88400 158369
rect 88640 158359 88720 158369
rect 87060 158280 87140 158290
rect 87210 158280 87290 158290
rect 87360 158280 87440 158290
rect 87140 158200 87150 158280
rect 87290 158200 87300 158280
rect 87440 158200 87450 158280
rect 87660 158279 87670 158359
rect 87980 158279 87990 158359
rect 88400 158279 88410 158359
rect 88720 158279 88730 158359
rect 89060 158280 89140 158290
rect 89210 158280 89290 158290
rect 87740 158199 87820 158209
rect 88060 158199 88140 158209
rect 88480 158199 88560 158209
rect 88800 158199 88880 158209
rect 89140 158200 89150 158280
rect 89290 158200 89300 158280
rect 87820 158119 87830 158199
rect 88140 158119 88150 158199
rect 88560 158119 88570 158199
rect 88880 158119 88890 158199
rect 87060 158100 87140 158110
rect 87210 158100 87290 158110
rect 87360 158100 87440 158110
rect 89060 158100 89140 158110
rect 89210 158100 89290 158110
rect 87140 158020 87150 158100
rect 87290 158020 87300 158100
rect 87440 158020 87450 158100
rect 87580 158039 87660 158049
rect 87900 158039 87980 158049
rect 88320 158039 88400 158049
rect 88640 158039 88720 158049
rect 87660 157959 87670 158039
rect 87980 157959 87990 158039
rect 88400 157959 88410 158039
rect 88720 157959 88730 158039
rect 89140 158020 89150 158100
rect 89290 158020 89300 158100
rect 87060 157920 87140 157930
rect 87210 157920 87290 157930
rect 87360 157920 87440 157930
rect 89060 157920 89140 157930
rect 89210 157920 89290 157930
rect 87140 157840 87150 157920
rect 87290 157840 87300 157920
rect 87440 157840 87450 157920
rect 87740 157879 87820 157889
rect 88060 157879 88140 157889
rect 88480 157879 88560 157889
rect 88800 157879 88880 157889
rect 87820 157799 87830 157879
rect 88140 157799 88150 157879
rect 88560 157799 88570 157879
rect 88880 157799 88890 157879
rect 89140 157840 89150 157920
rect 89290 157840 89300 157920
rect 87060 157740 87140 157750
rect 87210 157740 87290 157750
rect 87360 157740 87440 157750
rect 89060 157740 89140 157750
rect 89210 157740 89290 157750
rect 87140 157660 87150 157740
rect 87290 157660 87300 157740
rect 87440 157660 87450 157740
rect 87580 157719 87660 157729
rect 87900 157719 87980 157729
rect 88320 157719 88400 157729
rect 88640 157719 88720 157729
rect 87660 157639 87670 157719
rect 87980 157639 87990 157719
rect 88400 157639 88410 157719
rect 88720 157639 88730 157719
rect 89140 157660 89150 157740
rect 89290 157660 89300 157740
rect 87060 157560 87140 157570
rect 87210 157560 87290 157570
rect 87360 157560 87440 157570
rect 87140 157480 87150 157560
rect 87290 157480 87300 157560
rect 87440 157480 87450 157560
rect 87740 157559 87820 157569
rect 88060 157559 88140 157569
rect 88480 157559 88560 157569
rect 88800 157559 88880 157569
rect 89060 157560 89140 157570
rect 89210 157560 89290 157570
rect 87820 157479 87830 157559
rect 88140 157479 88150 157559
rect 88560 157479 88570 157559
rect 88880 157479 88890 157559
rect 89140 157480 89150 157560
rect 89290 157480 89300 157560
rect 87580 157399 87660 157409
rect 87900 157399 87980 157409
rect 88320 157399 88400 157409
rect 88640 157399 88720 157409
rect 87060 157380 87140 157390
rect 87210 157380 87290 157390
rect 87360 157380 87440 157390
rect 87140 157300 87150 157380
rect 87290 157300 87300 157380
rect 87440 157300 87450 157380
rect 87660 157319 87670 157399
rect 87980 157319 87990 157399
rect 88400 157319 88410 157399
rect 88720 157319 88730 157399
rect 89060 157380 89140 157390
rect 89210 157380 89290 157390
rect 89140 157300 89150 157380
rect 89290 157300 89300 157380
rect 87740 157239 87820 157249
rect 88060 157239 88140 157249
rect 88480 157239 88560 157249
rect 88800 157239 88880 157249
rect 87060 157200 87140 157210
rect 87210 157200 87290 157210
rect 87360 157200 87440 157210
rect 87140 157120 87150 157200
rect 87290 157120 87300 157200
rect 87440 157120 87450 157200
rect 87820 157159 87830 157239
rect 88140 157159 88150 157239
rect 88560 157159 88570 157239
rect 88880 157159 88890 157239
rect 89060 157200 89140 157210
rect 89210 157200 89290 157210
rect 89140 157120 89150 157200
rect 89290 157120 89300 157200
rect 87580 157079 87660 157089
rect 87900 157079 87980 157089
rect 88320 157079 88400 157089
rect 88640 157079 88720 157089
rect 87060 157020 87140 157030
rect 87210 157020 87290 157030
rect 87360 157020 87440 157030
rect 87140 156940 87150 157020
rect 87290 156940 87300 157020
rect 87440 156940 87450 157020
rect 87660 156999 87670 157079
rect 87980 156999 87990 157079
rect 88400 156999 88410 157079
rect 88720 156999 88730 157079
rect 89060 157020 89140 157030
rect 89210 157020 89290 157030
rect 89140 156940 89150 157020
rect 89290 156940 89300 157020
rect 87740 156919 87820 156929
rect 88060 156919 88140 156929
rect 88480 156919 88560 156929
rect 88800 156919 88880 156929
rect 87060 156840 87140 156850
rect 87210 156840 87290 156850
rect 87360 156840 87440 156850
rect 87140 156760 87150 156840
rect 87290 156760 87300 156840
rect 87440 156760 87450 156840
rect 87820 156839 87830 156919
rect 88140 156839 88150 156919
rect 88560 156839 88570 156919
rect 88880 156839 88890 156919
rect 89060 156840 89140 156850
rect 89210 156840 89290 156850
rect 87580 156759 87660 156769
rect 87900 156759 87980 156769
rect 88320 156759 88400 156769
rect 88640 156759 88720 156769
rect 89140 156760 89150 156840
rect 89290 156760 89300 156840
rect 87660 156679 87670 156759
rect 87980 156679 87990 156759
rect 88400 156679 88410 156759
rect 88720 156679 88730 156759
rect 87060 156660 87140 156670
rect 87210 156660 87290 156670
rect 87360 156660 87440 156670
rect 89060 156660 89140 156670
rect 89210 156660 89290 156670
rect 87140 156580 87150 156660
rect 87290 156580 87300 156660
rect 87440 156580 87450 156660
rect 87740 156599 87820 156609
rect 88060 156599 88140 156609
rect 88480 156599 88560 156609
rect 88800 156599 88880 156609
rect 87820 156519 87830 156599
rect 88140 156519 88150 156599
rect 88560 156519 88570 156599
rect 88880 156519 88890 156599
rect 89140 156580 89150 156660
rect 89290 156580 89300 156660
rect 87060 156480 87140 156490
rect 87210 156480 87290 156490
rect 87360 156480 87440 156490
rect 89060 156480 89140 156490
rect 89210 156480 89290 156490
rect 87140 156400 87150 156480
rect 87290 156400 87300 156480
rect 87440 156400 87450 156480
rect 87580 156439 87660 156449
rect 87900 156439 87980 156449
rect 88320 156439 88400 156449
rect 88640 156439 88720 156449
rect 87660 156359 87670 156439
rect 87980 156359 87990 156439
rect 88400 156359 88410 156439
rect 88720 156359 88730 156439
rect 89140 156400 89150 156480
rect 89290 156400 89300 156480
rect 87060 156300 87140 156310
rect 87210 156300 87290 156310
rect 87360 156300 87440 156310
rect 89060 156300 89140 156310
rect 89210 156300 89290 156310
rect 87140 156220 87150 156300
rect 87290 156220 87300 156300
rect 87440 156220 87450 156300
rect 87740 156279 87820 156289
rect 88060 156279 88140 156289
rect 88480 156279 88560 156289
rect 88800 156279 88880 156289
rect 87820 156199 87830 156279
rect 88140 156199 88150 156279
rect 88560 156199 88570 156279
rect 88880 156199 88890 156279
rect 89140 156220 89150 156300
rect 89290 156220 89300 156300
rect 87060 156120 87140 156130
rect 87210 156120 87290 156130
rect 87360 156120 87440 156130
rect 87140 156040 87150 156120
rect 87290 156040 87300 156120
rect 87440 156040 87450 156120
rect 87580 156119 87660 156129
rect 87900 156119 87980 156129
rect 88320 156119 88400 156129
rect 88640 156119 88720 156129
rect 89060 156120 89140 156130
rect 89210 156120 89290 156130
rect 87660 156039 87670 156119
rect 87980 156039 87990 156119
rect 88400 156039 88410 156119
rect 88720 156039 88730 156119
rect 89140 156040 89150 156120
rect 89290 156040 89300 156120
rect 87740 155959 87820 155969
rect 88060 155959 88140 155969
rect 88480 155959 88560 155969
rect 88800 155959 88880 155969
rect 87060 155940 87140 155950
rect 87210 155940 87290 155950
rect 87360 155940 87440 155950
rect 87140 155860 87150 155940
rect 87290 155860 87300 155940
rect 87440 155860 87450 155940
rect 87820 155879 87830 155959
rect 88140 155879 88150 155959
rect 88560 155879 88570 155959
rect 88880 155879 88890 155959
rect 89060 155940 89140 155950
rect 89210 155940 89290 155950
rect 89140 155860 89150 155940
rect 89290 155860 89300 155940
rect 87580 155799 87660 155809
rect 87900 155799 87980 155809
rect 88320 155799 88400 155809
rect 88640 155799 88720 155809
rect 87060 155760 87140 155770
rect 87210 155760 87290 155770
rect 87360 155760 87440 155770
rect 87140 155680 87150 155760
rect 87290 155680 87300 155760
rect 87440 155680 87450 155760
rect 87660 155719 87670 155799
rect 87980 155719 87990 155799
rect 88400 155719 88410 155799
rect 88720 155719 88730 155799
rect 89060 155760 89140 155770
rect 89210 155760 89290 155770
rect 89140 155680 89150 155760
rect 89290 155680 89300 155760
rect 87740 155639 87820 155649
rect 88060 155639 88140 155649
rect 88480 155639 88560 155649
rect 88800 155639 88880 155649
rect 87060 155580 87140 155590
rect 87210 155580 87290 155590
rect 87360 155580 87440 155590
rect 87140 155500 87150 155580
rect 87290 155500 87300 155580
rect 87440 155500 87450 155580
rect 87820 155559 87830 155639
rect 88140 155559 88150 155639
rect 88560 155559 88570 155639
rect 88880 155559 88890 155639
rect 89060 155580 89140 155590
rect 89210 155580 89290 155590
rect 89140 155500 89150 155580
rect 89290 155500 89300 155580
rect 87580 155479 87660 155489
rect 87900 155479 87980 155489
rect 88320 155479 88400 155489
rect 88640 155479 88720 155489
rect 87060 155400 87140 155410
rect 87210 155400 87290 155410
rect 87360 155400 87440 155410
rect 87140 155320 87150 155400
rect 87290 155320 87300 155400
rect 87440 155320 87450 155400
rect 87660 155399 87670 155479
rect 87980 155399 87990 155479
rect 88400 155399 88410 155479
rect 88720 155399 88730 155479
rect 89060 155400 89140 155410
rect 89210 155400 89290 155410
rect 87740 155319 87820 155329
rect 88060 155319 88140 155329
rect 88480 155319 88560 155329
rect 88800 155319 88880 155329
rect 89140 155320 89150 155400
rect 89290 155320 89300 155400
rect 87820 155239 87830 155319
rect 88140 155239 88150 155319
rect 88560 155239 88570 155319
rect 88880 155239 88890 155319
rect 87060 155220 87140 155230
rect 87210 155220 87290 155230
rect 87360 155220 87440 155230
rect 89060 155220 89140 155230
rect 89210 155220 89290 155230
rect 87140 155140 87150 155220
rect 87290 155140 87300 155220
rect 87440 155140 87450 155220
rect 87580 155159 87660 155169
rect 87900 155159 87980 155169
rect 88320 155159 88400 155169
rect 88640 155159 88720 155169
rect 87660 155079 87670 155159
rect 87980 155079 87990 155159
rect 88400 155079 88410 155159
rect 88720 155079 88730 155159
rect 89140 155140 89150 155220
rect 89290 155140 89300 155220
rect 87060 155040 87140 155050
rect 87210 155040 87290 155050
rect 87360 155040 87440 155050
rect 89060 155040 89140 155050
rect 89210 155040 89290 155050
rect 87140 154960 87150 155040
rect 87290 154960 87300 155040
rect 87440 154960 87450 155040
rect 87740 154999 87820 155009
rect 88060 154999 88140 155009
rect 88480 154999 88560 155009
rect 88800 154999 88880 155009
rect 87820 154919 87830 154999
rect 88140 154919 88150 154999
rect 88560 154919 88570 154999
rect 88880 154919 88890 154999
rect 89140 154960 89150 155040
rect 89290 154960 89300 155040
rect 87060 154860 87140 154870
rect 87210 154860 87290 154870
rect 87360 154860 87440 154870
rect 89060 154860 89140 154870
rect 89210 154860 89290 154870
rect 87140 154780 87150 154860
rect 87290 154780 87300 154860
rect 87440 154780 87450 154860
rect 87580 154839 87660 154849
rect 87900 154839 87980 154849
rect 88320 154839 88400 154849
rect 88640 154839 88720 154849
rect 87660 154759 87670 154839
rect 87980 154759 87990 154839
rect 88400 154759 88410 154839
rect 88720 154759 88730 154839
rect 89140 154780 89150 154860
rect 89290 154780 89300 154860
rect 87060 154680 87140 154690
rect 87210 154680 87290 154690
rect 87360 154680 87440 154690
rect 87140 154600 87150 154680
rect 87290 154600 87300 154680
rect 87440 154600 87450 154680
rect 87740 154679 87820 154689
rect 88060 154679 88140 154689
rect 88480 154679 88560 154689
rect 88800 154679 88880 154689
rect 89060 154680 89140 154690
rect 89210 154680 89290 154690
rect 87820 154599 87830 154679
rect 88140 154599 88150 154679
rect 88560 154599 88570 154679
rect 88880 154599 88890 154679
rect 89140 154600 89150 154680
rect 89290 154600 89300 154680
rect 87580 154519 87660 154529
rect 87900 154519 87980 154529
rect 88320 154519 88400 154529
rect 88640 154519 88720 154529
rect 87060 154500 87140 154510
rect 87210 154500 87290 154510
rect 87360 154500 87440 154510
rect 87140 154420 87150 154500
rect 87290 154420 87300 154500
rect 87440 154420 87450 154500
rect 87660 154439 87670 154519
rect 87980 154439 87990 154519
rect 88400 154439 88410 154519
rect 88720 154439 88730 154519
rect 89060 154500 89140 154510
rect 89210 154500 89290 154510
rect 89140 154420 89150 154500
rect 89290 154420 89300 154500
rect 87740 154359 87820 154369
rect 88060 154359 88140 154369
rect 88480 154359 88560 154369
rect 88800 154359 88880 154369
rect 87060 154320 87140 154330
rect 87210 154320 87290 154330
rect 87360 154320 87440 154330
rect 87140 154240 87150 154320
rect 87290 154240 87300 154320
rect 87440 154240 87450 154320
rect 87820 154279 87830 154359
rect 88140 154279 88150 154359
rect 88560 154279 88570 154359
rect 88880 154279 88890 154359
rect 89060 154320 89140 154330
rect 89210 154320 89290 154330
rect 89140 154240 89150 154320
rect 89290 154240 89300 154320
rect 87580 154199 87660 154209
rect 87900 154199 87980 154209
rect 88320 154199 88400 154209
rect 88640 154199 88720 154209
rect 87060 154140 87140 154150
rect 87210 154140 87290 154150
rect 87360 154140 87440 154150
rect 87140 154060 87150 154140
rect 87290 154060 87300 154140
rect 87440 154060 87450 154140
rect 87660 154119 87670 154199
rect 87980 154119 87990 154199
rect 88400 154119 88410 154199
rect 88720 154119 88730 154199
rect 89060 154140 89140 154150
rect 89210 154140 89290 154150
rect 89140 154060 89150 154140
rect 89290 154060 89300 154140
rect 87740 154039 87820 154049
rect 88060 154039 88140 154049
rect 88480 154039 88560 154049
rect 88800 154039 88880 154049
rect 87060 153960 87140 153970
rect 87210 153960 87290 153970
rect 87360 153960 87440 153970
rect 87140 153880 87150 153960
rect 87290 153880 87300 153960
rect 87440 153880 87450 153960
rect 87820 153959 87830 154039
rect 88140 153959 88150 154039
rect 88560 153959 88570 154039
rect 88880 153959 88890 154039
rect 89060 153960 89140 153970
rect 89210 153960 89290 153970
rect 87580 153879 87660 153889
rect 87900 153879 87980 153889
rect 88320 153879 88400 153889
rect 88640 153879 88720 153889
rect 89140 153880 89150 153960
rect 89290 153880 89300 153960
rect 87660 153799 87670 153879
rect 87980 153799 87990 153879
rect 88400 153799 88410 153879
rect 88720 153799 88730 153879
rect 87060 153780 87140 153790
rect 87210 153780 87290 153790
rect 87360 153780 87440 153790
rect 89060 153780 89140 153790
rect 89210 153780 89290 153790
rect 87140 153700 87150 153780
rect 87290 153700 87300 153780
rect 87440 153700 87450 153780
rect 87740 153719 87820 153729
rect 88060 153719 88140 153729
rect 88480 153719 88560 153729
rect 88800 153719 88880 153729
rect 87820 153639 87830 153719
rect 88140 153639 88150 153719
rect 88560 153639 88570 153719
rect 88880 153639 88890 153719
rect 89140 153700 89150 153780
rect 89290 153700 89300 153780
rect 87060 153600 87140 153610
rect 87210 153600 87290 153610
rect 87360 153600 87440 153610
rect 89060 153600 89140 153610
rect 89210 153600 89290 153610
rect 87140 153520 87150 153600
rect 87290 153520 87300 153600
rect 87440 153520 87450 153600
rect 87580 153559 87660 153569
rect 87900 153559 87980 153569
rect 88320 153559 88400 153569
rect 88640 153559 88720 153569
rect 87660 153479 87670 153559
rect 87980 153479 87990 153559
rect 88400 153479 88410 153559
rect 88720 153479 88730 153559
rect 89140 153520 89150 153600
rect 89290 153520 89300 153600
rect 87060 153420 87140 153430
rect 87210 153420 87290 153430
rect 87360 153420 87440 153430
rect 89060 153420 89140 153430
rect 89210 153420 89290 153430
rect 87140 153340 87150 153420
rect 87290 153340 87300 153420
rect 87440 153340 87450 153420
rect 87740 153399 87820 153409
rect 88060 153399 88140 153409
rect 88480 153399 88560 153409
rect 88800 153399 88880 153409
rect 87820 153319 87830 153399
rect 88140 153319 88150 153399
rect 88560 153319 88570 153399
rect 88880 153319 88890 153399
rect 89140 153340 89150 153420
rect 89290 153340 89300 153420
rect 87060 153240 87140 153250
rect 87210 153240 87290 153250
rect 87360 153240 87440 153250
rect 87140 153160 87150 153240
rect 87290 153160 87300 153240
rect 87440 153160 87450 153240
rect 87580 153239 87660 153249
rect 87900 153239 87980 153249
rect 88320 153239 88400 153249
rect 88640 153239 88720 153249
rect 89060 153240 89140 153250
rect 89210 153240 89290 153250
rect 87660 153159 87670 153239
rect 87980 153159 87990 153239
rect 88400 153159 88410 153239
rect 88720 153159 88730 153239
rect 89140 153160 89150 153240
rect 89290 153160 89300 153240
rect 87740 153079 87820 153089
rect 88060 153079 88140 153089
rect 88480 153079 88560 153089
rect 88800 153079 88880 153089
rect 87060 153060 87140 153070
rect 87210 153060 87290 153070
rect 87360 153060 87440 153070
rect 87140 152980 87150 153060
rect 87290 152980 87300 153060
rect 87440 152980 87450 153060
rect 87820 152999 87830 153079
rect 88140 152999 88150 153079
rect 88560 152999 88570 153079
rect 88880 152999 88890 153079
rect 89060 153060 89140 153070
rect 89210 153060 89290 153070
rect 89140 152980 89150 153060
rect 89290 152980 89300 153060
rect 87580 152919 87660 152929
rect 87900 152919 87980 152929
rect 88320 152919 88400 152929
rect 88640 152919 88720 152929
rect 75560 152880 75640 152890
rect 75710 152880 75790 152890
rect 87060 152880 87140 152890
rect 87210 152880 87290 152890
rect 87360 152880 87440 152890
rect 75640 152800 75650 152880
rect 75790 152800 75800 152880
rect 87140 152800 87150 152880
rect 87290 152800 87300 152880
rect 87440 152800 87450 152880
rect 87660 152839 87670 152919
rect 87980 152839 87990 152919
rect 88400 152839 88410 152919
rect 88720 152839 88730 152919
rect 100245 152900 100260 158990
rect 100640 158920 100650 159000
rect 100790 158920 100800 159000
rect 100940 158920 100950 159000
rect 101080 158999 101160 159009
rect 101400 158999 101480 159009
rect 101820 158999 101900 159009
rect 102140 158999 102220 159009
rect 114580 158999 114660 159009
rect 114900 158999 114980 159009
rect 115320 158999 115400 159009
rect 115640 158999 115720 159009
rect 116060 159000 116140 159010
rect 116210 159000 116290 159010
rect 127560 159000 127640 159010
rect 127710 159000 127790 159010
rect 127860 159000 127940 159010
rect 101160 158919 101170 158999
rect 101480 158919 101490 158999
rect 101900 158919 101910 158999
rect 102220 158919 102230 158999
rect 114660 158919 114670 158999
rect 114980 158919 114990 158999
rect 115400 158919 115410 158999
rect 115720 158919 115730 158999
rect 116140 158920 116150 159000
rect 116290 158920 116300 159000
rect 116740 158900 116755 158990
rect 101240 158839 101320 158849
rect 101560 158839 101640 158849
rect 101980 158839 102060 158849
rect 102300 158839 102380 158849
rect 114740 158839 114820 158849
rect 115060 158839 115140 158849
rect 115480 158839 115560 158849
rect 115800 158839 115880 158849
rect 100560 158820 100640 158830
rect 100710 158820 100790 158830
rect 100860 158820 100940 158830
rect 100640 158740 100650 158820
rect 100790 158740 100800 158820
rect 100940 158740 100950 158820
rect 101320 158759 101330 158839
rect 101640 158759 101650 158839
rect 102060 158759 102070 158839
rect 102380 158759 102390 158839
rect 114820 158759 114830 158839
rect 115140 158759 115150 158839
rect 115560 158759 115570 158839
rect 115880 158759 115890 158839
rect 116060 158820 116140 158830
rect 116210 158820 116290 158830
rect 116140 158740 116150 158820
rect 116290 158740 116300 158820
rect 101080 158679 101160 158689
rect 101400 158679 101480 158689
rect 101820 158679 101900 158689
rect 102140 158679 102220 158689
rect 114580 158679 114660 158689
rect 114900 158679 114980 158689
rect 115320 158679 115400 158689
rect 115640 158679 115720 158689
rect 100560 158640 100640 158650
rect 100710 158640 100790 158650
rect 100860 158640 100940 158650
rect 100640 158560 100650 158640
rect 100790 158560 100800 158640
rect 100940 158560 100950 158640
rect 101160 158599 101170 158679
rect 101480 158599 101490 158679
rect 101900 158599 101910 158679
rect 102220 158599 102230 158679
rect 114660 158599 114670 158679
rect 114980 158599 114990 158679
rect 115400 158599 115410 158679
rect 115720 158599 115730 158679
rect 116060 158640 116140 158650
rect 116210 158640 116290 158650
rect 116140 158560 116150 158640
rect 116290 158560 116300 158640
rect 101240 158519 101320 158529
rect 101560 158519 101640 158529
rect 101980 158519 102060 158529
rect 102300 158519 102380 158529
rect 114740 158519 114820 158529
rect 115060 158519 115140 158529
rect 115480 158519 115560 158529
rect 115800 158519 115880 158529
rect 100560 158460 100640 158470
rect 100710 158460 100790 158470
rect 100860 158460 100940 158470
rect 100640 158380 100650 158460
rect 100790 158380 100800 158460
rect 100940 158380 100950 158460
rect 101320 158439 101330 158519
rect 101640 158439 101650 158519
rect 102060 158439 102070 158519
rect 102380 158439 102390 158519
rect 114820 158439 114830 158519
rect 115140 158439 115150 158519
rect 115560 158439 115570 158519
rect 115880 158439 115890 158519
rect 116060 158460 116140 158470
rect 116210 158460 116290 158470
rect 116140 158380 116150 158460
rect 116290 158380 116300 158460
rect 101080 158359 101160 158369
rect 101400 158359 101480 158369
rect 101820 158359 101900 158369
rect 102140 158359 102220 158369
rect 114580 158359 114660 158369
rect 114900 158359 114980 158369
rect 115320 158359 115400 158369
rect 115640 158359 115720 158369
rect 100560 158280 100640 158290
rect 100710 158280 100790 158290
rect 100860 158280 100940 158290
rect 100640 158200 100650 158280
rect 100790 158200 100800 158280
rect 100940 158200 100950 158280
rect 101160 158279 101170 158359
rect 101480 158279 101490 158359
rect 101900 158279 101910 158359
rect 102220 158279 102230 158359
rect 114660 158279 114670 158359
rect 114980 158279 114990 158359
rect 115400 158279 115410 158359
rect 115720 158279 115730 158359
rect 116060 158280 116140 158290
rect 116210 158280 116290 158290
rect 101240 158199 101320 158209
rect 101560 158199 101640 158209
rect 101980 158199 102060 158209
rect 102300 158199 102380 158209
rect 114740 158199 114820 158209
rect 115060 158199 115140 158209
rect 115480 158199 115560 158209
rect 115800 158199 115880 158209
rect 116140 158200 116150 158280
rect 116290 158200 116300 158280
rect 101320 158119 101330 158199
rect 101640 158119 101650 158199
rect 102060 158119 102070 158199
rect 102380 158119 102390 158199
rect 114820 158119 114830 158199
rect 115140 158119 115150 158199
rect 115560 158119 115570 158199
rect 115880 158119 115890 158199
rect 100560 158100 100640 158110
rect 100710 158100 100790 158110
rect 100860 158100 100940 158110
rect 116060 158100 116140 158110
rect 116210 158100 116290 158110
rect 100640 158020 100650 158100
rect 100790 158020 100800 158100
rect 100940 158020 100950 158100
rect 101080 158039 101160 158049
rect 101400 158039 101480 158049
rect 101820 158039 101900 158049
rect 102140 158039 102220 158049
rect 114580 158039 114660 158049
rect 114900 158039 114980 158049
rect 115320 158039 115400 158049
rect 115640 158039 115720 158049
rect 101160 157959 101170 158039
rect 101480 157959 101490 158039
rect 101900 157959 101910 158039
rect 102220 157959 102230 158039
rect 114660 157959 114670 158039
rect 114980 157959 114990 158039
rect 115400 157959 115410 158039
rect 115720 157959 115730 158039
rect 116140 158020 116150 158100
rect 116290 158020 116300 158100
rect 100560 157920 100640 157930
rect 100710 157920 100790 157930
rect 100860 157920 100940 157930
rect 116060 157920 116140 157930
rect 116210 157920 116290 157930
rect 100640 157840 100650 157920
rect 100790 157840 100800 157920
rect 100940 157840 100950 157920
rect 101240 157879 101320 157889
rect 101560 157879 101640 157889
rect 101980 157879 102060 157889
rect 102300 157879 102380 157889
rect 114740 157879 114820 157889
rect 115060 157879 115140 157889
rect 115480 157879 115560 157889
rect 115800 157879 115880 157889
rect 101320 157799 101330 157879
rect 101640 157799 101650 157879
rect 102060 157799 102070 157879
rect 102380 157799 102390 157879
rect 114820 157799 114830 157879
rect 115140 157799 115150 157879
rect 115560 157799 115570 157879
rect 115880 157799 115890 157879
rect 116140 157840 116150 157920
rect 116290 157840 116300 157920
rect 100560 157740 100640 157750
rect 100710 157740 100790 157750
rect 100860 157740 100940 157750
rect 116060 157740 116140 157750
rect 116210 157740 116290 157750
rect 100640 157660 100650 157740
rect 100790 157660 100800 157740
rect 100940 157660 100950 157740
rect 101080 157719 101160 157729
rect 101400 157719 101480 157729
rect 101820 157719 101900 157729
rect 102140 157719 102220 157729
rect 114580 157719 114660 157729
rect 114900 157719 114980 157729
rect 115320 157719 115400 157729
rect 115640 157719 115720 157729
rect 101160 157639 101170 157719
rect 101480 157639 101490 157719
rect 101900 157639 101910 157719
rect 102220 157639 102230 157719
rect 114660 157639 114670 157719
rect 114980 157639 114990 157719
rect 115400 157639 115410 157719
rect 115720 157639 115730 157719
rect 116140 157660 116150 157740
rect 116290 157660 116300 157740
rect 100560 157560 100640 157570
rect 100710 157560 100790 157570
rect 100860 157560 100940 157570
rect 100640 157480 100650 157560
rect 100790 157480 100800 157560
rect 100940 157480 100950 157560
rect 101240 157559 101320 157569
rect 101560 157559 101640 157569
rect 101980 157559 102060 157569
rect 102300 157559 102380 157569
rect 114740 157559 114820 157569
rect 115060 157559 115140 157569
rect 115480 157559 115560 157569
rect 115800 157559 115880 157569
rect 116060 157560 116140 157570
rect 116210 157560 116290 157570
rect 101320 157479 101330 157559
rect 101640 157479 101650 157559
rect 102060 157479 102070 157559
rect 102380 157479 102390 157559
rect 114820 157479 114830 157559
rect 115140 157479 115150 157559
rect 115560 157479 115570 157559
rect 115880 157479 115890 157559
rect 116140 157480 116150 157560
rect 116290 157480 116300 157560
rect 101080 157399 101160 157409
rect 101400 157399 101480 157409
rect 101820 157399 101900 157409
rect 102140 157399 102220 157409
rect 114580 157399 114660 157409
rect 114900 157399 114980 157409
rect 115320 157399 115400 157409
rect 115640 157399 115720 157409
rect 100560 157380 100640 157390
rect 100710 157380 100790 157390
rect 100860 157380 100940 157390
rect 100640 157300 100650 157380
rect 100790 157300 100800 157380
rect 100940 157300 100950 157380
rect 101160 157319 101170 157399
rect 101480 157319 101490 157399
rect 101900 157319 101910 157399
rect 102220 157319 102230 157399
rect 114660 157319 114670 157399
rect 114980 157319 114990 157399
rect 115400 157319 115410 157399
rect 115720 157319 115730 157399
rect 116060 157380 116140 157390
rect 116210 157380 116290 157390
rect 116140 157300 116150 157380
rect 116290 157300 116300 157380
rect 101240 157239 101320 157249
rect 101560 157239 101640 157249
rect 101980 157239 102060 157249
rect 102300 157239 102380 157249
rect 114740 157239 114820 157249
rect 115060 157239 115140 157249
rect 115480 157239 115560 157249
rect 115800 157239 115880 157249
rect 100560 157200 100640 157210
rect 100710 157200 100790 157210
rect 100860 157200 100940 157210
rect 100640 157120 100650 157200
rect 100790 157120 100800 157200
rect 100940 157120 100950 157200
rect 101320 157159 101330 157239
rect 101640 157159 101650 157239
rect 102060 157159 102070 157239
rect 102380 157159 102390 157239
rect 114820 157159 114830 157239
rect 115140 157159 115150 157239
rect 115560 157159 115570 157239
rect 115880 157159 115890 157239
rect 116060 157200 116140 157210
rect 116210 157200 116290 157210
rect 116140 157120 116150 157200
rect 116290 157120 116300 157200
rect 101080 157079 101160 157089
rect 101400 157079 101480 157089
rect 101820 157079 101900 157089
rect 102140 157079 102220 157089
rect 114580 157079 114660 157089
rect 114900 157079 114980 157089
rect 115320 157079 115400 157089
rect 115640 157079 115720 157089
rect 100560 157020 100640 157030
rect 100710 157020 100790 157030
rect 100860 157020 100940 157030
rect 100640 156940 100650 157020
rect 100790 156940 100800 157020
rect 100940 156940 100950 157020
rect 101160 156999 101170 157079
rect 101480 156999 101490 157079
rect 101900 156999 101910 157079
rect 102220 156999 102230 157079
rect 114660 156999 114670 157079
rect 114980 156999 114990 157079
rect 115400 156999 115410 157079
rect 115720 156999 115730 157079
rect 116060 157020 116140 157030
rect 116210 157020 116290 157030
rect 116140 156940 116150 157020
rect 116290 156940 116300 157020
rect 101240 156919 101320 156929
rect 101560 156919 101640 156929
rect 101980 156919 102060 156929
rect 102300 156919 102380 156929
rect 114740 156919 114820 156929
rect 115060 156919 115140 156929
rect 115480 156919 115560 156929
rect 115800 156919 115880 156929
rect 100560 156840 100640 156850
rect 100710 156840 100790 156850
rect 100860 156840 100940 156850
rect 100640 156760 100650 156840
rect 100790 156760 100800 156840
rect 100940 156760 100950 156840
rect 101320 156839 101330 156919
rect 101640 156839 101650 156919
rect 102060 156839 102070 156919
rect 102380 156839 102390 156919
rect 114820 156839 114830 156919
rect 115140 156839 115150 156919
rect 115560 156839 115570 156919
rect 115880 156839 115890 156919
rect 116060 156840 116140 156850
rect 116210 156840 116290 156850
rect 101080 156759 101160 156769
rect 101400 156759 101480 156769
rect 101820 156759 101900 156769
rect 102140 156759 102220 156769
rect 114580 156759 114660 156769
rect 114900 156759 114980 156769
rect 115320 156759 115400 156769
rect 115640 156759 115720 156769
rect 116140 156760 116150 156840
rect 116290 156760 116300 156840
rect 101160 156679 101170 156759
rect 101480 156679 101490 156759
rect 101900 156679 101910 156759
rect 102220 156679 102230 156759
rect 114660 156679 114670 156759
rect 114980 156679 114990 156759
rect 115400 156679 115410 156759
rect 115720 156679 115730 156759
rect 100560 156660 100640 156670
rect 100710 156660 100790 156670
rect 100860 156660 100940 156670
rect 116060 156660 116140 156670
rect 116210 156660 116290 156670
rect 100640 156580 100650 156660
rect 100790 156580 100800 156660
rect 100940 156580 100950 156660
rect 101240 156599 101320 156609
rect 101560 156599 101640 156609
rect 101980 156599 102060 156609
rect 102300 156599 102380 156609
rect 114740 156599 114820 156609
rect 115060 156599 115140 156609
rect 115480 156599 115560 156609
rect 115800 156599 115880 156609
rect 101320 156519 101330 156599
rect 101640 156519 101650 156599
rect 102060 156519 102070 156599
rect 102380 156519 102390 156599
rect 114820 156519 114830 156599
rect 115140 156519 115150 156599
rect 115560 156519 115570 156599
rect 115880 156519 115890 156599
rect 116140 156580 116150 156660
rect 116290 156580 116300 156660
rect 100560 156480 100640 156490
rect 100710 156480 100790 156490
rect 100860 156480 100940 156490
rect 116060 156480 116140 156490
rect 116210 156480 116290 156490
rect 100640 156400 100650 156480
rect 100790 156400 100800 156480
rect 100940 156400 100950 156480
rect 101080 156439 101160 156449
rect 101400 156439 101480 156449
rect 101820 156439 101900 156449
rect 102140 156439 102220 156449
rect 114580 156439 114660 156449
rect 114900 156439 114980 156449
rect 115320 156439 115400 156449
rect 115640 156439 115720 156449
rect 101160 156359 101170 156439
rect 101480 156359 101490 156439
rect 101900 156359 101910 156439
rect 102220 156359 102230 156439
rect 114660 156359 114670 156439
rect 114980 156359 114990 156439
rect 115400 156359 115410 156439
rect 115720 156359 115730 156439
rect 116140 156400 116150 156480
rect 116290 156400 116300 156480
rect 100560 156300 100640 156310
rect 100710 156300 100790 156310
rect 100860 156300 100940 156310
rect 116060 156300 116140 156310
rect 116210 156300 116290 156310
rect 100640 156220 100650 156300
rect 100790 156220 100800 156300
rect 100940 156220 100950 156300
rect 101240 156279 101320 156289
rect 101560 156279 101640 156289
rect 101980 156279 102060 156289
rect 102300 156279 102380 156289
rect 114740 156279 114820 156289
rect 115060 156279 115140 156289
rect 115480 156279 115560 156289
rect 115800 156279 115880 156289
rect 101320 156199 101330 156279
rect 101640 156199 101650 156279
rect 102060 156199 102070 156279
rect 102380 156199 102390 156279
rect 114820 156199 114830 156279
rect 115140 156199 115150 156279
rect 115560 156199 115570 156279
rect 115880 156199 115890 156279
rect 116140 156220 116150 156300
rect 116290 156220 116300 156300
rect 100560 156120 100640 156130
rect 100710 156120 100790 156130
rect 100860 156120 100940 156130
rect 100640 156040 100650 156120
rect 100790 156040 100800 156120
rect 100940 156040 100950 156120
rect 101080 156119 101160 156129
rect 101400 156119 101480 156129
rect 101820 156119 101900 156129
rect 102140 156119 102220 156129
rect 114580 156119 114660 156129
rect 114900 156119 114980 156129
rect 115320 156119 115400 156129
rect 115640 156119 115720 156129
rect 116060 156120 116140 156130
rect 116210 156120 116290 156130
rect 101160 156039 101170 156119
rect 101480 156039 101490 156119
rect 101900 156039 101910 156119
rect 102220 156039 102230 156119
rect 114660 156039 114670 156119
rect 114980 156039 114990 156119
rect 115400 156039 115410 156119
rect 115720 156039 115730 156119
rect 116140 156040 116150 156120
rect 116290 156040 116300 156120
rect 101240 155959 101320 155969
rect 101560 155959 101640 155969
rect 101980 155959 102060 155969
rect 102300 155959 102380 155969
rect 114740 155959 114820 155969
rect 115060 155959 115140 155969
rect 115480 155959 115560 155969
rect 115800 155959 115880 155969
rect 100560 155940 100640 155950
rect 100710 155940 100790 155950
rect 100860 155940 100940 155950
rect 100640 155860 100650 155940
rect 100790 155860 100800 155940
rect 100940 155860 100950 155940
rect 101320 155879 101330 155959
rect 101640 155879 101650 155959
rect 102060 155879 102070 155959
rect 102380 155879 102390 155959
rect 114820 155879 114830 155959
rect 115140 155879 115150 155959
rect 115560 155879 115570 155959
rect 115880 155879 115890 155959
rect 116060 155940 116140 155950
rect 116210 155940 116290 155950
rect 116140 155860 116150 155940
rect 116290 155860 116300 155940
rect 101080 155799 101160 155809
rect 101400 155799 101480 155809
rect 101820 155799 101900 155809
rect 102140 155799 102220 155809
rect 114580 155799 114660 155809
rect 114900 155799 114980 155809
rect 115320 155799 115400 155809
rect 115640 155799 115720 155809
rect 100560 155760 100640 155770
rect 100710 155760 100790 155770
rect 100860 155760 100940 155770
rect 100640 155680 100650 155760
rect 100790 155680 100800 155760
rect 100940 155680 100950 155760
rect 101160 155719 101170 155799
rect 101480 155719 101490 155799
rect 101900 155719 101910 155799
rect 102220 155719 102230 155799
rect 114660 155719 114670 155799
rect 114980 155719 114990 155799
rect 115400 155719 115410 155799
rect 115720 155719 115730 155799
rect 116060 155760 116140 155770
rect 116210 155760 116290 155770
rect 116140 155680 116150 155760
rect 116290 155680 116300 155760
rect 101240 155639 101320 155649
rect 101560 155639 101640 155649
rect 101980 155639 102060 155649
rect 102300 155639 102380 155649
rect 114740 155639 114820 155649
rect 115060 155639 115140 155649
rect 115480 155639 115560 155649
rect 115800 155639 115880 155649
rect 100560 155580 100640 155590
rect 100710 155580 100790 155590
rect 100860 155580 100940 155590
rect 100640 155500 100650 155580
rect 100790 155500 100800 155580
rect 100940 155500 100950 155580
rect 101320 155559 101330 155639
rect 101640 155559 101650 155639
rect 102060 155559 102070 155639
rect 102380 155559 102390 155639
rect 114820 155559 114830 155639
rect 115140 155559 115150 155639
rect 115560 155559 115570 155639
rect 115880 155559 115890 155639
rect 116060 155580 116140 155590
rect 116210 155580 116290 155590
rect 116140 155500 116150 155580
rect 116290 155500 116300 155580
rect 101080 155479 101160 155489
rect 101400 155479 101480 155489
rect 101820 155479 101900 155489
rect 102140 155479 102220 155489
rect 114580 155479 114660 155489
rect 114900 155479 114980 155489
rect 115320 155479 115400 155489
rect 115640 155479 115720 155489
rect 100560 155400 100640 155410
rect 100710 155400 100790 155410
rect 100860 155400 100940 155410
rect 100640 155320 100650 155400
rect 100790 155320 100800 155400
rect 100940 155320 100950 155400
rect 101160 155399 101170 155479
rect 101480 155399 101490 155479
rect 101900 155399 101910 155479
rect 102220 155399 102230 155479
rect 114660 155399 114670 155479
rect 114980 155399 114990 155479
rect 115400 155399 115410 155479
rect 115720 155399 115730 155479
rect 116060 155400 116140 155410
rect 116210 155400 116290 155410
rect 101240 155319 101320 155329
rect 101560 155319 101640 155329
rect 101980 155319 102060 155329
rect 102300 155319 102380 155329
rect 114740 155319 114820 155329
rect 115060 155319 115140 155329
rect 115480 155319 115560 155329
rect 115800 155319 115880 155329
rect 116140 155320 116150 155400
rect 116290 155320 116300 155400
rect 101320 155239 101330 155319
rect 101640 155239 101650 155319
rect 102060 155239 102070 155319
rect 102380 155239 102390 155319
rect 114820 155239 114830 155319
rect 115140 155239 115150 155319
rect 115560 155239 115570 155319
rect 115880 155239 115890 155319
rect 100560 155220 100640 155230
rect 100710 155220 100790 155230
rect 100860 155220 100940 155230
rect 116060 155220 116140 155230
rect 116210 155220 116290 155230
rect 100640 155140 100650 155220
rect 100790 155140 100800 155220
rect 100940 155140 100950 155220
rect 101080 155159 101160 155169
rect 101400 155159 101480 155169
rect 101820 155159 101900 155169
rect 102140 155159 102220 155169
rect 114580 155159 114660 155169
rect 114900 155159 114980 155169
rect 115320 155159 115400 155169
rect 115640 155159 115720 155169
rect 101160 155079 101170 155159
rect 101480 155079 101490 155159
rect 101900 155079 101910 155159
rect 102220 155079 102230 155159
rect 114660 155079 114670 155159
rect 114980 155079 114990 155159
rect 115400 155079 115410 155159
rect 115720 155079 115730 155159
rect 116140 155140 116150 155220
rect 116290 155140 116300 155220
rect 100560 155040 100640 155050
rect 100710 155040 100790 155050
rect 100860 155040 100940 155050
rect 116060 155040 116140 155050
rect 116210 155040 116290 155050
rect 100640 154960 100650 155040
rect 100790 154960 100800 155040
rect 100940 154960 100950 155040
rect 101240 154999 101320 155009
rect 101560 154999 101640 155009
rect 101980 154999 102060 155009
rect 102300 154999 102380 155009
rect 114740 154999 114820 155009
rect 115060 154999 115140 155009
rect 115480 154999 115560 155009
rect 115800 154999 115880 155009
rect 101320 154919 101330 154999
rect 101640 154919 101650 154999
rect 102060 154919 102070 154999
rect 102380 154919 102390 154999
rect 114820 154919 114830 154999
rect 115140 154919 115150 154999
rect 115560 154919 115570 154999
rect 115880 154919 115890 154999
rect 116140 154960 116150 155040
rect 116290 154960 116300 155040
rect 100560 154860 100640 154870
rect 100710 154860 100790 154870
rect 100860 154860 100940 154870
rect 116060 154860 116140 154870
rect 116210 154860 116290 154870
rect 100640 154780 100650 154860
rect 100790 154780 100800 154860
rect 100940 154780 100950 154860
rect 101080 154839 101160 154849
rect 101400 154839 101480 154849
rect 101820 154839 101900 154849
rect 102140 154839 102220 154849
rect 114580 154839 114660 154849
rect 114900 154839 114980 154849
rect 115320 154839 115400 154849
rect 115640 154839 115720 154849
rect 101160 154759 101170 154839
rect 101480 154759 101490 154839
rect 101900 154759 101910 154839
rect 102220 154759 102230 154839
rect 114660 154759 114670 154839
rect 114980 154759 114990 154839
rect 115400 154759 115410 154839
rect 115720 154759 115730 154839
rect 116140 154780 116150 154860
rect 116290 154780 116300 154860
rect 100560 154680 100640 154690
rect 100710 154680 100790 154690
rect 100860 154680 100940 154690
rect 100640 154600 100650 154680
rect 100790 154600 100800 154680
rect 100940 154600 100950 154680
rect 101240 154679 101320 154689
rect 101560 154679 101640 154689
rect 101980 154679 102060 154689
rect 102300 154679 102380 154689
rect 114740 154679 114820 154689
rect 115060 154679 115140 154689
rect 115480 154679 115560 154689
rect 115800 154679 115880 154689
rect 116060 154680 116140 154690
rect 116210 154680 116290 154690
rect 101320 154599 101330 154679
rect 101640 154599 101650 154679
rect 102060 154599 102070 154679
rect 102380 154599 102390 154679
rect 114820 154599 114830 154679
rect 115140 154599 115150 154679
rect 115560 154599 115570 154679
rect 115880 154599 115890 154679
rect 116140 154600 116150 154680
rect 116290 154600 116300 154680
rect 101080 154519 101160 154529
rect 101400 154519 101480 154529
rect 101820 154519 101900 154529
rect 102140 154519 102220 154529
rect 114580 154519 114660 154529
rect 114900 154519 114980 154529
rect 115320 154519 115400 154529
rect 115640 154519 115720 154529
rect 100560 154500 100640 154510
rect 100710 154500 100790 154510
rect 100860 154500 100940 154510
rect 100640 154420 100650 154500
rect 100790 154420 100800 154500
rect 100940 154420 100950 154500
rect 101160 154439 101170 154519
rect 101480 154439 101490 154519
rect 101900 154439 101910 154519
rect 102220 154439 102230 154519
rect 114660 154439 114670 154519
rect 114980 154439 114990 154519
rect 115400 154439 115410 154519
rect 115720 154439 115730 154519
rect 116060 154500 116140 154510
rect 116210 154500 116290 154510
rect 116140 154420 116150 154500
rect 116290 154420 116300 154500
rect 101240 154359 101320 154369
rect 101560 154359 101640 154369
rect 101980 154359 102060 154369
rect 102300 154359 102380 154369
rect 114740 154359 114820 154369
rect 115060 154359 115140 154369
rect 115480 154359 115560 154369
rect 115800 154359 115880 154369
rect 100560 154320 100640 154330
rect 100710 154320 100790 154330
rect 100860 154320 100940 154330
rect 100640 154240 100650 154320
rect 100790 154240 100800 154320
rect 100940 154240 100950 154320
rect 101320 154279 101330 154359
rect 101640 154279 101650 154359
rect 102060 154279 102070 154359
rect 102380 154279 102390 154359
rect 114820 154279 114830 154359
rect 115140 154279 115150 154359
rect 115560 154279 115570 154359
rect 115880 154279 115890 154359
rect 116060 154320 116140 154330
rect 116210 154320 116290 154330
rect 116140 154240 116150 154320
rect 116290 154240 116300 154320
rect 101080 154199 101160 154209
rect 101400 154199 101480 154209
rect 101820 154199 101900 154209
rect 102140 154199 102220 154209
rect 114580 154199 114660 154209
rect 114900 154199 114980 154209
rect 115320 154199 115400 154209
rect 115640 154199 115720 154209
rect 100560 154140 100640 154150
rect 100710 154140 100790 154150
rect 100860 154140 100940 154150
rect 100640 154060 100650 154140
rect 100790 154060 100800 154140
rect 100940 154060 100950 154140
rect 101160 154119 101170 154199
rect 101480 154119 101490 154199
rect 101900 154119 101910 154199
rect 102220 154119 102230 154199
rect 114660 154119 114670 154199
rect 114980 154119 114990 154199
rect 115400 154119 115410 154199
rect 115720 154119 115730 154199
rect 116060 154140 116140 154150
rect 116210 154140 116290 154150
rect 116140 154060 116150 154140
rect 116290 154060 116300 154140
rect 101240 154039 101320 154049
rect 101560 154039 101640 154049
rect 101980 154039 102060 154049
rect 102300 154039 102380 154049
rect 114740 154039 114820 154049
rect 115060 154039 115140 154049
rect 115480 154039 115560 154049
rect 115800 154039 115880 154049
rect 100560 153960 100640 153970
rect 100710 153960 100790 153970
rect 100860 153960 100940 153970
rect 100640 153880 100650 153960
rect 100790 153880 100800 153960
rect 100940 153880 100950 153960
rect 101320 153959 101330 154039
rect 101640 153959 101650 154039
rect 102060 153959 102070 154039
rect 102380 153959 102390 154039
rect 114820 153959 114830 154039
rect 115140 153959 115150 154039
rect 115560 153959 115570 154039
rect 115880 153959 115890 154039
rect 116060 153960 116140 153970
rect 116210 153960 116290 153970
rect 101080 153879 101160 153889
rect 101400 153879 101480 153889
rect 101820 153879 101900 153889
rect 102140 153879 102220 153889
rect 114580 153879 114660 153889
rect 114900 153879 114980 153889
rect 115320 153879 115400 153889
rect 115640 153879 115720 153889
rect 116140 153880 116150 153960
rect 116290 153880 116300 153960
rect 101160 153799 101170 153879
rect 101480 153799 101490 153879
rect 101900 153799 101910 153879
rect 102220 153799 102230 153879
rect 114660 153799 114670 153879
rect 114980 153799 114990 153879
rect 115400 153799 115410 153879
rect 115720 153799 115730 153879
rect 100560 153780 100640 153790
rect 100710 153780 100790 153790
rect 100860 153780 100940 153790
rect 116060 153780 116140 153790
rect 116210 153780 116290 153790
rect 100640 153700 100650 153780
rect 100790 153700 100800 153780
rect 100940 153700 100950 153780
rect 101240 153719 101320 153729
rect 101560 153719 101640 153729
rect 101980 153719 102060 153729
rect 102300 153719 102380 153729
rect 114740 153719 114820 153729
rect 115060 153719 115140 153729
rect 115480 153719 115560 153729
rect 115800 153719 115880 153729
rect 101320 153639 101330 153719
rect 101640 153639 101650 153719
rect 102060 153639 102070 153719
rect 102380 153639 102390 153719
rect 114820 153639 114830 153719
rect 115140 153639 115150 153719
rect 115560 153639 115570 153719
rect 115880 153639 115890 153719
rect 116140 153700 116150 153780
rect 116290 153700 116300 153780
rect 100560 153600 100640 153610
rect 100710 153600 100790 153610
rect 100860 153600 100940 153610
rect 116060 153600 116140 153610
rect 116210 153600 116290 153610
rect 100640 153520 100650 153600
rect 100790 153520 100800 153600
rect 100940 153520 100950 153600
rect 101080 153559 101160 153569
rect 101400 153559 101480 153569
rect 101820 153559 101900 153569
rect 102140 153559 102220 153569
rect 114580 153559 114660 153569
rect 114900 153559 114980 153569
rect 115320 153559 115400 153569
rect 115640 153559 115720 153569
rect 101160 153479 101170 153559
rect 101480 153479 101490 153559
rect 101900 153479 101910 153559
rect 102220 153479 102230 153559
rect 114660 153479 114670 153559
rect 114980 153479 114990 153559
rect 115400 153479 115410 153559
rect 115720 153479 115730 153559
rect 116140 153520 116150 153600
rect 116290 153520 116300 153600
rect 100560 153420 100640 153430
rect 100710 153420 100790 153430
rect 100860 153420 100940 153430
rect 116060 153420 116140 153430
rect 116210 153420 116290 153430
rect 100640 153340 100650 153420
rect 100790 153340 100800 153420
rect 100940 153340 100950 153420
rect 101240 153399 101320 153409
rect 101560 153399 101640 153409
rect 101980 153399 102060 153409
rect 102300 153399 102380 153409
rect 114740 153399 114820 153409
rect 115060 153399 115140 153409
rect 115480 153399 115560 153409
rect 115800 153399 115880 153409
rect 101320 153319 101330 153399
rect 101640 153319 101650 153399
rect 102060 153319 102070 153399
rect 102380 153319 102390 153399
rect 114820 153319 114830 153399
rect 115140 153319 115150 153399
rect 115560 153319 115570 153399
rect 115880 153319 115890 153399
rect 116140 153340 116150 153420
rect 116290 153340 116300 153420
rect 100560 153240 100640 153250
rect 100710 153240 100790 153250
rect 100860 153240 100940 153250
rect 100640 153160 100650 153240
rect 100790 153160 100800 153240
rect 100940 153160 100950 153240
rect 101080 153239 101160 153249
rect 101400 153239 101480 153249
rect 101820 153239 101900 153249
rect 102140 153239 102220 153249
rect 114580 153239 114660 153249
rect 114900 153239 114980 153249
rect 115320 153239 115400 153249
rect 115640 153239 115720 153249
rect 116060 153240 116140 153250
rect 116210 153240 116290 153250
rect 101160 153159 101170 153239
rect 101480 153159 101490 153239
rect 101900 153159 101910 153239
rect 102220 153159 102230 153239
rect 114660 153159 114670 153239
rect 114980 153159 114990 153239
rect 115400 153159 115410 153239
rect 115720 153159 115730 153239
rect 116140 153160 116150 153240
rect 116290 153160 116300 153240
rect 101240 153079 101320 153089
rect 101560 153079 101640 153089
rect 101980 153079 102060 153089
rect 102300 153079 102380 153089
rect 114740 153079 114820 153089
rect 115060 153079 115140 153089
rect 115480 153079 115560 153089
rect 115800 153079 115880 153089
rect 100560 153060 100640 153070
rect 100710 153060 100790 153070
rect 100860 153060 100940 153070
rect 100640 152980 100650 153060
rect 100790 152980 100800 153060
rect 100940 152980 100950 153060
rect 101320 152999 101330 153079
rect 101640 152999 101650 153079
rect 102060 152999 102070 153079
rect 102380 152999 102390 153079
rect 114820 152999 114830 153079
rect 115140 152999 115150 153079
rect 115560 152999 115570 153079
rect 115880 152999 115890 153079
rect 116060 153060 116140 153070
rect 116210 153060 116290 153070
rect 116140 152980 116150 153060
rect 116290 152980 116300 153060
rect 101080 152919 101160 152929
rect 101400 152919 101480 152929
rect 101820 152919 101900 152929
rect 102140 152919 102220 152929
rect 114580 152919 114660 152929
rect 114900 152919 114980 152929
rect 115320 152919 115400 152929
rect 115640 152919 115720 152929
rect 89060 152880 89140 152890
rect 89210 152880 89290 152890
rect 100560 152880 100640 152890
rect 100710 152880 100790 152890
rect 100860 152880 100940 152890
rect 89140 152800 89150 152880
rect 89290 152800 89300 152880
rect 100640 152800 100650 152880
rect 100790 152800 100800 152880
rect 100940 152800 100950 152880
rect 101160 152839 101170 152919
rect 101480 152839 101490 152919
rect 101900 152839 101910 152919
rect 102220 152839 102230 152919
rect 114660 152839 114670 152919
rect 114980 152839 114990 152919
rect 115400 152839 115410 152919
rect 115720 152839 115730 152919
rect 127245 152900 127260 158990
rect 127640 158920 127650 159000
rect 127790 158920 127800 159000
rect 127940 158920 127950 159000
rect 128080 158999 128160 159009
rect 128400 158999 128480 159009
rect 128820 158999 128900 159009
rect 129140 158999 129220 159009
rect 129560 159000 129640 159010
rect 129710 159000 129790 159010
rect 141060 159000 141140 159010
rect 141210 159000 141290 159010
rect 141360 159000 141440 159010
rect 141545 159000 141625 159010
rect 141865 159000 141945 159010
rect 142185 159000 142200 159010
rect 145385 159000 145465 159010
rect 145705 159000 145785 159010
rect 146025 159000 146105 159010
rect 128160 158919 128170 158999
rect 128480 158919 128490 158999
rect 128900 158919 128910 158999
rect 129220 158919 129230 158999
rect 129640 158920 129650 159000
rect 129790 158920 129800 159000
rect 130240 158900 130255 158990
rect 128240 158839 128320 158849
rect 128560 158839 128640 158849
rect 128980 158839 129060 158849
rect 129300 158839 129380 158849
rect 127560 158820 127640 158830
rect 127710 158820 127790 158830
rect 127860 158820 127940 158830
rect 127640 158740 127650 158820
rect 127790 158740 127800 158820
rect 127940 158740 127950 158820
rect 128320 158759 128330 158839
rect 128640 158759 128650 158839
rect 129060 158759 129070 158839
rect 129380 158759 129390 158839
rect 129560 158820 129640 158830
rect 129710 158820 129790 158830
rect 129640 158740 129650 158820
rect 129790 158740 129800 158820
rect 128080 158679 128160 158689
rect 128400 158679 128480 158689
rect 128820 158679 128900 158689
rect 129140 158679 129220 158689
rect 127560 158640 127640 158650
rect 127710 158640 127790 158650
rect 127860 158640 127940 158650
rect 127640 158560 127650 158640
rect 127790 158560 127800 158640
rect 127940 158560 127950 158640
rect 128160 158599 128170 158679
rect 128480 158599 128490 158679
rect 128900 158599 128910 158679
rect 129220 158599 129230 158679
rect 129560 158640 129640 158650
rect 129710 158640 129790 158650
rect 129640 158560 129650 158640
rect 129790 158560 129800 158640
rect 128240 158519 128320 158529
rect 128560 158519 128640 158529
rect 128980 158519 129060 158529
rect 129300 158519 129380 158529
rect 127560 158460 127640 158470
rect 127710 158460 127790 158470
rect 127860 158460 127940 158470
rect 127640 158380 127650 158460
rect 127790 158380 127800 158460
rect 127940 158380 127950 158460
rect 128320 158439 128330 158519
rect 128640 158439 128650 158519
rect 129060 158439 129070 158519
rect 129380 158439 129390 158519
rect 129560 158460 129640 158470
rect 129710 158460 129790 158470
rect 129640 158380 129650 158460
rect 129790 158380 129800 158460
rect 128080 158359 128160 158369
rect 128400 158359 128480 158369
rect 128820 158359 128900 158369
rect 129140 158359 129220 158369
rect 127560 158280 127640 158290
rect 127710 158280 127790 158290
rect 127860 158280 127940 158290
rect 127640 158200 127650 158280
rect 127790 158200 127800 158280
rect 127940 158200 127950 158280
rect 128160 158279 128170 158359
rect 128480 158279 128490 158359
rect 128900 158279 128910 158359
rect 129220 158279 129230 158359
rect 129560 158280 129640 158290
rect 129710 158280 129790 158290
rect 128240 158199 128320 158209
rect 128560 158199 128640 158209
rect 128980 158199 129060 158209
rect 129300 158199 129380 158209
rect 129640 158200 129650 158280
rect 129790 158200 129800 158280
rect 128320 158119 128330 158199
rect 128640 158119 128650 158199
rect 129060 158119 129070 158199
rect 129380 158119 129390 158199
rect 127560 158100 127640 158110
rect 127710 158100 127790 158110
rect 127860 158100 127940 158110
rect 129560 158100 129640 158110
rect 129710 158100 129790 158110
rect 127640 158020 127650 158100
rect 127790 158020 127800 158100
rect 127940 158020 127950 158100
rect 128080 158039 128160 158049
rect 128400 158039 128480 158049
rect 128820 158039 128900 158049
rect 129140 158039 129220 158049
rect 128160 157959 128170 158039
rect 128480 157959 128490 158039
rect 128900 157959 128910 158039
rect 129220 157959 129230 158039
rect 129640 158020 129650 158100
rect 129790 158020 129800 158100
rect 127560 157920 127640 157930
rect 127710 157920 127790 157930
rect 127860 157920 127940 157930
rect 129560 157920 129640 157930
rect 129710 157920 129790 157930
rect 127640 157840 127650 157920
rect 127790 157840 127800 157920
rect 127940 157840 127950 157920
rect 128240 157879 128320 157889
rect 128560 157879 128640 157889
rect 128980 157879 129060 157889
rect 129300 157879 129380 157889
rect 128320 157799 128330 157879
rect 128640 157799 128650 157879
rect 129060 157799 129070 157879
rect 129380 157799 129390 157879
rect 129640 157840 129650 157920
rect 129790 157840 129800 157920
rect 127560 157740 127640 157750
rect 127710 157740 127790 157750
rect 127860 157740 127940 157750
rect 129560 157740 129640 157750
rect 129710 157740 129790 157750
rect 127640 157660 127650 157740
rect 127790 157660 127800 157740
rect 127940 157660 127950 157740
rect 128080 157719 128160 157729
rect 128400 157719 128480 157729
rect 128820 157719 128900 157729
rect 129140 157719 129220 157729
rect 128160 157639 128170 157719
rect 128480 157639 128490 157719
rect 128900 157639 128910 157719
rect 129220 157639 129230 157719
rect 129640 157660 129650 157740
rect 129790 157660 129800 157740
rect 127560 157560 127640 157570
rect 127710 157560 127790 157570
rect 127860 157560 127940 157570
rect 127640 157480 127650 157560
rect 127790 157480 127800 157560
rect 127940 157480 127950 157560
rect 128240 157559 128320 157569
rect 128560 157559 128640 157569
rect 128980 157559 129060 157569
rect 129300 157559 129380 157569
rect 129560 157560 129640 157570
rect 129710 157560 129790 157570
rect 128320 157479 128330 157559
rect 128640 157479 128650 157559
rect 129060 157479 129070 157559
rect 129380 157479 129390 157559
rect 129640 157480 129650 157560
rect 129790 157480 129800 157560
rect 128080 157399 128160 157409
rect 128400 157399 128480 157409
rect 128820 157399 128900 157409
rect 129140 157399 129220 157409
rect 127560 157380 127640 157390
rect 127710 157380 127790 157390
rect 127860 157380 127940 157390
rect 127640 157300 127650 157380
rect 127790 157300 127800 157380
rect 127940 157300 127950 157380
rect 128160 157319 128170 157399
rect 128480 157319 128490 157399
rect 128900 157319 128910 157399
rect 129220 157319 129230 157399
rect 129560 157380 129640 157390
rect 129710 157380 129790 157390
rect 129640 157300 129650 157380
rect 129790 157300 129800 157380
rect 128240 157239 128320 157249
rect 128560 157239 128640 157249
rect 128980 157239 129060 157249
rect 129300 157239 129380 157249
rect 127560 157200 127640 157210
rect 127710 157200 127790 157210
rect 127860 157200 127940 157210
rect 127640 157120 127650 157200
rect 127790 157120 127800 157200
rect 127940 157120 127950 157200
rect 128320 157159 128330 157239
rect 128640 157159 128650 157239
rect 129060 157159 129070 157239
rect 129380 157159 129390 157239
rect 129560 157200 129640 157210
rect 129710 157200 129790 157210
rect 129640 157120 129650 157200
rect 129790 157120 129800 157200
rect 128080 157079 128160 157089
rect 128400 157079 128480 157089
rect 128820 157079 128900 157089
rect 129140 157079 129220 157089
rect 127560 157020 127640 157030
rect 127710 157020 127790 157030
rect 127860 157020 127940 157030
rect 127640 156940 127650 157020
rect 127790 156940 127800 157020
rect 127940 156940 127950 157020
rect 128160 156999 128170 157079
rect 128480 156999 128490 157079
rect 128900 156999 128910 157079
rect 129220 156999 129230 157079
rect 129560 157020 129640 157030
rect 129710 157020 129790 157030
rect 129640 156940 129650 157020
rect 129790 156940 129800 157020
rect 128240 156919 128320 156929
rect 128560 156919 128640 156929
rect 128980 156919 129060 156929
rect 129300 156919 129380 156929
rect 127560 156840 127640 156850
rect 127710 156840 127790 156850
rect 127860 156840 127940 156850
rect 127640 156760 127650 156840
rect 127790 156760 127800 156840
rect 127940 156760 127950 156840
rect 128320 156839 128330 156919
rect 128640 156839 128650 156919
rect 129060 156839 129070 156919
rect 129380 156839 129390 156919
rect 129560 156840 129640 156850
rect 129710 156840 129790 156850
rect 128080 156759 128160 156769
rect 128400 156759 128480 156769
rect 128820 156759 128900 156769
rect 129140 156759 129220 156769
rect 129640 156760 129650 156840
rect 129790 156760 129800 156840
rect 128160 156679 128170 156759
rect 128480 156679 128490 156759
rect 128900 156679 128910 156759
rect 129220 156679 129230 156759
rect 127560 156660 127640 156670
rect 127710 156660 127790 156670
rect 127860 156660 127940 156670
rect 129560 156660 129640 156670
rect 129710 156660 129790 156670
rect 127640 156580 127650 156660
rect 127790 156580 127800 156660
rect 127940 156580 127950 156660
rect 128240 156599 128320 156609
rect 128560 156599 128640 156609
rect 128980 156599 129060 156609
rect 129300 156599 129380 156609
rect 128320 156519 128330 156599
rect 128640 156519 128650 156599
rect 129060 156519 129070 156599
rect 129380 156519 129390 156599
rect 129640 156580 129650 156660
rect 129790 156580 129800 156660
rect 127560 156480 127640 156490
rect 127710 156480 127790 156490
rect 127860 156480 127940 156490
rect 129560 156480 129640 156490
rect 129710 156480 129790 156490
rect 127640 156400 127650 156480
rect 127790 156400 127800 156480
rect 127940 156400 127950 156480
rect 128080 156439 128160 156449
rect 128400 156439 128480 156449
rect 128820 156439 128900 156449
rect 129140 156439 129220 156449
rect 128160 156359 128170 156439
rect 128480 156359 128490 156439
rect 128900 156359 128910 156439
rect 129220 156359 129230 156439
rect 129640 156400 129650 156480
rect 129790 156400 129800 156480
rect 127560 156300 127640 156310
rect 127710 156300 127790 156310
rect 127860 156300 127940 156310
rect 129560 156300 129640 156310
rect 129710 156300 129790 156310
rect 127640 156220 127650 156300
rect 127790 156220 127800 156300
rect 127940 156220 127950 156300
rect 128240 156279 128320 156289
rect 128560 156279 128640 156289
rect 128980 156279 129060 156289
rect 129300 156279 129380 156289
rect 128320 156199 128330 156279
rect 128640 156199 128650 156279
rect 129060 156199 129070 156279
rect 129380 156199 129390 156279
rect 129640 156220 129650 156300
rect 129790 156220 129800 156300
rect 127560 156120 127640 156130
rect 127710 156120 127790 156130
rect 127860 156120 127940 156130
rect 127640 156040 127650 156120
rect 127790 156040 127800 156120
rect 127940 156040 127950 156120
rect 128080 156119 128160 156129
rect 128400 156119 128480 156129
rect 128820 156119 128900 156129
rect 129140 156119 129220 156129
rect 129560 156120 129640 156130
rect 129710 156120 129790 156130
rect 128160 156039 128170 156119
rect 128480 156039 128490 156119
rect 128900 156039 128910 156119
rect 129220 156039 129230 156119
rect 129640 156040 129650 156120
rect 129790 156040 129800 156120
rect 128240 155959 128320 155969
rect 128560 155959 128640 155969
rect 128980 155959 129060 155969
rect 129300 155959 129380 155969
rect 127560 155940 127640 155950
rect 127710 155940 127790 155950
rect 127860 155940 127940 155950
rect 127640 155860 127650 155940
rect 127790 155860 127800 155940
rect 127940 155860 127950 155940
rect 128320 155879 128330 155959
rect 128640 155879 128650 155959
rect 129060 155879 129070 155959
rect 129380 155879 129390 155959
rect 129560 155940 129640 155950
rect 129710 155940 129790 155950
rect 129640 155860 129650 155940
rect 129790 155860 129800 155940
rect 128080 155799 128160 155809
rect 128400 155799 128480 155809
rect 128820 155799 128900 155809
rect 129140 155799 129220 155809
rect 127560 155760 127640 155770
rect 127710 155760 127790 155770
rect 127860 155760 127940 155770
rect 127640 155680 127650 155760
rect 127790 155680 127800 155760
rect 127940 155680 127950 155760
rect 128160 155719 128170 155799
rect 128480 155719 128490 155799
rect 128900 155719 128910 155799
rect 129220 155719 129230 155799
rect 129560 155760 129640 155770
rect 129710 155760 129790 155770
rect 129640 155680 129650 155760
rect 129790 155680 129800 155760
rect 128240 155639 128320 155649
rect 128560 155639 128640 155649
rect 128980 155639 129060 155649
rect 129300 155639 129380 155649
rect 127560 155580 127640 155590
rect 127710 155580 127790 155590
rect 127860 155580 127940 155590
rect 127640 155500 127650 155580
rect 127790 155500 127800 155580
rect 127940 155500 127950 155580
rect 128320 155559 128330 155639
rect 128640 155559 128650 155639
rect 129060 155559 129070 155639
rect 129380 155559 129390 155639
rect 129560 155580 129640 155590
rect 129710 155580 129790 155590
rect 129640 155500 129650 155580
rect 129790 155500 129800 155580
rect 128080 155479 128160 155489
rect 128400 155479 128480 155489
rect 128820 155479 128900 155489
rect 129140 155479 129220 155489
rect 127560 155400 127640 155410
rect 127710 155400 127790 155410
rect 127860 155400 127940 155410
rect 127640 155320 127650 155400
rect 127790 155320 127800 155400
rect 127940 155320 127950 155400
rect 128160 155399 128170 155479
rect 128480 155399 128490 155479
rect 128900 155399 128910 155479
rect 129220 155399 129230 155479
rect 129560 155400 129640 155410
rect 129710 155400 129790 155410
rect 128240 155319 128320 155329
rect 128560 155319 128640 155329
rect 128980 155319 129060 155329
rect 129300 155319 129380 155329
rect 129640 155320 129650 155400
rect 129790 155320 129800 155400
rect 128320 155239 128330 155319
rect 128640 155239 128650 155319
rect 129060 155239 129070 155319
rect 129380 155239 129390 155319
rect 127560 155220 127640 155230
rect 127710 155220 127790 155230
rect 127860 155220 127940 155230
rect 129560 155220 129640 155230
rect 129710 155220 129790 155230
rect 127640 155140 127650 155220
rect 127790 155140 127800 155220
rect 127940 155140 127950 155220
rect 128080 155159 128160 155169
rect 128400 155159 128480 155169
rect 128820 155159 128900 155169
rect 129140 155159 129220 155169
rect 128160 155079 128170 155159
rect 128480 155079 128490 155159
rect 128900 155079 128910 155159
rect 129220 155079 129230 155159
rect 129640 155140 129650 155220
rect 129790 155140 129800 155220
rect 127560 155040 127640 155050
rect 127710 155040 127790 155050
rect 127860 155040 127940 155050
rect 129560 155040 129640 155050
rect 129710 155040 129790 155050
rect 127640 154960 127650 155040
rect 127790 154960 127800 155040
rect 127940 154960 127950 155040
rect 128240 154999 128320 155009
rect 128560 154999 128640 155009
rect 128980 154999 129060 155009
rect 129300 154999 129380 155009
rect 128320 154919 128330 154999
rect 128640 154919 128650 154999
rect 129060 154919 129070 154999
rect 129380 154919 129390 154999
rect 129640 154960 129650 155040
rect 129790 154960 129800 155040
rect 127560 154860 127640 154870
rect 127710 154860 127790 154870
rect 127860 154860 127940 154870
rect 129560 154860 129640 154870
rect 129710 154860 129790 154870
rect 127640 154780 127650 154860
rect 127790 154780 127800 154860
rect 127940 154780 127950 154860
rect 128080 154839 128160 154849
rect 128400 154839 128480 154849
rect 128820 154839 128900 154849
rect 129140 154839 129220 154849
rect 128160 154759 128170 154839
rect 128480 154759 128490 154839
rect 128900 154759 128910 154839
rect 129220 154759 129230 154839
rect 129640 154780 129650 154860
rect 129790 154780 129800 154860
rect 127560 154680 127640 154690
rect 127710 154680 127790 154690
rect 127860 154680 127940 154690
rect 127640 154600 127650 154680
rect 127790 154600 127800 154680
rect 127940 154600 127950 154680
rect 128240 154679 128320 154689
rect 128560 154679 128640 154689
rect 128980 154679 129060 154689
rect 129300 154679 129380 154689
rect 129560 154680 129640 154690
rect 129710 154680 129790 154690
rect 128320 154599 128330 154679
rect 128640 154599 128650 154679
rect 129060 154599 129070 154679
rect 129380 154599 129390 154679
rect 129640 154600 129650 154680
rect 129790 154600 129800 154680
rect 128080 154519 128160 154529
rect 128400 154519 128480 154529
rect 128820 154519 128900 154529
rect 129140 154519 129220 154529
rect 127560 154500 127640 154510
rect 127710 154500 127790 154510
rect 127860 154500 127940 154510
rect 127640 154420 127650 154500
rect 127790 154420 127800 154500
rect 127940 154420 127950 154500
rect 128160 154439 128170 154519
rect 128480 154439 128490 154519
rect 128900 154439 128910 154519
rect 129220 154439 129230 154519
rect 129560 154500 129640 154510
rect 129710 154500 129790 154510
rect 129640 154420 129650 154500
rect 129790 154420 129800 154500
rect 128240 154359 128320 154369
rect 128560 154359 128640 154369
rect 128980 154359 129060 154369
rect 129300 154359 129380 154369
rect 127560 154320 127640 154330
rect 127710 154320 127790 154330
rect 127860 154320 127940 154330
rect 127640 154240 127650 154320
rect 127790 154240 127800 154320
rect 127940 154240 127950 154320
rect 128320 154279 128330 154359
rect 128640 154279 128650 154359
rect 129060 154279 129070 154359
rect 129380 154279 129390 154359
rect 129560 154320 129640 154330
rect 129710 154320 129790 154330
rect 129640 154240 129650 154320
rect 129790 154240 129800 154320
rect 128080 154199 128160 154209
rect 128400 154199 128480 154209
rect 128820 154199 128900 154209
rect 129140 154199 129220 154209
rect 127560 154140 127640 154150
rect 127710 154140 127790 154150
rect 127860 154140 127940 154150
rect 127640 154060 127650 154140
rect 127790 154060 127800 154140
rect 127940 154060 127950 154140
rect 128160 154119 128170 154199
rect 128480 154119 128490 154199
rect 128900 154119 128910 154199
rect 129220 154119 129230 154199
rect 129560 154140 129640 154150
rect 129710 154140 129790 154150
rect 129640 154060 129650 154140
rect 129790 154060 129800 154140
rect 128240 154039 128320 154049
rect 128560 154039 128640 154049
rect 128980 154039 129060 154049
rect 129300 154039 129380 154049
rect 127560 153960 127640 153970
rect 127710 153960 127790 153970
rect 127860 153960 127940 153970
rect 127640 153880 127650 153960
rect 127790 153880 127800 153960
rect 127940 153880 127950 153960
rect 128320 153959 128330 154039
rect 128640 153959 128650 154039
rect 129060 153959 129070 154039
rect 129380 153959 129390 154039
rect 129560 153960 129640 153970
rect 129710 153960 129790 153970
rect 128080 153879 128160 153889
rect 128400 153879 128480 153889
rect 128820 153879 128900 153889
rect 129140 153879 129220 153889
rect 129640 153880 129650 153960
rect 129790 153880 129800 153960
rect 128160 153799 128170 153879
rect 128480 153799 128490 153879
rect 128900 153799 128910 153879
rect 129220 153799 129230 153879
rect 127560 153780 127640 153790
rect 127710 153780 127790 153790
rect 127860 153780 127940 153790
rect 129560 153780 129640 153790
rect 129710 153780 129790 153790
rect 127640 153700 127650 153780
rect 127790 153700 127800 153780
rect 127940 153700 127950 153780
rect 128240 153719 128320 153729
rect 128560 153719 128640 153729
rect 128980 153719 129060 153729
rect 129300 153719 129380 153729
rect 128320 153639 128330 153719
rect 128640 153639 128650 153719
rect 129060 153639 129070 153719
rect 129380 153639 129390 153719
rect 129640 153700 129650 153780
rect 129790 153700 129800 153780
rect 127560 153600 127640 153610
rect 127710 153600 127790 153610
rect 127860 153600 127940 153610
rect 129560 153600 129640 153610
rect 129710 153600 129790 153610
rect 127640 153520 127650 153600
rect 127790 153520 127800 153600
rect 127940 153520 127950 153600
rect 128080 153559 128160 153569
rect 128400 153559 128480 153569
rect 128820 153559 128900 153569
rect 129140 153559 129220 153569
rect 128160 153479 128170 153559
rect 128480 153479 128490 153559
rect 128900 153479 128910 153559
rect 129220 153479 129230 153559
rect 129640 153520 129650 153600
rect 129790 153520 129800 153600
rect 127560 153420 127640 153430
rect 127710 153420 127790 153430
rect 127860 153420 127940 153430
rect 129560 153420 129640 153430
rect 129710 153420 129790 153430
rect 127640 153340 127650 153420
rect 127790 153340 127800 153420
rect 127940 153340 127950 153420
rect 128240 153399 128320 153409
rect 128560 153399 128640 153409
rect 128980 153399 129060 153409
rect 129300 153399 129380 153409
rect 128320 153319 128330 153399
rect 128640 153319 128650 153399
rect 129060 153319 129070 153399
rect 129380 153319 129390 153399
rect 129640 153340 129650 153420
rect 129790 153340 129800 153420
rect 127560 153240 127640 153250
rect 127710 153240 127790 153250
rect 127860 153240 127940 153250
rect 127640 153160 127650 153240
rect 127790 153160 127800 153240
rect 127940 153160 127950 153240
rect 128080 153239 128160 153249
rect 128400 153239 128480 153249
rect 128820 153239 128900 153249
rect 129140 153239 129220 153249
rect 129560 153240 129640 153250
rect 129710 153240 129790 153250
rect 128160 153159 128170 153239
rect 128480 153159 128490 153239
rect 128900 153159 128910 153239
rect 129220 153159 129230 153239
rect 129640 153160 129650 153240
rect 129790 153160 129800 153240
rect 128240 153079 128320 153089
rect 128560 153079 128640 153089
rect 128980 153079 129060 153089
rect 129300 153079 129380 153089
rect 127560 153060 127640 153070
rect 127710 153060 127790 153070
rect 127860 153060 127940 153070
rect 127640 152980 127650 153060
rect 127790 152980 127800 153060
rect 127940 152980 127950 153060
rect 128320 152999 128330 153079
rect 128640 152999 128650 153079
rect 129060 152999 129070 153079
rect 129380 152999 129390 153079
rect 129560 153060 129640 153070
rect 129710 153060 129790 153070
rect 129640 152980 129650 153060
rect 129790 152980 129800 153060
rect 128080 152919 128160 152929
rect 128400 152919 128480 152929
rect 128820 152919 128900 152929
rect 129140 152919 129220 152929
rect 116060 152880 116140 152890
rect 116210 152880 116290 152890
rect 127560 152880 127640 152890
rect 127710 152880 127790 152890
rect 127860 152880 127940 152890
rect 116140 152800 116150 152880
rect 116290 152800 116300 152880
rect 127640 152800 127650 152880
rect 127790 152800 127800 152880
rect 127940 152800 127950 152880
rect 128160 152839 128170 152919
rect 128480 152839 128490 152919
rect 128900 152839 128910 152919
rect 129220 152839 129230 152919
rect 140710 152900 140760 158990
rect 141140 158920 141150 159000
rect 141290 158920 141300 159000
rect 141440 158920 141450 159000
rect 141625 158920 141635 159000
rect 141945 158920 141955 159000
rect 145465 158920 145475 159000
rect 145785 158920 145795 159000
rect 146105 158920 146115 159000
rect 146700 158940 146780 158950
rect 146780 158860 146790 158940
rect 141705 158840 141785 158850
rect 142025 158840 142105 158850
rect 145225 158840 145305 158850
rect 145545 158840 145625 158850
rect 145865 158840 145945 158850
rect 141060 158820 141140 158830
rect 141210 158820 141290 158830
rect 141360 158820 141440 158830
rect 141140 158740 141150 158820
rect 141290 158740 141300 158820
rect 141440 158740 141450 158820
rect 141785 158760 141795 158840
rect 142105 158760 142115 158840
rect 145305 158760 145315 158840
rect 145625 158760 145635 158840
rect 145945 158760 145955 158840
rect 146540 158780 146620 158790
rect 146860 158780 146940 158790
rect 146620 158700 146630 158780
rect 146940 158700 146950 158780
rect 141545 158680 141625 158690
rect 141865 158680 141945 158690
rect 142185 158680 142200 158690
rect 145385 158680 145465 158690
rect 145705 158680 145785 158690
rect 146025 158680 146105 158690
rect 141060 158640 141140 158650
rect 141210 158640 141290 158650
rect 141360 158640 141440 158650
rect 141140 158560 141150 158640
rect 141290 158560 141300 158640
rect 141440 158560 141450 158640
rect 141625 158600 141635 158680
rect 141945 158600 141955 158680
rect 145465 158600 145475 158680
rect 145785 158600 145795 158680
rect 146105 158600 146115 158680
rect 146700 158620 146780 158630
rect 146780 158540 146790 158620
rect 141705 158520 141785 158530
rect 142025 158520 142105 158530
rect 145225 158520 145305 158530
rect 145545 158520 145625 158530
rect 145865 158520 145945 158530
rect 141060 158460 141140 158470
rect 141210 158460 141290 158470
rect 141360 158460 141440 158470
rect 141140 158380 141150 158460
rect 141290 158380 141300 158460
rect 141440 158380 141450 158460
rect 141785 158440 141795 158520
rect 142105 158440 142115 158520
rect 145305 158440 145315 158520
rect 145625 158440 145635 158520
rect 145945 158440 145955 158520
rect 146540 158460 146620 158470
rect 146860 158460 146940 158470
rect 146620 158380 146630 158460
rect 146940 158380 146950 158460
rect 141545 158360 141625 158370
rect 141865 158360 141945 158370
rect 142185 158360 142200 158370
rect 145385 158360 145465 158370
rect 145705 158360 145785 158370
rect 146025 158360 146105 158370
rect 141060 158280 141140 158290
rect 141210 158280 141290 158290
rect 141360 158280 141440 158290
rect 141625 158280 141635 158360
rect 141945 158280 141955 158360
rect 145465 158280 145475 158360
rect 145785 158280 145795 158360
rect 146105 158280 146115 158360
rect 146700 158300 146780 158310
rect 141140 158200 141150 158280
rect 141290 158200 141300 158280
rect 141440 158200 141450 158280
rect 146780 158220 146790 158300
rect 141705 158200 141785 158210
rect 142025 158200 142105 158210
rect 145225 158200 145305 158210
rect 145545 158200 145625 158210
rect 145865 158200 145945 158210
rect 141785 158120 141795 158200
rect 142105 158120 142115 158200
rect 145305 158120 145315 158200
rect 145625 158120 145635 158200
rect 145945 158120 145955 158200
rect 146540 158140 146620 158150
rect 146860 158140 146940 158150
rect 141060 158100 141140 158110
rect 141210 158100 141290 158110
rect 141360 158100 141440 158110
rect 141140 158020 141150 158100
rect 141290 158020 141300 158100
rect 141440 158020 141450 158100
rect 146620 158060 146630 158140
rect 146940 158060 146950 158140
rect 141545 158040 141625 158050
rect 141865 158040 141945 158050
rect 142185 158040 142200 158050
rect 145385 158040 145465 158050
rect 145705 158040 145785 158050
rect 146025 158040 146105 158050
rect 141625 157960 141635 158040
rect 141945 157960 141955 158040
rect 145465 157960 145475 158040
rect 145785 157960 145795 158040
rect 146105 157960 146115 158040
rect 146700 157980 146780 157990
rect 141060 157920 141140 157930
rect 141210 157920 141290 157930
rect 141360 157920 141440 157930
rect 141140 157840 141150 157920
rect 141290 157840 141300 157920
rect 141440 157840 141450 157920
rect 146780 157900 146790 157980
rect 141705 157880 141785 157890
rect 142025 157880 142105 157890
rect 145225 157880 145305 157890
rect 145545 157880 145625 157890
rect 145865 157880 145945 157890
rect 141785 157800 141795 157880
rect 142105 157800 142115 157880
rect 145305 157800 145315 157880
rect 145625 157800 145635 157880
rect 145945 157800 145955 157880
rect 146540 157820 146620 157830
rect 146860 157820 146940 157830
rect 141060 157740 141140 157750
rect 141210 157740 141290 157750
rect 141360 157740 141440 157750
rect 146620 157740 146630 157820
rect 146940 157740 146950 157820
rect 141140 157660 141150 157740
rect 141290 157660 141300 157740
rect 141440 157660 141450 157740
rect 141545 157720 141625 157730
rect 141865 157720 141945 157730
rect 142185 157720 142200 157730
rect 145385 157720 145465 157730
rect 145705 157720 145785 157730
rect 146025 157720 146105 157730
rect 141625 157640 141635 157720
rect 141945 157640 141955 157720
rect 145465 157640 145475 157720
rect 145785 157640 145795 157720
rect 146105 157640 146115 157720
rect 146700 157660 146780 157670
rect 146780 157580 146790 157660
rect 141060 157560 141140 157570
rect 141210 157560 141290 157570
rect 141360 157560 141440 157570
rect 141705 157560 141785 157570
rect 142025 157560 142105 157570
rect 145225 157560 145305 157570
rect 145545 157560 145625 157570
rect 145865 157560 145945 157570
rect 141140 157480 141150 157560
rect 141290 157480 141300 157560
rect 141440 157480 141450 157560
rect 141785 157480 141795 157560
rect 142105 157480 142115 157560
rect 145305 157480 145315 157560
rect 145625 157480 145635 157560
rect 145945 157480 145955 157560
rect 146540 157500 146620 157510
rect 146860 157500 146940 157510
rect 146620 157420 146630 157500
rect 146940 157420 146950 157500
rect 141545 157400 141625 157410
rect 141865 157400 141945 157410
rect 142185 157400 142200 157410
rect 145385 157400 145465 157410
rect 145705 157400 145785 157410
rect 146025 157400 146105 157410
rect 141060 157380 141140 157390
rect 141210 157380 141290 157390
rect 141360 157380 141440 157390
rect 141140 157300 141150 157380
rect 141290 157300 141300 157380
rect 141440 157300 141450 157380
rect 141625 157320 141635 157400
rect 141945 157320 141955 157400
rect 145465 157320 145475 157400
rect 145785 157320 145795 157400
rect 146105 157320 146115 157400
rect 146700 157340 146780 157350
rect 146780 157260 146790 157340
rect 141705 157240 141785 157250
rect 142025 157240 142105 157250
rect 145225 157240 145305 157250
rect 145545 157240 145625 157250
rect 145865 157240 145945 157250
rect 141060 157200 141140 157210
rect 141210 157200 141290 157210
rect 141360 157200 141440 157210
rect 141140 157120 141150 157200
rect 141290 157120 141300 157200
rect 141440 157120 141450 157200
rect 141785 157160 141795 157240
rect 142105 157160 142115 157240
rect 145305 157160 145315 157240
rect 145625 157160 145635 157240
rect 145945 157160 145955 157240
rect 146540 157180 146620 157190
rect 146860 157180 146940 157190
rect 146620 157100 146630 157180
rect 146940 157100 146950 157180
rect 141545 157080 141625 157090
rect 141865 157080 141945 157090
rect 142185 157080 142200 157090
rect 145385 157080 145465 157090
rect 145705 157080 145785 157090
rect 146025 157080 146105 157090
rect 141060 157020 141140 157030
rect 141210 157020 141290 157030
rect 141360 157020 141440 157030
rect 141140 156940 141150 157020
rect 141290 156940 141300 157020
rect 141440 156940 141450 157020
rect 141625 157000 141635 157080
rect 141945 157000 141955 157080
rect 145465 157000 145475 157080
rect 145785 157000 145795 157080
rect 146105 157000 146115 157080
rect 146700 157020 146780 157030
rect 146780 156940 146790 157020
rect 141705 156920 141785 156930
rect 142025 156920 142105 156930
rect 145225 156920 145305 156930
rect 145545 156920 145625 156930
rect 145865 156920 145945 156930
rect 141060 156840 141140 156850
rect 141210 156840 141290 156850
rect 141360 156840 141440 156850
rect 141785 156840 141795 156920
rect 142105 156840 142115 156920
rect 145305 156840 145315 156920
rect 145625 156840 145635 156920
rect 145945 156840 145955 156920
rect 146540 156860 146620 156870
rect 146860 156860 146940 156870
rect 141140 156760 141150 156840
rect 141290 156760 141300 156840
rect 141440 156760 141450 156840
rect 146620 156780 146630 156860
rect 146940 156780 146950 156860
rect 141545 156760 141625 156770
rect 141865 156760 141945 156770
rect 142185 156760 142200 156770
rect 145385 156760 145465 156770
rect 145705 156760 145785 156770
rect 146025 156760 146105 156770
rect 141625 156680 141635 156760
rect 141945 156680 141955 156760
rect 145465 156680 145475 156760
rect 145785 156680 145795 156760
rect 146105 156680 146115 156760
rect 146700 156700 146780 156710
rect 141060 156660 141140 156670
rect 141210 156660 141290 156670
rect 141360 156660 141440 156670
rect 141140 156580 141150 156660
rect 141290 156580 141300 156660
rect 141440 156580 141450 156660
rect 146780 156620 146790 156700
rect 141705 156600 141785 156610
rect 142025 156600 142105 156610
rect 145225 156600 145305 156610
rect 145545 156600 145625 156610
rect 145865 156600 145945 156610
rect 141785 156520 141795 156600
rect 142105 156520 142115 156600
rect 145305 156520 145315 156600
rect 145625 156520 145635 156600
rect 145945 156520 145955 156600
rect 146540 156540 146620 156550
rect 146860 156540 146940 156550
rect 141060 156480 141140 156490
rect 141210 156480 141290 156490
rect 141360 156480 141440 156490
rect 141140 156400 141150 156480
rect 141290 156400 141300 156480
rect 141440 156400 141450 156480
rect 146620 156460 146630 156540
rect 146940 156460 146950 156540
rect 141545 156440 141625 156450
rect 141865 156440 141945 156450
rect 142185 156440 142200 156450
rect 145385 156440 145465 156450
rect 145705 156440 145785 156450
rect 146025 156440 146105 156450
rect 141625 156360 141635 156440
rect 141945 156360 141955 156440
rect 145465 156360 145475 156440
rect 145785 156360 145795 156440
rect 146105 156360 146115 156440
rect 146700 156380 146780 156390
rect 141060 156300 141140 156310
rect 141210 156300 141290 156310
rect 141360 156300 141440 156310
rect 146780 156300 146790 156380
rect 141140 156220 141150 156300
rect 141290 156220 141300 156300
rect 141440 156220 141450 156300
rect 141705 156280 141785 156290
rect 142025 156280 142105 156290
rect 145225 156280 145305 156290
rect 145545 156280 145625 156290
rect 145865 156280 145945 156290
rect 141785 156200 141795 156280
rect 142105 156200 142115 156280
rect 145305 156200 145315 156280
rect 145625 156200 145635 156280
rect 145945 156200 145955 156280
rect 146540 156220 146620 156230
rect 146860 156220 146940 156230
rect 146620 156140 146630 156220
rect 146940 156140 146950 156220
rect 141060 156120 141140 156130
rect 141210 156120 141290 156130
rect 141360 156120 141440 156130
rect 141545 156120 141625 156130
rect 141865 156120 141945 156130
rect 142185 156120 142200 156130
rect 145385 156120 145465 156130
rect 145705 156120 145785 156130
rect 146025 156120 146105 156130
rect 141140 156040 141150 156120
rect 141290 156040 141300 156120
rect 141440 156040 141450 156120
rect 141625 156040 141635 156120
rect 141945 156040 141955 156120
rect 145465 156040 145475 156120
rect 145785 156040 145795 156120
rect 146105 156040 146115 156120
rect 146700 156060 146780 156070
rect 146780 155980 146790 156060
rect 147100 155980 147110 156000
rect 147420 155980 147430 156000
rect 147740 155980 147750 156000
rect 148060 155980 148070 156000
rect 148380 155980 148390 156000
rect 148700 155980 148710 156000
rect 149020 155980 149030 156000
rect 149340 155980 149350 156000
rect 149660 155980 149670 156000
rect 149980 155980 149990 156000
rect 150300 155980 150310 156000
rect 150620 155980 150630 156000
rect 150940 155980 150950 156000
rect 151260 155980 151270 156000
rect 151580 155980 151590 156000
rect 151900 155980 151910 156000
rect 152220 155980 152230 156000
rect 152540 155980 152550 156000
rect 152860 155980 152870 156000
rect 153180 155980 153190 156000
rect 153500 155980 153510 156000
rect 153820 155980 153830 156000
rect 154140 155980 154150 156000
rect 154460 155980 154470 156000
rect 154780 155980 154790 156000
rect 155100 155980 155110 156000
rect 155420 155980 155430 156000
rect 155740 155980 155750 156000
rect 141705 155960 141785 155970
rect 142025 155960 142105 155970
rect 145225 155960 145305 155970
rect 145545 155960 145625 155970
rect 145865 155960 145945 155970
rect 141060 155940 141140 155950
rect 141210 155940 141290 155950
rect 141360 155940 141440 155950
rect 141140 155860 141150 155940
rect 141290 155860 141300 155940
rect 141440 155860 141450 155940
rect 141785 155880 141795 155960
rect 142105 155880 142115 155960
rect 145305 155880 145315 155960
rect 145625 155880 145635 155960
rect 145945 155880 145955 155960
rect 146540 155900 146620 155910
rect 146860 155900 146940 155910
rect 147180 155900 147260 155910
rect 147500 155900 147580 155910
rect 147820 155900 147900 155910
rect 148140 155900 148220 155910
rect 148460 155900 148540 155910
rect 148780 155900 148860 155910
rect 149100 155900 149180 155910
rect 149420 155900 149500 155910
rect 149740 155900 149820 155910
rect 150060 155900 150140 155910
rect 150380 155900 150460 155910
rect 150700 155900 150780 155910
rect 151020 155900 151100 155910
rect 151340 155900 151420 155910
rect 151660 155900 151740 155910
rect 151980 155900 152060 155910
rect 152300 155900 152380 155910
rect 152620 155900 152700 155910
rect 152940 155900 153020 155910
rect 153260 155900 153340 155910
rect 153580 155900 153660 155910
rect 153900 155900 153980 155910
rect 154220 155900 154300 155910
rect 154540 155900 154620 155910
rect 154860 155900 154940 155910
rect 155180 155900 155260 155910
rect 155500 155900 155580 155910
rect 155820 155900 155900 155910
rect 146620 155820 146630 155900
rect 146940 155820 146950 155900
rect 147260 155820 147270 155900
rect 147580 155820 147590 155900
rect 147900 155820 147910 155900
rect 148220 155820 148230 155900
rect 148540 155820 148550 155900
rect 148860 155820 148870 155900
rect 149180 155820 149190 155900
rect 149500 155820 149510 155900
rect 149820 155820 149830 155900
rect 150140 155820 150150 155900
rect 150460 155820 150470 155900
rect 150780 155820 150790 155900
rect 151100 155820 151110 155900
rect 151420 155820 151430 155900
rect 151740 155820 151750 155900
rect 152060 155820 152070 155900
rect 152380 155820 152390 155900
rect 152700 155820 152710 155900
rect 153020 155820 153030 155900
rect 153340 155820 153350 155900
rect 153660 155820 153670 155900
rect 153980 155820 153990 155900
rect 154300 155820 154310 155900
rect 154620 155820 154630 155900
rect 154940 155820 154950 155900
rect 155260 155820 155270 155900
rect 155580 155820 155590 155900
rect 155900 155820 155910 155900
rect 141545 155800 141625 155810
rect 141865 155800 141945 155810
rect 142185 155800 142200 155810
rect 145385 155800 145465 155810
rect 145705 155800 145785 155810
rect 146025 155800 146105 155810
rect 141060 155760 141140 155770
rect 141210 155760 141290 155770
rect 141360 155760 141440 155770
rect 141140 155680 141150 155760
rect 141290 155680 141300 155760
rect 141440 155680 141450 155760
rect 141625 155720 141635 155800
rect 141945 155720 141955 155800
rect 145465 155720 145475 155800
rect 145785 155720 145795 155800
rect 146105 155720 146115 155800
rect 146700 155740 146780 155750
rect 147020 155740 147100 155750
rect 147340 155740 147420 155750
rect 147660 155740 147740 155750
rect 147980 155740 148060 155750
rect 148300 155740 148380 155750
rect 148620 155740 148700 155750
rect 148940 155740 149020 155750
rect 149260 155740 149340 155750
rect 149580 155740 149660 155750
rect 149900 155740 149980 155750
rect 150220 155740 150300 155750
rect 150540 155740 150620 155750
rect 150860 155740 150940 155750
rect 151180 155740 151260 155750
rect 151500 155740 151580 155750
rect 151820 155740 151900 155750
rect 152140 155740 152220 155750
rect 152460 155740 152540 155750
rect 152780 155740 152860 155750
rect 153100 155740 153180 155750
rect 153420 155740 153500 155750
rect 153740 155740 153820 155750
rect 154060 155740 154140 155750
rect 154380 155740 154460 155750
rect 154700 155740 154780 155750
rect 155020 155740 155100 155750
rect 155340 155740 155420 155750
rect 155660 155740 155740 155750
rect 155980 155740 156000 155750
rect 146780 155660 146790 155740
rect 147100 155660 147110 155740
rect 147420 155660 147430 155740
rect 147740 155660 147750 155740
rect 148060 155660 148070 155740
rect 148380 155660 148390 155740
rect 148700 155660 148710 155740
rect 149020 155660 149030 155740
rect 149340 155660 149350 155740
rect 149660 155660 149670 155740
rect 149980 155660 149990 155740
rect 150300 155660 150310 155740
rect 150620 155660 150630 155740
rect 150940 155660 150950 155740
rect 151260 155660 151270 155740
rect 151580 155660 151590 155740
rect 151900 155660 151910 155740
rect 152220 155660 152230 155740
rect 152540 155660 152550 155740
rect 152860 155660 152870 155740
rect 153180 155660 153190 155740
rect 153500 155660 153510 155740
rect 153820 155660 153830 155740
rect 154140 155660 154150 155740
rect 154460 155660 154470 155740
rect 154780 155660 154790 155740
rect 155100 155660 155110 155740
rect 155420 155660 155430 155740
rect 155740 155660 155750 155740
rect 141705 155640 141785 155650
rect 142025 155640 142105 155650
rect 145225 155640 145305 155650
rect 145545 155640 145625 155650
rect 145865 155640 145945 155650
rect 141060 155580 141140 155590
rect 141210 155580 141290 155590
rect 141360 155580 141440 155590
rect 141140 155500 141150 155580
rect 141290 155500 141300 155580
rect 141440 155500 141450 155580
rect 141785 155560 141795 155640
rect 142105 155560 142115 155640
rect 145305 155560 145315 155640
rect 145625 155560 145635 155640
rect 145945 155560 145955 155640
rect 146540 155580 146620 155590
rect 146860 155580 146940 155590
rect 147180 155580 147260 155590
rect 147500 155580 147580 155590
rect 147820 155580 147900 155590
rect 148140 155580 148220 155590
rect 148460 155580 148540 155590
rect 148780 155580 148860 155590
rect 149100 155580 149180 155590
rect 149420 155580 149500 155590
rect 149740 155580 149820 155590
rect 150060 155580 150140 155590
rect 150380 155580 150460 155590
rect 150700 155580 150780 155590
rect 151020 155580 151100 155590
rect 151340 155580 151420 155590
rect 151660 155580 151740 155590
rect 151980 155580 152060 155590
rect 152300 155580 152380 155590
rect 152620 155580 152700 155590
rect 152940 155580 153020 155590
rect 153260 155580 153340 155590
rect 153580 155580 153660 155590
rect 153900 155580 153980 155590
rect 154220 155580 154300 155590
rect 154540 155580 154620 155590
rect 154860 155580 154940 155590
rect 155180 155580 155260 155590
rect 155500 155580 155580 155590
rect 155820 155580 155900 155590
rect 146620 155500 146630 155580
rect 146940 155500 146950 155580
rect 147260 155500 147270 155580
rect 147580 155500 147590 155580
rect 147900 155500 147910 155580
rect 148220 155500 148230 155580
rect 148540 155500 148550 155580
rect 148860 155500 148870 155580
rect 149180 155500 149190 155580
rect 149500 155500 149510 155580
rect 149820 155500 149830 155580
rect 150140 155500 150150 155580
rect 150460 155500 150470 155580
rect 150780 155500 150790 155580
rect 151100 155500 151110 155580
rect 151420 155500 151430 155580
rect 151740 155500 151750 155580
rect 152060 155500 152070 155580
rect 152380 155500 152390 155580
rect 152700 155500 152710 155580
rect 153020 155500 153030 155580
rect 153340 155500 153350 155580
rect 153660 155500 153670 155580
rect 153980 155500 153990 155580
rect 154300 155500 154310 155580
rect 154620 155500 154630 155580
rect 154940 155500 154950 155580
rect 155260 155500 155270 155580
rect 155580 155500 155590 155580
rect 155900 155500 155910 155580
rect 141545 155480 141625 155490
rect 141865 155480 141945 155490
rect 142185 155480 142200 155490
rect 145385 155480 145465 155490
rect 145705 155480 145785 155490
rect 146025 155480 146105 155490
rect 141060 155400 141140 155410
rect 141210 155400 141290 155410
rect 141360 155400 141440 155410
rect 141625 155400 141635 155480
rect 141945 155400 141955 155480
rect 145465 155400 145475 155480
rect 145785 155400 145795 155480
rect 146105 155400 146115 155480
rect 146700 155420 146780 155430
rect 147020 155420 147100 155430
rect 147340 155420 147420 155430
rect 147660 155420 147740 155430
rect 147980 155420 148060 155430
rect 148300 155420 148380 155430
rect 148620 155420 148700 155430
rect 148940 155420 149020 155430
rect 149260 155420 149340 155430
rect 149580 155420 149660 155430
rect 149900 155420 149980 155430
rect 150220 155420 150300 155430
rect 150540 155420 150620 155430
rect 150860 155420 150940 155430
rect 151180 155420 151260 155430
rect 151500 155420 151580 155430
rect 151820 155420 151900 155430
rect 152140 155420 152220 155430
rect 152460 155420 152540 155430
rect 152780 155420 152860 155430
rect 153100 155420 153180 155430
rect 153420 155420 153500 155430
rect 153740 155420 153820 155430
rect 154060 155420 154140 155430
rect 154380 155420 154460 155430
rect 154700 155420 154780 155430
rect 155020 155420 155100 155430
rect 155340 155420 155420 155430
rect 155660 155420 155740 155430
rect 155980 155420 156000 155430
rect 141140 155320 141150 155400
rect 141290 155320 141300 155400
rect 141440 155320 141450 155400
rect 146780 155340 146790 155420
rect 147100 155340 147110 155420
rect 147420 155340 147430 155420
rect 147740 155340 147750 155420
rect 148060 155340 148070 155420
rect 148380 155340 148390 155420
rect 148700 155340 148710 155420
rect 149020 155340 149030 155420
rect 149340 155340 149350 155420
rect 149660 155340 149670 155420
rect 149980 155340 149990 155420
rect 150300 155340 150310 155420
rect 150620 155340 150630 155420
rect 150940 155340 150950 155420
rect 151260 155340 151270 155420
rect 151580 155340 151590 155420
rect 151900 155340 151910 155420
rect 152220 155340 152230 155420
rect 152540 155340 152550 155420
rect 152860 155340 152870 155420
rect 153180 155340 153190 155420
rect 153500 155340 153510 155420
rect 153820 155340 153830 155420
rect 154140 155340 154150 155420
rect 154460 155340 154470 155420
rect 154780 155340 154790 155420
rect 155100 155340 155110 155420
rect 155420 155340 155430 155420
rect 155740 155340 155750 155420
rect 141705 155320 141785 155330
rect 142025 155320 142105 155330
rect 145225 155320 145305 155330
rect 145545 155320 145625 155330
rect 145865 155320 145945 155330
rect 141785 155240 141795 155320
rect 142105 155240 142115 155320
rect 145305 155240 145315 155320
rect 145625 155240 145635 155320
rect 145945 155240 145955 155320
rect 146540 155260 146620 155270
rect 146860 155260 146940 155270
rect 147180 155260 147260 155270
rect 147500 155260 147580 155270
rect 147820 155260 147900 155270
rect 148140 155260 148220 155270
rect 148460 155260 148540 155270
rect 148780 155260 148860 155270
rect 149100 155260 149180 155270
rect 149420 155260 149500 155270
rect 149740 155260 149820 155270
rect 150060 155260 150140 155270
rect 150380 155260 150460 155270
rect 150700 155260 150780 155270
rect 151020 155260 151100 155270
rect 151340 155260 151420 155270
rect 151660 155260 151740 155270
rect 151980 155260 152060 155270
rect 152300 155260 152380 155270
rect 152620 155260 152700 155270
rect 152940 155260 153020 155270
rect 153260 155260 153340 155270
rect 153580 155260 153660 155270
rect 153900 155260 153980 155270
rect 154220 155260 154300 155270
rect 154540 155260 154620 155270
rect 154860 155260 154940 155270
rect 155180 155260 155260 155270
rect 155500 155260 155580 155270
rect 155820 155260 155900 155270
rect 141060 155220 141140 155230
rect 141210 155220 141290 155230
rect 141360 155220 141440 155230
rect 141140 155140 141150 155220
rect 141290 155140 141300 155220
rect 141440 155140 141450 155220
rect 146620 155180 146630 155260
rect 146940 155180 146950 155260
rect 147260 155180 147270 155260
rect 147580 155180 147590 155260
rect 147900 155180 147910 155260
rect 148220 155180 148230 155260
rect 148540 155180 148550 155260
rect 148860 155180 148870 155260
rect 149180 155180 149190 155260
rect 149500 155180 149510 155260
rect 149820 155180 149830 155260
rect 150140 155180 150150 155260
rect 150460 155180 150470 155260
rect 150780 155180 150790 155260
rect 151100 155180 151110 155260
rect 151420 155180 151430 155260
rect 151740 155180 151750 155260
rect 152060 155180 152070 155260
rect 152380 155180 152390 155260
rect 152700 155180 152710 155260
rect 153020 155180 153030 155260
rect 153340 155180 153350 155260
rect 153660 155180 153670 155260
rect 153980 155180 153990 155260
rect 154300 155180 154310 155260
rect 154620 155180 154630 155260
rect 154940 155180 154950 155260
rect 155260 155180 155270 155260
rect 155580 155180 155590 155260
rect 155900 155180 155910 155260
rect 141545 155160 141625 155170
rect 141865 155160 141945 155170
rect 142185 155160 142200 155170
rect 145385 155160 145465 155170
rect 145705 155160 145785 155170
rect 146025 155160 146105 155170
rect 141625 155080 141635 155160
rect 141945 155080 141955 155160
rect 145465 155080 145475 155160
rect 145785 155080 145795 155160
rect 146105 155080 146115 155160
rect 146700 155100 146780 155110
rect 147020 155100 147100 155110
rect 147340 155100 147420 155110
rect 147660 155100 147740 155110
rect 147980 155100 148060 155110
rect 148300 155100 148380 155110
rect 148620 155100 148700 155110
rect 148940 155100 149020 155110
rect 149260 155100 149340 155110
rect 149580 155100 149660 155110
rect 149900 155100 149980 155110
rect 150220 155100 150300 155110
rect 150540 155100 150620 155110
rect 150860 155100 150940 155110
rect 151180 155100 151260 155110
rect 151500 155100 151580 155110
rect 151820 155100 151900 155110
rect 152140 155100 152220 155110
rect 152460 155100 152540 155110
rect 152780 155100 152860 155110
rect 153100 155100 153180 155110
rect 153420 155100 153500 155110
rect 153740 155100 153820 155110
rect 154060 155100 154140 155110
rect 154380 155100 154460 155110
rect 154700 155100 154780 155110
rect 155020 155100 155100 155110
rect 155340 155100 155420 155110
rect 155660 155100 155740 155110
rect 155980 155100 156000 155110
rect 141060 155040 141140 155050
rect 141210 155040 141290 155050
rect 141360 155040 141440 155050
rect 141140 154960 141150 155040
rect 141290 154960 141300 155040
rect 141440 154960 141450 155040
rect 146780 155020 146790 155100
rect 147100 155020 147110 155100
rect 147420 155020 147430 155100
rect 147740 155020 147750 155100
rect 148060 155020 148070 155100
rect 148380 155020 148390 155100
rect 148700 155020 148710 155100
rect 149020 155020 149030 155100
rect 149340 155020 149350 155100
rect 149660 155020 149670 155100
rect 149980 155020 149990 155100
rect 150300 155020 150310 155100
rect 150620 155020 150630 155100
rect 150940 155020 150950 155100
rect 151260 155020 151270 155100
rect 151580 155020 151590 155100
rect 151900 155020 151910 155100
rect 152220 155020 152230 155100
rect 152540 155020 152550 155100
rect 152860 155020 152870 155100
rect 153180 155020 153190 155100
rect 153500 155020 153510 155100
rect 153820 155020 153830 155100
rect 154140 155020 154150 155100
rect 154460 155020 154470 155100
rect 154780 155020 154790 155100
rect 155100 155020 155110 155100
rect 155420 155020 155430 155100
rect 155740 155020 155750 155100
rect 141705 155000 141785 155010
rect 142025 155000 142105 155010
rect 145225 155000 145305 155010
rect 145545 155000 145625 155010
rect 145865 155000 145945 155010
rect 141785 154920 141795 155000
rect 142105 154920 142115 155000
rect 145305 154920 145315 155000
rect 145625 154920 145635 155000
rect 145945 154920 145955 155000
rect 146540 154940 146620 154950
rect 146860 154940 146940 154950
rect 147180 154940 147260 154950
rect 147500 154940 147580 154950
rect 147820 154940 147900 154950
rect 148140 154940 148220 154950
rect 148460 154940 148540 154950
rect 148780 154940 148860 154950
rect 149100 154940 149180 154950
rect 149420 154940 149500 154950
rect 149740 154940 149820 154950
rect 150060 154940 150140 154950
rect 150380 154940 150460 154950
rect 150700 154940 150780 154950
rect 151020 154940 151100 154950
rect 151340 154940 151420 154950
rect 151660 154940 151740 154950
rect 151980 154940 152060 154950
rect 152300 154940 152380 154950
rect 152620 154940 152700 154950
rect 152940 154940 153020 154950
rect 153260 154940 153340 154950
rect 153580 154940 153660 154950
rect 153900 154940 153980 154950
rect 154220 154940 154300 154950
rect 154540 154940 154620 154950
rect 154860 154940 154940 154950
rect 155180 154940 155260 154950
rect 155500 154940 155580 154950
rect 155820 154940 155900 154950
rect 141060 154860 141140 154870
rect 141210 154860 141290 154870
rect 141360 154860 141440 154870
rect 146620 154860 146630 154940
rect 146940 154860 146950 154940
rect 147260 154860 147270 154940
rect 147580 154860 147590 154940
rect 147900 154860 147910 154940
rect 148220 154860 148230 154940
rect 148540 154860 148550 154940
rect 148860 154860 148870 154940
rect 149180 154860 149190 154940
rect 149500 154860 149510 154940
rect 149820 154860 149830 154940
rect 150140 154860 150150 154940
rect 150460 154860 150470 154940
rect 150780 154860 150790 154940
rect 151100 154860 151110 154940
rect 151420 154860 151430 154940
rect 151740 154860 151750 154940
rect 152060 154860 152070 154940
rect 152380 154860 152390 154940
rect 152700 154860 152710 154940
rect 153020 154860 153030 154940
rect 153340 154860 153350 154940
rect 153660 154860 153670 154940
rect 153980 154860 153990 154940
rect 154300 154860 154310 154940
rect 154620 154860 154630 154940
rect 154940 154860 154950 154940
rect 155260 154860 155270 154940
rect 155580 154860 155590 154940
rect 155900 154860 155910 154940
rect 141140 154780 141150 154860
rect 141290 154780 141300 154860
rect 141440 154780 141450 154860
rect 141545 154840 141625 154850
rect 141865 154840 141945 154850
rect 142185 154840 142200 154850
rect 145385 154840 145465 154850
rect 145705 154840 145785 154850
rect 146025 154840 146105 154850
rect 141625 154760 141635 154840
rect 141945 154760 141955 154840
rect 145465 154760 145475 154840
rect 145785 154760 145795 154840
rect 146105 154760 146115 154840
rect 146700 154780 146780 154790
rect 147020 154780 147100 154790
rect 147340 154780 147420 154790
rect 147660 154780 147740 154790
rect 147980 154780 148060 154790
rect 148300 154780 148380 154790
rect 148620 154780 148700 154790
rect 148940 154780 149020 154790
rect 149260 154780 149340 154790
rect 149580 154780 149660 154790
rect 149900 154780 149980 154790
rect 150220 154780 150300 154790
rect 150540 154780 150620 154790
rect 150860 154780 150940 154790
rect 151180 154780 151260 154790
rect 151500 154780 151580 154790
rect 151820 154780 151900 154790
rect 152140 154780 152220 154790
rect 152460 154780 152540 154790
rect 152780 154780 152860 154790
rect 153100 154780 153180 154790
rect 153420 154780 153500 154790
rect 153740 154780 153820 154790
rect 154060 154780 154140 154790
rect 154380 154780 154460 154790
rect 154700 154780 154780 154790
rect 155020 154780 155100 154790
rect 155340 154780 155420 154790
rect 155660 154780 155740 154790
rect 155980 154780 156000 154790
rect 146780 154700 146790 154780
rect 147100 154700 147110 154780
rect 147420 154700 147430 154780
rect 147740 154700 147750 154780
rect 148060 154700 148070 154780
rect 148380 154700 148390 154780
rect 148700 154700 148710 154780
rect 149020 154700 149030 154780
rect 149340 154700 149350 154780
rect 149660 154700 149670 154780
rect 149980 154700 149990 154780
rect 150300 154700 150310 154780
rect 150620 154700 150630 154780
rect 150940 154700 150950 154780
rect 151260 154700 151270 154780
rect 151580 154700 151590 154780
rect 151900 154700 151910 154780
rect 152220 154700 152230 154780
rect 152540 154700 152550 154780
rect 152860 154700 152870 154780
rect 153180 154700 153190 154780
rect 153500 154700 153510 154780
rect 153820 154700 153830 154780
rect 154140 154700 154150 154780
rect 154460 154700 154470 154780
rect 154780 154700 154790 154780
rect 155100 154700 155110 154780
rect 155420 154700 155430 154780
rect 155740 154700 155750 154780
rect 141060 154680 141140 154690
rect 141210 154680 141290 154690
rect 141360 154680 141440 154690
rect 141705 154680 141785 154690
rect 142025 154680 142105 154690
rect 145225 154680 145305 154690
rect 145545 154680 145625 154690
rect 145865 154680 145945 154690
rect 141140 154600 141150 154680
rect 141290 154600 141300 154680
rect 141440 154600 141450 154680
rect 141785 154600 141795 154680
rect 142105 154600 142115 154680
rect 145305 154600 145315 154680
rect 145625 154600 145635 154680
rect 145945 154600 145955 154680
rect 146540 154620 146620 154630
rect 146860 154620 146940 154630
rect 147180 154620 147260 154630
rect 147500 154620 147580 154630
rect 147820 154620 147900 154630
rect 148140 154620 148220 154630
rect 148460 154620 148540 154630
rect 148780 154620 148860 154630
rect 149100 154620 149180 154630
rect 149420 154620 149500 154630
rect 149740 154620 149820 154630
rect 150060 154620 150140 154630
rect 150380 154620 150460 154630
rect 150700 154620 150780 154630
rect 151020 154620 151100 154630
rect 151340 154620 151420 154630
rect 151660 154620 151740 154630
rect 151980 154620 152060 154630
rect 152300 154620 152380 154630
rect 152620 154620 152700 154630
rect 152940 154620 153020 154630
rect 153260 154620 153340 154630
rect 153580 154620 153660 154630
rect 153900 154620 153980 154630
rect 154220 154620 154300 154630
rect 154540 154620 154620 154630
rect 154860 154620 154940 154630
rect 155180 154620 155260 154630
rect 155500 154620 155580 154630
rect 155820 154620 155900 154630
rect 146620 154540 146630 154620
rect 146940 154540 146950 154620
rect 147260 154540 147270 154620
rect 147580 154540 147590 154620
rect 147900 154540 147910 154620
rect 148220 154540 148230 154620
rect 148540 154540 148550 154620
rect 148860 154540 148870 154620
rect 149180 154540 149190 154620
rect 149500 154540 149510 154620
rect 149820 154540 149830 154620
rect 150140 154540 150150 154620
rect 150460 154540 150470 154620
rect 150780 154540 150790 154620
rect 151100 154540 151110 154620
rect 151420 154540 151430 154620
rect 151740 154540 151750 154620
rect 152060 154540 152070 154620
rect 152380 154540 152390 154620
rect 152700 154540 152710 154620
rect 153020 154540 153030 154620
rect 153340 154540 153350 154620
rect 153660 154540 153670 154620
rect 153980 154540 153990 154620
rect 154300 154540 154310 154620
rect 154620 154540 154630 154620
rect 154940 154540 154950 154620
rect 155260 154540 155270 154620
rect 155580 154540 155590 154620
rect 155900 154540 155910 154620
rect 141545 154520 141625 154530
rect 141865 154520 141945 154530
rect 142185 154520 142200 154530
rect 145385 154520 145465 154530
rect 145705 154520 145785 154530
rect 146025 154520 146105 154530
rect 141060 154500 141140 154510
rect 141210 154500 141290 154510
rect 141360 154500 141440 154510
rect 141140 154420 141150 154500
rect 141290 154420 141300 154500
rect 141440 154420 141450 154500
rect 141625 154440 141635 154520
rect 141945 154440 141955 154520
rect 145465 154440 145475 154520
rect 145785 154440 145795 154520
rect 146105 154440 146115 154520
rect 146700 154460 146780 154470
rect 147020 154460 147100 154470
rect 147340 154460 147420 154470
rect 147660 154460 147740 154470
rect 147980 154460 148060 154470
rect 148300 154460 148380 154470
rect 148620 154460 148700 154470
rect 148940 154460 149020 154470
rect 149260 154460 149340 154470
rect 149580 154460 149660 154470
rect 149900 154460 149980 154470
rect 150220 154460 150300 154470
rect 150540 154460 150620 154470
rect 150860 154460 150940 154470
rect 151180 154460 151260 154470
rect 151500 154460 151580 154470
rect 151820 154460 151900 154470
rect 152140 154460 152220 154470
rect 152460 154460 152540 154470
rect 152780 154460 152860 154470
rect 153100 154460 153180 154470
rect 153420 154460 153500 154470
rect 153740 154460 153820 154470
rect 154060 154460 154140 154470
rect 154380 154460 154460 154470
rect 154700 154460 154780 154470
rect 155020 154460 155100 154470
rect 155340 154460 155420 154470
rect 155660 154460 155740 154470
rect 155980 154460 156000 154470
rect 146780 154380 146790 154460
rect 147100 154380 147110 154460
rect 147420 154380 147430 154460
rect 147740 154380 147750 154460
rect 148060 154380 148070 154460
rect 148380 154380 148390 154460
rect 148700 154380 148710 154460
rect 149020 154380 149030 154460
rect 149340 154380 149350 154460
rect 149660 154380 149670 154460
rect 149980 154380 149990 154460
rect 150300 154380 150310 154460
rect 150620 154380 150630 154460
rect 150940 154380 150950 154460
rect 151260 154380 151270 154460
rect 151580 154380 151590 154460
rect 151900 154380 151910 154460
rect 152220 154380 152230 154460
rect 152540 154380 152550 154460
rect 152860 154380 152870 154460
rect 153180 154380 153190 154460
rect 153500 154380 153510 154460
rect 153820 154380 153830 154460
rect 154140 154380 154150 154460
rect 154460 154380 154470 154460
rect 154780 154380 154790 154460
rect 155100 154380 155110 154460
rect 155420 154380 155430 154460
rect 155740 154380 155750 154460
rect 141705 154360 141785 154370
rect 142025 154360 142105 154370
rect 145225 154360 145305 154370
rect 145545 154360 145625 154370
rect 145865 154360 145945 154370
rect 141060 154320 141140 154330
rect 141210 154320 141290 154330
rect 141360 154320 141440 154330
rect 141140 154240 141150 154320
rect 141290 154240 141300 154320
rect 141440 154240 141450 154320
rect 141785 154280 141795 154360
rect 142105 154280 142115 154360
rect 145305 154280 145315 154360
rect 145625 154280 145635 154360
rect 145945 154280 145955 154360
rect 146540 154300 146620 154310
rect 146860 154300 146940 154310
rect 147180 154300 147260 154310
rect 147500 154300 147580 154310
rect 147820 154300 147900 154310
rect 148140 154300 148220 154310
rect 148460 154300 148540 154310
rect 148780 154300 148860 154310
rect 149100 154300 149180 154310
rect 149420 154300 149500 154310
rect 149740 154300 149820 154310
rect 150060 154300 150140 154310
rect 150380 154300 150460 154310
rect 150700 154300 150780 154310
rect 151020 154300 151100 154310
rect 151340 154300 151420 154310
rect 151660 154300 151740 154310
rect 151980 154300 152060 154310
rect 152300 154300 152380 154310
rect 152620 154300 152700 154310
rect 152940 154300 153020 154310
rect 153260 154300 153340 154310
rect 153580 154300 153660 154310
rect 153900 154300 153980 154310
rect 154220 154300 154300 154310
rect 154540 154300 154620 154310
rect 154860 154300 154940 154310
rect 155180 154300 155260 154310
rect 155500 154300 155580 154310
rect 155820 154300 155900 154310
rect 146620 154220 146630 154300
rect 146940 154220 146950 154300
rect 147260 154220 147270 154300
rect 147580 154220 147590 154300
rect 147900 154220 147910 154300
rect 148220 154220 148230 154300
rect 148540 154220 148550 154300
rect 148860 154220 148870 154300
rect 149180 154220 149190 154300
rect 149500 154220 149510 154300
rect 149820 154220 149830 154300
rect 150140 154220 150150 154300
rect 150460 154220 150470 154300
rect 150780 154220 150790 154300
rect 151100 154220 151110 154300
rect 151420 154220 151430 154300
rect 151740 154220 151750 154300
rect 152060 154220 152070 154300
rect 152380 154220 152390 154300
rect 152700 154220 152710 154300
rect 153020 154220 153030 154300
rect 153340 154220 153350 154300
rect 153660 154220 153670 154300
rect 153980 154220 153990 154300
rect 154300 154220 154310 154300
rect 154620 154220 154630 154300
rect 154940 154220 154950 154300
rect 155260 154220 155270 154300
rect 155580 154220 155590 154300
rect 155900 154220 155910 154300
rect 141545 154200 141625 154210
rect 141865 154200 141945 154210
rect 142185 154200 142200 154210
rect 145385 154200 145465 154210
rect 145705 154200 145785 154210
rect 146025 154200 146105 154210
rect 141060 154140 141140 154150
rect 141210 154140 141290 154150
rect 141360 154140 141440 154150
rect 141140 154060 141150 154140
rect 141290 154060 141300 154140
rect 141440 154060 141450 154140
rect 141625 154120 141635 154200
rect 141945 154120 141955 154200
rect 145465 154120 145475 154200
rect 145785 154120 145795 154200
rect 146105 154120 146115 154200
rect 146700 154140 146780 154150
rect 147020 154140 147100 154150
rect 147340 154140 147420 154150
rect 147660 154140 147740 154150
rect 147980 154140 148060 154150
rect 148300 154140 148380 154150
rect 148620 154140 148700 154150
rect 148940 154140 149020 154150
rect 149260 154140 149340 154150
rect 149580 154140 149660 154150
rect 149900 154140 149980 154150
rect 150220 154140 150300 154150
rect 150540 154140 150620 154150
rect 150860 154140 150940 154150
rect 151180 154140 151260 154150
rect 151500 154140 151580 154150
rect 151820 154140 151900 154150
rect 152140 154140 152220 154150
rect 152460 154140 152540 154150
rect 152780 154140 152860 154150
rect 153100 154140 153180 154150
rect 153420 154140 153500 154150
rect 153740 154140 153820 154150
rect 154060 154140 154140 154150
rect 154380 154140 154460 154150
rect 154700 154140 154780 154150
rect 155020 154140 155100 154150
rect 155340 154140 155420 154150
rect 155660 154140 155740 154150
rect 155980 154140 156000 154150
rect 146780 154060 146790 154140
rect 147100 154060 147110 154140
rect 147420 154060 147430 154140
rect 147740 154060 147750 154140
rect 148060 154060 148070 154140
rect 148380 154060 148390 154140
rect 148700 154060 148710 154140
rect 149020 154060 149030 154140
rect 149340 154060 149350 154140
rect 149660 154060 149670 154140
rect 149980 154060 149990 154140
rect 150300 154060 150310 154140
rect 150620 154060 150630 154140
rect 150940 154060 150950 154140
rect 151260 154060 151270 154140
rect 151580 154060 151590 154140
rect 151900 154060 151910 154140
rect 152220 154060 152230 154140
rect 152540 154060 152550 154140
rect 152860 154060 152870 154140
rect 153180 154060 153190 154140
rect 153500 154060 153510 154140
rect 153820 154060 153830 154140
rect 154140 154060 154150 154140
rect 154460 154060 154470 154140
rect 154780 154060 154790 154140
rect 155100 154060 155110 154140
rect 155420 154060 155430 154140
rect 155740 154060 155750 154140
rect 141705 154040 141785 154050
rect 142025 154040 142105 154050
rect 145225 154040 145305 154050
rect 145545 154040 145625 154050
rect 145865 154040 145945 154050
rect 141060 153960 141140 153970
rect 141210 153960 141290 153970
rect 141360 153960 141440 153970
rect 141785 153960 141795 154040
rect 142105 153960 142115 154040
rect 145305 153960 145315 154040
rect 145625 153960 145635 154040
rect 145945 153960 145955 154040
rect 146540 153980 146620 153990
rect 146860 153980 146940 153990
rect 147180 153980 147260 153990
rect 147500 153980 147580 153990
rect 147820 153980 147900 153990
rect 148140 153980 148220 153990
rect 148460 153980 148540 153990
rect 148780 153980 148860 153990
rect 149100 153980 149180 153990
rect 149420 153980 149500 153990
rect 149740 153980 149820 153990
rect 150060 153980 150140 153990
rect 150380 153980 150460 153990
rect 150700 153980 150780 153990
rect 151020 153980 151100 153990
rect 151340 153980 151420 153990
rect 151660 153980 151740 153990
rect 151980 153980 152060 153990
rect 152300 153980 152380 153990
rect 152620 153980 152700 153990
rect 152940 153980 153020 153990
rect 153260 153980 153340 153990
rect 153580 153980 153660 153990
rect 153900 153980 153980 153990
rect 154220 153980 154300 153990
rect 154540 153980 154620 153990
rect 154860 153980 154940 153990
rect 155180 153980 155260 153990
rect 155500 153980 155580 153990
rect 155820 153980 155900 153990
rect 141140 153880 141150 153960
rect 141290 153880 141300 153960
rect 141440 153880 141450 153960
rect 146620 153900 146630 153980
rect 146940 153900 146950 153980
rect 147260 153900 147270 153980
rect 147580 153900 147590 153980
rect 147900 153900 147910 153980
rect 148220 153900 148230 153980
rect 148540 153900 148550 153980
rect 148860 153900 148870 153980
rect 149180 153900 149190 153980
rect 149500 153900 149510 153980
rect 149820 153900 149830 153980
rect 150140 153900 150150 153980
rect 150460 153900 150470 153980
rect 150780 153900 150790 153980
rect 151100 153900 151110 153980
rect 151420 153900 151430 153980
rect 151740 153900 151750 153980
rect 152060 153900 152070 153980
rect 152380 153900 152390 153980
rect 152700 153900 152710 153980
rect 153020 153900 153030 153980
rect 153340 153900 153350 153980
rect 153660 153900 153670 153980
rect 153980 153900 153990 153980
rect 154300 153900 154310 153980
rect 154620 153900 154630 153980
rect 154940 153900 154950 153980
rect 155260 153900 155270 153980
rect 155580 153900 155590 153980
rect 155900 153900 155910 153980
rect 141545 153880 141625 153890
rect 141865 153880 141945 153890
rect 142185 153880 142200 153890
rect 145385 153880 145465 153890
rect 145705 153880 145785 153890
rect 146025 153880 146105 153890
rect 141625 153800 141635 153880
rect 141945 153800 141955 153880
rect 145465 153800 145475 153880
rect 145785 153800 145795 153880
rect 146105 153800 146115 153880
rect 146700 153820 146780 153830
rect 147020 153820 147100 153830
rect 147340 153820 147420 153830
rect 147660 153820 147740 153830
rect 147980 153820 148060 153830
rect 148300 153820 148380 153830
rect 148620 153820 148700 153830
rect 148940 153820 149020 153830
rect 149260 153820 149340 153830
rect 149580 153820 149660 153830
rect 149900 153820 149980 153830
rect 150220 153820 150300 153830
rect 150540 153820 150620 153830
rect 150860 153820 150940 153830
rect 151180 153820 151260 153830
rect 151500 153820 151580 153830
rect 151820 153820 151900 153830
rect 152140 153820 152220 153830
rect 152460 153820 152540 153830
rect 152780 153820 152860 153830
rect 153100 153820 153180 153830
rect 153420 153820 153500 153830
rect 153740 153820 153820 153830
rect 154060 153820 154140 153830
rect 154380 153820 154460 153830
rect 154700 153820 154780 153830
rect 155020 153820 155100 153830
rect 155340 153820 155420 153830
rect 155660 153820 155740 153830
rect 155980 153820 156000 153830
rect 141060 153780 141140 153790
rect 141210 153780 141290 153790
rect 141360 153780 141440 153790
rect 141140 153700 141150 153780
rect 141290 153700 141300 153780
rect 141440 153700 141450 153780
rect 146780 153740 146790 153820
rect 147100 153740 147110 153820
rect 147420 153740 147430 153820
rect 147740 153740 147750 153820
rect 148060 153740 148070 153820
rect 148380 153740 148390 153820
rect 148700 153740 148710 153820
rect 149020 153740 149030 153820
rect 149340 153740 149350 153820
rect 149660 153740 149670 153820
rect 149980 153740 149990 153820
rect 150300 153740 150310 153820
rect 150620 153740 150630 153820
rect 150940 153740 150950 153820
rect 151260 153740 151270 153820
rect 151580 153740 151590 153820
rect 151900 153740 151910 153820
rect 152220 153740 152230 153820
rect 152540 153740 152550 153820
rect 152860 153740 152870 153820
rect 153180 153740 153190 153820
rect 153500 153740 153510 153820
rect 153820 153740 153830 153820
rect 154140 153740 154150 153820
rect 154460 153740 154470 153820
rect 154780 153740 154790 153820
rect 155100 153740 155110 153820
rect 155420 153740 155430 153820
rect 155740 153740 155750 153820
rect 141705 153720 141785 153730
rect 142025 153720 142105 153730
rect 145225 153720 145305 153730
rect 145545 153720 145625 153730
rect 145865 153720 145945 153730
rect 141785 153640 141795 153720
rect 142105 153640 142115 153720
rect 145305 153640 145315 153720
rect 145625 153640 145635 153720
rect 145945 153640 145955 153720
rect 146540 153660 146620 153670
rect 146860 153660 146940 153670
rect 147180 153660 147260 153670
rect 147500 153660 147580 153670
rect 147820 153660 147900 153670
rect 148140 153660 148220 153670
rect 148460 153660 148540 153670
rect 148780 153660 148860 153670
rect 149100 153660 149180 153670
rect 149420 153660 149500 153670
rect 149740 153660 149820 153670
rect 150060 153660 150140 153670
rect 150380 153660 150460 153670
rect 150700 153660 150780 153670
rect 151020 153660 151100 153670
rect 151340 153660 151420 153670
rect 151660 153660 151740 153670
rect 151980 153660 152060 153670
rect 152300 153660 152380 153670
rect 152620 153660 152700 153670
rect 152940 153660 153020 153670
rect 153260 153660 153340 153670
rect 153580 153660 153660 153670
rect 153900 153660 153980 153670
rect 154220 153660 154300 153670
rect 154540 153660 154620 153670
rect 154860 153660 154940 153670
rect 155180 153660 155260 153670
rect 155500 153660 155580 153670
rect 155820 153660 155900 153670
rect 141060 153600 141140 153610
rect 141210 153600 141290 153610
rect 141360 153600 141440 153610
rect 141140 153520 141150 153600
rect 141290 153520 141300 153600
rect 141440 153520 141450 153600
rect 146620 153580 146630 153660
rect 146940 153580 146950 153660
rect 147260 153580 147270 153660
rect 147580 153580 147590 153660
rect 147900 153580 147910 153660
rect 148220 153580 148230 153660
rect 148540 153580 148550 153660
rect 148860 153580 148870 153660
rect 149180 153580 149190 153660
rect 149500 153580 149510 153660
rect 149820 153580 149830 153660
rect 150140 153580 150150 153660
rect 150460 153580 150470 153660
rect 150780 153580 150790 153660
rect 151100 153580 151110 153660
rect 151420 153580 151430 153660
rect 151740 153580 151750 153660
rect 152060 153580 152070 153660
rect 152380 153580 152390 153660
rect 152700 153580 152710 153660
rect 153020 153580 153030 153660
rect 153340 153580 153350 153660
rect 153660 153580 153670 153660
rect 153980 153580 153990 153660
rect 154300 153580 154310 153660
rect 154620 153580 154630 153660
rect 154940 153580 154950 153660
rect 155260 153580 155270 153660
rect 155580 153580 155590 153660
rect 155900 153580 155910 153660
rect 141545 153560 141625 153570
rect 141865 153560 141945 153570
rect 142185 153560 142200 153570
rect 145385 153560 145465 153570
rect 145705 153560 145785 153570
rect 146025 153560 146105 153570
rect 141625 153480 141635 153560
rect 141945 153480 141955 153560
rect 145465 153480 145475 153560
rect 145785 153480 145795 153560
rect 146105 153480 146115 153560
rect 146700 153500 146780 153510
rect 147020 153500 147100 153510
rect 147340 153500 147420 153510
rect 147660 153500 147740 153510
rect 147980 153500 148060 153510
rect 148300 153500 148380 153510
rect 148620 153500 148700 153510
rect 148940 153500 149020 153510
rect 149260 153500 149340 153510
rect 149580 153500 149660 153510
rect 149900 153500 149980 153510
rect 150220 153500 150300 153510
rect 150540 153500 150620 153510
rect 150860 153500 150940 153510
rect 151180 153500 151260 153510
rect 151500 153500 151580 153510
rect 151820 153500 151900 153510
rect 152140 153500 152220 153510
rect 152460 153500 152540 153510
rect 152780 153500 152860 153510
rect 153100 153500 153180 153510
rect 153420 153500 153500 153510
rect 153740 153500 153820 153510
rect 154060 153500 154140 153510
rect 154380 153500 154460 153510
rect 154700 153500 154780 153510
rect 155020 153500 155100 153510
rect 155340 153500 155420 153510
rect 155660 153500 155740 153510
rect 155980 153500 156000 153510
rect 141060 153420 141140 153430
rect 141210 153420 141290 153430
rect 141360 153420 141440 153430
rect 146780 153420 146790 153500
rect 147100 153420 147110 153500
rect 147420 153420 147430 153500
rect 147740 153420 147750 153500
rect 148060 153420 148070 153500
rect 148380 153420 148390 153500
rect 148700 153420 148710 153500
rect 149020 153420 149030 153500
rect 149340 153420 149350 153500
rect 149660 153420 149670 153500
rect 149980 153420 149990 153500
rect 150300 153420 150310 153500
rect 150620 153420 150630 153500
rect 150940 153420 150950 153500
rect 151260 153420 151270 153500
rect 151580 153420 151590 153500
rect 151900 153420 151910 153500
rect 152220 153420 152230 153500
rect 152540 153420 152550 153500
rect 152860 153420 152870 153500
rect 153180 153420 153190 153500
rect 153500 153420 153510 153500
rect 153820 153420 153830 153500
rect 154140 153420 154150 153500
rect 154460 153420 154470 153500
rect 154780 153420 154790 153500
rect 155100 153420 155110 153500
rect 155420 153420 155430 153500
rect 155740 153420 155750 153500
rect 141140 153340 141150 153420
rect 141290 153340 141300 153420
rect 141440 153340 141450 153420
rect 141705 153400 141785 153410
rect 142025 153400 142105 153410
rect 145225 153400 145305 153410
rect 145545 153400 145625 153410
rect 145865 153400 145945 153410
rect 141785 153320 141795 153400
rect 142105 153320 142115 153400
rect 145305 153320 145315 153400
rect 145625 153320 145635 153400
rect 145945 153320 145955 153400
rect 146540 153340 146620 153350
rect 146860 153340 146940 153350
rect 147180 153340 147260 153350
rect 147500 153340 147580 153350
rect 147820 153340 147900 153350
rect 148140 153340 148220 153350
rect 148460 153340 148540 153350
rect 148780 153340 148860 153350
rect 149100 153340 149180 153350
rect 149420 153340 149500 153350
rect 149740 153340 149820 153350
rect 150060 153340 150140 153350
rect 150380 153340 150460 153350
rect 150700 153340 150780 153350
rect 151020 153340 151100 153350
rect 151340 153340 151420 153350
rect 151660 153340 151740 153350
rect 151980 153340 152060 153350
rect 152300 153340 152380 153350
rect 152620 153340 152700 153350
rect 152940 153340 153020 153350
rect 153260 153340 153340 153350
rect 153580 153340 153660 153350
rect 153900 153340 153980 153350
rect 154220 153340 154300 153350
rect 154540 153340 154620 153350
rect 154860 153340 154940 153350
rect 155180 153340 155260 153350
rect 155500 153340 155580 153350
rect 155820 153340 155900 153350
rect 146620 153260 146630 153340
rect 146940 153260 146950 153340
rect 147260 153260 147270 153340
rect 147580 153260 147590 153340
rect 147900 153260 147910 153340
rect 148220 153260 148230 153340
rect 148540 153260 148550 153340
rect 148860 153260 148870 153340
rect 149180 153260 149190 153340
rect 149500 153260 149510 153340
rect 149820 153260 149830 153340
rect 150140 153260 150150 153340
rect 150460 153260 150470 153340
rect 150780 153260 150790 153340
rect 151100 153260 151110 153340
rect 151420 153260 151430 153340
rect 151740 153260 151750 153340
rect 152060 153260 152070 153340
rect 152380 153260 152390 153340
rect 152700 153260 152710 153340
rect 153020 153260 153030 153340
rect 153340 153260 153350 153340
rect 153660 153260 153670 153340
rect 153980 153260 153990 153340
rect 154300 153260 154310 153340
rect 154620 153260 154630 153340
rect 154940 153260 154950 153340
rect 155260 153260 155270 153340
rect 155580 153260 155590 153340
rect 155900 153260 155910 153340
rect 141060 153240 141140 153250
rect 141210 153240 141290 153250
rect 141360 153240 141440 153250
rect 141545 153240 141625 153250
rect 141865 153240 141945 153250
rect 142185 153240 142200 153250
rect 145385 153240 145465 153250
rect 145705 153240 145785 153250
rect 146025 153240 146105 153250
rect 141140 153160 141150 153240
rect 141290 153160 141300 153240
rect 141440 153160 141450 153240
rect 141625 153160 141635 153240
rect 141945 153160 141955 153240
rect 145465 153160 145475 153240
rect 145785 153160 145795 153240
rect 146105 153160 146115 153240
rect 146700 153180 146780 153190
rect 147020 153180 147100 153190
rect 147340 153180 147420 153190
rect 147660 153180 147740 153190
rect 147980 153180 148060 153190
rect 148300 153180 148380 153190
rect 148620 153180 148700 153190
rect 148940 153180 149020 153190
rect 149260 153180 149340 153190
rect 149580 153180 149660 153190
rect 149900 153180 149980 153190
rect 150220 153180 150300 153190
rect 150540 153180 150620 153190
rect 150860 153180 150940 153190
rect 151180 153180 151260 153190
rect 151500 153180 151580 153190
rect 151820 153180 151900 153190
rect 152140 153180 152220 153190
rect 152460 153180 152540 153190
rect 152780 153180 152860 153190
rect 153100 153180 153180 153190
rect 153420 153180 153500 153190
rect 153740 153180 153820 153190
rect 154060 153180 154140 153190
rect 154380 153180 154460 153190
rect 154700 153180 154780 153190
rect 155020 153180 155100 153190
rect 155340 153180 155420 153190
rect 155660 153180 155740 153190
rect 155980 153180 156000 153190
rect 146780 153100 146790 153180
rect 147100 153100 147110 153180
rect 147420 153100 147430 153180
rect 147740 153100 147750 153180
rect 148060 153100 148070 153180
rect 148380 153100 148390 153180
rect 148700 153100 148710 153180
rect 149020 153100 149030 153180
rect 149340 153100 149350 153180
rect 149660 153100 149670 153180
rect 149980 153100 149990 153180
rect 150300 153100 150310 153180
rect 150620 153100 150630 153180
rect 150940 153100 150950 153180
rect 151260 153100 151270 153180
rect 151580 153100 151590 153180
rect 151900 153100 151910 153180
rect 152220 153100 152230 153180
rect 152540 153100 152550 153180
rect 152860 153100 152870 153180
rect 153180 153100 153190 153180
rect 153500 153100 153510 153180
rect 153820 153100 153830 153180
rect 154140 153100 154150 153180
rect 154460 153100 154470 153180
rect 154780 153100 154790 153180
rect 155100 153100 155110 153180
rect 155420 153100 155430 153180
rect 155740 153100 155750 153180
rect 141705 153080 141785 153090
rect 142025 153080 142105 153090
rect 145225 153080 145305 153090
rect 145545 153080 145625 153090
rect 145865 153080 145945 153090
rect 141060 153060 141140 153070
rect 141210 153060 141290 153070
rect 141360 153060 141440 153070
rect 141140 152980 141150 153060
rect 141290 152980 141300 153060
rect 141440 152980 141450 153060
rect 141785 153000 141795 153080
rect 142105 153000 142115 153080
rect 145305 153000 145315 153080
rect 145625 153000 145635 153080
rect 145945 153000 145955 153080
rect 146540 153020 146620 153030
rect 146860 153020 146940 153030
rect 147180 153020 147260 153030
rect 147500 153020 147580 153030
rect 147820 153020 147900 153030
rect 148140 153020 148220 153030
rect 148460 153020 148540 153030
rect 148780 153020 148860 153030
rect 149100 153020 149180 153030
rect 149420 153020 149500 153030
rect 149740 153020 149820 153030
rect 150060 153020 150140 153030
rect 150380 153020 150460 153030
rect 150700 153020 150780 153030
rect 151020 153020 151100 153030
rect 151340 153020 151420 153030
rect 151660 153020 151740 153030
rect 151980 153020 152060 153030
rect 152300 153020 152380 153030
rect 152620 153020 152700 153030
rect 152940 153020 153020 153030
rect 153260 153020 153340 153030
rect 153580 153020 153660 153030
rect 153900 153020 153980 153030
rect 154220 153020 154300 153030
rect 154540 153020 154620 153030
rect 154860 153020 154940 153030
rect 155180 153020 155260 153030
rect 155500 153020 155580 153030
rect 155820 153020 155900 153030
rect 146620 152940 146630 153020
rect 146940 152940 146950 153020
rect 147260 152940 147270 153020
rect 147580 152940 147590 153020
rect 147900 152940 147910 153020
rect 148220 152940 148230 153020
rect 148540 152940 148550 153020
rect 148860 152940 148870 153020
rect 149180 152940 149190 153020
rect 149500 152940 149510 153020
rect 149820 152940 149830 153020
rect 150140 152940 150150 153020
rect 150460 152940 150470 153020
rect 150780 152940 150790 153020
rect 151100 152940 151110 153020
rect 151420 152940 151430 153020
rect 151740 152940 151750 153020
rect 152060 152940 152070 153020
rect 152380 152940 152390 153020
rect 152700 152940 152710 153020
rect 153020 152940 153030 153020
rect 153340 152940 153350 153020
rect 153660 152940 153670 153020
rect 153980 152940 153990 153020
rect 154300 152940 154310 153020
rect 154620 152940 154630 153020
rect 154940 152940 154950 153020
rect 155260 152940 155270 153020
rect 155580 152940 155590 153020
rect 155900 152940 155910 153020
rect 141545 152920 141625 152930
rect 141865 152920 141945 152930
rect 142185 152920 142200 152930
rect 145385 152920 145465 152930
rect 145705 152920 145785 152930
rect 146025 152920 146105 152930
rect 129560 152880 129640 152890
rect 129710 152880 129790 152890
rect 141060 152880 141140 152890
rect 141210 152880 141290 152890
rect 141360 152880 141440 152890
rect 129640 152800 129650 152880
rect 129790 152800 129800 152880
rect 141140 152800 141150 152880
rect 141290 152800 141300 152880
rect 141440 152800 141450 152880
rect 141625 152840 141635 152920
rect 141945 152840 141955 152920
rect 145465 152840 145475 152920
rect 145785 152840 145795 152920
rect 146105 152840 146115 152920
rect 146700 152860 146780 152870
rect 147020 152860 147100 152870
rect 147340 152860 147420 152870
rect 147660 152860 147740 152870
rect 147980 152860 148060 152870
rect 148300 152860 148380 152870
rect 148620 152860 148700 152870
rect 148940 152860 149020 152870
rect 149260 152860 149340 152870
rect 149580 152860 149660 152870
rect 149900 152860 149980 152870
rect 150220 152860 150300 152870
rect 150540 152860 150620 152870
rect 150860 152860 150940 152870
rect 151180 152860 151260 152870
rect 151500 152860 151580 152870
rect 151820 152860 151900 152870
rect 152140 152860 152220 152870
rect 152460 152860 152540 152870
rect 152780 152860 152860 152870
rect 153100 152860 153180 152870
rect 153420 152860 153500 152870
rect 153740 152860 153820 152870
rect 154060 152860 154140 152870
rect 154380 152860 154460 152870
rect 154700 152860 154780 152870
rect 155020 152860 155100 152870
rect 155340 152860 155420 152870
rect 155660 152860 155740 152870
rect 155980 152860 156000 152870
rect 146780 152780 146790 152860
rect 147100 152780 147110 152860
rect 147420 152780 147430 152860
rect 147740 152780 147750 152860
rect 148060 152780 148070 152860
rect 148380 152780 148390 152860
rect 148700 152780 148710 152860
rect 149020 152780 149030 152860
rect 149340 152780 149350 152860
rect 149660 152780 149670 152860
rect 149980 152780 149990 152860
rect 150300 152780 150310 152860
rect 150620 152780 150630 152860
rect 150940 152780 150950 152860
rect 151260 152780 151270 152860
rect 151580 152780 151590 152860
rect 151900 152780 151910 152860
rect 152220 152780 152230 152860
rect 152540 152780 152550 152860
rect 152860 152780 152870 152860
rect 153180 152780 153190 152860
rect 153500 152780 153510 152860
rect 153820 152780 153830 152860
rect 154140 152780 154150 152860
rect 154460 152780 154470 152860
rect 154780 152780 154790 152860
rect 155100 152780 155110 152860
rect 155420 152780 155430 152860
rect 155740 152780 155750 152860
rect 60740 152759 60820 152769
rect 61060 152759 61140 152769
rect 61480 152759 61560 152769
rect 61800 152759 61880 152769
rect 74240 152759 74320 152769
rect 74560 152759 74640 152769
rect 74980 152759 75060 152769
rect 75300 152759 75380 152769
rect 87740 152759 87820 152769
rect 88060 152759 88140 152769
rect 88480 152759 88560 152769
rect 88800 152759 88880 152769
rect 101240 152759 101320 152769
rect 101560 152759 101640 152769
rect 101980 152759 102060 152769
rect 102300 152759 102380 152769
rect 114740 152759 114820 152769
rect 115060 152759 115140 152769
rect 115480 152759 115560 152769
rect 115800 152759 115880 152769
rect 128240 152759 128320 152769
rect 128560 152759 128640 152769
rect 128980 152759 129060 152769
rect 129300 152759 129380 152769
rect 141705 152760 141785 152770
rect 142025 152760 142105 152770
rect 145225 152760 145305 152770
rect 145545 152760 145625 152770
rect 145865 152760 145945 152770
rect 50070 152740 50150 152750
rect 50230 152740 50310 152750
rect 48500 152700 48640 152710
rect 48710 152700 48790 152710
rect 43785 152600 43865 152610
rect 44105 152600 44185 152610
rect 44425 152600 44505 152610
rect 44745 152600 44825 152610
rect 45065 152600 45145 152610
rect 45385 152600 45465 152610
rect 45705 152600 45785 152610
rect 46025 152600 46105 152610
rect 46345 152600 46425 152610
rect 46665 152600 46745 152610
rect 46985 152600 47065 152610
rect 47305 152600 47385 152610
rect 47625 152600 47705 152610
rect 47945 152600 48025 152610
rect 48265 152600 48345 152610
rect 36180 152540 36260 152550
rect 36500 152540 36580 152550
rect 36820 152540 36900 152550
rect 37140 152540 37220 152550
rect 37460 152540 37540 152550
rect 37780 152540 37860 152550
rect 38100 152540 38180 152550
rect 38420 152540 38500 152550
rect 38740 152540 38820 152550
rect 39060 152540 39140 152550
rect 39380 152540 39460 152550
rect 39700 152540 39780 152550
rect 40020 152540 40100 152550
rect 40340 152540 40420 152550
rect 40660 152540 40740 152550
rect 40980 152540 41060 152550
rect 41300 152540 41380 152550
rect 41620 152540 41700 152550
rect 41940 152540 42020 152550
rect 42260 152540 42340 152550
rect 42580 152540 42660 152550
rect 42900 152540 42980 152550
rect 43220 152540 43300 152550
rect 36260 152460 36270 152540
rect 36580 152460 36590 152540
rect 36900 152460 36910 152540
rect 37220 152460 37230 152540
rect 37540 152460 37550 152540
rect 37860 152460 37870 152540
rect 38180 152460 38190 152540
rect 38500 152460 38510 152540
rect 38820 152460 38830 152540
rect 39140 152460 39150 152540
rect 39460 152460 39470 152540
rect 39780 152460 39790 152540
rect 40100 152460 40110 152540
rect 40420 152460 40430 152540
rect 40740 152460 40750 152540
rect 41060 152460 41070 152540
rect 41380 152460 41390 152540
rect 41700 152460 41710 152540
rect 42020 152460 42030 152540
rect 42340 152460 42350 152540
rect 42660 152460 42670 152540
rect 42980 152460 42990 152540
rect 43300 152460 43310 152540
rect 43865 152520 43875 152600
rect 44185 152520 44195 152600
rect 44505 152520 44515 152600
rect 44825 152520 44835 152600
rect 45145 152520 45155 152600
rect 45465 152520 45475 152600
rect 45785 152520 45795 152600
rect 46105 152520 46115 152600
rect 46425 152520 46435 152600
rect 46745 152520 46755 152600
rect 47065 152520 47075 152600
rect 47385 152520 47395 152600
rect 47705 152520 47715 152600
rect 48025 152520 48035 152600
rect 48345 152520 48355 152600
rect 48500 152530 48605 152700
rect 48640 152620 48650 152700
rect 48790 152620 48800 152700
rect 50150 152660 50160 152740
rect 50230 152660 50240 152740
rect 50310 152660 50320 152740
rect 60060 152700 60140 152710
rect 60210 152700 60290 152710
rect 60360 152700 60440 152710
rect 60140 152620 60150 152700
rect 60290 152620 60300 152700
rect 60440 152620 60450 152700
rect 60820 152679 60830 152759
rect 61140 152679 61150 152759
rect 61560 152679 61570 152759
rect 61880 152679 61890 152759
rect 62060 152700 62140 152710
rect 62210 152700 62290 152710
rect 73560 152700 73640 152710
rect 73710 152700 73790 152710
rect 73860 152700 73940 152710
rect 62140 152620 62150 152700
rect 62290 152620 62300 152700
rect 73640 152620 73650 152700
rect 73790 152620 73800 152700
rect 73940 152620 73950 152700
rect 74320 152679 74330 152759
rect 74640 152679 74650 152759
rect 75060 152679 75070 152759
rect 75380 152679 75390 152759
rect 75560 152700 75640 152710
rect 75710 152700 75790 152710
rect 87060 152700 87140 152710
rect 87210 152700 87290 152710
rect 87360 152700 87440 152710
rect 75640 152620 75650 152700
rect 75790 152620 75800 152700
rect 87140 152620 87150 152700
rect 87290 152620 87300 152700
rect 87440 152620 87450 152700
rect 87820 152679 87830 152759
rect 88140 152679 88150 152759
rect 88560 152679 88570 152759
rect 88880 152679 88890 152759
rect 89060 152700 89140 152710
rect 89210 152700 89290 152710
rect 100560 152700 100640 152710
rect 100710 152700 100790 152710
rect 100860 152700 100940 152710
rect 89140 152620 89150 152700
rect 89290 152620 89300 152700
rect 100640 152620 100650 152700
rect 100790 152620 100800 152700
rect 100940 152620 100950 152700
rect 101320 152679 101330 152759
rect 101640 152679 101650 152759
rect 102060 152679 102070 152759
rect 102380 152679 102390 152759
rect 114820 152679 114830 152759
rect 115140 152679 115150 152759
rect 115560 152679 115570 152759
rect 115880 152679 115890 152759
rect 116060 152700 116140 152710
rect 116210 152700 116290 152710
rect 127560 152700 127640 152710
rect 127710 152700 127790 152710
rect 127860 152700 127940 152710
rect 116140 152620 116150 152700
rect 116290 152620 116300 152700
rect 127640 152620 127650 152700
rect 127790 152620 127800 152700
rect 127940 152620 127950 152700
rect 128320 152679 128330 152759
rect 128640 152679 128650 152759
rect 129060 152679 129070 152759
rect 129380 152679 129390 152759
rect 129560 152700 129640 152710
rect 129710 152700 129790 152710
rect 141060 152700 141140 152710
rect 141210 152700 141290 152710
rect 141360 152700 141440 152710
rect 129640 152620 129650 152700
rect 129790 152620 129800 152700
rect 141140 152620 141150 152700
rect 141290 152620 141300 152700
rect 141440 152620 141450 152700
rect 141785 152680 141795 152760
rect 142105 152680 142115 152760
rect 145305 152680 145315 152760
rect 145625 152680 145635 152760
rect 145945 152680 145955 152760
rect 146540 152700 146620 152710
rect 146860 152700 146940 152710
rect 147180 152700 147260 152710
rect 147500 152700 147580 152710
rect 147820 152700 147900 152710
rect 148140 152700 148220 152710
rect 148460 152700 148540 152710
rect 148780 152700 148860 152710
rect 149100 152700 149180 152710
rect 149420 152700 149500 152710
rect 149740 152700 149820 152710
rect 150060 152700 150140 152710
rect 150380 152700 150460 152710
rect 150700 152700 150780 152710
rect 151020 152700 151100 152710
rect 151340 152700 151420 152710
rect 151660 152700 151740 152710
rect 151980 152700 152060 152710
rect 152300 152700 152380 152710
rect 152620 152700 152700 152710
rect 152940 152700 153020 152710
rect 153260 152700 153340 152710
rect 153580 152700 153660 152710
rect 153900 152700 153980 152710
rect 154220 152700 154300 152710
rect 154540 152700 154620 152710
rect 154860 152700 154940 152710
rect 155180 152700 155260 152710
rect 155500 152700 155580 152710
rect 155820 152700 155900 152710
rect 146620 152620 146630 152700
rect 146940 152620 146950 152700
rect 147260 152620 147270 152700
rect 147580 152620 147590 152700
rect 147900 152620 147910 152700
rect 148220 152620 148230 152700
rect 148540 152620 148550 152700
rect 148860 152620 148870 152700
rect 149180 152620 149190 152700
rect 149500 152620 149510 152700
rect 149820 152620 149830 152700
rect 150140 152620 150150 152700
rect 150460 152620 150470 152700
rect 150780 152620 150790 152700
rect 151100 152620 151110 152700
rect 151420 152620 151430 152700
rect 151740 152620 151750 152700
rect 152060 152620 152070 152700
rect 152380 152620 152390 152700
rect 152700 152620 152710 152700
rect 153020 152620 153030 152700
rect 153340 152620 153350 152700
rect 153660 152620 153670 152700
rect 153980 152620 153990 152700
rect 154300 152620 154310 152700
rect 154620 152620 154630 152700
rect 154940 152620 154950 152700
rect 155260 152620 155270 152700
rect 155580 152620 155590 152700
rect 155900 152620 155910 152700
rect 60580 152599 60660 152609
rect 60900 152599 60980 152609
rect 61320 152599 61400 152609
rect 61640 152599 61720 152609
rect 74080 152599 74160 152609
rect 74400 152599 74480 152609
rect 74820 152599 74900 152609
rect 75140 152599 75220 152609
rect 87580 152599 87660 152609
rect 87900 152599 87980 152609
rect 88320 152599 88400 152609
rect 88640 152599 88720 152609
rect 101080 152599 101160 152609
rect 101400 152599 101480 152609
rect 101820 152599 101900 152609
rect 102140 152599 102220 152609
rect 114580 152599 114660 152609
rect 114900 152599 114980 152609
rect 115320 152599 115400 152609
rect 115640 152599 115720 152609
rect 128080 152599 128160 152609
rect 128400 152599 128480 152609
rect 128820 152599 128900 152609
rect 129140 152599 129220 152609
rect 141545 152600 141625 152610
rect 141865 152600 141945 152610
rect 142185 152600 142200 152610
rect 145385 152600 145465 152610
rect 145705 152600 145785 152610
rect 146025 152600 146105 152610
rect 48500 152520 48640 152530
rect 48710 152520 48790 152530
rect 60060 152520 60140 152530
rect 60210 152520 60290 152530
rect 60360 152520 60440 152530
rect 43945 152440 44025 152450
rect 44265 152440 44345 152450
rect 44585 152440 44665 152450
rect 44905 152440 44985 152450
rect 45225 152440 45305 152450
rect 45545 152440 45625 152450
rect 45865 152440 45945 152450
rect 46185 152440 46265 152450
rect 46505 152440 46585 152450
rect 46825 152440 46905 152450
rect 47145 152440 47225 152450
rect 47465 152440 47545 152450
rect 47785 152440 47865 152450
rect 48105 152440 48185 152450
rect 36020 152380 36100 152390
rect 36340 152380 36420 152390
rect 36660 152380 36740 152390
rect 36980 152380 37060 152390
rect 37300 152380 37380 152390
rect 37620 152380 37700 152390
rect 37940 152380 38020 152390
rect 38260 152380 38340 152390
rect 38580 152380 38660 152390
rect 38900 152380 38980 152390
rect 39220 152380 39300 152390
rect 39540 152380 39620 152390
rect 39860 152380 39940 152390
rect 40180 152380 40260 152390
rect 40500 152380 40580 152390
rect 40820 152380 40900 152390
rect 41140 152380 41220 152390
rect 41460 152380 41540 152390
rect 41780 152380 41860 152390
rect 42100 152380 42180 152390
rect 42420 152380 42500 152390
rect 42740 152380 42820 152390
rect 43060 152380 43140 152390
rect 43380 152380 43460 152390
rect 36100 152300 36110 152380
rect 36420 152300 36430 152380
rect 36740 152300 36750 152380
rect 37060 152300 37070 152380
rect 37380 152300 37390 152380
rect 37700 152300 37710 152380
rect 38020 152300 38030 152380
rect 38340 152300 38350 152380
rect 38660 152300 38670 152380
rect 38980 152300 38990 152380
rect 39300 152300 39310 152380
rect 39620 152300 39630 152380
rect 39940 152300 39950 152380
rect 40260 152300 40270 152380
rect 40580 152300 40590 152380
rect 40900 152300 40910 152380
rect 41220 152300 41230 152380
rect 41540 152300 41550 152380
rect 41860 152300 41870 152380
rect 42180 152300 42190 152380
rect 42500 152300 42510 152380
rect 42820 152300 42830 152380
rect 43140 152300 43150 152380
rect 43460 152300 43470 152380
rect 44025 152360 44035 152440
rect 44345 152360 44355 152440
rect 44665 152360 44675 152440
rect 44985 152360 44995 152440
rect 45305 152360 45315 152440
rect 45625 152360 45635 152440
rect 45945 152360 45955 152440
rect 46265 152360 46275 152440
rect 46585 152360 46595 152440
rect 46905 152360 46915 152440
rect 47225 152360 47235 152440
rect 47545 152360 47555 152440
rect 47865 152360 47875 152440
rect 48185 152360 48195 152440
rect 48500 152350 48605 152520
rect 48640 152440 48650 152520
rect 48790 152440 48800 152520
rect 60140 152440 60150 152520
rect 60290 152440 60300 152520
rect 60440 152440 60450 152520
rect 60660 152519 60670 152599
rect 60980 152519 60990 152599
rect 61400 152519 61410 152599
rect 61720 152519 61730 152599
rect 62060 152520 62140 152530
rect 62210 152520 62290 152530
rect 73560 152520 73640 152530
rect 73710 152520 73790 152530
rect 73860 152520 73940 152530
rect 60740 152439 60820 152449
rect 61060 152439 61140 152449
rect 61480 152439 61560 152449
rect 61800 152439 61880 152449
rect 62140 152440 62150 152520
rect 62290 152440 62300 152520
rect 73640 152440 73650 152520
rect 73790 152440 73800 152520
rect 73940 152440 73950 152520
rect 74160 152519 74170 152599
rect 74480 152519 74490 152599
rect 74900 152519 74910 152599
rect 75220 152519 75230 152599
rect 75560 152520 75640 152530
rect 75710 152520 75790 152530
rect 87060 152520 87140 152530
rect 87210 152520 87290 152530
rect 87360 152520 87440 152530
rect 74240 152439 74320 152449
rect 74560 152439 74640 152449
rect 74980 152439 75060 152449
rect 75300 152439 75380 152449
rect 75640 152440 75650 152520
rect 75790 152440 75800 152520
rect 87140 152440 87150 152520
rect 87290 152440 87300 152520
rect 87440 152440 87450 152520
rect 87660 152519 87670 152599
rect 87980 152519 87990 152599
rect 88400 152519 88410 152599
rect 88720 152519 88730 152599
rect 89060 152520 89140 152530
rect 89210 152520 89290 152530
rect 100560 152520 100640 152530
rect 100710 152520 100790 152530
rect 100860 152520 100940 152530
rect 87740 152439 87820 152449
rect 88060 152439 88140 152449
rect 88480 152439 88560 152449
rect 88800 152439 88880 152449
rect 89140 152440 89150 152520
rect 89290 152440 89300 152520
rect 100640 152440 100650 152520
rect 100790 152440 100800 152520
rect 100940 152440 100950 152520
rect 101160 152519 101170 152599
rect 101480 152519 101490 152599
rect 101900 152519 101910 152599
rect 102220 152519 102230 152599
rect 114660 152519 114670 152599
rect 114980 152519 114990 152599
rect 115400 152519 115410 152599
rect 115720 152519 115730 152599
rect 116060 152520 116140 152530
rect 116210 152520 116290 152530
rect 127560 152520 127640 152530
rect 127710 152520 127790 152530
rect 127860 152520 127940 152530
rect 101240 152439 101320 152449
rect 101560 152439 101640 152449
rect 101980 152439 102060 152449
rect 102300 152439 102380 152449
rect 114740 152439 114820 152449
rect 115060 152439 115140 152449
rect 115480 152439 115560 152449
rect 115800 152439 115880 152449
rect 116140 152440 116150 152520
rect 116290 152440 116300 152520
rect 127640 152440 127650 152520
rect 127790 152440 127800 152520
rect 127940 152440 127950 152520
rect 128160 152519 128170 152599
rect 128480 152519 128490 152599
rect 128900 152519 128910 152599
rect 129220 152519 129230 152599
rect 129560 152520 129640 152530
rect 129710 152520 129790 152530
rect 141060 152520 141140 152530
rect 141210 152520 141290 152530
rect 141360 152520 141440 152530
rect 141625 152520 141635 152600
rect 141945 152520 141955 152600
rect 145465 152520 145475 152600
rect 145785 152520 145795 152600
rect 146105 152520 146115 152600
rect 146700 152540 146780 152550
rect 147020 152540 147100 152550
rect 147340 152540 147420 152550
rect 147660 152540 147740 152550
rect 147980 152540 148060 152550
rect 148300 152540 148380 152550
rect 148620 152540 148700 152550
rect 148940 152540 149020 152550
rect 149260 152540 149340 152550
rect 149580 152540 149660 152550
rect 149900 152540 149980 152550
rect 150220 152540 150300 152550
rect 150540 152540 150620 152550
rect 150860 152540 150940 152550
rect 151180 152540 151260 152550
rect 151500 152540 151580 152550
rect 151820 152540 151900 152550
rect 152140 152540 152220 152550
rect 152460 152540 152540 152550
rect 152780 152540 152860 152550
rect 153100 152540 153180 152550
rect 153420 152540 153500 152550
rect 153740 152540 153820 152550
rect 154060 152540 154140 152550
rect 154380 152540 154460 152550
rect 154700 152540 154780 152550
rect 155020 152540 155100 152550
rect 155340 152540 155420 152550
rect 155660 152540 155740 152550
rect 155980 152540 156000 152550
rect 128240 152439 128320 152449
rect 128560 152439 128640 152449
rect 128980 152439 129060 152449
rect 129300 152439 129380 152449
rect 129640 152440 129650 152520
rect 129790 152440 129800 152520
rect 141140 152440 141150 152520
rect 141290 152440 141300 152520
rect 141440 152440 141450 152520
rect 146780 152460 146790 152540
rect 147100 152460 147110 152540
rect 147420 152460 147430 152540
rect 147740 152460 147750 152540
rect 148060 152460 148070 152540
rect 148380 152460 148390 152540
rect 148700 152460 148710 152540
rect 149020 152460 149030 152540
rect 149340 152460 149350 152540
rect 149660 152460 149670 152540
rect 149980 152460 149990 152540
rect 150300 152460 150310 152540
rect 150620 152460 150630 152540
rect 150940 152460 150950 152540
rect 151260 152460 151270 152540
rect 151580 152460 151590 152540
rect 151900 152460 151910 152540
rect 152220 152460 152230 152540
rect 152540 152460 152550 152540
rect 152860 152460 152870 152540
rect 153180 152460 153190 152540
rect 153500 152460 153510 152540
rect 153820 152460 153830 152540
rect 154140 152460 154150 152540
rect 154460 152460 154470 152540
rect 154780 152460 154790 152540
rect 155100 152460 155110 152540
rect 155420 152460 155430 152540
rect 155740 152460 155750 152540
rect 141705 152440 141785 152450
rect 142025 152440 142105 152450
rect 145225 152440 145305 152450
rect 145545 152440 145625 152450
rect 145865 152440 145945 152450
rect 49180 152370 49210 152400
rect 49300 152370 49330 152400
rect 49420 152370 49450 152400
rect 49540 152370 49570 152400
rect 49660 152370 49690 152400
rect 49780 152370 49810 152400
rect 49900 152370 49930 152400
rect 50020 152370 50050 152400
rect 50140 152370 50170 152400
rect 50260 152370 50290 152400
rect 50380 152370 50410 152400
rect 50500 152370 50530 152400
rect 50620 152370 50650 152400
rect 50740 152370 50770 152400
rect 50860 152370 50890 152400
rect 50980 152370 51010 152400
rect 51100 152370 51130 152400
rect 51220 152370 51250 152400
rect 51340 152370 51370 152400
rect 51460 152370 51490 152400
rect 51580 152370 51610 152400
rect 51700 152370 51730 152400
rect 51820 152370 51850 152400
rect 51940 152370 51970 152400
rect 52060 152370 52090 152400
rect 52180 152370 52210 152400
rect 52300 152370 52330 152400
rect 52420 152370 52450 152400
rect 52540 152370 52570 152400
rect 52660 152370 52690 152400
rect 52780 152370 52810 152400
rect 52900 152370 52930 152400
rect 53020 152370 53050 152400
rect 53140 152370 53170 152400
rect 53260 152370 53290 152400
rect 53380 152370 53410 152400
rect 53500 152370 53530 152400
rect 53620 152370 53650 152400
rect 53740 152370 53770 152400
rect 53860 152370 53890 152400
rect 53980 152370 54010 152400
rect 54100 152370 54130 152400
rect 54220 152370 54250 152400
rect 54340 152370 54370 152400
rect 54460 152370 54490 152400
rect 54580 152370 54610 152400
rect 54700 152370 54730 152400
rect 54820 152370 54850 152400
rect 54940 152370 54970 152400
rect 55060 152370 55090 152400
rect 55180 152370 55210 152400
rect 55300 152370 55330 152400
rect 55420 152370 55450 152400
rect 55540 152370 55570 152400
rect 55660 152370 55690 152400
rect 55780 152370 55810 152400
rect 55900 152370 55930 152400
rect 56020 152370 56050 152400
rect 56140 152370 56170 152400
rect 56260 152370 56290 152400
rect 56380 152370 56410 152400
rect 56500 152370 56530 152400
rect 56620 152370 56650 152400
rect 56740 152370 56770 152400
rect 56860 152370 56890 152400
rect 56980 152370 57010 152400
rect 57100 152370 57130 152400
rect 57220 152370 57250 152400
rect 57340 152370 57370 152400
rect 57460 152370 57490 152400
rect 57580 152370 57610 152400
rect 57700 152370 57730 152400
rect 57820 152370 57850 152400
rect 57940 152370 57970 152400
rect 58060 152370 58090 152400
rect 58180 152370 58210 152400
rect 58300 152370 58330 152400
rect 58420 152370 58450 152400
rect 58540 152370 58570 152400
rect 58660 152370 58690 152400
rect 58780 152370 58810 152400
rect 58900 152370 58930 152400
rect 59020 152370 59050 152400
rect 59140 152370 59170 152400
rect 59260 152370 59290 152400
rect 59380 152370 59410 152400
rect 59500 152370 59530 152400
rect 59620 152370 59650 152400
rect 59740 152370 59770 152400
rect 59860 152370 59890 152400
rect 48500 152340 48640 152350
rect 48710 152340 48790 152350
rect 49060 152340 49120 152370
rect 49180 152340 49240 152370
rect 49300 152340 49360 152370
rect 49420 152340 49480 152370
rect 49540 152340 49600 152370
rect 49660 152340 49720 152370
rect 49780 152340 49840 152370
rect 49900 152340 49960 152370
rect 50020 152340 50080 152370
rect 50140 152340 50200 152370
rect 50260 152340 50320 152370
rect 50380 152340 50440 152370
rect 50500 152340 50560 152370
rect 50620 152340 50680 152370
rect 50740 152340 50800 152370
rect 50860 152340 50920 152370
rect 50980 152340 51040 152370
rect 51100 152340 51160 152370
rect 51220 152340 51280 152370
rect 51340 152340 51400 152370
rect 51460 152340 51520 152370
rect 51580 152340 51640 152370
rect 51700 152340 51760 152370
rect 51820 152340 51880 152370
rect 51940 152340 52000 152370
rect 52060 152340 52120 152370
rect 52180 152340 52240 152370
rect 52300 152340 52360 152370
rect 52420 152340 52480 152370
rect 52540 152340 52600 152370
rect 52660 152340 52720 152370
rect 52780 152340 52840 152370
rect 52900 152340 52960 152370
rect 53020 152340 53080 152370
rect 53140 152340 53200 152370
rect 53260 152340 53320 152370
rect 53380 152340 53440 152370
rect 53500 152340 53560 152370
rect 53620 152340 53680 152370
rect 53740 152340 53800 152370
rect 53860 152340 53920 152370
rect 53980 152340 54040 152370
rect 54100 152340 54160 152370
rect 54220 152340 54280 152370
rect 54340 152340 54400 152370
rect 54460 152340 54520 152370
rect 54580 152340 54640 152370
rect 54700 152340 54760 152370
rect 54820 152340 54880 152370
rect 54940 152340 55000 152370
rect 55060 152340 55120 152370
rect 55180 152340 55240 152370
rect 55300 152340 55360 152370
rect 55420 152340 55480 152370
rect 55540 152340 55600 152370
rect 55660 152340 55720 152370
rect 55780 152340 55840 152370
rect 55900 152340 55960 152370
rect 56020 152340 56080 152370
rect 56140 152340 56200 152370
rect 56260 152340 56320 152370
rect 56380 152340 56440 152370
rect 56500 152340 56560 152370
rect 56620 152340 56680 152370
rect 56740 152340 56800 152370
rect 56860 152340 56920 152370
rect 56980 152340 57040 152370
rect 57100 152340 57160 152370
rect 57220 152340 57280 152370
rect 57340 152340 57400 152370
rect 57460 152340 57520 152370
rect 57580 152340 57640 152370
rect 57700 152340 57760 152370
rect 57820 152340 57880 152370
rect 57940 152340 58000 152370
rect 58060 152340 58120 152370
rect 58180 152340 58240 152370
rect 58300 152340 58360 152370
rect 58420 152340 58480 152370
rect 58540 152340 58600 152370
rect 58660 152340 58720 152370
rect 58780 152340 58840 152370
rect 58900 152340 58960 152370
rect 59020 152340 59080 152370
rect 59140 152340 59200 152370
rect 59260 152340 59320 152370
rect 59380 152340 59440 152370
rect 59500 152340 59560 152370
rect 59620 152340 59680 152370
rect 59740 152340 59800 152370
rect 59860 152340 59920 152370
rect 60820 152359 60830 152439
rect 61140 152359 61150 152439
rect 61560 152359 61570 152439
rect 61880 152359 61890 152439
rect 62680 152370 62710 152400
rect 73245 152370 73270 152400
rect 73360 152370 73390 152400
rect 60060 152340 60140 152350
rect 60210 152340 60290 152350
rect 60360 152340 60440 152350
rect 62060 152340 62140 152350
rect 62210 152340 62290 152350
rect 62560 152340 62620 152370
rect 62680 152340 62740 152370
rect 73245 152340 73300 152370
rect 73360 152340 73420 152370
rect 74320 152359 74330 152439
rect 74640 152359 74650 152439
rect 75060 152359 75070 152439
rect 75380 152359 75390 152439
rect 76180 152370 76210 152400
rect 86745 152370 86770 152400
rect 86860 152370 86890 152400
rect 73560 152340 73640 152350
rect 73710 152340 73790 152350
rect 73860 152340 73940 152350
rect 75560 152340 75640 152350
rect 75710 152340 75790 152350
rect 76060 152340 76120 152370
rect 76180 152340 76240 152370
rect 86745 152340 86800 152370
rect 86860 152340 86920 152370
rect 87820 152359 87830 152439
rect 88140 152359 88150 152439
rect 88560 152359 88570 152439
rect 88880 152359 88890 152439
rect 89680 152370 89710 152400
rect 100245 152370 100270 152400
rect 100360 152370 100390 152400
rect 87060 152340 87140 152350
rect 87210 152340 87290 152350
rect 87360 152340 87440 152350
rect 89060 152340 89140 152350
rect 89210 152340 89290 152350
rect 89560 152340 89620 152370
rect 89680 152340 89740 152370
rect 100245 152340 100300 152370
rect 100360 152340 100420 152370
rect 101320 152359 101330 152439
rect 101640 152359 101650 152439
rect 102060 152359 102070 152439
rect 102380 152359 102390 152439
rect 114820 152359 114830 152439
rect 115140 152359 115150 152439
rect 115560 152359 115570 152439
rect 115880 152359 115890 152439
rect 116680 152370 116710 152400
rect 127245 152370 127270 152400
rect 127360 152370 127390 152400
rect 100560 152340 100640 152350
rect 100710 152340 100790 152350
rect 100860 152340 100940 152350
rect 116060 152340 116140 152350
rect 116210 152340 116290 152350
rect 116560 152340 116620 152370
rect 116680 152340 116740 152370
rect 127245 152340 127300 152370
rect 127360 152340 127420 152370
rect 128320 152359 128330 152439
rect 128640 152359 128650 152439
rect 129060 152359 129070 152439
rect 129380 152359 129390 152439
rect 130180 152370 130210 152400
rect 140740 152370 140770 152400
rect 140860 152370 140890 152400
rect 127560 152340 127640 152350
rect 127710 152340 127790 152350
rect 127860 152340 127940 152350
rect 129560 152340 129640 152350
rect 129710 152340 129790 152350
rect 130060 152340 130120 152370
rect 130180 152340 130240 152370
rect 140740 152340 140800 152370
rect 140860 152340 140920 152370
rect 141785 152360 141795 152440
rect 142105 152360 142115 152440
rect 145305 152360 145315 152440
rect 145625 152360 145635 152440
rect 145945 152360 145955 152440
rect 146540 152380 146620 152390
rect 146860 152380 146940 152390
rect 147180 152380 147260 152390
rect 147500 152380 147580 152390
rect 147820 152380 147900 152390
rect 148140 152380 148220 152390
rect 148460 152380 148540 152390
rect 148780 152380 148860 152390
rect 149100 152380 149180 152390
rect 149420 152380 149500 152390
rect 149740 152380 149820 152390
rect 150060 152380 150140 152390
rect 150380 152380 150460 152390
rect 150700 152380 150780 152390
rect 151020 152380 151100 152390
rect 151340 152380 151420 152390
rect 151660 152380 151740 152390
rect 151980 152380 152060 152390
rect 152300 152380 152380 152390
rect 152620 152380 152700 152390
rect 152940 152380 153020 152390
rect 153260 152380 153340 152390
rect 153580 152380 153660 152390
rect 153900 152380 153980 152390
rect 154220 152380 154300 152390
rect 154540 152380 154620 152390
rect 154860 152380 154940 152390
rect 155180 152380 155260 152390
rect 155500 152380 155580 152390
rect 155820 152380 155900 152390
rect 141060 152340 141140 152350
rect 141210 152340 141290 152350
rect 141360 152340 141440 152350
rect 43785 152280 43865 152290
rect 44105 152280 44185 152290
rect 44425 152280 44505 152290
rect 44745 152280 44825 152290
rect 45065 152280 45145 152290
rect 45385 152280 45465 152290
rect 45705 152280 45785 152290
rect 46025 152280 46105 152290
rect 46345 152280 46425 152290
rect 46665 152280 46745 152290
rect 46985 152280 47065 152290
rect 47305 152280 47385 152290
rect 47625 152280 47705 152290
rect 47945 152280 48025 152290
rect 48265 152280 48345 152290
rect 36180 152220 36260 152230
rect 36500 152220 36580 152230
rect 36820 152220 36900 152230
rect 37140 152220 37220 152230
rect 37460 152220 37540 152230
rect 37780 152220 37860 152230
rect 38100 152220 38180 152230
rect 38420 152220 38500 152230
rect 38740 152220 38820 152230
rect 39060 152220 39140 152230
rect 39380 152220 39460 152230
rect 39700 152220 39780 152230
rect 36260 152140 36270 152220
rect 36580 152140 36590 152220
rect 36900 152140 36910 152220
rect 37220 152140 37230 152220
rect 37540 152140 37550 152220
rect 37860 152140 37870 152220
rect 38180 152140 38190 152220
rect 38500 152140 38510 152220
rect 38820 152140 38830 152220
rect 39140 152140 39150 152220
rect 39460 152140 39470 152220
rect 39780 152140 39790 152220
rect 43865 152200 43875 152280
rect 44185 152200 44195 152280
rect 44505 152200 44515 152280
rect 44825 152200 44835 152280
rect 45145 152200 45155 152280
rect 45465 152200 45475 152280
rect 45785 152200 45795 152280
rect 46105 152200 46115 152280
rect 46425 152200 46435 152280
rect 46745 152200 46755 152280
rect 47065 152200 47075 152280
rect 47385 152200 47395 152280
rect 47705 152200 47715 152280
rect 48025 152200 48035 152280
rect 48345 152200 48355 152280
rect 48500 152170 48605 152340
rect 48640 152260 48650 152340
rect 48790 152260 48800 152340
rect 49180 152250 49210 152280
rect 49300 152250 49330 152280
rect 49420 152250 49450 152280
rect 49540 152250 49570 152280
rect 49660 152250 49690 152280
rect 49780 152250 49810 152280
rect 49900 152250 49930 152280
rect 50020 152250 50050 152280
rect 50140 152250 50170 152280
rect 50260 152250 50290 152280
rect 50380 152250 50410 152280
rect 50500 152250 50530 152280
rect 50620 152250 50650 152280
rect 50740 152250 50770 152280
rect 50860 152250 50890 152280
rect 50980 152250 51010 152280
rect 51100 152250 51130 152280
rect 51220 152250 51250 152280
rect 51340 152250 51370 152280
rect 51460 152250 51490 152280
rect 51580 152250 51610 152280
rect 51700 152250 51730 152280
rect 51820 152250 51850 152280
rect 51940 152250 51970 152280
rect 52060 152250 52090 152280
rect 52180 152250 52210 152280
rect 52300 152250 52330 152280
rect 52420 152250 52450 152280
rect 52540 152250 52570 152280
rect 52660 152250 52690 152280
rect 52780 152250 52810 152280
rect 52900 152250 52930 152280
rect 53020 152250 53050 152280
rect 53140 152250 53170 152280
rect 53260 152250 53290 152280
rect 53380 152250 53410 152280
rect 53500 152250 53530 152280
rect 53620 152250 53650 152280
rect 53740 152250 53770 152280
rect 53860 152250 53890 152280
rect 53980 152250 54010 152280
rect 54100 152250 54130 152280
rect 54220 152250 54250 152280
rect 54340 152250 54370 152280
rect 54460 152250 54490 152280
rect 54580 152250 54610 152280
rect 54700 152250 54730 152280
rect 54820 152250 54850 152280
rect 54940 152250 54970 152280
rect 55060 152250 55090 152280
rect 55180 152250 55210 152280
rect 55300 152250 55330 152280
rect 55420 152250 55450 152280
rect 55540 152250 55570 152280
rect 55660 152250 55690 152280
rect 55780 152250 55810 152280
rect 55900 152250 55930 152280
rect 56020 152250 56050 152280
rect 56140 152250 56170 152280
rect 56260 152250 56290 152280
rect 56380 152250 56410 152280
rect 56500 152250 56530 152280
rect 56620 152250 56650 152280
rect 56740 152250 56770 152280
rect 56860 152250 56890 152280
rect 56980 152250 57010 152280
rect 57100 152250 57130 152280
rect 57220 152250 57250 152280
rect 57340 152250 57370 152280
rect 57460 152250 57490 152280
rect 57580 152250 57610 152280
rect 57700 152250 57730 152280
rect 57820 152250 57850 152280
rect 57940 152250 57970 152280
rect 58060 152250 58090 152280
rect 58180 152250 58210 152280
rect 58300 152250 58330 152280
rect 58420 152250 58450 152280
rect 58540 152250 58570 152280
rect 58660 152250 58690 152280
rect 58780 152250 58810 152280
rect 58900 152250 58930 152280
rect 59020 152250 59050 152280
rect 59140 152250 59170 152280
rect 59260 152250 59290 152280
rect 59380 152250 59410 152280
rect 59500 152250 59530 152280
rect 59620 152250 59650 152280
rect 59740 152250 59770 152280
rect 59860 152250 59890 152280
rect 60140 152260 60150 152340
rect 60290 152260 60300 152340
rect 60440 152260 60450 152340
rect 60580 152279 60660 152289
rect 60900 152279 60980 152289
rect 61320 152279 61400 152289
rect 61640 152279 61720 152289
rect 49060 152220 49120 152250
rect 49180 152220 49240 152250
rect 49300 152220 49360 152250
rect 49420 152220 49480 152250
rect 49540 152220 49600 152250
rect 49660 152220 49720 152250
rect 49780 152220 49840 152250
rect 49900 152220 49960 152250
rect 50020 152220 50080 152250
rect 50140 152220 50200 152250
rect 50260 152220 50320 152250
rect 50380 152220 50440 152250
rect 50500 152220 50560 152250
rect 50620 152220 50680 152250
rect 50740 152220 50800 152250
rect 50860 152220 50920 152250
rect 50980 152220 51040 152250
rect 51100 152220 51160 152250
rect 51220 152220 51280 152250
rect 51340 152220 51400 152250
rect 51460 152220 51520 152250
rect 51580 152220 51640 152250
rect 51700 152220 51760 152250
rect 51820 152220 51880 152250
rect 51940 152220 52000 152250
rect 52060 152220 52120 152250
rect 52180 152220 52240 152250
rect 52300 152220 52360 152250
rect 52420 152220 52480 152250
rect 52540 152220 52600 152250
rect 52660 152220 52720 152250
rect 52780 152220 52840 152250
rect 52900 152220 52960 152250
rect 53020 152220 53080 152250
rect 53140 152220 53200 152250
rect 53260 152220 53320 152250
rect 53380 152220 53440 152250
rect 53500 152220 53560 152250
rect 53620 152220 53680 152250
rect 53740 152220 53800 152250
rect 53860 152220 53920 152250
rect 53980 152220 54040 152250
rect 54100 152220 54160 152250
rect 54220 152220 54280 152250
rect 54340 152220 54400 152250
rect 54460 152220 54520 152250
rect 54580 152220 54640 152250
rect 54700 152220 54760 152250
rect 54820 152220 54880 152250
rect 54940 152220 55000 152250
rect 55060 152220 55120 152250
rect 55180 152220 55240 152250
rect 55300 152220 55360 152250
rect 55420 152220 55480 152250
rect 55540 152220 55600 152250
rect 55660 152220 55720 152250
rect 55780 152220 55840 152250
rect 55900 152220 55960 152250
rect 56020 152220 56080 152250
rect 56140 152220 56200 152250
rect 56260 152220 56320 152250
rect 56380 152220 56440 152250
rect 56500 152220 56560 152250
rect 56620 152220 56680 152250
rect 56740 152220 56800 152250
rect 56860 152220 56920 152250
rect 56980 152220 57040 152250
rect 57100 152220 57160 152250
rect 57220 152220 57280 152250
rect 57340 152220 57400 152250
rect 57460 152220 57520 152250
rect 57580 152220 57640 152250
rect 57700 152220 57760 152250
rect 57820 152220 57880 152250
rect 57940 152220 58000 152250
rect 58060 152220 58120 152250
rect 58180 152220 58240 152250
rect 58300 152220 58360 152250
rect 58420 152220 58480 152250
rect 58540 152220 58600 152250
rect 58660 152220 58720 152250
rect 58780 152220 58840 152250
rect 58900 152220 58960 152250
rect 59020 152220 59080 152250
rect 59140 152220 59200 152250
rect 59260 152220 59320 152250
rect 59380 152220 59440 152250
rect 59500 152220 59560 152250
rect 59620 152220 59680 152250
rect 59740 152220 59800 152250
rect 59860 152220 59920 152250
rect 60660 152199 60670 152279
rect 60980 152199 60990 152279
rect 61400 152199 61410 152279
rect 61720 152199 61730 152279
rect 62140 152260 62150 152340
rect 62290 152260 62300 152340
rect 62680 152250 62710 152280
rect 73245 152250 73270 152280
rect 73360 152250 73390 152280
rect 73640 152260 73650 152340
rect 73790 152260 73800 152340
rect 73940 152260 73950 152340
rect 74080 152279 74160 152289
rect 74400 152279 74480 152289
rect 74820 152279 74900 152289
rect 75140 152279 75220 152289
rect 62560 152220 62620 152250
rect 62680 152220 62740 152250
rect 73245 152220 73300 152250
rect 73360 152220 73420 152250
rect 74160 152199 74170 152279
rect 74480 152199 74490 152279
rect 74900 152199 74910 152279
rect 75220 152199 75230 152279
rect 75640 152260 75650 152340
rect 75790 152260 75800 152340
rect 76180 152250 76210 152280
rect 86745 152250 86770 152280
rect 86860 152250 86890 152280
rect 87140 152260 87150 152340
rect 87290 152260 87300 152340
rect 87440 152260 87450 152340
rect 87580 152279 87660 152289
rect 87900 152279 87980 152289
rect 88320 152279 88400 152289
rect 88640 152279 88720 152289
rect 76060 152220 76120 152250
rect 76180 152220 76240 152250
rect 86745 152220 86800 152250
rect 86860 152220 86920 152250
rect 87660 152199 87670 152279
rect 87980 152199 87990 152279
rect 88400 152199 88410 152279
rect 88720 152199 88730 152279
rect 89140 152260 89150 152340
rect 89290 152260 89300 152340
rect 89680 152250 89710 152280
rect 100245 152250 100270 152280
rect 100360 152250 100390 152280
rect 100640 152260 100650 152340
rect 100790 152260 100800 152340
rect 100940 152260 100950 152340
rect 101080 152279 101160 152289
rect 101400 152279 101480 152289
rect 101820 152279 101900 152289
rect 102140 152279 102220 152289
rect 114580 152279 114660 152289
rect 114900 152279 114980 152289
rect 115320 152279 115400 152289
rect 115640 152279 115720 152289
rect 89560 152220 89620 152250
rect 89680 152220 89740 152250
rect 100245 152220 100300 152250
rect 100360 152220 100420 152250
rect 101160 152199 101170 152279
rect 101480 152199 101490 152279
rect 101900 152199 101910 152279
rect 102220 152199 102230 152279
rect 114660 152199 114670 152279
rect 114980 152199 114990 152279
rect 115400 152199 115410 152279
rect 115720 152199 115730 152279
rect 116140 152260 116150 152340
rect 116290 152260 116300 152340
rect 116680 152250 116710 152280
rect 127245 152250 127270 152280
rect 127360 152250 127390 152280
rect 127640 152260 127650 152340
rect 127790 152260 127800 152340
rect 127940 152260 127950 152340
rect 128080 152279 128160 152289
rect 128400 152279 128480 152289
rect 128820 152279 128900 152289
rect 129140 152279 129220 152289
rect 116560 152220 116620 152250
rect 116680 152220 116740 152250
rect 127245 152220 127300 152250
rect 127360 152220 127420 152250
rect 128160 152199 128170 152279
rect 128480 152199 128490 152279
rect 128900 152199 128910 152279
rect 129220 152199 129230 152279
rect 129640 152260 129650 152340
rect 129790 152260 129800 152340
rect 130180 152250 130210 152280
rect 140740 152250 140770 152280
rect 140860 152250 140890 152280
rect 141140 152260 141150 152340
rect 141290 152260 141300 152340
rect 141440 152260 141450 152340
rect 146620 152300 146630 152380
rect 146940 152300 146950 152380
rect 147260 152300 147270 152380
rect 147580 152300 147590 152380
rect 147900 152300 147910 152380
rect 148220 152300 148230 152380
rect 148540 152300 148550 152380
rect 148860 152300 148870 152380
rect 149180 152300 149190 152380
rect 149500 152300 149510 152380
rect 149820 152300 149830 152380
rect 150140 152300 150150 152380
rect 150460 152300 150470 152380
rect 150780 152300 150790 152380
rect 151100 152300 151110 152380
rect 151420 152300 151430 152380
rect 151740 152300 151750 152380
rect 152060 152300 152070 152380
rect 152380 152300 152390 152380
rect 152700 152300 152710 152380
rect 153020 152300 153030 152380
rect 153340 152300 153350 152380
rect 153660 152300 153670 152380
rect 153980 152300 153990 152380
rect 154300 152300 154310 152380
rect 154620 152300 154630 152380
rect 154940 152300 154950 152380
rect 155260 152300 155270 152380
rect 155580 152300 155590 152380
rect 155900 152300 155910 152380
rect 141545 152280 141625 152290
rect 141865 152280 141945 152290
rect 142185 152280 142200 152290
rect 145385 152280 145465 152290
rect 145705 152280 145785 152290
rect 146025 152280 146105 152290
rect 130060 152220 130120 152250
rect 130180 152220 130240 152250
rect 140740 152220 140800 152250
rect 140860 152220 140920 152250
rect 141625 152200 141635 152280
rect 141945 152200 141955 152280
rect 145465 152200 145475 152280
rect 145785 152200 145795 152280
rect 146105 152200 146115 152280
rect 150220 152220 150300 152230
rect 150540 152220 150620 152230
rect 150860 152220 150940 152230
rect 151180 152220 151260 152230
rect 151500 152220 151580 152230
rect 151820 152220 151900 152230
rect 152140 152220 152220 152230
rect 152460 152220 152540 152230
rect 152780 152220 152860 152230
rect 153100 152220 153180 152230
rect 153420 152220 153500 152230
rect 153740 152220 153820 152230
rect 154060 152220 154140 152230
rect 154380 152220 154460 152230
rect 154700 152220 154780 152230
rect 155020 152220 155100 152230
rect 155340 152220 155420 152230
rect 155660 152220 155740 152230
rect 155980 152220 156000 152230
rect 48500 152160 48640 152170
rect 48710 152160 48790 152170
rect 60060 152160 60140 152170
rect 60210 152160 60290 152170
rect 60360 152160 60440 152170
rect 62060 152160 62140 152170
rect 62210 152160 62290 152170
rect 73560 152160 73640 152170
rect 73710 152160 73790 152170
rect 73860 152160 73940 152170
rect 75560 152160 75640 152170
rect 75710 152160 75790 152170
rect 87060 152160 87140 152170
rect 87210 152160 87290 152170
rect 87360 152160 87440 152170
rect 89060 152160 89140 152170
rect 89210 152160 89290 152170
rect 100560 152160 100640 152170
rect 100710 152160 100790 152170
rect 100860 152160 100940 152170
rect 116060 152160 116140 152170
rect 116210 152160 116290 152170
rect 127560 152160 127640 152170
rect 127710 152160 127790 152170
rect 127860 152160 127940 152170
rect 129560 152160 129640 152170
rect 129710 152160 129790 152170
rect 141060 152160 141140 152170
rect 141210 152160 141290 152170
rect 141360 152160 141440 152170
rect 36020 152060 36100 152070
rect 36340 152060 36420 152070
rect 36660 152060 36740 152070
rect 36980 152060 37060 152070
rect 37300 152060 37380 152070
rect 37620 152060 37700 152070
rect 37940 152060 38020 152070
rect 38260 152060 38340 152070
rect 38580 152060 38660 152070
rect 38900 152060 38980 152070
rect 39220 152060 39300 152070
rect 39540 152060 39620 152070
rect 36100 151980 36110 152060
rect 36420 151980 36430 152060
rect 36740 151980 36750 152060
rect 37060 151980 37070 152060
rect 37380 151980 37390 152060
rect 37700 151980 37710 152060
rect 38020 151980 38030 152060
rect 38340 151980 38350 152060
rect 38660 151980 38670 152060
rect 38980 151980 38990 152060
rect 39300 151980 39310 152060
rect 39620 151980 39630 152060
rect 48500 152000 48605 152160
rect 48640 152080 48650 152160
rect 48790 152080 48800 152160
rect 49180 152100 49210 152160
rect 49300 152100 49330 152160
rect 49420 152100 49450 152160
rect 49540 152100 49570 152160
rect 49660 152100 49690 152160
rect 49780 152100 49810 152160
rect 49900 152100 49930 152160
rect 50020 152100 50050 152160
rect 50140 152100 50170 152160
rect 50260 152100 50290 152160
rect 50380 152100 50410 152160
rect 50500 152100 50530 152160
rect 50620 152100 50650 152160
rect 50740 152100 50770 152160
rect 50860 152100 50890 152160
rect 50980 152100 51010 152160
rect 51100 152100 51130 152160
rect 51220 152100 51250 152160
rect 51340 152100 51370 152160
rect 51460 152100 51490 152160
rect 51580 152100 51610 152160
rect 51700 152100 51730 152160
rect 51820 152100 51850 152160
rect 51940 152100 51970 152160
rect 52060 152100 52090 152160
rect 52180 152100 52210 152160
rect 52300 152100 52330 152160
rect 52420 152100 52450 152160
rect 52540 152100 52570 152160
rect 52660 152100 52690 152160
rect 52780 152100 52810 152160
rect 52900 152100 52930 152160
rect 53020 152100 53050 152160
rect 53140 152100 53170 152160
rect 53260 152100 53290 152160
rect 53380 152100 53410 152160
rect 53500 152100 53530 152160
rect 53620 152100 53650 152160
rect 53740 152100 53770 152160
rect 53860 152100 53890 152160
rect 53980 152100 54010 152160
rect 54100 152100 54130 152160
rect 54220 152100 54250 152160
rect 54340 152100 54370 152160
rect 54460 152100 54490 152160
rect 54580 152100 54610 152160
rect 54700 152100 54730 152160
rect 54820 152100 54850 152160
rect 54940 152100 54970 152160
rect 55060 152100 55090 152160
rect 55180 152100 55210 152160
rect 55300 152100 55330 152160
rect 55420 152100 55450 152160
rect 55540 152100 55570 152160
rect 55660 152100 55690 152160
rect 55780 152100 55810 152160
rect 55900 152100 55930 152160
rect 56020 152100 56050 152160
rect 56140 152100 56170 152160
rect 56260 152100 56290 152160
rect 56380 152100 56410 152160
rect 56500 152100 56530 152160
rect 56620 152100 56650 152160
rect 56740 152100 56770 152160
rect 56860 152100 56890 152160
rect 56980 152100 57010 152160
rect 57100 152100 57130 152160
rect 57220 152100 57250 152160
rect 57340 152100 57370 152160
rect 57460 152100 57490 152160
rect 57580 152100 57610 152160
rect 57700 152100 57730 152160
rect 57820 152100 57850 152160
rect 57940 152100 57970 152160
rect 58060 152100 58090 152160
rect 58180 152100 58210 152160
rect 58300 152100 58330 152160
rect 58420 152100 58450 152160
rect 58540 152100 58570 152160
rect 58660 152100 58690 152160
rect 58780 152100 58810 152160
rect 58900 152100 58930 152160
rect 59020 152100 59050 152160
rect 59140 152100 59170 152160
rect 59260 152100 59290 152160
rect 59380 152100 59410 152160
rect 59500 152100 59530 152160
rect 59620 152100 59650 152160
rect 59740 152100 59770 152160
rect 59860 152100 59890 152160
rect 60140 152080 60150 152160
rect 60290 152080 60300 152160
rect 60440 152080 60450 152160
rect 62140 152080 62150 152160
rect 62290 152080 62300 152160
rect 62680 152100 62710 152160
rect 73245 152100 73270 152160
rect 73360 152100 73390 152160
rect 73640 152080 73650 152160
rect 73790 152080 73800 152160
rect 73940 152080 73950 152160
rect 75640 152080 75650 152160
rect 75790 152080 75800 152160
rect 76180 152100 76210 152160
rect 86745 152100 86770 152160
rect 86860 152100 86890 152160
rect 87140 152080 87150 152160
rect 87290 152080 87300 152160
rect 87440 152080 87450 152160
rect 89140 152080 89150 152160
rect 89290 152080 89300 152160
rect 89680 152100 89710 152160
rect 100245 152100 100270 152160
rect 100360 152100 100390 152160
rect 100640 152080 100650 152160
rect 100790 152080 100800 152160
rect 100940 152080 100950 152160
rect 116140 152080 116150 152160
rect 116290 152080 116300 152160
rect 116680 152100 116710 152160
rect 127245 152100 127270 152160
rect 127360 152100 127390 152160
rect 127640 152080 127650 152160
rect 127790 152080 127800 152160
rect 127940 152080 127950 152160
rect 129640 152080 129650 152160
rect 129790 152080 129800 152160
rect 130180 152100 130210 152160
rect 140740 152100 140770 152160
rect 140860 152100 140890 152160
rect 141140 152080 141150 152160
rect 141290 152080 141300 152160
rect 141440 152080 141450 152160
rect 150300 152140 150310 152220
rect 150620 152140 150630 152220
rect 150940 152140 150950 152220
rect 151260 152140 151270 152220
rect 151580 152140 151590 152220
rect 151900 152140 151910 152220
rect 152220 152140 152230 152220
rect 152540 152140 152550 152220
rect 152860 152140 152870 152220
rect 153180 152140 153190 152220
rect 153500 152140 153510 152220
rect 153820 152140 153830 152220
rect 154140 152140 154150 152220
rect 154460 152140 154470 152220
rect 154780 152140 154790 152220
rect 155100 152140 155110 152220
rect 155420 152140 155430 152220
rect 155740 152140 155750 152220
rect 150380 152060 150460 152070
rect 150700 152060 150780 152070
rect 151020 152060 151100 152070
rect 151340 152060 151420 152070
rect 151660 152060 151740 152070
rect 151980 152060 152060 152070
rect 152300 152060 152380 152070
rect 152620 152060 152700 152070
rect 152940 152060 153020 152070
rect 153260 152060 153340 152070
rect 153580 152060 153660 152070
rect 153900 152060 153980 152070
rect 154220 152060 154300 152070
rect 154540 152060 154620 152070
rect 154860 152060 154940 152070
rect 155180 152060 155260 152070
rect 155500 152060 155580 152070
rect 155820 152060 155900 152070
rect 150460 151980 150470 152060
rect 150780 151980 150790 152060
rect 151100 151980 151110 152060
rect 151420 151980 151430 152060
rect 151740 151980 151750 152060
rect 152060 151980 152070 152060
rect 152380 151980 152390 152060
rect 152700 151980 152710 152060
rect 153020 151980 153030 152060
rect 153340 151980 153350 152060
rect 153660 151980 153670 152060
rect 153980 151980 153990 152060
rect 154300 151980 154310 152060
rect 154620 151980 154630 152060
rect 154940 151980 154950 152060
rect 155260 151980 155270 152060
rect 155580 151980 155590 152060
rect 155900 151980 155910 152060
rect 36180 151900 36260 151910
rect 36500 151900 36580 151910
rect 36820 151900 36900 151910
rect 37140 151900 37220 151910
rect 37460 151900 37540 151910
rect 37780 151900 37860 151910
rect 38100 151900 38180 151910
rect 38420 151900 38500 151910
rect 38740 151900 38820 151910
rect 39060 151900 39140 151910
rect 39380 151900 39460 151910
rect 150540 151900 150620 151910
rect 150860 151900 150940 151910
rect 151180 151900 151260 151910
rect 151500 151900 151580 151910
rect 151820 151900 151900 151910
rect 152140 151900 152220 151910
rect 152460 151900 152540 151910
rect 152780 151900 152860 151910
rect 153100 151900 153180 151910
rect 153420 151900 153500 151910
rect 153740 151900 153820 151910
rect 154060 151900 154140 151910
rect 154380 151900 154460 151910
rect 154700 151900 154780 151910
rect 155020 151900 155100 151910
rect 155340 151900 155420 151910
rect 155660 151900 155740 151910
rect 155980 151900 156000 151910
rect 36260 151820 36270 151900
rect 36580 151820 36590 151900
rect 36900 151820 36910 151900
rect 37220 151820 37230 151900
rect 37540 151820 37550 151900
rect 37860 151820 37870 151900
rect 38180 151820 38190 151900
rect 38500 151820 38510 151900
rect 38820 151820 38830 151900
rect 39140 151820 39150 151900
rect 39460 151820 39470 151900
rect 150620 151820 150630 151900
rect 150940 151820 150950 151900
rect 151260 151820 151270 151900
rect 151580 151820 151590 151900
rect 151900 151820 151910 151900
rect 152220 151820 152230 151900
rect 152540 151820 152550 151900
rect 152860 151820 152870 151900
rect 153180 151820 153190 151900
rect 153500 151820 153510 151900
rect 153820 151820 153830 151900
rect 154140 151820 154150 151900
rect 154460 151820 154470 151900
rect 154780 151820 154790 151900
rect 155100 151820 155110 151900
rect 155420 151820 155430 151900
rect 155740 151820 155750 151900
rect 36020 151740 36100 151750
rect 36340 151740 36420 151750
rect 36660 151740 36740 151750
rect 36980 151740 37060 151750
rect 37300 151740 37380 151750
rect 37620 151740 37700 151750
rect 37940 151740 38020 151750
rect 38260 151740 38340 151750
rect 38580 151740 38660 151750
rect 38900 151740 38980 151750
rect 39220 151740 39300 151750
rect 150700 151740 150780 151750
rect 151020 151740 151100 151750
rect 151340 151740 151420 151750
rect 151660 151740 151740 151750
rect 151980 151740 152060 151750
rect 152300 151740 152380 151750
rect 152620 151740 152700 151750
rect 152940 151740 153020 151750
rect 153260 151740 153340 151750
rect 153580 151740 153660 151750
rect 153900 151740 153980 151750
rect 154220 151740 154300 151750
rect 154540 151740 154620 151750
rect 154860 151740 154940 151750
rect 155180 151740 155260 151750
rect 155500 151740 155580 151750
rect 155820 151740 155900 151750
rect 36100 151660 36110 151740
rect 36420 151660 36430 151740
rect 36740 151660 36750 151740
rect 37060 151660 37070 151740
rect 37380 151660 37390 151740
rect 37700 151660 37710 151740
rect 38020 151660 38030 151740
rect 38340 151660 38350 151740
rect 38660 151660 38670 151740
rect 38980 151660 38990 151740
rect 39300 151660 39310 151740
rect 150780 151660 150790 151740
rect 151100 151660 151110 151740
rect 151420 151660 151430 151740
rect 151740 151660 151750 151740
rect 152060 151660 152070 151740
rect 152380 151660 152390 151740
rect 152700 151660 152710 151740
rect 153020 151660 153030 151740
rect 153340 151660 153350 151740
rect 153660 151660 153670 151740
rect 153980 151660 153990 151740
rect 154300 151660 154310 151740
rect 154620 151660 154630 151740
rect 154940 151660 154950 151740
rect 155260 151660 155270 151740
rect 155580 151660 155590 151740
rect 155900 151660 155910 151740
rect 36180 151580 36260 151590
rect 36500 151580 36580 151590
rect 36820 151580 36900 151590
rect 37140 151580 37220 151590
rect 37460 151580 37540 151590
rect 37780 151580 37860 151590
rect 38100 151580 38180 151590
rect 38420 151580 38500 151590
rect 38740 151580 38820 151590
rect 39060 151580 39140 151590
rect 150860 151580 150940 151590
rect 151180 151580 151260 151590
rect 151500 151580 151580 151590
rect 151820 151580 151900 151590
rect 152140 151580 152220 151590
rect 152460 151580 152540 151590
rect 152780 151580 152860 151590
rect 153100 151580 153180 151590
rect 153420 151580 153500 151590
rect 153740 151580 153820 151590
rect 154060 151580 154140 151590
rect 154380 151580 154460 151590
rect 154700 151580 154780 151590
rect 155020 151580 155100 151590
rect 155340 151580 155420 151590
rect 155660 151580 155740 151590
rect 155980 151580 156000 151590
rect 36260 151500 36270 151580
rect 36580 151500 36590 151580
rect 36900 151500 36910 151580
rect 37220 151500 37230 151580
rect 37540 151500 37550 151580
rect 37860 151500 37870 151580
rect 38180 151500 38190 151580
rect 38500 151500 38510 151580
rect 38820 151500 38830 151580
rect 39140 151500 39150 151580
rect 150940 151500 150950 151580
rect 151260 151500 151270 151580
rect 151580 151500 151590 151580
rect 151900 151500 151910 151580
rect 152220 151500 152230 151580
rect 152540 151500 152550 151580
rect 152860 151500 152870 151580
rect 153180 151500 153190 151580
rect 153500 151500 153510 151580
rect 153820 151500 153830 151580
rect 154140 151500 154150 151580
rect 154460 151500 154470 151580
rect 154780 151500 154790 151580
rect 155100 151500 155110 151580
rect 155420 151500 155430 151580
rect 155740 151500 155750 151580
rect 36020 151420 36100 151430
rect 36340 151420 36420 151430
rect 36660 151420 36740 151430
rect 36980 151420 37060 151430
rect 37300 151420 37380 151430
rect 37620 151420 37700 151430
rect 37940 151420 38020 151430
rect 38260 151420 38340 151430
rect 38580 151420 38660 151430
rect 38900 151420 38980 151430
rect 151020 151420 151100 151430
rect 151340 151420 151420 151430
rect 151660 151420 151740 151430
rect 151980 151420 152060 151430
rect 152300 151420 152380 151430
rect 152620 151420 152700 151430
rect 152940 151420 153020 151430
rect 153260 151420 153340 151430
rect 153580 151420 153660 151430
rect 153900 151420 153980 151430
rect 154220 151420 154300 151430
rect 154540 151420 154620 151430
rect 154860 151420 154940 151430
rect 155180 151420 155260 151430
rect 155500 151420 155580 151430
rect 155820 151420 155900 151430
rect 36100 151340 36110 151420
rect 36420 151340 36430 151420
rect 36740 151340 36750 151420
rect 37060 151340 37070 151420
rect 37380 151340 37390 151420
rect 37700 151340 37710 151420
rect 38020 151340 38030 151420
rect 38340 151340 38350 151420
rect 38660 151340 38670 151420
rect 38980 151340 38990 151420
rect 151100 151340 151110 151420
rect 151420 151340 151430 151420
rect 151740 151340 151750 151420
rect 152060 151340 152070 151420
rect 152380 151340 152390 151420
rect 152700 151340 152710 151420
rect 153020 151340 153030 151420
rect 153340 151340 153350 151420
rect 153660 151340 153670 151420
rect 153980 151340 153990 151420
rect 154300 151340 154310 151420
rect 154620 151340 154630 151420
rect 154940 151340 154950 151420
rect 155260 151340 155270 151420
rect 155580 151340 155590 151420
rect 155900 151340 155910 151420
rect 36180 151260 36260 151270
rect 36500 151260 36580 151270
rect 36820 151260 36900 151270
rect 37140 151260 37220 151270
rect 37460 151260 37540 151270
rect 37780 151260 37860 151270
rect 38100 151260 38180 151270
rect 38420 151260 38500 151270
rect 38740 151260 38820 151270
rect 151180 151260 151260 151270
rect 151500 151260 151580 151270
rect 151820 151260 151900 151270
rect 152140 151260 152220 151270
rect 152460 151260 152540 151270
rect 152780 151260 152860 151270
rect 153100 151260 153180 151270
rect 153420 151260 153500 151270
rect 153740 151260 153820 151270
rect 154060 151260 154140 151270
rect 154380 151260 154460 151270
rect 154700 151260 154780 151270
rect 155020 151260 155100 151270
rect 155340 151260 155420 151270
rect 155660 151260 155740 151270
rect 155980 151260 156000 151270
rect 36260 151180 36270 151260
rect 36580 151180 36590 151260
rect 36900 151180 36910 151260
rect 37220 151180 37230 151260
rect 37540 151180 37550 151260
rect 37860 151180 37870 151260
rect 38180 151180 38190 151260
rect 38500 151180 38510 151260
rect 38820 151180 38830 151260
rect 151260 151180 151270 151260
rect 151580 151180 151590 151260
rect 151900 151180 151910 151260
rect 152220 151180 152230 151260
rect 152540 151180 152550 151260
rect 152860 151180 152870 151260
rect 153180 151180 153190 151260
rect 153500 151180 153510 151260
rect 153820 151180 153830 151260
rect 154140 151180 154150 151260
rect 154460 151180 154470 151260
rect 154780 151180 154790 151260
rect 155100 151180 155110 151260
rect 155420 151180 155430 151260
rect 155740 151180 155750 151260
rect 36020 151100 36100 151110
rect 36340 151100 36420 151110
rect 36660 151100 36740 151110
rect 36980 151100 37060 151110
rect 37300 151100 37380 151110
rect 37620 151100 37700 151110
rect 37940 151100 38020 151110
rect 38260 151100 38340 151110
rect 38580 151100 38660 151110
rect 151340 151100 151420 151110
rect 151660 151100 151740 151110
rect 151980 151100 152060 151110
rect 152300 151100 152380 151110
rect 152620 151100 152700 151110
rect 152940 151100 153020 151110
rect 153260 151100 153340 151110
rect 153580 151100 153660 151110
rect 153900 151100 153980 151110
rect 154220 151100 154300 151110
rect 154540 151100 154620 151110
rect 154860 151100 154940 151110
rect 155180 151100 155260 151110
rect 155500 151100 155580 151110
rect 155820 151100 155900 151110
rect 36100 151020 36110 151100
rect 36420 151020 36430 151100
rect 36740 151020 36750 151100
rect 37060 151020 37070 151100
rect 37380 151020 37390 151100
rect 37700 151020 37710 151100
rect 38020 151020 38030 151100
rect 38340 151020 38350 151100
rect 38660 151020 38670 151100
rect 151420 151020 151430 151100
rect 151740 151020 151750 151100
rect 152060 151020 152070 151100
rect 152380 151020 152390 151100
rect 152700 151020 152710 151100
rect 153020 151020 153030 151100
rect 153340 151020 153350 151100
rect 153660 151020 153670 151100
rect 153980 151020 153990 151100
rect 154300 151020 154310 151100
rect 154620 151020 154630 151100
rect 154940 151020 154950 151100
rect 155260 151020 155270 151100
rect 155580 151020 155590 151100
rect 155900 151020 155910 151100
rect 36180 150940 36260 150950
rect 36500 150940 36580 150950
rect 36820 150940 36900 150950
rect 37140 150940 37220 150950
rect 37460 150940 37540 150950
rect 37780 150940 37860 150950
rect 38100 150940 38180 150950
rect 38420 150940 38500 150950
rect 151500 150940 151580 150950
rect 151820 150940 151900 150950
rect 152140 150940 152220 150950
rect 152460 150940 152540 150950
rect 152780 150940 152860 150950
rect 153100 150940 153180 150950
rect 153420 150940 153500 150950
rect 153740 150940 153820 150950
rect 154060 150940 154140 150950
rect 154380 150940 154460 150950
rect 154700 150940 154780 150950
rect 155020 150940 155100 150950
rect 155340 150940 155420 150950
rect 155660 150940 155740 150950
rect 155980 150940 156000 150950
rect 36260 150860 36270 150940
rect 36580 150860 36590 150940
rect 36900 150860 36910 150940
rect 37220 150860 37230 150940
rect 37540 150860 37550 150940
rect 37860 150860 37870 150940
rect 38180 150860 38190 150940
rect 38500 150860 38510 150940
rect 151580 150860 151590 150940
rect 151900 150860 151910 150940
rect 152220 150860 152230 150940
rect 152540 150860 152550 150940
rect 152860 150860 152870 150940
rect 153180 150860 153190 150940
rect 153500 150860 153510 150940
rect 153820 150860 153830 150940
rect 154140 150860 154150 150940
rect 154460 150860 154470 150940
rect 154780 150860 154790 150940
rect 155100 150860 155110 150940
rect 155420 150860 155430 150940
rect 155740 150860 155750 150940
rect 36020 150780 36100 150790
rect 36340 150780 36420 150790
rect 36660 150780 36740 150790
rect 36980 150780 37060 150790
rect 37300 150780 37380 150790
rect 37620 150780 37700 150790
rect 37940 150780 38020 150790
rect 38260 150780 38340 150790
rect 151660 150780 151740 150790
rect 151980 150780 152060 150790
rect 152300 150780 152380 150790
rect 152620 150780 152700 150790
rect 152940 150780 153020 150790
rect 153260 150780 153340 150790
rect 153580 150780 153660 150790
rect 153900 150780 153980 150790
rect 154220 150780 154300 150790
rect 154540 150780 154620 150790
rect 154860 150780 154940 150790
rect 155180 150780 155260 150790
rect 155500 150780 155580 150790
rect 155820 150780 155900 150790
rect 36100 150700 36110 150780
rect 36420 150700 36430 150780
rect 36740 150700 36750 150780
rect 37060 150700 37070 150780
rect 37380 150700 37390 150780
rect 37700 150700 37710 150780
rect 38020 150700 38030 150780
rect 38340 150700 38350 150780
rect 151740 150700 151750 150780
rect 152060 150700 152070 150780
rect 152380 150700 152390 150780
rect 152700 150700 152710 150780
rect 153020 150700 153030 150780
rect 153340 150700 153350 150780
rect 153660 150700 153670 150780
rect 153980 150700 153990 150780
rect 154300 150700 154310 150780
rect 154620 150700 154630 150780
rect 154940 150700 154950 150780
rect 155260 150700 155270 150780
rect 155580 150700 155590 150780
rect 155900 150700 155910 150780
rect 36180 150620 36260 150630
rect 36500 150620 36580 150630
rect 36820 150620 36900 150630
rect 37140 150620 37220 150630
rect 37460 150620 37540 150630
rect 37780 150620 37860 150630
rect 38100 150620 38180 150630
rect 151820 150620 151900 150630
rect 152140 150620 152220 150630
rect 152460 150620 152540 150630
rect 152780 150620 152860 150630
rect 153100 150620 153180 150630
rect 153420 150620 153500 150630
rect 153740 150620 153820 150630
rect 154060 150620 154140 150630
rect 154380 150620 154460 150630
rect 154700 150620 154780 150630
rect 155020 150620 155100 150630
rect 155340 150620 155420 150630
rect 155660 150620 155740 150630
rect 155980 150620 156000 150630
rect 36260 150540 36270 150620
rect 36580 150540 36590 150620
rect 36900 150540 36910 150620
rect 37220 150540 37230 150620
rect 37540 150540 37550 150620
rect 37860 150540 37870 150620
rect 38180 150540 38190 150620
rect 151900 150540 151910 150620
rect 152220 150540 152230 150620
rect 152540 150540 152550 150620
rect 152860 150540 152870 150620
rect 153180 150540 153190 150620
rect 153500 150540 153510 150620
rect 153820 150540 153830 150620
rect 154140 150540 154150 150620
rect 154460 150540 154470 150620
rect 154780 150540 154790 150620
rect 155100 150540 155110 150620
rect 155420 150540 155430 150620
rect 155740 150540 155750 150620
rect 36020 150460 36100 150470
rect 36340 150460 36420 150470
rect 36660 150460 36740 150470
rect 36980 150460 37060 150470
rect 37300 150460 37380 150470
rect 37620 150460 37700 150470
rect 37940 150460 38020 150470
rect 151980 150460 152060 150470
rect 152300 150460 152380 150470
rect 152620 150460 152700 150470
rect 152940 150460 153020 150470
rect 153260 150460 153340 150470
rect 153580 150460 153660 150470
rect 153900 150460 153980 150470
rect 154220 150460 154300 150470
rect 154540 150460 154620 150470
rect 154860 150460 154940 150470
rect 155180 150460 155260 150470
rect 155500 150460 155580 150470
rect 155820 150460 155900 150470
rect 36100 150380 36110 150460
rect 36420 150380 36430 150460
rect 36740 150380 36750 150460
rect 37060 150380 37070 150460
rect 37380 150380 37390 150460
rect 37700 150380 37710 150460
rect 38020 150380 38030 150460
rect 152060 150380 152070 150460
rect 152380 150380 152390 150460
rect 152700 150380 152710 150460
rect 153020 150380 153030 150460
rect 153340 150380 153350 150460
rect 153660 150380 153670 150460
rect 153980 150380 153990 150460
rect 154300 150380 154310 150460
rect 154620 150380 154630 150460
rect 154940 150380 154950 150460
rect 155260 150380 155270 150460
rect 155580 150380 155590 150460
rect 155900 150380 155910 150460
rect 36180 150300 36260 150310
rect 36500 150300 36580 150310
rect 36820 150300 36900 150310
rect 37140 150300 37220 150310
rect 37460 150300 37540 150310
rect 37780 150300 37860 150310
rect 152140 150300 152220 150310
rect 152460 150300 152540 150310
rect 152780 150300 152860 150310
rect 153100 150300 153180 150310
rect 153420 150300 153500 150310
rect 153740 150300 153820 150310
rect 154060 150300 154140 150310
rect 154380 150300 154460 150310
rect 154700 150300 154780 150310
rect 155020 150300 155100 150310
rect 155340 150300 155420 150310
rect 155660 150300 155740 150310
rect 155980 150300 156000 150310
rect 36260 150220 36270 150300
rect 36580 150220 36590 150300
rect 36900 150220 36910 150300
rect 37220 150220 37230 150300
rect 37540 150220 37550 150300
rect 37860 150220 37870 150300
rect 152220 150220 152230 150300
rect 152540 150220 152550 150300
rect 152860 150220 152870 150300
rect 153180 150220 153190 150300
rect 153500 150220 153510 150300
rect 153820 150220 153830 150300
rect 154140 150220 154150 150300
rect 154460 150220 154470 150300
rect 154780 150220 154790 150300
rect 155100 150220 155110 150300
rect 155420 150220 155430 150300
rect 155740 150220 155750 150300
rect 36020 150140 36100 150150
rect 36340 150140 36420 150150
rect 36660 150140 36740 150150
rect 36980 150140 37060 150150
rect 37300 150140 37380 150150
rect 37620 150140 37700 150150
rect 152300 150140 152380 150150
rect 152620 150140 152700 150150
rect 152940 150140 153020 150150
rect 153260 150140 153340 150150
rect 153580 150140 153660 150150
rect 153900 150140 153980 150150
rect 154220 150140 154300 150150
rect 154540 150140 154620 150150
rect 154860 150140 154940 150150
rect 155180 150140 155260 150150
rect 155500 150140 155580 150150
rect 155820 150140 155900 150150
rect 36100 150060 36110 150140
rect 36420 150060 36430 150140
rect 36740 150060 36750 150140
rect 37060 150060 37070 150140
rect 37380 150060 37390 150140
rect 37700 150060 37710 150140
rect 152380 150060 152390 150140
rect 152700 150060 152710 150140
rect 153020 150060 153030 150140
rect 153340 150060 153350 150140
rect 153660 150060 153670 150140
rect 153980 150060 153990 150140
rect 154300 150060 154310 150140
rect 154620 150060 154630 150140
rect 154940 150060 154950 150140
rect 155260 150060 155270 150140
rect 155580 150060 155590 150140
rect 155900 150060 155910 150140
rect 36180 149980 36260 149990
rect 36500 149980 36580 149990
rect 36820 149980 36900 149990
rect 37140 149980 37220 149990
rect 37460 149980 37540 149990
rect 36260 149900 36270 149980
rect 36580 149900 36590 149980
rect 36900 149900 36910 149980
rect 37220 149900 37230 149980
rect 37540 149900 37550 149980
rect 48500 149950 48605 150000
rect 51775 149999 60500 150000
rect 73245 149999 74000 150000
rect 86745 149999 87500 150000
rect 100245 149999 101000 150000
rect 127245 149999 128000 150000
rect 48500 149940 48640 149950
rect 51775 149940 60570 149999
rect 62060 149940 62140 149950
rect 36020 149820 36100 149830
rect 36340 149820 36420 149830
rect 36660 149820 36740 149830
rect 36980 149820 37060 149830
rect 37300 149820 37380 149830
rect 37620 149820 37700 149830
rect 41460 149820 41540 149830
rect 41780 149820 41860 149830
rect 42100 149820 42180 149830
rect 42420 149820 42500 149830
rect 42740 149820 42820 149830
rect 43060 149820 43140 149830
rect 43380 149820 43460 149830
rect 43785 149820 43865 149830
rect 44105 149820 44185 149830
rect 44425 149820 44505 149830
rect 44745 149820 44825 149830
rect 45065 149820 45145 149830
rect 45385 149820 45465 149830
rect 45705 149820 45785 149830
rect 46025 149820 46105 149830
rect 46345 149820 46425 149830
rect 46665 149820 46745 149830
rect 46985 149820 47065 149830
rect 47305 149820 47385 149830
rect 47625 149820 47705 149830
rect 47945 149820 48025 149830
rect 48265 149820 48345 149830
rect 36100 149740 36110 149820
rect 36420 149740 36430 149820
rect 36740 149740 36750 149820
rect 37060 149740 37070 149820
rect 37380 149740 37390 149820
rect 37700 149740 37710 149820
rect 41540 149740 41550 149820
rect 41860 149740 41870 149820
rect 42180 149740 42190 149820
rect 42500 149740 42510 149820
rect 42820 149740 42830 149820
rect 43140 149740 43150 149820
rect 43460 149740 43470 149820
rect 43865 149740 43875 149820
rect 44185 149740 44195 149820
rect 44505 149740 44515 149820
rect 44825 149740 44835 149820
rect 45145 149740 45155 149820
rect 45465 149740 45475 149820
rect 45785 149740 45795 149820
rect 46105 149740 46115 149820
rect 46425 149740 46435 149820
rect 46745 149740 46755 149820
rect 47065 149740 47075 149820
rect 47385 149740 47395 149820
rect 47705 149740 47715 149820
rect 48025 149740 48035 149820
rect 48345 149740 48355 149820
rect 48500 149810 48605 149940
rect 48640 149860 48650 149940
rect 48870 149880 48900 149940
rect 48990 149880 49020 149940
rect 49110 149880 49140 149940
rect 49230 149880 49260 149940
rect 49350 149880 49380 149940
rect 49470 149880 49500 149940
rect 49590 149880 49620 149940
rect 49710 149880 49740 149940
rect 49830 149880 49860 149940
rect 49950 149880 49980 149940
rect 50070 149880 50100 149940
rect 50190 149880 50220 149940
rect 50310 149880 50340 149940
rect 50430 149880 50460 149940
rect 50550 149880 50580 149940
rect 50670 149880 50700 149940
rect 50790 149880 50820 149940
rect 50910 149880 50940 149940
rect 51030 149880 51060 149940
rect 51150 149880 51180 149940
rect 51270 149880 51300 149940
rect 51390 149880 51420 149940
rect 51510 149880 51540 149940
rect 51630 149880 51660 149940
rect 51750 149880 60570 149940
rect 48970 149820 51150 149830
rect 51775 149820 60570 149880
rect 62140 149860 62150 149940
rect 62370 149880 62400 149940
rect 62490 149880 62520 149940
rect 62610 149880 62640 149940
rect 62730 149880 62755 149940
rect 48500 149800 48640 149810
rect 48500 149670 48605 149800
rect 48640 149720 48650 149800
rect 36180 149660 36260 149670
rect 36500 149660 36580 149670
rect 36820 149660 36900 149670
rect 37140 149660 37220 149670
rect 37460 149660 37540 149670
rect 41300 149660 41380 149670
rect 41620 149660 41700 149670
rect 41940 149660 42020 149670
rect 42260 149660 42340 149670
rect 42580 149660 42660 149670
rect 42900 149660 42980 149670
rect 43220 149660 43300 149670
rect 43945 149660 44025 149670
rect 44265 149660 44345 149670
rect 44585 149660 44665 149670
rect 44905 149660 44985 149670
rect 45225 149660 45305 149670
rect 45545 149660 45625 149670
rect 45865 149660 45945 149670
rect 46185 149660 46265 149670
rect 46505 149660 46585 149670
rect 46825 149660 46905 149670
rect 47145 149660 47225 149670
rect 47465 149660 47545 149670
rect 47785 149660 47865 149670
rect 48105 149660 48185 149670
rect 48500 149660 48640 149670
rect 36260 149580 36270 149660
rect 36580 149580 36590 149660
rect 36900 149580 36910 149660
rect 37220 149580 37230 149660
rect 37540 149580 37550 149660
rect 41380 149580 41390 149660
rect 41700 149580 41710 149660
rect 42020 149580 42030 149660
rect 42340 149580 42350 149660
rect 42660 149580 42670 149660
rect 42980 149580 42990 149660
rect 43300 149580 43310 149660
rect 44025 149580 44035 149660
rect 44345 149580 44355 149660
rect 44665 149580 44675 149660
rect 44985 149580 44995 149660
rect 45305 149580 45315 149660
rect 45625 149580 45635 149660
rect 45945 149580 45955 149660
rect 46265 149580 46275 149660
rect 46585 149580 46595 149660
rect 46905 149580 46915 149660
rect 47225 149580 47235 149660
rect 47545 149580 47555 149660
rect 47865 149580 47875 149660
rect 48185 149580 48195 149660
rect 48500 149530 48605 149660
rect 48640 149580 48650 149660
rect 49260 149620 49660 149630
rect 49860 149620 50260 149630
rect 50460 149620 50860 149630
rect 48980 149530 51140 149620
rect 48500 149520 48640 149530
rect 36020 149500 36100 149510
rect 36340 149500 36420 149510
rect 36660 149500 36740 149510
rect 36980 149500 37060 149510
rect 37300 149500 37380 149510
rect 37620 149500 37700 149510
rect 41140 149500 41220 149510
rect 41460 149500 41540 149510
rect 41780 149500 41860 149510
rect 42100 149500 42180 149510
rect 42420 149500 42500 149510
rect 42740 149500 42820 149510
rect 43060 149500 43140 149510
rect 43380 149500 43460 149510
rect 43785 149500 43865 149510
rect 44105 149500 44185 149510
rect 44425 149500 44505 149510
rect 44745 149500 44825 149510
rect 45065 149500 45145 149510
rect 45385 149500 45465 149510
rect 45705 149500 45785 149510
rect 46025 149500 46105 149510
rect 46345 149500 46425 149510
rect 46665 149500 46745 149510
rect 46985 149500 47065 149510
rect 47305 149500 47385 149510
rect 47625 149500 47705 149510
rect 47945 149500 48025 149510
rect 48265 149500 48345 149510
rect 36100 149420 36110 149500
rect 36420 149420 36430 149500
rect 36740 149420 36750 149500
rect 37060 149420 37070 149500
rect 37380 149420 37390 149500
rect 37700 149420 37710 149500
rect 41220 149420 41230 149500
rect 41540 149420 41550 149500
rect 41860 149420 41870 149500
rect 42180 149420 42190 149500
rect 42500 149420 42510 149500
rect 42820 149420 42830 149500
rect 43140 149420 43150 149500
rect 43460 149420 43470 149500
rect 43865 149420 43875 149500
rect 44185 149420 44195 149500
rect 44505 149420 44515 149500
rect 44825 149420 44835 149500
rect 45145 149420 45155 149500
rect 45465 149420 45475 149500
rect 45785 149420 45795 149500
rect 46105 149420 46115 149500
rect 46425 149420 46435 149500
rect 46745 149420 46755 149500
rect 47065 149420 47075 149500
rect 47385 149420 47395 149500
rect 47705 149420 47715 149500
rect 48025 149420 48035 149500
rect 48345 149420 48355 149500
rect 48500 149390 48605 149520
rect 48640 149440 48650 149520
rect 48500 149380 48640 149390
rect 36180 149340 36260 149350
rect 36500 149340 36580 149350
rect 36820 149340 36900 149350
rect 37140 149340 37220 149350
rect 37460 149340 37540 149350
rect 40980 149340 41060 149350
rect 41300 149340 41380 149350
rect 41620 149340 41700 149350
rect 41940 149340 42020 149350
rect 42260 149340 42340 149350
rect 42580 149340 42660 149350
rect 42900 149340 42980 149350
rect 43220 149340 43300 149350
rect 43945 149340 44025 149350
rect 44265 149340 44345 149350
rect 44585 149340 44665 149350
rect 44905 149340 44985 149350
rect 45225 149340 45305 149350
rect 45545 149340 45625 149350
rect 45865 149340 45945 149350
rect 46185 149340 46265 149350
rect 46505 149340 46585 149350
rect 46825 149340 46905 149350
rect 47145 149340 47225 149350
rect 47465 149340 47545 149350
rect 47785 149340 47865 149350
rect 48105 149340 48185 149350
rect 36260 149260 36270 149340
rect 36580 149260 36590 149340
rect 36900 149260 36910 149340
rect 37220 149260 37230 149340
rect 37540 149260 37550 149340
rect 41060 149260 41070 149340
rect 41380 149260 41390 149340
rect 41700 149260 41710 149340
rect 42020 149260 42030 149340
rect 42340 149260 42350 149340
rect 42660 149260 42670 149340
rect 42980 149260 42990 149340
rect 43300 149260 43310 149340
rect 44025 149260 44035 149340
rect 44345 149260 44355 149340
rect 44665 149260 44675 149340
rect 44985 149260 44995 149340
rect 45305 149260 45315 149340
rect 45625 149260 45635 149340
rect 45945 149260 45955 149340
rect 46265 149260 46275 149340
rect 46585 149260 46595 149340
rect 46905 149260 46915 149340
rect 47225 149260 47235 149340
rect 47545 149260 47555 149340
rect 47865 149260 47875 149340
rect 48185 149260 48195 149340
rect 48500 149250 48605 149380
rect 48640 149300 48650 149380
rect 49100 149350 49220 149410
rect 49255 149350 49285 149530
rect 48500 149240 48640 149250
rect 49220 149240 49285 149350
rect 36020 149180 36100 149190
rect 36340 149180 36420 149190
rect 36660 149180 36740 149190
rect 36980 149180 37060 149190
rect 37300 149180 37380 149190
rect 37620 149180 37700 149190
rect 40820 149180 40900 149190
rect 41140 149180 41220 149190
rect 41460 149180 41540 149190
rect 41780 149180 41860 149190
rect 42100 149180 42180 149190
rect 42420 149180 42500 149190
rect 42740 149180 42820 149190
rect 43060 149180 43140 149190
rect 43380 149180 43460 149190
rect 43785 149180 43865 149190
rect 44105 149180 44185 149190
rect 44425 149180 44505 149190
rect 44745 149180 44825 149190
rect 45065 149180 45145 149190
rect 45385 149180 45465 149190
rect 45705 149180 45785 149190
rect 46025 149180 46105 149190
rect 46345 149180 46425 149190
rect 46665 149180 46745 149190
rect 46985 149180 47065 149190
rect 47305 149180 47385 149190
rect 47625 149180 47705 149190
rect 47945 149180 48025 149190
rect 48265 149180 48345 149190
rect 36100 149100 36110 149180
rect 36420 149100 36430 149180
rect 36740 149100 36750 149180
rect 37060 149100 37070 149180
rect 37380 149100 37390 149180
rect 37700 149100 37710 149180
rect 40900 149100 40910 149180
rect 41220 149100 41230 149180
rect 41540 149100 41550 149180
rect 41860 149100 41870 149180
rect 42180 149100 42190 149180
rect 42500 149100 42510 149180
rect 42820 149100 42830 149180
rect 43140 149100 43150 149180
rect 43460 149100 43470 149180
rect 43865 149100 43875 149180
rect 44185 149100 44195 149180
rect 44505 149100 44515 149180
rect 44825 149100 44835 149180
rect 45145 149100 45155 149180
rect 45465 149100 45475 149180
rect 45785 149100 45795 149180
rect 46105 149100 46115 149180
rect 46425 149100 46435 149180
rect 46745 149100 46755 149180
rect 47065 149100 47075 149180
rect 47385 149100 47395 149180
rect 47705 149100 47715 149180
rect 48025 149100 48035 149180
rect 48345 149100 48355 149180
rect 48500 149110 48605 149240
rect 48640 149160 48650 149240
rect 49100 149230 49285 149240
rect 48500 149100 48640 149110
rect 36180 149020 36260 149030
rect 36500 149020 36580 149030
rect 36820 149020 36900 149030
rect 37140 149020 37220 149030
rect 37460 149020 37540 149030
rect 40660 149020 40740 149030
rect 40980 149020 41060 149030
rect 41300 149020 41380 149030
rect 41620 149020 41700 149030
rect 41940 149020 42020 149030
rect 42260 149020 42340 149030
rect 42580 149020 42660 149030
rect 42900 149020 42980 149030
rect 43220 149020 43300 149030
rect 43945 149020 44025 149030
rect 44265 149020 44345 149030
rect 44585 149020 44665 149030
rect 44905 149020 44985 149030
rect 45225 149020 45305 149030
rect 45545 149020 45625 149030
rect 45865 149020 45945 149030
rect 46185 149020 46265 149030
rect 46505 149020 46585 149030
rect 46825 149020 46905 149030
rect 47145 149020 47225 149030
rect 47465 149020 47545 149030
rect 47785 149020 47865 149030
rect 48105 149020 48185 149030
rect 36260 148940 36270 149020
rect 36580 148940 36590 149020
rect 36900 148940 36910 149020
rect 37220 148940 37230 149020
rect 37540 148940 37550 149020
rect 40740 148940 40750 149020
rect 41060 148940 41070 149020
rect 41380 148940 41390 149020
rect 41700 148940 41710 149020
rect 42020 148940 42030 149020
rect 42340 148940 42350 149020
rect 42660 148940 42670 149020
rect 42980 148940 42990 149020
rect 43300 148940 43310 149020
rect 44025 148940 44035 149020
rect 44345 148940 44355 149020
rect 44665 148940 44675 149020
rect 44985 148940 44995 149020
rect 45305 148940 45315 149020
rect 45625 148940 45635 149020
rect 45945 148940 45955 149020
rect 46265 148940 46275 149020
rect 46585 148940 46595 149020
rect 46905 148940 46915 149020
rect 47225 148940 47235 149020
rect 47545 148940 47555 149020
rect 47865 148940 47875 149020
rect 48185 148940 48195 149020
rect 48500 148970 48605 149100
rect 48640 149020 48650 149100
rect 49100 149070 49220 149130
rect 49255 149070 49285 149230
rect 48500 148960 48640 148970
rect 36020 148860 36100 148870
rect 36340 148860 36420 148870
rect 36660 148860 36740 148870
rect 36980 148860 37060 148870
rect 37300 148860 37380 148870
rect 37620 148860 37700 148870
rect 40500 148860 40580 148870
rect 40820 148860 40900 148870
rect 41140 148860 41220 148870
rect 41460 148860 41540 148870
rect 41780 148860 41860 148870
rect 42100 148860 42180 148870
rect 42420 148860 42500 148870
rect 42740 148860 42820 148870
rect 43060 148860 43140 148870
rect 43380 148860 43460 148870
rect 43785 148860 43865 148870
rect 44105 148860 44185 148870
rect 44425 148860 44505 148870
rect 44745 148860 44825 148870
rect 45065 148860 45145 148870
rect 45385 148860 45465 148870
rect 45705 148860 45785 148870
rect 46025 148860 46105 148870
rect 46345 148860 46425 148870
rect 46665 148860 46745 148870
rect 46985 148860 47065 148870
rect 47305 148860 47385 148870
rect 47625 148860 47705 148870
rect 47945 148860 48025 148870
rect 48265 148860 48345 148870
rect 36100 148780 36110 148860
rect 36420 148780 36430 148860
rect 36740 148780 36750 148860
rect 37060 148780 37070 148860
rect 37380 148780 37390 148860
rect 37700 148780 37710 148860
rect 40580 148780 40590 148860
rect 40900 148780 40910 148860
rect 41220 148780 41230 148860
rect 41540 148780 41550 148860
rect 41860 148780 41870 148860
rect 42180 148780 42190 148860
rect 42500 148780 42510 148860
rect 42820 148780 42830 148860
rect 43140 148780 43150 148860
rect 43460 148780 43470 148860
rect 43865 148780 43875 148860
rect 44185 148780 44195 148860
rect 44505 148780 44515 148860
rect 44825 148780 44835 148860
rect 45145 148780 45155 148860
rect 45465 148780 45475 148860
rect 45785 148780 45795 148860
rect 46105 148780 46115 148860
rect 46425 148780 46435 148860
rect 46745 148780 46755 148860
rect 47065 148780 47075 148860
rect 47385 148780 47395 148860
rect 47705 148780 47715 148860
rect 48025 148780 48035 148860
rect 48345 148780 48355 148860
rect 48500 148830 48605 148960
rect 48640 148880 48650 148960
rect 49220 148950 49285 149070
rect 49255 148910 49285 148950
rect 49335 148910 49365 149530
rect 49420 149470 49500 149480
rect 49500 149410 49510 149470
rect 49400 149350 49520 149410
rect 49555 149350 49585 149530
rect 49420 149330 49500 149340
rect 49500 149250 49510 149330
rect 49520 149230 49585 149350
rect 49420 149190 49500 149200
rect 49500 149130 49510 149190
rect 49400 149070 49520 149130
rect 49555 149070 49585 149230
rect 49420 149050 49500 149060
rect 49500 148970 49510 149050
rect 49520 148950 49585 149070
rect 49555 148910 49585 148950
rect 49635 148910 49665 149530
rect 49700 149350 49820 149410
rect 49855 149350 49885 149530
rect 49820 149240 49885 149350
rect 49700 149230 49885 149240
rect 49700 149070 49820 149130
rect 49855 149070 49885 149230
rect 49820 148950 49885 149070
rect 49855 148910 49885 148950
rect 49935 148910 49965 149530
rect 50020 149470 50100 149480
rect 50100 149410 50110 149470
rect 50000 149350 50120 149410
rect 50155 149350 50185 149530
rect 50020 149330 50100 149340
rect 50100 149250 50110 149330
rect 50120 149230 50185 149350
rect 50020 149190 50100 149200
rect 50100 149130 50110 149190
rect 50000 149070 50120 149130
rect 50155 149070 50185 149230
rect 50020 149050 50100 149060
rect 50100 148970 50110 149050
rect 50120 148950 50185 149070
rect 50155 148910 50185 148950
rect 50235 148910 50265 149530
rect 50300 149350 50420 149410
rect 50455 149350 50485 149530
rect 50420 149240 50485 149350
rect 50300 149230 50485 149240
rect 50300 149070 50420 149130
rect 50455 149070 50485 149230
rect 50420 148950 50485 149070
rect 50455 148910 50485 148950
rect 50535 148910 50565 149530
rect 50620 149470 50700 149480
rect 50700 149410 50710 149470
rect 50600 149350 50720 149410
rect 50755 149350 50785 149530
rect 50620 149330 50700 149340
rect 50700 149250 50710 149330
rect 50720 149230 50785 149350
rect 50620 149190 50700 149200
rect 50700 149130 50710 149190
rect 50600 149070 50720 149130
rect 50755 149070 50785 149230
rect 50620 149050 50700 149060
rect 50700 148970 50710 149050
rect 50720 148950 50785 149070
rect 50755 148910 50785 148950
rect 50835 148910 50865 149530
rect 50920 149470 51000 149480
rect 51000 149410 51010 149470
rect 50900 149350 51020 149410
rect 51050 149350 51140 149530
rect 51020 149230 51140 149350
rect 50920 149190 51000 149200
rect 51000 149130 51010 149190
rect 50900 149070 51020 149130
rect 51050 149070 51140 149230
rect 51020 148950 51140 149070
rect 51050 148910 51140 148950
rect 49335 148830 49345 148910
rect 49350 148900 49360 148910
rect 49635 148830 49645 148910
rect 49650 148900 49660 148910
rect 49935 148830 49945 148910
rect 50235 148830 50245 148910
rect 50250 148900 50260 148910
rect 50535 148830 50545 148910
rect 50835 148830 50845 148910
rect 50850 148900 50860 148910
rect 48500 148820 48640 148830
rect 36180 148700 36260 148710
rect 36500 148700 36580 148710
rect 36820 148700 36900 148710
rect 37140 148700 37220 148710
rect 37460 148700 37540 148710
rect 40340 148700 40420 148710
rect 40660 148700 40740 148710
rect 40980 148700 41060 148710
rect 41300 148700 41380 148710
rect 41620 148700 41700 148710
rect 41940 148700 42020 148710
rect 36260 148620 36270 148700
rect 36580 148620 36590 148700
rect 36900 148620 36910 148700
rect 37220 148620 37230 148700
rect 37540 148620 37550 148700
rect 40420 148620 40430 148700
rect 40740 148620 40750 148700
rect 41060 148620 41070 148700
rect 41380 148620 41390 148700
rect 41700 148620 41710 148700
rect 42020 148620 42030 148700
rect 48500 148690 48605 148820
rect 48640 148740 48650 148820
rect 49250 148770 49370 148830
rect 49550 148770 49670 148830
rect 49850 148770 49970 148830
rect 50150 148770 50270 148830
rect 50450 148770 50570 148830
rect 50750 148770 50870 148830
rect 60300 148790 60570 149820
rect 60580 149819 60660 149829
rect 60900 149819 60980 149829
rect 61320 149819 61400 149829
rect 61640 149819 61720 149829
rect 62470 149820 62755 149830
rect 73245 149820 74070 149999
rect 75560 149940 75640 149950
rect 75640 149860 75650 149940
rect 75870 149880 75900 149940
rect 75990 149880 76020 149940
rect 76110 149880 76140 149940
rect 76230 149880 76255 149940
rect 60660 149739 60670 149819
rect 60980 149739 60990 149819
rect 61400 149739 61410 149819
rect 61720 149739 61730 149819
rect 62060 149800 62140 149810
rect 62140 149720 62150 149800
rect 60740 149659 60820 149669
rect 61060 149659 61140 149669
rect 61480 149659 61560 149669
rect 61800 149659 61880 149669
rect 62060 149660 62140 149670
rect 60820 149579 60830 149659
rect 61140 149579 61150 149659
rect 61560 149579 61570 149659
rect 61880 149579 61890 149659
rect 62140 149580 62150 149660
rect 62480 149530 62755 149620
rect 62060 149520 62140 149530
rect 60580 149499 60660 149509
rect 60900 149499 60980 149509
rect 61320 149499 61400 149509
rect 61640 149499 61720 149509
rect 60660 149419 60670 149499
rect 60980 149419 60990 149499
rect 61400 149419 61410 149499
rect 61720 149419 61730 149499
rect 62140 149440 62150 149520
rect 62060 149380 62140 149390
rect 60740 149339 60820 149349
rect 61060 149339 61140 149349
rect 61480 149339 61560 149349
rect 61800 149339 61880 149349
rect 60820 149259 60830 149339
rect 61140 149259 61150 149339
rect 61560 149259 61570 149339
rect 61880 149259 61890 149339
rect 62140 149300 62150 149380
rect 62600 149350 62720 149410
rect 62060 149240 62140 149250
rect 62720 149240 62755 149350
rect 60580 149179 60660 149189
rect 60900 149179 60980 149189
rect 61320 149179 61400 149189
rect 61640 149179 61720 149189
rect 60660 149099 60670 149179
rect 60980 149099 60990 149179
rect 61400 149099 61410 149179
rect 61720 149099 61730 149179
rect 62140 149160 62150 149240
rect 62600 149230 62755 149240
rect 62060 149100 62140 149110
rect 60740 149019 60820 149029
rect 61060 149019 61140 149029
rect 61480 149019 61560 149029
rect 61800 149019 61880 149029
rect 62140 149020 62150 149100
rect 62600 149070 62720 149130
rect 60820 148939 60830 149019
rect 61140 148939 61150 149019
rect 61560 148939 61570 149019
rect 61880 148939 61890 149019
rect 62060 148960 62140 148970
rect 62140 148880 62150 148960
rect 62720 148950 62755 149070
rect 60580 148859 60660 148869
rect 60900 148859 60980 148869
rect 61320 148859 61400 148869
rect 61640 148859 61720 148869
rect 49370 148750 49430 148770
rect 49670 148750 49730 148770
rect 49970 148750 50030 148770
rect 50270 148750 50330 148770
rect 50570 148750 50630 148770
rect 49370 148740 49500 148750
rect 49670 148740 49800 148750
rect 49970 148740 50100 148750
rect 50270 148740 50400 148750
rect 50570 148740 50710 148750
rect 48500 148680 48640 148690
rect 36020 148540 36100 148550
rect 36340 148540 36420 148550
rect 36660 148540 36740 148550
rect 36980 148540 37060 148550
rect 37300 148540 37380 148550
rect 37620 148540 37700 148550
rect 40180 148540 40260 148550
rect 40500 148540 40580 148550
rect 40820 148540 40900 148550
rect 41140 148540 41220 148550
rect 41460 148540 41540 148550
rect 41780 148540 41860 148550
rect 36100 148460 36110 148540
rect 36420 148460 36430 148540
rect 36740 148460 36750 148540
rect 37060 148460 37070 148540
rect 37380 148460 37390 148540
rect 37700 148460 37710 148540
rect 40260 148460 40270 148540
rect 40580 148460 40590 148540
rect 40900 148460 40910 148540
rect 41220 148460 41230 148540
rect 41540 148460 41550 148540
rect 41860 148460 41870 148540
rect 36180 148380 36260 148390
rect 36500 148380 36580 148390
rect 36820 148380 36900 148390
rect 37140 148380 37220 148390
rect 37460 148380 37540 148390
rect 40340 148380 40420 148390
rect 40660 148380 40740 148390
rect 40980 148380 41060 148390
rect 41300 148380 41380 148390
rect 41620 148380 41700 148390
rect 36260 148300 36270 148380
rect 36580 148300 36590 148380
rect 36900 148300 36910 148380
rect 37220 148300 37230 148380
rect 37540 148300 37550 148380
rect 40420 148300 40430 148380
rect 40740 148300 40750 148380
rect 41060 148300 41070 148380
rect 41380 148300 41390 148380
rect 41700 148300 41710 148380
rect 48500 148340 48605 148680
rect 48640 148600 48650 148680
rect 49370 148650 49430 148740
rect 49500 148660 49510 148740
rect 49670 148650 49730 148740
rect 49800 148660 49810 148740
rect 49970 148650 50030 148740
rect 50100 148660 50110 148740
rect 50270 148650 50330 148740
rect 50400 148660 50410 148740
rect 50570 148650 50630 148740
rect 50710 148660 50720 148740
rect 50870 148650 50930 148770
rect 49220 148600 50900 148610
rect 52045 148520 60570 148790
rect 60660 148779 60670 148859
rect 60980 148779 60990 148859
rect 61400 148779 61410 148859
rect 61720 148779 61730 148859
rect 62060 148820 62140 148830
rect 62140 148740 62150 148820
rect 62750 148770 62755 148830
rect 73800 148790 74070 149820
rect 74080 149819 74160 149829
rect 74400 149819 74480 149829
rect 74820 149819 74900 149829
rect 75140 149819 75220 149829
rect 75970 149820 76255 149830
rect 86745 149820 87570 149999
rect 89060 149940 89140 149950
rect 89140 149860 89150 149940
rect 89370 149880 89400 149940
rect 89490 149880 89520 149940
rect 89610 149880 89640 149940
rect 89730 149880 89755 149940
rect 74160 149739 74170 149819
rect 74480 149739 74490 149819
rect 74900 149739 74910 149819
rect 75220 149739 75230 149819
rect 75560 149800 75640 149810
rect 75640 149720 75650 149800
rect 74240 149659 74320 149669
rect 74560 149659 74640 149669
rect 74980 149659 75060 149669
rect 75300 149659 75380 149669
rect 75560 149660 75640 149670
rect 74320 149579 74330 149659
rect 74640 149579 74650 149659
rect 75060 149579 75070 149659
rect 75380 149579 75390 149659
rect 75640 149580 75650 149660
rect 75980 149530 76255 149620
rect 75560 149520 75640 149530
rect 74080 149499 74160 149509
rect 74400 149499 74480 149509
rect 74820 149499 74900 149509
rect 75140 149499 75220 149509
rect 74160 149419 74170 149499
rect 74480 149419 74490 149499
rect 74900 149419 74910 149499
rect 75220 149419 75230 149499
rect 75640 149440 75650 149520
rect 75560 149380 75640 149390
rect 74240 149339 74320 149349
rect 74560 149339 74640 149349
rect 74980 149339 75060 149349
rect 75300 149339 75380 149349
rect 74320 149259 74330 149339
rect 74640 149259 74650 149339
rect 75060 149259 75070 149339
rect 75380 149259 75390 149339
rect 75640 149300 75650 149380
rect 76100 149350 76220 149410
rect 75560 149240 75640 149250
rect 76220 149240 76255 149350
rect 74080 149179 74160 149189
rect 74400 149179 74480 149189
rect 74820 149179 74900 149189
rect 75140 149179 75220 149189
rect 74160 149099 74170 149179
rect 74480 149099 74490 149179
rect 74900 149099 74910 149179
rect 75220 149099 75230 149179
rect 75640 149160 75650 149240
rect 76100 149230 76255 149240
rect 75560 149100 75640 149110
rect 74240 149019 74320 149029
rect 74560 149019 74640 149029
rect 74980 149019 75060 149029
rect 75300 149019 75380 149029
rect 75640 149020 75650 149100
rect 76100 149070 76220 149130
rect 74320 148939 74330 149019
rect 74640 148939 74650 149019
rect 75060 148939 75070 149019
rect 75380 148939 75390 149019
rect 75560 148960 75640 148970
rect 75640 148880 75650 148960
rect 76220 148950 76255 149070
rect 74080 148859 74160 148869
rect 74400 148859 74480 148869
rect 74820 148859 74900 148869
rect 75140 148859 75220 148869
rect 62060 148680 62140 148690
rect 62140 148600 62150 148680
rect 62720 148600 62755 148610
rect 73245 148520 74070 148790
rect 74160 148779 74170 148859
rect 74480 148779 74490 148859
rect 74900 148779 74910 148859
rect 75220 148779 75230 148859
rect 75560 148820 75640 148830
rect 75640 148740 75650 148820
rect 76250 148770 76255 148830
rect 87300 148790 87570 149820
rect 87580 149819 87660 149829
rect 87900 149819 87980 149829
rect 88320 149819 88400 149829
rect 88640 149819 88720 149829
rect 89470 149820 89755 149830
rect 100245 149820 101070 149999
rect 116060 149940 116140 149950
rect 116140 149860 116150 149940
rect 116370 149880 116400 149940
rect 116490 149880 116520 149940
rect 116610 149880 116640 149940
rect 116730 149880 116755 149940
rect 87660 149739 87670 149819
rect 87980 149739 87990 149819
rect 88400 149739 88410 149819
rect 88720 149739 88730 149819
rect 89060 149800 89140 149810
rect 89140 149720 89150 149800
rect 87740 149659 87820 149669
rect 88060 149659 88140 149669
rect 88480 149659 88560 149669
rect 88800 149659 88880 149669
rect 89060 149660 89140 149670
rect 87820 149579 87830 149659
rect 88140 149579 88150 149659
rect 88560 149579 88570 149659
rect 88880 149579 88890 149659
rect 89140 149580 89150 149660
rect 89480 149530 89755 149620
rect 89060 149520 89140 149530
rect 87580 149499 87660 149509
rect 87900 149499 87980 149509
rect 88320 149499 88400 149509
rect 88640 149499 88720 149509
rect 87660 149419 87670 149499
rect 87980 149419 87990 149499
rect 88400 149419 88410 149499
rect 88720 149419 88730 149499
rect 89140 149440 89150 149520
rect 89060 149380 89140 149390
rect 87740 149339 87820 149349
rect 88060 149339 88140 149349
rect 88480 149339 88560 149349
rect 88800 149339 88880 149349
rect 87820 149259 87830 149339
rect 88140 149259 88150 149339
rect 88560 149259 88570 149339
rect 88880 149259 88890 149339
rect 89140 149300 89150 149380
rect 89600 149350 89720 149410
rect 89060 149240 89140 149250
rect 89720 149240 89755 149350
rect 87580 149179 87660 149189
rect 87900 149179 87980 149189
rect 88320 149179 88400 149189
rect 88640 149179 88720 149189
rect 87660 149099 87670 149179
rect 87980 149099 87990 149179
rect 88400 149099 88410 149179
rect 88720 149099 88730 149179
rect 89140 149160 89150 149240
rect 89600 149230 89755 149240
rect 89060 149100 89140 149110
rect 87740 149019 87820 149029
rect 88060 149019 88140 149029
rect 88480 149019 88560 149029
rect 88800 149019 88880 149029
rect 89140 149020 89150 149100
rect 89600 149070 89720 149130
rect 87820 148939 87830 149019
rect 88140 148939 88150 149019
rect 88560 148939 88570 149019
rect 88880 148939 88890 149019
rect 89060 148960 89140 148970
rect 89140 148880 89150 148960
rect 89720 148950 89755 149070
rect 87580 148859 87660 148869
rect 87900 148859 87980 148869
rect 88320 148859 88400 148869
rect 88640 148859 88720 148869
rect 75560 148680 75640 148690
rect 75640 148600 75650 148680
rect 76220 148600 76255 148610
rect 86745 148520 87570 148790
rect 87660 148779 87670 148859
rect 87980 148779 87990 148859
rect 88400 148779 88410 148859
rect 88720 148779 88730 148859
rect 89060 148820 89140 148830
rect 89140 148740 89150 148820
rect 89750 148770 89755 148830
rect 100800 148790 101070 149820
rect 101080 149819 101160 149829
rect 101400 149819 101480 149829
rect 101820 149819 101900 149829
rect 102140 149819 102220 149829
rect 114580 149819 114660 149829
rect 114900 149819 114980 149829
rect 115320 149819 115400 149829
rect 115640 149819 115720 149829
rect 116470 149820 116755 149830
rect 127245 149820 128070 149999
rect 129560 149940 129640 149950
rect 129640 149860 129650 149940
rect 129870 149880 129900 149940
rect 129990 149880 130020 149940
rect 130110 149880 130140 149940
rect 130230 149880 130255 149940
rect 140710 149830 141570 150000
rect 152460 149980 152540 149990
rect 152780 149980 152860 149990
rect 153100 149980 153180 149990
rect 153420 149980 153500 149990
rect 153740 149980 153820 149990
rect 154060 149980 154140 149990
rect 154380 149980 154460 149990
rect 154700 149980 154780 149990
rect 155020 149980 155100 149990
rect 155340 149980 155420 149990
rect 155660 149980 155740 149990
rect 155980 149980 156000 149990
rect 152540 149900 152550 149980
rect 152860 149900 152870 149980
rect 153180 149900 153190 149980
rect 153500 149900 153510 149980
rect 153820 149900 153830 149980
rect 154140 149900 154150 149980
rect 154460 149900 154470 149980
rect 154780 149900 154790 149980
rect 155100 149900 155110 149980
rect 155420 149900 155430 149980
rect 155740 149900 155750 149980
rect 101160 149739 101170 149819
rect 101480 149739 101490 149819
rect 101900 149739 101910 149819
rect 102220 149739 102230 149819
rect 114660 149739 114670 149819
rect 114980 149739 114990 149819
rect 115400 149739 115410 149819
rect 115720 149739 115730 149819
rect 116060 149800 116140 149810
rect 116140 149720 116150 149800
rect 101240 149659 101320 149669
rect 101560 149659 101640 149669
rect 101980 149659 102060 149669
rect 102300 149659 102380 149669
rect 114740 149659 114820 149669
rect 115060 149659 115140 149669
rect 115480 149659 115560 149669
rect 115800 149659 115880 149669
rect 116060 149660 116140 149670
rect 101320 149579 101330 149659
rect 101640 149579 101650 149659
rect 102060 149579 102070 149659
rect 102380 149579 102390 149659
rect 114820 149579 114830 149659
rect 115140 149579 115150 149659
rect 115560 149579 115570 149659
rect 115880 149579 115890 149659
rect 116140 149580 116150 149660
rect 116480 149530 116755 149620
rect 116060 149520 116140 149530
rect 101080 149499 101160 149509
rect 101400 149499 101480 149509
rect 101820 149499 101900 149509
rect 102140 149499 102220 149509
rect 114580 149499 114660 149509
rect 114900 149499 114980 149509
rect 115320 149499 115400 149509
rect 115640 149499 115720 149509
rect 101160 149419 101170 149499
rect 101480 149419 101490 149499
rect 101900 149419 101910 149499
rect 102220 149419 102230 149499
rect 114660 149419 114670 149499
rect 114980 149419 114990 149499
rect 115400 149419 115410 149499
rect 115720 149419 115730 149499
rect 116140 149440 116150 149520
rect 116060 149380 116140 149390
rect 101240 149339 101320 149349
rect 101560 149339 101640 149349
rect 101980 149339 102060 149349
rect 102300 149339 102380 149349
rect 114740 149339 114820 149349
rect 115060 149339 115140 149349
rect 115480 149339 115560 149349
rect 115800 149339 115880 149349
rect 101320 149259 101330 149339
rect 101640 149259 101650 149339
rect 102060 149259 102070 149339
rect 102380 149259 102390 149339
rect 114820 149259 114830 149339
rect 115140 149259 115150 149339
rect 115560 149259 115570 149339
rect 115880 149259 115890 149339
rect 116140 149300 116150 149380
rect 116600 149350 116720 149410
rect 116060 149240 116140 149250
rect 116720 149240 116755 149350
rect 101080 149179 101160 149189
rect 101400 149179 101480 149189
rect 101820 149179 101900 149189
rect 102140 149179 102220 149189
rect 114580 149179 114660 149189
rect 114900 149179 114980 149189
rect 115320 149179 115400 149189
rect 115640 149179 115720 149189
rect 101160 149099 101170 149179
rect 101480 149099 101490 149179
rect 101900 149099 101910 149179
rect 102220 149099 102230 149179
rect 114660 149099 114670 149179
rect 114980 149099 114990 149179
rect 115400 149099 115410 149179
rect 115720 149099 115730 149179
rect 116140 149160 116150 149240
rect 116600 149230 116755 149240
rect 116060 149100 116140 149110
rect 101240 149019 101320 149029
rect 101560 149019 101640 149029
rect 101980 149019 102060 149029
rect 102300 149019 102380 149029
rect 114740 149019 114820 149029
rect 115060 149019 115140 149029
rect 115480 149019 115560 149029
rect 115800 149019 115880 149029
rect 116140 149020 116150 149100
rect 116600 149070 116720 149130
rect 101320 148939 101330 149019
rect 101640 148939 101650 149019
rect 102060 148939 102070 149019
rect 102380 148939 102390 149019
rect 114820 148939 114830 149019
rect 115140 148939 115150 149019
rect 115560 148939 115570 149019
rect 115880 148939 115890 149019
rect 116060 148960 116140 148970
rect 116140 148880 116150 148960
rect 116720 148950 116755 149070
rect 101080 148859 101160 148869
rect 101400 148859 101480 148869
rect 101820 148859 101900 148869
rect 102140 148859 102220 148869
rect 114580 148859 114660 148869
rect 114900 148859 114980 148869
rect 115320 148859 115400 148869
rect 115640 148859 115720 148869
rect 89060 148680 89140 148690
rect 89140 148600 89150 148680
rect 89720 148600 89755 148610
rect 100245 148520 101070 148790
rect 101160 148779 101170 148859
rect 101480 148779 101490 148859
rect 101900 148779 101910 148859
rect 102220 148779 102230 148859
rect 114660 148779 114670 148859
rect 114980 148779 114990 148859
rect 115400 148779 115410 148859
rect 115720 148779 115730 148859
rect 116060 148820 116140 148830
rect 116140 148740 116150 148820
rect 116750 148770 116755 148830
rect 127800 148790 128070 149820
rect 128080 149819 128160 149829
rect 128400 149819 128480 149829
rect 128820 149819 128900 149829
rect 129140 149819 129220 149829
rect 129970 149820 130255 149830
rect 140710 149820 141625 149830
rect 141865 149820 141945 149830
rect 142185 149820 142200 149830
rect 145385 149820 145465 149830
rect 145705 149820 145785 149830
rect 146025 149820 146105 149830
rect 146540 149820 146620 149830
rect 146860 149820 146940 149830
rect 147180 149820 147260 149830
rect 147500 149820 147580 149830
rect 147820 149820 147900 149830
rect 148140 149820 148220 149830
rect 148460 149820 148540 149830
rect 152300 149820 152380 149830
rect 152620 149820 152700 149830
rect 152940 149820 153020 149830
rect 153260 149820 153340 149830
rect 153580 149820 153660 149830
rect 153900 149820 153980 149830
rect 154220 149820 154300 149830
rect 154540 149820 154620 149830
rect 154860 149820 154940 149830
rect 155180 149820 155260 149830
rect 155500 149820 155580 149830
rect 155820 149820 155900 149830
rect 128160 149739 128170 149819
rect 128480 149739 128490 149819
rect 128900 149739 128910 149819
rect 129220 149739 129230 149819
rect 129560 149800 129640 149810
rect 129640 149720 129650 149800
rect 128240 149659 128320 149669
rect 128560 149659 128640 149669
rect 128980 149659 129060 149669
rect 129300 149659 129380 149669
rect 129560 149660 129640 149670
rect 128320 149579 128330 149659
rect 128640 149579 128650 149659
rect 129060 149579 129070 149659
rect 129380 149579 129390 149659
rect 129640 149580 129650 149660
rect 129980 149530 130255 149620
rect 129560 149520 129640 149530
rect 128080 149499 128160 149509
rect 128400 149499 128480 149509
rect 128820 149499 128900 149509
rect 129140 149499 129220 149509
rect 128160 149419 128170 149499
rect 128480 149419 128490 149499
rect 128900 149419 128910 149499
rect 129220 149419 129230 149499
rect 129640 149440 129650 149520
rect 141300 149510 141570 149820
rect 141625 149740 141635 149820
rect 141945 149740 141955 149820
rect 145465 149740 145475 149820
rect 145785 149740 145795 149820
rect 146105 149740 146115 149820
rect 146620 149740 146630 149820
rect 146940 149740 146950 149820
rect 147260 149740 147270 149820
rect 147580 149740 147590 149820
rect 147900 149740 147910 149820
rect 148220 149740 148230 149820
rect 148540 149740 148550 149820
rect 152380 149740 152390 149820
rect 152700 149740 152710 149820
rect 153020 149740 153030 149820
rect 153340 149740 153350 149820
rect 153660 149740 153670 149820
rect 153980 149740 153990 149820
rect 154300 149740 154310 149820
rect 154620 149740 154630 149820
rect 154940 149740 154950 149820
rect 155260 149740 155270 149820
rect 155580 149740 155590 149820
rect 155900 149740 155910 149820
rect 141705 149660 141785 149670
rect 142025 149660 142105 149670
rect 145225 149660 145305 149670
rect 145545 149660 145625 149670
rect 145865 149660 145945 149670
rect 146700 149660 146780 149670
rect 147020 149660 147100 149670
rect 147340 149660 147420 149670
rect 147660 149660 147740 149670
rect 147980 149660 148060 149670
rect 148300 149660 148380 149670
rect 148620 149660 148700 149670
rect 152460 149660 152540 149670
rect 152780 149660 152860 149670
rect 153100 149660 153180 149670
rect 153420 149660 153500 149670
rect 153740 149660 153820 149670
rect 154060 149660 154140 149670
rect 154380 149660 154460 149670
rect 154700 149660 154780 149670
rect 155020 149660 155100 149670
rect 155340 149660 155420 149670
rect 155660 149660 155740 149670
rect 155980 149660 156000 149670
rect 141785 149580 141795 149660
rect 142105 149580 142115 149660
rect 145305 149580 145315 149660
rect 145625 149580 145635 149660
rect 145945 149580 145955 149660
rect 146780 149580 146790 149660
rect 147100 149580 147110 149660
rect 147420 149580 147430 149660
rect 147740 149580 147750 149660
rect 148060 149580 148070 149660
rect 148380 149580 148390 149660
rect 148700 149580 148710 149660
rect 152540 149580 152550 149660
rect 152860 149580 152870 149660
rect 153180 149580 153190 149660
rect 153500 149580 153510 149660
rect 153820 149580 153830 149660
rect 154140 149580 154150 149660
rect 154460 149580 154470 149660
rect 154780 149580 154790 149660
rect 155100 149580 155110 149660
rect 155420 149580 155430 149660
rect 155740 149580 155750 149660
rect 141300 149500 141625 149510
rect 141865 149500 141945 149510
rect 142185 149500 142200 149510
rect 145385 149500 145465 149510
rect 145705 149500 145785 149510
rect 146025 149500 146105 149510
rect 146540 149500 146620 149510
rect 146860 149500 146940 149510
rect 147180 149500 147260 149510
rect 147500 149500 147580 149510
rect 147820 149500 147900 149510
rect 148140 149500 148220 149510
rect 148460 149500 148540 149510
rect 148780 149500 148860 149510
rect 152300 149500 152380 149510
rect 152620 149500 152700 149510
rect 152940 149500 153020 149510
rect 153260 149500 153340 149510
rect 153580 149500 153660 149510
rect 153900 149500 153980 149510
rect 154220 149500 154300 149510
rect 154540 149500 154620 149510
rect 154860 149500 154940 149510
rect 155180 149500 155260 149510
rect 155500 149500 155580 149510
rect 155820 149500 155900 149510
rect 129560 149380 129640 149390
rect 128240 149339 128320 149349
rect 128560 149339 128640 149349
rect 128980 149339 129060 149349
rect 129300 149339 129380 149349
rect 128320 149259 128330 149339
rect 128640 149259 128650 149339
rect 129060 149259 129070 149339
rect 129380 149259 129390 149339
rect 129640 149300 129650 149380
rect 130100 149350 130220 149410
rect 129560 149240 129640 149250
rect 130220 149240 130255 149350
rect 128080 149179 128160 149189
rect 128400 149179 128480 149189
rect 128820 149179 128900 149189
rect 129140 149179 129220 149189
rect 128160 149099 128170 149179
rect 128480 149099 128490 149179
rect 128900 149099 128910 149179
rect 129220 149099 129230 149179
rect 129640 149160 129650 149240
rect 130100 149230 130255 149240
rect 141300 149190 141570 149500
rect 141625 149420 141635 149500
rect 141945 149420 141955 149500
rect 145465 149420 145475 149500
rect 145785 149420 145795 149500
rect 146105 149420 146115 149500
rect 146620 149420 146630 149500
rect 146940 149420 146950 149500
rect 147260 149420 147270 149500
rect 147580 149420 147590 149500
rect 147900 149420 147910 149500
rect 148220 149420 148230 149500
rect 148540 149420 148550 149500
rect 148860 149420 148870 149500
rect 152380 149420 152390 149500
rect 152700 149420 152710 149500
rect 153020 149420 153030 149500
rect 153340 149420 153350 149500
rect 153660 149420 153670 149500
rect 153980 149420 153990 149500
rect 154300 149420 154310 149500
rect 154620 149420 154630 149500
rect 154940 149420 154950 149500
rect 155260 149420 155270 149500
rect 155580 149420 155590 149500
rect 155900 149420 155910 149500
rect 141705 149340 141785 149350
rect 142025 149340 142105 149350
rect 145225 149340 145305 149350
rect 145545 149340 145625 149350
rect 145865 149340 145945 149350
rect 146700 149340 146780 149350
rect 147020 149340 147100 149350
rect 147340 149340 147420 149350
rect 147660 149340 147740 149350
rect 147980 149340 148060 149350
rect 148300 149340 148380 149350
rect 148620 149340 148700 149350
rect 148940 149340 149020 149350
rect 152460 149340 152540 149350
rect 152780 149340 152860 149350
rect 153100 149340 153180 149350
rect 153420 149340 153500 149350
rect 153740 149340 153820 149350
rect 154060 149340 154140 149350
rect 154380 149340 154460 149350
rect 154700 149340 154780 149350
rect 155020 149340 155100 149350
rect 155340 149340 155420 149350
rect 155660 149340 155740 149350
rect 155980 149340 156000 149350
rect 141785 149260 141795 149340
rect 142105 149260 142115 149340
rect 145305 149260 145315 149340
rect 145625 149260 145635 149340
rect 145945 149260 145955 149340
rect 146780 149260 146790 149340
rect 147100 149260 147110 149340
rect 147420 149260 147430 149340
rect 147740 149260 147750 149340
rect 148060 149260 148070 149340
rect 148380 149260 148390 149340
rect 148700 149260 148710 149340
rect 149020 149260 149030 149340
rect 152540 149260 152550 149340
rect 152860 149260 152870 149340
rect 153180 149260 153190 149340
rect 153500 149260 153510 149340
rect 153820 149260 153830 149340
rect 154140 149260 154150 149340
rect 154460 149260 154470 149340
rect 154780 149260 154790 149340
rect 155100 149260 155110 149340
rect 155420 149260 155430 149340
rect 155740 149260 155750 149340
rect 141300 149180 141625 149190
rect 141865 149180 141945 149190
rect 142185 149180 142200 149190
rect 145385 149180 145465 149190
rect 145705 149180 145785 149190
rect 146025 149180 146105 149190
rect 146540 149180 146620 149190
rect 146860 149180 146940 149190
rect 147180 149180 147260 149190
rect 147500 149180 147580 149190
rect 147820 149180 147900 149190
rect 148140 149180 148220 149190
rect 148460 149180 148540 149190
rect 148780 149180 148860 149190
rect 149100 149180 149180 149190
rect 152300 149180 152380 149190
rect 152620 149180 152700 149190
rect 152940 149180 153020 149190
rect 153260 149180 153340 149190
rect 153580 149180 153660 149190
rect 153900 149180 153980 149190
rect 154220 149180 154300 149190
rect 154540 149180 154620 149190
rect 154860 149180 154940 149190
rect 155180 149180 155260 149190
rect 155500 149180 155580 149190
rect 155820 149180 155900 149190
rect 129560 149100 129640 149110
rect 128240 149019 128320 149029
rect 128560 149019 128640 149029
rect 128980 149019 129060 149029
rect 129300 149019 129380 149029
rect 129640 149020 129650 149100
rect 130100 149070 130220 149130
rect 128320 148939 128330 149019
rect 128640 148939 128650 149019
rect 129060 148939 129070 149019
rect 129380 148939 129390 149019
rect 129560 148960 129640 148970
rect 129640 148880 129650 148960
rect 130220 148950 130255 149070
rect 141300 148870 141570 149180
rect 141625 149100 141635 149180
rect 141945 149100 141955 149180
rect 145465 149100 145475 149180
rect 145785 149100 145795 149180
rect 146105 149100 146115 149180
rect 146620 149100 146630 149180
rect 146940 149100 146950 149180
rect 147260 149100 147270 149180
rect 147580 149100 147590 149180
rect 147900 149100 147910 149180
rect 148220 149100 148230 149180
rect 148540 149100 148550 149180
rect 148860 149100 148870 149180
rect 149180 149100 149190 149180
rect 152380 149100 152390 149180
rect 152700 149100 152710 149180
rect 153020 149100 153030 149180
rect 153340 149100 153350 149180
rect 153660 149100 153670 149180
rect 153980 149100 153990 149180
rect 154300 149100 154310 149180
rect 154620 149100 154630 149180
rect 154940 149100 154950 149180
rect 155260 149100 155270 149180
rect 155580 149100 155590 149180
rect 155900 149100 155910 149180
rect 141705 149020 141785 149030
rect 142025 149020 142105 149030
rect 145225 149020 145305 149030
rect 145545 149020 145625 149030
rect 145865 149020 145945 149030
rect 146700 149020 146780 149030
rect 147020 149020 147100 149030
rect 147340 149020 147420 149030
rect 147660 149020 147740 149030
rect 147980 149020 148060 149030
rect 148300 149020 148380 149030
rect 148620 149020 148700 149030
rect 148940 149020 149020 149030
rect 149260 149020 149340 149030
rect 152460 149020 152540 149030
rect 152780 149020 152860 149030
rect 153100 149020 153180 149030
rect 153420 149020 153500 149030
rect 153740 149020 153820 149030
rect 154060 149020 154140 149030
rect 154380 149020 154460 149030
rect 154700 149020 154780 149030
rect 155020 149020 155100 149030
rect 155340 149020 155420 149030
rect 155660 149020 155740 149030
rect 155980 149020 156000 149030
rect 141785 148940 141795 149020
rect 142105 148940 142115 149020
rect 145305 148940 145315 149020
rect 145625 148940 145635 149020
rect 145945 148940 145955 149020
rect 146780 148940 146790 149020
rect 147100 148940 147110 149020
rect 147420 148940 147430 149020
rect 147740 148940 147750 149020
rect 148060 148940 148070 149020
rect 148380 148940 148390 149020
rect 148700 148940 148710 149020
rect 149020 148940 149030 149020
rect 149340 148940 149350 149020
rect 152540 148940 152550 149020
rect 152860 148940 152870 149020
rect 153180 148940 153190 149020
rect 153500 148940 153510 149020
rect 153820 148940 153830 149020
rect 154140 148940 154150 149020
rect 154460 148940 154470 149020
rect 154780 148940 154790 149020
rect 155100 148940 155110 149020
rect 155420 148940 155430 149020
rect 155740 148940 155750 149020
rect 128080 148859 128160 148869
rect 128400 148859 128480 148869
rect 128820 148859 128900 148869
rect 129140 148859 129220 148869
rect 141300 148860 141625 148870
rect 141865 148860 141945 148870
rect 142185 148860 142200 148870
rect 145385 148860 145465 148870
rect 145705 148860 145785 148870
rect 146025 148860 146105 148870
rect 146540 148860 146620 148870
rect 146860 148860 146940 148870
rect 147180 148860 147260 148870
rect 147500 148860 147580 148870
rect 147820 148860 147900 148870
rect 148140 148860 148220 148870
rect 148460 148860 148540 148870
rect 148780 148860 148860 148870
rect 149100 148860 149180 148870
rect 149420 148860 149500 148870
rect 152300 148860 152380 148870
rect 152620 148860 152700 148870
rect 152940 148860 153020 148870
rect 153260 148860 153340 148870
rect 153580 148860 153660 148870
rect 153900 148860 153980 148870
rect 154220 148860 154300 148870
rect 154540 148860 154620 148870
rect 154860 148860 154940 148870
rect 155180 148860 155260 148870
rect 155500 148860 155580 148870
rect 155820 148860 155900 148870
rect 116060 148680 116140 148690
rect 116140 148600 116150 148680
rect 116720 148600 116755 148610
rect 127245 148520 128070 148790
rect 128160 148779 128170 148859
rect 128480 148779 128490 148859
rect 128900 148779 128910 148859
rect 129220 148779 129230 148859
rect 129560 148820 129640 148830
rect 129640 148740 129650 148820
rect 130250 148770 130255 148830
rect 141300 148790 141570 148860
rect 129560 148680 129640 148690
rect 129640 148600 129650 148680
rect 130220 148600 130255 148610
rect 140710 148520 141570 148790
rect 141625 148780 141635 148860
rect 141945 148780 141955 148860
rect 145465 148780 145475 148860
rect 145785 148780 145795 148860
rect 146105 148780 146115 148860
rect 146620 148780 146630 148860
rect 146940 148780 146950 148860
rect 147260 148780 147270 148860
rect 147580 148780 147590 148860
rect 147900 148780 147910 148860
rect 148220 148780 148230 148860
rect 148540 148780 148550 148860
rect 148860 148780 148870 148860
rect 149180 148780 149190 148860
rect 149500 148780 149510 148860
rect 152380 148780 152390 148860
rect 152700 148780 152710 148860
rect 153020 148780 153030 148860
rect 153340 148780 153350 148860
rect 153660 148780 153670 148860
rect 153980 148780 153990 148860
rect 154300 148780 154310 148860
rect 154620 148780 154630 148860
rect 154940 148780 154950 148860
rect 155260 148780 155270 148860
rect 155580 148780 155590 148860
rect 155900 148780 155910 148860
rect 147980 148700 148060 148710
rect 148300 148700 148380 148710
rect 148620 148700 148700 148710
rect 148940 148700 149020 148710
rect 149260 148700 149340 148710
rect 149580 148700 149660 148710
rect 152460 148700 152540 148710
rect 152780 148700 152860 148710
rect 153100 148700 153180 148710
rect 153420 148700 153500 148710
rect 153740 148700 153820 148710
rect 154060 148700 154140 148710
rect 154380 148700 154460 148710
rect 154700 148700 154780 148710
rect 155020 148700 155100 148710
rect 155340 148700 155420 148710
rect 155660 148700 155740 148710
rect 155980 148700 156000 148710
rect 148060 148620 148070 148700
rect 148380 148620 148390 148700
rect 148700 148620 148710 148700
rect 149020 148620 149030 148700
rect 149340 148620 149350 148700
rect 149660 148620 149670 148700
rect 152540 148620 152550 148700
rect 152860 148620 152870 148700
rect 153180 148620 153190 148700
rect 153500 148620 153510 148700
rect 153820 148620 153830 148700
rect 154140 148620 154150 148700
rect 154460 148620 154470 148700
rect 154780 148620 154790 148700
rect 155100 148620 155110 148700
rect 155420 148620 155430 148700
rect 155740 148620 155750 148700
rect 148140 148540 148220 148550
rect 148460 148540 148540 148550
rect 148780 148540 148860 148550
rect 149100 148540 149180 148550
rect 149420 148540 149500 148550
rect 149740 148540 149820 148550
rect 152300 148540 152380 148550
rect 152620 148540 152700 148550
rect 152940 148540 153020 148550
rect 153260 148540 153340 148550
rect 153580 148540 153660 148550
rect 153900 148540 153980 148550
rect 154220 148540 154300 148550
rect 154540 148540 154620 148550
rect 154860 148540 154940 148550
rect 155180 148540 155260 148550
rect 155500 148540 155580 148550
rect 155820 148540 155900 148550
rect 148220 148460 148230 148540
rect 148540 148460 148550 148540
rect 148860 148460 148870 148540
rect 149180 148460 149190 148540
rect 149500 148460 149510 148540
rect 149820 148460 149830 148540
rect 152380 148460 152390 148540
rect 152700 148460 152710 148540
rect 153020 148460 153030 148540
rect 153340 148460 153350 148540
rect 153660 148460 153670 148540
rect 153980 148460 153990 148540
rect 154300 148460 154310 148540
rect 154620 148460 154630 148540
rect 154940 148460 154950 148540
rect 155260 148460 155270 148540
rect 155580 148460 155590 148540
rect 155900 148460 155910 148540
rect 48870 148400 48900 148460
rect 48990 148400 49020 148460
rect 49110 148400 49140 148460
rect 49230 148400 49260 148460
rect 49350 148400 49380 148460
rect 49470 148400 49500 148460
rect 49590 148400 49620 148460
rect 49710 148400 49740 148460
rect 49830 148400 49860 148460
rect 49950 148400 49980 148460
rect 50070 148400 50100 148460
rect 50190 148400 50220 148460
rect 50310 148400 50340 148460
rect 50430 148400 50460 148460
rect 50550 148400 50580 148460
rect 50670 148400 50700 148460
rect 50790 148400 50820 148460
rect 50910 148400 50940 148460
rect 51030 148400 51060 148460
rect 51150 148400 51180 148460
rect 51270 148400 51300 148460
rect 51390 148400 51420 148460
rect 51510 148400 51540 148460
rect 51630 148400 51660 148460
rect 51750 148400 51780 148460
rect 51870 148400 51900 148460
rect 51990 148400 52020 148460
rect 52110 148400 52140 148460
rect 52230 148400 52260 148460
rect 52350 148400 52380 148460
rect 52470 148400 52500 148460
rect 52590 148400 52620 148460
rect 52710 148400 52740 148460
rect 52830 148400 52860 148460
rect 52950 148400 52980 148460
rect 53070 148400 53100 148460
rect 53190 148400 53220 148460
rect 53310 148400 53340 148460
rect 53430 148400 53460 148460
rect 53550 148400 53580 148460
rect 53670 148400 53700 148460
rect 53790 148400 53820 148460
rect 53910 148400 53940 148460
rect 54030 148400 54060 148460
rect 54150 148400 54180 148460
rect 54270 148400 54300 148460
rect 54390 148400 54420 148460
rect 54510 148400 54540 148460
rect 54630 148400 54660 148460
rect 54750 148400 54780 148460
rect 54870 148400 54900 148460
rect 54990 148400 55020 148460
rect 55110 148400 55140 148460
rect 55230 148400 55260 148460
rect 55350 148400 55380 148460
rect 55470 148400 55500 148460
rect 55590 148400 55620 148460
rect 55710 148400 55740 148460
rect 55830 148400 55860 148460
rect 55950 148400 55980 148460
rect 56070 148400 56100 148460
rect 56190 148400 56220 148460
rect 56310 148400 56340 148460
rect 56430 148400 56460 148460
rect 56550 148400 56580 148460
rect 56670 148400 56700 148460
rect 56790 148400 56820 148460
rect 56910 148400 56940 148460
rect 57030 148400 57060 148460
rect 57150 148400 57180 148460
rect 57270 148400 57300 148460
rect 57390 148400 57420 148460
rect 57510 148400 57540 148460
rect 57630 148400 57660 148460
rect 57750 148400 57780 148460
rect 57870 148400 57900 148460
rect 57990 148400 58020 148460
rect 58110 148400 58140 148460
rect 58230 148400 58260 148460
rect 58350 148400 58380 148460
rect 58470 148400 58500 148460
rect 58590 148400 58620 148460
rect 58710 148400 58740 148460
rect 58830 148400 58860 148460
rect 58950 148400 58980 148460
rect 59070 148400 59100 148460
rect 59190 148400 59220 148460
rect 59310 148400 59340 148460
rect 59430 148400 59460 148460
rect 59550 148400 59580 148460
rect 59670 148400 59700 148460
rect 59790 148400 59820 148460
rect 59910 148400 59940 148460
rect 60030 148400 60060 148460
rect 60150 148400 60180 148460
rect 62370 148400 62400 148460
rect 62490 148400 62520 148460
rect 62610 148400 62640 148460
rect 62730 148400 62755 148460
rect 73290 148400 73320 148460
rect 73410 148400 73440 148460
rect 73530 148400 73560 148460
rect 73650 148400 73680 148460
rect 75870 148400 75900 148460
rect 75990 148400 76020 148460
rect 76110 148400 76140 148460
rect 76230 148400 76255 148460
rect 86790 148400 86820 148460
rect 86910 148400 86940 148460
rect 87030 148400 87060 148460
rect 87150 148400 87180 148460
rect 89370 148400 89400 148460
rect 89490 148400 89520 148460
rect 89610 148400 89640 148460
rect 89730 148400 89755 148460
rect 100290 148400 100320 148460
rect 100410 148400 100440 148460
rect 100530 148400 100560 148460
rect 100650 148400 100680 148460
rect 116370 148400 116400 148460
rect 116490 148400 116520 148460
rect 116610 148400 116640 148460
rect 116730 148400 116755 148460
rect 127290 148400 127320 148460
rect 127410 148400 127440 148460
rect 127530 148400 127560 148460
rect 127650 148400 127680 148460
rect 129870 148400 129900 148460
rect 129990 148400 130020 148460
rect 130110 148400 130140 148460
rect 130230 148400 130255 148460
rect 140790 148400 140820 148460
rect 140910 148400 140940 148460
rect 141030 148400 141060 148460
rect 141150 148400 141180 148460
rect 148300 148380 148380 148390
rect 148620 148380 148700 148390
rect 148940 148380 149020 148390
rect 149260 148380 149340 148390
rect 149580 148380 149660 148390
rect 152460 148380 152540 148390
rect 152780 148380 152860 148390
rect 153100 148380 153180 148390
rect 153420 148380 153500 148390
rect 153740 148380 153820 148390
rect 154060 148380 154140 148390
rect 154380 148380 154460 148390
rect 154700 148380 154780 148390
rect 155020 148380 155100 148390
rect 155340 148380 155420 148390
rect 155660 148380 155740 148390
rect 155980 148380 156000 148390
rect 148380 148300 148390 148380
rect 148700 148300 148710 148380
rect 149020 148300 149030 148380
rect 149340 148300 149350 148380
rect 149660 148300 149670 148380
rect 152540 148300 152550 148380
rect 152860 148300 152870 148380
rect 153180 148300 153190 148380
rect 153500 148300 153510 148380
rect 153820 148300 153830 148380
rect 154140 148300 154150 148380
rect 154460 148300 154470 148380
rect 154780 148300 154790 148380
rect 155100 148300 155110 148380
rect 155420 148300 155430 148380
rect 155740 148300 155750 148380
rect 36020 148220 36100 148230
rect 36340 148220 36420 148230
rect 36660 148220 36740 148230
rect 36980 148220 37060 148230
rect 37300 148220 37380 148230
rect 37620 148220 37700 148230
rect 40180 148220 40260 148230
rect 40500 148220 40580 148230
rect 40820 148220 40900 148230
rect 41140 148220 41220 148230
rect 41460 148220 41540 148230
rect 148460 148220 148540 148230
rect 148780 148220 148860 148230
rect 149100 148220 149180 148230
rect 149420 148220 149500 148230
rect 149740 148220 149820 148230
rect 152300 148220 152380 148230
rect 152620 148220 152700 148230
rect 152940 148220 153020 148230
rect 153260 148220 153340 148230
rect 153580 148220 153660 148230
rect 153900 148220 153980 148230
rect 154220 148220 154300 148230
rect 154540 148220 154620 148230
rect 154860 148220 154940 148230
rect 155180 148220 155260 148230
rect 155500 148220 155580 148230
rect 155820 148220 155900 148230
rect 36100 148140 36110 148220
rect 36420 148140 36430 148220
rect 36740 148140 36750 148220
rect 37060 148140 37070 148220
rect 37380 148140 37390 148220
rect 37700 148140 37710 148220
rect 40260 148140 40270 148220
rect 40580 148140 40590 148220
rect 40900 148140 40910 148220
rect 41220 148140 41230 148220
rect 41540 148140 41550 148220
rect 148540 148140 148550 148220
rect 148860 148140 148870 148220
rect 149180 148140 149190 148220
rect 149500 148140 149510 148220
rect 149820 148140 149830 148220
rect 152380 148140 152390 148220
rect 152700 148140 152710 148220
rect 153020 148140 153030 148220
rect 153340 148140 153350 148220
rect 153660 148140 153670 148220
rect 153980 148140 153990 148220
rect 154300 148140 154310 148220
rect 154620 148140 154630 148220
rect 154940 148140 154950 148220
rect 155260 148140 155270 148220
rect 155580 148140 155590 148220
rect 155900 148140 155910 148220
rect 36180 148060 36260 148070
rect 36500 148060 36580 148070
rect 36820 148060 36900 148070
rect 37140 148060 37220 148070
rect 37460 148060 37540 148070
rect 40340 148060 40420 148070
rect 40660 148060 40740 148070
rect 40980 148060 41060 148070
rect 41300 148060 41380 148070
rect 148620 148060 148700 148070
rect 148940 148060 149020 148070
rect 149260 148060 149340 148070
rect 149580 148060 149660 148070
rect 152460 148060 152540 148070
rect 152780 148060 152860 148070
rect 153100 148060 153180 148070
rect 153420 148060 153500 148070
rect 153740 148060 153820 148070
rect 154060 148060 154140 148070
rect 154380 148060 154460 148070
rect 154700 148060 154780 148070
rect 155020 148060 155100 148070
rect 155340 148060 155420 148070
rect 155660 148060 155740 148070
rect 155980 148060 156000 148070
rect 36260 147980 36270 148060
rect 36580 147980 36590 148060
rect 36900 147980 36910 148060
rect 37220 147980 37230 148060
rect 37540 147980 37550 148060
rect 40420 147980 40430 148060
rect 40740 147980 40750 148060
rect 41060 147980 41070 148060
rect 41380 147980 41390 148060
rect 148700 147980 148710 148060
rect 149020 147980 149030 148060
rect 149340 147980 149350 148060
rect 149660 147980 149670 148060
rect 152540 147980 152550 148060
rect 152860 147980 152870 148060
rect 153180 147980 153190 148060
rect 153500 147980 153510 148060
rect 153820 147980 153830 148060
rect 154140 147980 154150 148060
rect 154460 147980 154470 148060
rect 154780 147980 154790 148060
rect 155100 147980 155110 148060
rect 155420 147980 155430 148060
rect 155740 147980 155750 148060
rect 36020 147900 36100 147910
rect 36340 147900 36420 147910
rect 36660 147900 36740 147910
rect 36980 147900 37060 147910
rect 37300 147900 37380 147910
rect 37620 147900 37700 147910
rect 40180 147900 40260 147910
rect 40500 147900 40580 147910
rect 40820 147900 40900 147910
rect 41140 147900 41220 147910
rect 148780 147900 148860 147910
rect 149100 147900 149180 147910
rect 149420 147900 149500 147910
rect 149740 147900 149820 147910
rect 152300 147900 152380 147910
rect 152620 147900 152700 147910
rect 152940 147900 153020 147910
rect 153260 147900 153340 147910
rect 153580 147900 153660 147910
rect 153900 147900 153980 147910
rect 154220 147900 154300 147910
rect 154540 147900 154620 147910
rect 154860 147900 154940 147910
rect 155180 147900 155260 147910
rect 155500 147900 155580 147910
rect 155820 147900 155900 147910
rect 36100 147820 36110 147900
rect 36420 147820 36430 147900
rect 36740 147820 36750 147900
rect 37060 147820 37070 147900
rect 37380 147820 37390 147900
rect 37700 147820 37710 147900
rect 40260 147820 40270 147900
rect 40580 147820 40590 147900
rect 40900 147820 40910 147900
rect 41220 147820 41230 147900
rect 148860 147820 148870 147900
rect 149180 147820 149190 147900
rect 149500 147820 149510 147900
rect 149820 147820 149830 147900
rect 152380 147820 152390 147900
rect 152700 147820 152710 147900
rect 153020 147820 153030 147900
rect 153340 147820 153350 147900
rect 153660 147820 153670 147900
rect 153980 147820 153990 147900
rect 154300 147820 154310 147900
rect 154620 147820 154630 147900
rect 154940 147820 154950 147900
rect 155260 147820 155270 147900
rect 155580 147820 155590 147900
rect 155900 147820 155910 147900
rect 36180 147740 36260 147750
rect 36500 147740 36580 147750
rect 36820 147740 36900 147750
rect 37140 147740 37220 147750
rect 37460 147740 37540 147750
rect 40340 147740 40420 147750
rect 40660 147740 40740 147750
rect 40980 147740 41060 147750
rect 148940 147740 149020 147750
rect 149260 147740 149340 147750
rect 149580 147740 149660 147750
rect 152460 147740 152540 147750
rect 152780 147740 152860 147750
rect 153100 147740 153180 147750
rect 153420 147740 153500 147750
rect 153740 147740 153820 147750
rect 154060 147740 154140 147750
rect 154380 147740 154460 147750
rect 154700 147740 154780 147750
rect 155020 147740 155100 147750
rect 155340 147740 155420 147750
rect 155660 147740 155740 147750
rect 155980 147740 156000 147750
rect 36260 147660 36270 147740
rect 36580 147660 36590 147740
rect 36900 147660 36910 147740
rect 37220 147660 37230 147740
rect 37540 147660 37550 147740
rect 40420 147660 40430 147740
rect 40740 147660 40750 147740
rect 41060 147660 41070 147740
rect 48500 147650 48605 147700
rect 149020 147660 149030 147740
rect 149340 147660 149350 147740
rect 149660 147660 149670 147740
rect 152540 147660 152550 147740
rect 152860 147660 152870 147740
rect 153180 147660 153190 147740
rect 153500 147660 153510 147740
rect 153820 147660 153830 147740
rect 154140 147660 154150 147740
rect 154460 147660 154470 147740
rect 154780 147660 154790 147740
rect 155100 147660 155110 147740
rect 155420 147660 155430 147740
rect 155740 147660 155750 147740
rect 48500 147640 48640 147650
rect 60360 147640 60440 147650
rect 62060 147640 62140 147650
rect 73860 147640 73940 147650
rect 75560 147640 75640 147650
rect 87360 147640 87440 147650
rect 89060 147640 89140 147650
rect 100860 147640 100940 147650
rect 116060 147640 116140 147650
rect 127860 147640 127940 147650
rect 129560 147640 129640 147650
rect 141360 147640 141440 147650
rect 36020 147580 36100 147590
rect 36340 147580 36420 147590
rect 36660 147580 36740 147590
rect 36980 147580 37060 147590
rect 37300 147580 37380 147590
rect 37620 147580 37700 147590
rect 40180 147580 40260 147590
rect 40500 147580 40580 147590
rect 40820 147580 40900 147590
rect 41140 147580 41220 147590
rect 43060 147580 43140 147590
rect 43380 147580 43460 147590
rect 43700 147580 43780 147590
rect 36100 147500 36110 147580
rect 36420 147500 36430 147580
rect 36740 147500 36750 147580
rect 37060 147500 37070 147580
rect 37380 147500 37390 147580
rect 37700 147500 37710 147580
rect 40260 147500 40270 147580
rect 40580 147500 40590 147580
rect 40900 147500 40910 147580
rect 41220 147500 41230 147580
rect 43140 147500 43150 147580
rect 43460 147500 43470 147580
rect 43780 147530 43790 147580
rect 43700 147500 43790 147530
rect 48500 147510 48605 147640
rect 48640 147560 48650 147640
rect 48870 147580 48900 147640
rect 48990 147580 49020 147640
rect 49110 147580 49140 147640
rect 49230 147580 49260 147640
rect 49350 147580 49380 147640
rect 49470 147580 49500 147640
rect 49590 147580 49620 147640
rect 49710 147580 49740 147640
rect 49830 147580 49860 147640
rect 49950 147580 49980 147640
rect 50070 147580 50100 147640
rect 50190 147580 50220 147640
rect 50310 147580 50340 147640
rect 50430 147580 50460 147640
rect 50550 147580 50580 147640
rect 50670 147580 50700 147640
rect 50790 147580 50820 147640
rect 50910 147580 50940 147640
rect 51030 147580 51060 147640
rect 51150 147580 51180 147640
rect 51270 147580 51300 147640
rect 51390 147580 51420 147640
rect 51510 147580 51540 147640
rect 51630 147580 51660 147640
rect 51750 147580 51780 147640
rect 51870 147580 51900 147640
rect 51990 147580 52020 147640
rect 52110 147580 52140 147640
rect 52230 147580 52260 147640
rect 52350 147580 52380 147640
rect 52470 147580 52500 147640
rect 52590 147580 52620 147640
rect 52710 147580 52740 147640
rect 52830 147580 52860 147640
rect 52950 147580 52980 147640
rect 53070 147580 53100 147640
rect 53190 147580 53220 147640
rect 53310 147580 53340 147640
rect 53430 147580 53460 147640
rect 53550 147580 53580 147640
rect 53670 147580 53700 147640
rect 53790 147580 53820 147640
rect 53910 147580 53940 147640
rect 54030 147580 54060 147640
rect 54150 147580 54180 147640
rect 54270 147580 54300 147640
rect 54390 147580 54420 147640
rect 54510 147580 54540 147640
rect 54630 147580 54660 147640
rect 54750 147580 54780 147640
rect 54870 147580 54900 147640
rect 54990 147580 55020 147640
rect 55110 147580 55140 147640
rect 55230 147580 55260 147640
rect 55350 147580 55380 147640
rect 55470 147580 55500 147640
rect 55590 147580 55620 147640
rect 55710 147580 55740 147640
rect 55830 147580 55860 147640
rect 55950 147580 55980 147640
rect 56070 147580 56100 147640
rect 56190 147580 56220 147640
rect 56310 147580 56340 147640
rect 56430 147580 56460 147640
rect 56550 147580 56580 147640
rect 56670 147580 56700 147640
rect 56790 147580 56820 147640
rect 56910 147580 56940 147640
rect 57030 147580 57060 147640
rect 57150 147580 57180 147640
rect 57270 147580 57300 147640
rect 57390 147580 57420 147640
rect 57510 147580 57540 147640
rect 57630 147580 57660 147640
rect 57750 147580 57780 147640
rect 57870 147580 57900 147640
rect 57990 147580 58020 147640
rect 58110 147580 58140 147640
rect 58230 147580 58260 147640
rect 58350 147580 58380 147640
rect 58470 147580 58500 147640
rect 58590 147580 58620 147640
rect 58710 147580 58740 147640
rect 58830 147580 58860 147640
rect 58950 147580 58980 147640
rect 59070 147580 59100 147640
rect 59190 147580 59220 147640
rect 59310 147580 59340 147640
rect 59430 147580 59460 147640
rect 59550 147580 59580 147640
rect 59670 147580 59700 147640
rect 59790 147580 59820 147640
rect 59910 147580 59940 147640
rect 60030 147580 60060 147640
rect 60150 147580 60180 147640
rect 60440 147560 60450 147640
rect 62140 147560 62150 147640
rect 62370 147580 62400 147640
rect 62490 147580 62520 147640
rect 62610 147580 62640 147640
rect 62730 147580 62755 147640
rect 73290 147580 73320 147640
rect 73410 147580 73440 147640
rect 73530 147580 73560 147640
rect 73650 147580 73680 147640
rect 73940 147560 73950 147640
rect 75640 147560 75650 147640
rect 75870 147580 75900 147640
rect 75990 147580 76020 147640
rect 76110 147580 76140 147640
rect 76230 147580 76255 147640
rect 86790 147580 86820 147640
rect 86910 147580 86940 147640
rect 87030 147580 87060 147640
rect 87150 147580 87180 147640
rect 87440 147560 87450 147640
rect 89140 147560 89150 147640
rect 89370 147580 89400 147640
rect 89490 147580 89520 147640
rect 89610 147580 89640 147640
rect 89730 147580 89755 147640
rect 100290 147580 100320 147640
rect 100410 147580 100440 147640
rect 100530 147580 100560 147640
rect 100650 147580 100680 147640
rect 100940 147560 100950 147640
rect 116140 147560 116150 147640
rect 116370 147580 116400 147640
rect 116490 147580 116520 147640
rect 116610 147580 116640 147640
rect 116730 147580 116755 147640
rect 127290 147580 127320 147640
rect 127410 147580 127440 147640
rect 127530 147580 127560 147640
rect 127650 147580 127680 147640
rect 127940 147560 127950 147640
rect 129640 147560 129650 147640
rect 129870 147580 129900 147640
rect 129990 147580 130020 147640
rect 130110 147580 130140 147640
rect 130230 147580 130255 147640
rect 140790 147580 140820 147640
rect 140910 147580 140940 147640
rect 141030 147580 141060 147640
rect 141150 147580 141180 147640
rect 141440 147560 141450 147640
rect 146220 147580 146300 147590
rect 146540 147580 146620 147590
rect 146860 147580 146940 147590
rect 148780 147580 148860 147590
rect 149100 147580 149180 147590
rect 149420 147580 149500 147590
rect 149740 147580 149820 147590
rect 152300 147580 152380 147590
rect 152620 147580 152700 147590
rect 152940 147580 153020 147590
rect 153260 147580 153340 147590
rect 153580 147580 153660 147590
rect 153900 147580 153980 147590
rect 154220 147580 154300 147590
rect 154540 147580 154620 147590
rect 154860 147580 154940 147590
rect 155180 147580 155260 147590
rect 155500 147580 155580 147590
rect 155820 147580 155900 147590
rect 49430 147520 50970 147530
rect 48500 147500 48640 147510
rect 60360 147500 60440 147510
rect 62060 147500 62140 147510
rect 73860 147500 73940 147510
rect 75560 147500 75640 147510
rect 87360 147500 87440 147510
rect 89060 147500 89140 147510
rect 100860 147500 100940 147510
rect 116060 147500 116140 147510
rect 127860 147500 127940 147510
rect 129560 147500 129640 147510
rect 141360 147500 141440 147510
rect 146300 147500 146310 147580
rect 146620 147500 146630 147580
rect 146940 147500 146950 147580
rect 148860 147500 148870 147580
rect 149180 147500 149190 147580
rect 149500 147500 149510 147580
rect 149820 147500 149830 147580
rect 152380 147500 152390 147580
rect 152700 147500 152710 147580
rect 153020 147500 153030 147580
rect 153340 147500 153350 147580
rect 153660 147500 153670 147580
rect 153980 147500 153990 147580
rect 154300 147500 154310 147580
rect 154620 147500 154630 147580
rect 154940 147500 154950 147580
rect 155260 147500 155270 147580
rect 155580 147500 155590 147580
rect 155900 147500 155910 147580
rect 43785 147440 43865 147450
rect 44105 147440 44185 147450
rect 44425 147440 44505 147450
rect 44745 147440 44825 147450
rect 45065 147440 45145 147450
rect 45385 147440 45465 147450
rect 45705 147440 45785 147450
rect 46025 147440 46105 147450
rect 46345 147440 46425 147450
rect 46665 147440 46745 147450
rect 46985 147440 47065 147450
rect 47305 147440 47385 147450
rect 47625 147440 47705 147450
rect 47945 147440 48025 147450
rect 48265 147440 48345 147450
rect 36180 147420 36260 147430
rect 36500 147420 36580 147430
rect 36820 147420 36900 147430
rect 37140 147420 37220 147430
rect 37460 147420 37540 147430
rect 40340 147420 40420 147430
rect 40660 147420 40740 147430
rect 40980 147420 41060 147430
rect 42900 147420 42980 147430
rect 43220 147420 43300 147430
rect 43540 147420 43620 147430
rect 36260 147340 36270 147420
rect 36580 147340 36590 147420
rect 36900 147340 36910 147420
rect 37220 147340 37230 147420
rect 37540 147340 37550 147420
rect 40420 147340 40430 147420
rect 40740 147340 40750 147420
rect 41060 147340 41070 147420
rect 42980 147340 42990 147420
rect 43300 147340 43310 147420
rect 43620 147340 43630 147420
rect 43865 147360 43875 147440
rect 44185 147360 44195 147440
rect 44505 147360 44515 147440
rect 44825 147360 44835 147440
rect 45145 147360 45155 147440
rect 45465 147360 45475 147440
rect 45785 147360 45795 147440
rect 46105 147360 46115 147440
rect 46425 147360 46435 147440
rect 46745 147360 46755 147440
rect 47065 147360 47075 147440
rect 47385 147360 47395 147440
rect 47705 147360 47715 147440
rect 48025 147360 48035 147440
rect 48345 147360 48355 147440
rect 48500 147370 48605 147500
rect 48640 147420 48650 147500
rect 49550 147390 49670 147450
rect 50140 147390 50260 147450
rect 50730 147390 50850 147450
rect 60440 147420 60450 147500
rect 60580 147439 60660 147449
rect 60900 147439 60980 147449
rect 61320 147439 61400 147449
rect 61640 147439 61720 147449
rect 48500 147360 48640 147370
rect 43945 147280 44025 147290
rect 44265 147280 44345 147290
rect 44585 147280 44665 147290
rect 44905 147280 44985 147290
rect 45225 147280 45305 147290
rect 45545 147280 45625 147290
rect 45865 147280 45945 147290
rect 46185 147280 46265 147290
rect 46505 147280 46585 147290
rect 46825 147280 46905 147290
rect 47145 147280 47225 147290
rect 47465 147280 47545 147290
rect 47785 147280 47865 147290
rect 48105 147280 48185 147290
rect 36020 147260 36100 147270
rect 36340 147260 36420 147270
rect 36660 147260 36740 147270
rect 36980 147260 37060 147270
rect 37300 147260 37380 147270
rect 37620 147260 37700 147270
rect 40180 147260 40260 147270
rect 40500 147260 40580 147270
rect 40820 147260 40900 147270
rect 41140 147260 41220 147270
rect 42740 147260 42820 147270
rect 43060 147260 43140 147270
rect 43380 147260 43460 147270
rect 43700 147260 43780 147270
rect 36100 147180 36110 147260
rect 36420 147180 36430 147260
rect 36740 147180 36750 147260
rect 37060 147180 37070 147260
rect 37380 147180 37390 147260
rect 37700 147180 37710 147260
rect 40260 147180 40270 147260
rect 40580 147180 40590 147260
rect 40900 147180 40910 147260
rect 41220 147180 41230 147260
rect 42820 147180 42830 147260
rect 43140 147180 43150 147260
rect 43460 147180 43470 147260
rect 43780 147210 43790 147260
rect 43700 147180 43790 147210
rect 44025 147200 44035 147280
rect 44345 147200 44355 147280
rect 44665 147200 44675 147280
rect 44985 147200 44995 147280
rect 45305 147200 45315 147280
rect 45625 147200 45635 147280
rect 45945 147200 45955 147280
rect 46265 147200 46275 147280
rect 46585 147200 46595 147280
rect 46905 147200 46915 147280
rect 47225 147200 47235 147280
rect 47545 147200 47555 147280
rect 47865 147200 47875 147280
rect 48185 147200 48195 147280
rect 48500 147230 48605 147360
rect 48640 147280 48650 147360
rect 49670 147270 49730 147390
rect 49760 147380 49840 147390
rect 49940 147380 50020 147390
rect 49840 147300 49850 147380
rect 50020 147300 50030 147380
rect 50260 147270 50320 147390
rect 50360 147380 50440 147390
rect 50540 147380 50620 147390
rect 50440 147300 50450 147380
rect 50620 147300 50630 147380
rect 50850 147270 50910 147390
rect 60360 147360 60440 147370
rect 60440 147280 60450 147360
rect 60660 147359 60670 147439
rect 60980 147359 60990 147439
rect 61400 147359 61410 147439
rect 61720 147359 61730 147439
rect 62140 147420 62150 147500
rect 73940 147420 73950 147500
rect 74080 147439 74160 147449
rect 74400 147439 74480 147449
rect 74820 147439 74900 147449
rect 75140 147439 75220 147449
rect 62060 147360 62140 147370
rect 73860 147360 73940 147370
rect 60740 147279 60820 147289
rect 61060 147279 61140 147289
rect 61480 147279 61560 147289
rect 61800 147279 61880 147289
rect 62140 147280 62150 147360
rect 73940 147280 73950 147360
rect 74160 147359 74170 147439
rect 74480 147359 74490 147439
rect 74900 147359 74910 147439
rect 75220 147359 75230 147439
rect 75640 147420 75650 147500
rect 87440 147420 87450 147500
rect 87580 147439 87660 147449
rect 87900 147439 87980 147449
rect 88320 147439 88400 147449
rect 88640 147439 88720 147449
rect 75560 147360 75640 147370
rect 87360 147360 87440 147370
rect 74240 147279 74320 147289
rect 74560 147279 74640 147289
rect 74980 147279 75060 147289
rect 75300 147279 75380 147289
rect 75640 147280 75650 147360
rect 87440 147280 87450 147360
rect 87660 147359 87670 147439
rect 87980 147359 87990 147439
rect 88400 147359 88410 147439
rect 88720 147359 88730 147439
rect 89140 147420 89150 147500
rect 100940 147420 100950 147500
rect 101080 147439 101160 147449
rect 101400 147439 101480 147449
rect 101820 147439 101900 147449
rect 102140 147439 102220 147449
rect 114580 147439 114660 147449
rect 114900 147439 114980 147449
rect 115320 147439 115400 147449
rect 115640 147439 115720 147449
rect 89060 147360 89140 147370
rect 100860 147360 100940 147370
rect 87740 147279 87820 147289
rect 88060 147279 88140 147289
rect 88480 147279 88560 147289
rect 88800 147279 88880 147289
rect 89140 147280 89150 147360
rect 100940 147280 100950 147360
rect 101160 147359 101170 147439
rect 101480 147359 101490 147439
rect 101900 147359 101910 147439
rect 102220 147359 102230 147439
rect 114660 147359 114670 147439
rect 114980 147359 114990 147439
rect 115400 147359 115410 147439
rect 115720 147359 115730 147439
rect 116140 147420 116150 147500
rect 127940 147420 127950 147500
rect 128080 147439 128160 147449
rect 128400 147439 128480 147449
rect 128820 147439 128900 147449
rect 129140 147439 129220 147449
rect 116060 147360 116140 147370
rect 127860 147360 127940 147370
rect 101240 147279 101320 147289
rect 101560 147279 101640 147289
rect 101980 147279 102060 147289
rect 102300 147279 102380 147289
rect 114740 147279 114820 147289
rect 115060 147279 115140 147289
rect 115480 147279 115560 147289
rect 115800 147279 115880 147289
rect 116140 147280 116150 147360
rect 127940 147280 127950 147360
rect 128160 147359 128170 147439
rect 128480 147359 128490 147439
rect 128900 147359 128910 147439
rect 129220 147359 129230 147439
rect 129640 147420 129650 147500
rect 141440 147420 141450 147500
rect 141545 147440 141625 147450
rect 141865 147440 141945 147450
rect 142185 147440 142200 147450
rect 145385 147440 145465 147450
rect 145705 147440 145785 147450
rect 146025 147440 146105 147450
rect 129560 147360 129640 147370
rect 141360 147360 141440 147370
rect 141625 147360 141635 147440
rect 141945 147360 141955 147440
rect 145465 147360 145475 147440
rect 145785 147360 145795 147440
rect 146105 147360 146115 147440
rect 146380 147420 146460 147430
rect 146700 147420 146780 147430
rect 147020 147420 147100 147430
rect 148940 147420 149020 147430
rect 149260 147420 149340 147430
rect 149580 147420 149660 147430
rect 152460 147420 152540 147430
rect 152780 147420 152860 147430
rect 153100 147420 153180 147430
rect 153420 147420 153500 147430
rect 153740 147420 153820 147430
rect 154060 147420 154140 147430
rect 154380 147420 154460 147430
rect 154700 147420 154780 147430
rect 155020 147420 155100 147430
rect 155340 147420 155420 147430
rect 155660 147420 155740 147430
rect 155980 147420 156000 147430
rect 128240 147279 128320 147289
rect 128560 147279 128640 147289
rect 128980 147279 129060 147289
rect 129300 147279 129380 147289
rect 129640 147280 129650 147360
rect 141440 147280 141450 147360
rect 146460 147340 146470 147420
rect 146780 147340 146790 147420
rect 147100 147340 147110 147420
rect 149020 147340 149030 147420
rect 149340 147340 149350 147420
rect 149660 147340 149670 147420
rect 152540 147340 152550 147420
rect 152860 147340 152870 147420
rect 153180 147340 153190 147420
rect 153500 147340 153510 147420
rect 153820 147340 153830 147420
rect 154140 147340 154150 147420
rect 154460 147340 154470 147420
rect 154780 147340 154790 147420
rect 155100 147340 155110 147420
rect 155420 147340 155430 147420
rect 155740 147340 155750 147420
rect 141705 147280 141785 147290
rect 142025 147280 142105 147290
rect 145225 147280 145305 147290
rect 145545 147280 145625 147290
rect 145865 147280 145945 147290
rect 49635 147230 49645 147250
rect 50225 147230 50235 147250
rect 50815 147230 50825 147250
rect 48500 147220 48640 147230
rect 49520 147220 50880 147230
rect 60360 147220 60440 147230
rect 43785 147120 43865 147130
rect 44105 147120 44185 147130
rect 44425 147120 44505 147130
rect 44745 147120 44825 147130
rect 45065 147120 45145 147130
rect 45385 147120 45465 147130
rect 45705 147120 45785 147130
rect 46025 147120 46105 147130
rect 46345 147120 46425 147130
rect 46665 147120 46745 147130
rect 46985 147120 47065 147130
rect 47305 147120 47385 147130
rect 47625 147120 47705 147130
rect 47945 147120 48025 147130
rect 48265 147120 48345 147130
rect 36180 147100 36260 147110
rect 36500 147100 36580 147110
rect 36820 147100 36900 147110
rect 37140 147100 37220 147110
rect 37460 147100 37540 147110
rect 40340 147100 40420 147110
rect 40660 147100 40740 147110
rect 40980 147100 41060 147110
rect 42580 147100 42660 147110
rect 42900 147100 42980 147110
rect 43220 147100 43300 147110
rect 43540 147100 43620 147110
rect 19300 147020 19310 147050
rect 19620 147020 19630 147050
rect 19940 147020 19950 147050
rect 20260 147020 20270 147050
rect 20580 147020 20590 147050
rect 20900 147020 20910 147050
rect 21220 147020 21230 147050
rect 21540 147020 21550 147050
rect 21860 147020 21870 147050
rect 22180 147020 22190 147050
rect 22500 147020 22510 147050
rect 22820 147020 22830 147050
rect 23140 147020 23150 147050
rect 23460 147020 23470 147050
rect 23780 147020 23790 147050
rect 24100 147020 24110 147050
rect 24420 147020 24430 147050
rect 24740 147020 24750 147050
rect 25060 147020 25070 147050
rect 25380 147020 25390 147050
rect 25700 147020 25710 147050
rect 26020 147020 26030 147050
rect 26340 147020 26350 147050
rect 30500 147020 30510 147050
rect 30820 147020 30830 147050
rect 31140 147020 31150 147050
rect 31460 147020 31470 147050
rect 31780 147020 31790 147050
rect 32100 147020 32110 147050
rect 32420 147020 32430 147050
rect 32740 147020 32750 147050
rect 33060 147020 33070 147050
rect 33380 147020 33390 147050
rect 33700 147020 33710 147050
rect 34020 147020 34030 147050
rect 34340 147020 34350 147050
rect 34660 147020 34670 147050
rect 34980 147020 34990 147050
rect 35300 147020 35310 147050
rect 35620 147020 35630 147050
rect 35940 147020 35950 147050
rect 36260 147020 36270 147100
rect 36580 147020 36590 147100
rect 36900 147020 36910 147100
rect 37220 147020 37230 147100
rect 37540 147020 37550 147100
rect 40420 147020 40430 147100
rect 40740 147020 40750 147100
rect 41060 147020 41070 147100
rect 42660 147020 42670 147100
rect 42980 147020 42990 147100
rect 43300 147020 43310 147100
rect 43620 147020 43630 147100
rect 43865 147040 43875 147120
rect 44185 147040 44195 147120
rect 44505 147040 44515 147120
rect 44825 147040 44835 147120
rect 45145 147040 45155 147120
rect 45465 147040 45475 147120
rect 45785 147040 45795 147120
rect 46105 147040 46115 147120
rect 46425 147040 46435 147120
rect 46745 147040 46755 147120
rect 47065 147040 47075 147120
rect 47385 147040 47395 147120
rect 47705 147040 47715 147120
rect 48025 147040 48035 147120
rect 48345 147040 48355 147120
rect 48500 147090 48605 147220
rect 48640 147140 48650 147220
rect 49400 147090 49520 147150
rect 48500 147080 48640 147090
rect 43945 146960 44025 146970
rect 44265 146960 44345 146970
rect 44585 146960 44665 146970
rect 44905 146960 44985 146970
rect 45225 146960 45305 146970
rect 45545 146960 45625 146970
rect 45865 146960 45945 146970
rect 46185 146960 46265 146970
rect 46505 146960 46585 146970
rect 46825 146960 46905 146970
rect 47145 146960 47225 146970
rect 47465 146960 47545 146970
rect 47785 146960 47865 146970
rect 48105 146960 48185 146970
rect 19060 146940 19140 146950
rect 19380 146940 19460 146950
rect 19700 146940 19780 146950
rect 20020 146940 20100 146950
rect 20340 146940 20420 146950
rect 20660 146940 20740 146950
rect 20980 146940 21060 146950
rect 21300 146940 21380 146950
rect 21620 146940 21700 146950
rect 21940 146940 22020 146950
rect 22260 146940 22340 146950
rect 22580 146940 22660 146950
rect 22900 146940 22980 146950
rect 23220 146940 23300 146950
rect 23540 146940 23620 146950
rect 23860 146940 23940 146950
rect 24180 146940 24260 146950
rect 24500 146940 24580 146950
rect 24820 146940 24900 146950
rect 25140 146940 25220 146950
rect 25460 146940 25540 146950
rect 25780 146940 25860 146950
rect 26100 146940 26180 146950
rect 26420 146940 26500 146950
rect 30580 146940 30660 146950
rect 30900 146940 30980 146950
rect 31220 146940 31300 146950
rect 31540 146940 31620 146950
rect 31860 146940 31940 146950
rect 32180 146940 32260 146950
rect 32500 146940 32580 146950
rect 32820 146940 32900 146950
rect 33140 146940 33220 146950
rect 33460 146940 33540 146950
rect 33780 146940 33860 146950
rect 34100 146940 34180 146950
rect 34420 146940 34500 146950
rect 34740 146940 34820 146950
rect 35060 146940 35140 146950
rect 35380 146940 35460 146950
rect 35700 146940 35780 146950
rect 36020 146940 36100 146950
rect 36340 146940 36420 146950
rect 36660 146940 36740 146950
rect 36980 146940 37060 146950
rect 37300 146940 37380 146950
rect 37620 146940 37700 146950
rect 40180 146940 40260 146950
rect 40500 146940 40580 146950
rect 40820 146940 40900 146950
rect 41140 146940 41220 146950
rect 42420 146940 42500 146950
rect 42740 146940 42820 146950
rect 43060 146940 43140 146950
rect 43380 146940 43460 146950
rect 43700 146940 43780 146950
rect 19140 146860 19150 146940
rect 19460 146860 19470 146940
rect 19780 146860 19790 146940
rect 20100 146860 20110 146940
rect 20420 146860 20430 146940
rect 20740 146860 20750 146940
rect 21060 146860 21070 146940
rect 21380 146860 21390 146940
rect 21700 146860 21710 146940
rect 22020 146860 22030 146940
rect 22340 146860 22350 146940
rect 22660 146860 22670 146940
rect 22980 146860 22990 146940
rect 23300 146860 23310 146940
rect 23620 146860 23630 146940
rect 23940 146860 23950 146940
rect 24260 146860 24270 146940
rect 24580 146860 24590 146940
rect 24900 146860 24910 146940
rect 25220 146860 25230 146940
rect 25540 146860 25550 146940
rect 25860 146860 25870 146940
rect 26180 146860 26190 146940
rect 26500 146860 26510 146940
rect 30660 146860 30670 146940
rect 30980 146860 30990 146940
rect 31300 146860 31310 146940
rect 31620 146860 31630 146940
rect 31940 146860 31950 146940
rect 32260 146860 32270 146940
rect 32580 146860 32590 146940
rect 32900 146860 32910 146940
rect 33220 146860 33230 146940
rect 33540 146860 33550 146940
rect 33860 146860 33870 146940
rect 34180 146860 34190 146940
rect 34500 146860 34510 146940
rect 34820 146860 34830 146940
rect 35140 146860 35150 146940
rect 35460 146860 35470 146940
rect 35780 146860 35790 146940
rect 36100 146860 36110 146940
rect 36420 146860 36430 146940
rect 36740 146860 36750 146940
rect 37060 146860 37070 146940
rect 37380 146860 37390 146940
rect 37700 146860 37710 146940
rect 40260 146860 40270 146940
rect 40580 146860 40590 146940
rect 40900 146860 40910 146940
rect 41220 146860 41230 146940
rect 42500 146860 42510 146940
rect 42820 146860 42830 146940
rect 43140 146860 43150 146940
rect 43460 146860 43470 146940
rect 43780 146890 43790 146940
rect 43700 146860 43790 146890
rect 44025 146880 44035 146960
rect 44345 146880 44355 146960
rect 44665 146880 44675 146960
rect 44985 146880 44995 146960
rect 45305 146880 45315 146960
rect 45625 146880 45635 146960
rect 45945 146880 45955 146960
rect 46265 146880 46275 146960
rect 46585 146880 46595 146960
rect 46905 146880 46915 146960
rect 47225 146880 47235 146960
rect 47545 146880 47555 146960
rect 47865 146880 47875 146960
rect 48185 146880 48195 146960
rect 48500 146950 48605 147080
rect 48640 147000 48650 147080
rect 49420 147070 49500 147080
rect 49500 146990 49510 147070
rect 49520 146970 49580 147090
rect 48500 146940 48640 146950
rect 48500 146810 48605 146940
rect 48640 146860 48650 146940
rect 49420 146930 49500 146940
rect 49500 146870 49510 146930
rect 49400 146810 49520 146870
rect 43785 146800 43865 146810
rect 44105 146800 44185 146810
rect 44425 146800 44505 146810
rect 44745 146800 44825 146810
rect 45065 146800 45145 146810
rect 45385 146800 45465 146810
rect 45705 146800 45785 146810
rect 46025 146800 46105 146810
rect 46345 146800 46425 146810
rect 46665 146800 46745 146810
rect 46985 146800 47065 146810
rect 47305 146800 47385 146810
rect 47625 146800 47705 146810
rect 47945 146800 48025 146810
rect 48265 146800 48345 146810
rect 48500 146800 48640 146810
rect 19220 146780 19300 146790
rect 19540 146780 19620 146790
rect 19860 146780 19940 146790
rect 20180 146780 20260 146790
rect 20500 146780 20580 146790
rect 20820 146780 20900 146790
rect 21140 146780 21220 146790
rect 21460 146780 21540 146790
rect 21780 146780 21860 146790
rect 22100 146780 22180 146790
rect 22420 146780 22500 146790
rect 22740 146780 22820 146790
rect 23060 146780 23140 146790
rect 23380 146780 23460 146790
rect 23700 146780 23780 146790
rect 24020 146780 24100 146790
rect 24340 146780 24420 146790
rect 24660 146780 24740 146790
rect 24980 146780 25060 146790
rect 25300 146780 25380 146790
rect 25620 146780 25700 146790
rect 25940 146780 26020 146790
rect 26260 146780 26340 146790
rect 30420 146780 30500 146790
rect 30740 146780 30820 146790
rect 31060 146780 31140 146790
rect 31380 146780 31460 146790
rect 31700 146780 31780 146790
rect 32020 146780 32100 146790
rect 32340 146780 32420 146790
rect 32660 146780 32740 146790
rect 32980 146780 33060 146790
rect 33300 146780 33380 146790
rect 33620 146780 33700 146790
rect 33940 146780 34020 146790
rect 34260 146780 34340 146790
rect 34580 146780 34660 146790
rect 34900 146780 34980 146790
rect 35220 146780 35300 146790
rect 35540 146780 35620 146790
rect 35860 146780 35940 146790
rect 36180 146780 36260 146790
rect 36500 146780 36580 146790
rect 36820 146780 36900 146790
rect 37140 146780 37220 146790
rect 37460 146780 37540 146790
rect 40340 146780 40420 146790
rect 40660 146780 40740 146790
rect 40980 146780 41060 146790
rect 42580 146780 42660 146790
rect 42900 146780 42980 146790
rect 43220 146780 43300 146790
rect 43540 146780 43620 146790
rect 19300 146700 19310 146780
rect 19620 146700 19630 146780
rect 19940 146700 19950 146780
rect 20260 146700 20270 146780
rect 20580 146700 20590 146780
rect 20900 146700 20910 146780
rect 21220 146700 21230 146780
rect 21540 146700 21550 146780
rect 21860 146700 21870 146780
rect 22180 146700 22190 146780
rect 22500 146700 22510 146780
rect 22820 146700 22830 146780
rect 23140 146700 23150 146780
rect 23460 146700 23470 146780
rect 23780 146700 23790 146780
rect 24100 146700 24110 146780
rect 24420 146700 24430 146780
rect 24740 146700 24750 146780
rect 25060 146700 25070 146780
rect 25380 146700 25390 146780
rect 25700 146700 25710 146780
rect 26020 146700 26030 146780
rect 26340 146700 26350 146780
rect 30500 146700 30510 146780
rect 30820 146700 30830 146780
rect 31140 146700 31150 146780
rect 31460 146700 31470 146780
rect 31780 146700 31790 146780
rect 32100 146700 32110 146780
rect 32420 146700 32430 146780
rect 32740 146700 32750 146780
rect 33060 146700 33070 146780
rect 33380 146700 33390 146780
rect 33700 146700 33710 146780
rect 34020 146700 34030 146780
rect 34340 146700 34350 146780
rect 34660 146700 34670 146780
rect 34980 146700 34990 146780
rect 35300 146700 35310 146780
rect 35620 146700 35630 146780
rect 35940 146700 35950 146780
rect 36260 146700 36270 146780
rect 36580 146700 36590 146780
rect 36900 146700 36910 146780
rect 37220 146700 37230 146780
rect 37540 146700 37550 146780
rect 40420 146700 40430 146780
rect 40740 146700 40750 146780
rect 41060 146700 41070 146780
rect 42660 146700 42670 146780
rect 42980 146700 42990 146780
rect 43300 146700 43310 146780
rect 43620 146700 43630 146780
rect 43865 146720 43875 146800
rect 44185 146720 44195 146800
rect 44505 146720 44515 146800
rect 44825 146720 44835 146800
rect 45145 146720 45155 146800
rect 45465 146720 45475 146800
rect 45785 146720 45795 146800
rect 46105 146720 46115 146800
rect 46425 146720 46435 146800
rect 46745 146720 46755 146800
rect 47065 146720 47075 146800
rect 47385 146720 47395 146800
rect 47705 146720 47715 146800
rect 48025 146720 48035 146800
rect 48345 146720 48355 146800
rect 48500 146670 48605 146800
rect 48640 146720 48650 146800
rect 49420 146790 49500 146800
rect 49500 146710 49510 146790
rect 49520 146690 49580 146810
rect 48500 146660 48640 146670
rect 43945 146640 44025 146650
rect 44265 146640 44345 146650
rect 44585 146640 44665 146650
rect 44905 146640 44985 146650
rect 45225 146640 45305 146650
rect 45545 146640 45625 146650
rect 45865 146640 45945 146650
rect 46185 146640 46265 146650
rect 46505 146640 46585 146650
rect 46825 146640 46905 146650
rect 47145 146640 47225 146650
rect 47465 146640 47545 146650
rect 47785 146640 47865 146650
rect 48105 146640 48185 146650
rect 19060 146620 19140 146630
rect 19380 146620 19460 146630
rect 19700 146620 19780 146630
rect 20020 146620 20100 146630
rect 20340 146620 20420 146630
rect 20660 146620 20740 146630
rect 20980 146620 21060 146630
rect 21300 146620 21380 146630
rect 21620 146620 21700 146630
rect 21940 146620 22020 146630
rect 22260 146620 22340 146630
rect 22580 146620 22660 146630
rect 22900 146620 22980 146630
rect 23220 146620 23300 146630
rect 23540 146620 23620 146630
rect 23860 146620 23940 146630
rect 24180 146620 24260 146630
rect 24500 146620 24580 146630
rect 24820 146620 24900 146630
rect 25140 146620 25220 146630
rect 25460 146620 25540 146630
rect 25780 146620 25860 146630
rect 26100 146620 26180 146630
rect 26420 146620 26500 146630
rect 30580 146620 30660 146630
rect 30900 146620 30980 146630
rect 31220 146620 31300 146630
rect 31540 146620 31620 146630
rect 31860 146620 31940 146630
rect 32180 146620 32260 146630
rect 32500 146620 32580 146630
rect 32820 146620 32900 146630
rect 33140 146620 33220 146630
rect 33460 146620 33540 146630
rect 33780 146620 33860 146630
rect 34100 146620 34180 146630
rect 34420 146620 34500 146630
rect 34740 146620 34820 146630
rect 35060 146620 35140 146630
rect 35380 146620 35460 146630
rect 35700 146620 35780 146630
rect 36020 146620 36100 146630
rect 36340 146620 36420 146630
rect 36660 146620 36740 146630
rect 36980 146620 37060 146630
rect 37300 146620 37380 146630
rect 37620 146620 37700 146630
rect 40180 146620 40260 146630
rect 40500 146620 40580 146630
rect 40820 146620 40900 146630
rect 41140 146620 41220 146630
rect 42420 146620 42500 146630
rect 42740 146620 42820 146630
rect 43060 146620 43140 146630
rect 43380 146620 43460 146630
rect 43700 146620 43780 146630
rect 19140 146540 19150 146620
rect 19460 146540 19470 146620
rect 19780 146540 19790 146620
rect 20100 146540 20110 146620
rect 20420 146540 20430 146620
rect 20740 146540 20750 146620
rect 21060 146540 21070 146620
rect 21380 146540 21390 146620
rect 21700 146540 21710 146620
rect 22020 146540 22030 146620
rect 22340 146540 22350 146620
rect 22660 146540 22670 146620
rect 22980 146540 22990 146620
rect 23300 146540 23310 146620
rect 23620 146540 23630 146620
rect 23940 146540 23950 146620
rect 24260 146540 24270 146620
rect 24580 146540 24590 146620
rect 24900 146540 24910 146620
rect 25220 146540 25230 146620
rect 25540 146540 25550 146620
rect 25860 146540 25870 146620
rect 26180 146540 26190 146620
rect 26500 146540 26510 146620
rect 30660 146540 30670 146620
rect 30980 146540 30990 146620
rect 31300 146540 31310 146620
rect 31620 146540 31630 146620
rect 31940 146540 31950 146620
rect 32260 146540 32270 146620
rect 32580 146540 32590 146620
rect 32900 146540 32910 146620
rect 33220 146540 33230 146620
rect 33540 146540 33550 146620
rect 33860 146540 33870 146620
rect 34180 146540 34190 146620
rect 34500 146540 34510 146620
rect 34820 146540 34830 146620
rect 35140 146540 35150 146620
rect 35460 146540 35470 146620
rect 35780 146540 35790 146620
rect 36100 146540 36110 146620
rect 36420 146540 36430 146620
rect 36740 146540 36750 146620
rect 37060 146540 37070 146620
rect 37380 146540 37390 146620
rect 37700 146540 37710 146620
rect 40260 146540 40270 146620
rect 40580 146540 40590 146620
rect 40900 146540 40910 146620
rect 41220 146540 41230 146620
rect 42500 146540 42510 146620
rect 42820 146540 42830 146620
rect 43140 146540 43150 146620
rect 43460 146540 43470 146620
rect 43780 146570 43790 146620
rect 43700 146540 43790 146570
rect 44025 146560 44035 146640
rect 44345 146560 44355 146640
rect 44665 146560 44675 146640
rect 44985 146560 44995 146640
rect 45305 146560 45315 146640
rect 45625 146560 45635 146640
rect 45945 146560 45955 146640
rect 46265 146560 46275 146640
rect 46585 146560 46595 146640
rect 46905 146560 46915 146640
rect 47225 146560 47235 146640
rect 47545 146560 47555 146640
rect 47865 146560 47875 146640
rect 48185 146560 48195 146640
rect 48500 146530 48605 146660
rect 48640 146580 48650 146660
rect 49420 146650 49500 146660
rect 49500 146570 49510 146650
rect 48500 146520 48640 146530
rect 43785 146480 43865 146490
rect 44105 146480 44185 146490
rect 44425 146480 44505 146490
rect 44745 146480 44825 146490
rect 45065 146480 45145 146490
rect 45385 146480 45465 146490
rect 45705 146480 45785 146490
rect 46025 146480 46105 146490
rect 46345 146480 46425 146490
rect 46665 146480 46745 146490
rect 46985 146480 47065 146490
rect 47305 146480 47385 146490
rect 47625 146480 47705 146490
rect 47945 146480 48025 146490
rect 48265 146480 48345 146490
rect 42580 146460 42660 146470
rect 42900 146460 42980 146470
rect 43220 146460 43300 146470
rect 43540 146460 43620 146470
rect 42660 146380 42670 146460
rect 42980 146380 42990 146460
rect 43300 146380 43310 146460
rect 43620 146380 43630 146460
rect 43865 146400 43875 146480
rect 44185 146400 44195 146480
rect 44505 146400 44515 146480
rect 44825 146400 44835 146480
rect 45145 146400 45155 146480
rect 45465 146400 45475 146480
rect 45785 146400 45795 146480
rect 46105 146400 46115 146480
rect 46425 146400 46435 146480
rect 46745 146400 46755 146480
rect 47065 146400 47075 146480
rect 47385 146400 47395 146480
rect 47705 146400 47715 146480
rect 48025 146400 48035 146480
rect 48345 146400 48355 146480
rect 48500 146390 48605 146520
rect 48640 146440 48650 146520
rect 49635 146460 49645 147220
rect 49650 146500 49660 147140
rect 49700 147090 49820 147150
rect 49820 146980 49880 147090
rect 49700 146970 49880 146980
rect 49700 146810 49820 146870
rect 49820 146700 49880 146810
rect 49700 146690 49880 146700
rect 49960 146510 49970 147130
rect 49990 147090 50110 147150
rect 50010 147070 50090 147080
rect 50090 146990 50100 147070
rect 50110 146970 50170 147090
rect 50010 146930 50090 146940
rect 50090 146870 50100 146930
rect 49990 146810 50110 146870
rect 50010 146790 50090 146800
rect 50090 146710 50100 146790
rect 50110 146690 50170 146810
rect 50010 146650 50090 146660
rect 50090 146570 50100 146650
rect 49950 146500 50160 146510
rect 50225 146460 50235 147220
rect 50240 146500 50250 147140
rect 50290 147090 50410 147150
rect 50410 146980 50470 147090
rect 50290 146970 50470 146980
rect 50290 146810 50410 146870
rect 50410 146700 50470 146810
rect 50290 146690 50470 146700
rect 50550 146510 50560 147130
rect 50580 147090 50700 147150
rect 50600 147070 50680 147080
rect 50680 146990 50690 147070
rect 50700 146970 50760 147090
rect 50600 146930 50680 146940
rect 50680 146870 50690 146930
rect 50580 146810 50700 146870
rect 50600 146790 50680 146800
rect 50680 146710 50690 146790
rect 50700 146690 50760 146810
rect 50600 146650 50680 146660
rect 50680 146570 50690 146650
rect 50540 146500 50750 146510
rect 50815 146460 50825 147220
rect 50830 146500 50840 147140
rect 50880 147090 51000 147150
rect 60440 147140 60450 147220
rect 60820 147199 60830 147279
rect 61140 147199 61150 147279
rect 61560 147199 61570 147279
rect 61880 147199 61890 147279
rect 62060 147220 62140 147230
rect 73860 147220 73940 147230
rect 62140 147140 62150 147220
rect 73940 147140 73950 147220
rect 74320 147199 74330 147279
rect 74640 147199 74650 147279
rect 75060 147199 75070 147279
rect 75380 147199 75390 147279
rect 75560 147220 75640 147230
rect 87360 147220 87440 147230
rect 75640 147140 75650 147220
rect 87440 147140 87450 147220
rect 87820 147199 87830 147279
rect 88140 147199 88150 147279
rect 88560 147199 88570 147279
rect 88880 147199 88890 147279
rect 89060 147220 89140 147230
rect 100860 147220 100940 147230
rect 89140 147140 89150 147220
rect 100940 147140 100950 147220
rect 101320 147199 101330 147279
rect 101640 147199 101650 147279
rect 102060 147199 102070 147279
rect 102380 147199 102390 147279
rect 103990 147140 104000 147200
rect 104170 147140 104180 147200
rect 104350 147140 104360 147200
rect 104530 147140 104540 147200
rect 104710 147140 104720 147200
rect 104890 147140 104900 147200
rect 105070 147140 105080 147200
rect 105250 147140 105260 147200
rect 105430 147140 105440 147200
rect 105610 147140 105620 147200
rect 105790 147140 105800 147200
rect 105970 147140 105980 147200
rect 106150 147140 106160 147200
rect 106330 147140 106340 147200
rect 106510 147140 106520 147200
rect 106690 147140 106700 147200
rect 106870 147140 106880 147200
rect 107050 147140 107060 147200
rect 107230 147140 107240 147200
rect 107410 147140 107420 147200
rect 107590 147140 107600 147200
rect 107770 147140 107780 147200
rect 107950 147140 107960 147200
rect 108130 147140 108140 147200
rect 108310 147140 108320 147200
rect 108490 147140 108500 147200
rect 108670 147140 108680 147200
rect 108850 147140 108860 147200
rect 109030 147140 109040 147200
rect 109210 147140 109220 147200
rect 109390 147140 109400 147200
rect 109570 147140 109580 147200
rect 109750 147140 109760 147200
rect 109930 147140 109940 147200
rect 110110 147140 110120 147200
rect 110290 147140 110300 147200
rect 110470 147140 110480 147200
rect 110650 147140 110660 147200
rect 110830 147140 110840 147200
rect 111010 147140 111020 147200
rect 111190 147140 111200 147200
rect 111370 147140 111380 147200
rect 111550 147140 111560 147200
rect 111730 147140 111740 147200
rect 111910 147140 111920 147200
rect 112090 147140 112100 147200
rect 112270 147140 112280 147200
rect 112450 147140 112460 147200
rect 112630 147140 112640 147200
rect 112810 147140 112820 147200
rect 112990 147140 113000 147200
rect 114820 147199 114830 147279
rect 115140 147199 115150 147279
rect 115560 147199 115570 147279
rect 115880 147199 115890 147279
rect 116060 147220 116140 147230
rect 127860 147220 127940 147230
rect 116140 147140 116150 147220
rect 60580 147119 60660 147129
rect 60900 147119 60980 147129
rect 61320 147119 61400 147129
rect 61640 147119 61720 147129
rect 51000 146970 51060 147090
rect 60360 147080 60440 147090
rect 60440 147000 60450 147080
rect 60660 147039 60670 147119
rect 60980 147039 60990 147119
rect 61400 147039 61410 147119
rect 61720 147039 61730 147119
rect 62900 147090 63020 147140
rect 62060 147080 62140 147090
rect 62140 147000 62150 147080
rect 62920 147070 63000 147080
rect 63000 146990 63010 147070
rect 63020 146970 63080 147090
rect 60740 146959 60820 146969
rect 61060 146959 61140 146969
rect 61480 146959 61560 146969
rect 61800 146959 61880 146969
rect 60360 146940 60440 146950
rect 50900 146930 50980 146940
rect 50980 146870 50990 146930
rect 50880 146810 51000 146870
rect 60440 146860 60450 146940
rect 60820 146879 60830 146959
rect 61140 146879 61150 146959
rect 61560 146879 61570 146959
rect 61880 146879 61890 146959
rect 62060 146940 62140 146950
rect 62140 146860 62150 146940
rect 62920 146930 63000 146940
rect 63000 146870 63010 146930
rect 62900 146810 63020 146870
rect 51000 146690 51060 146810
rect 60360 146800 60440 146810
rect 60440 146720 60450 146800
rect 60580 146799 60660 146809
rect 60900 146799 60980 146809
rect 61320 146799 61400 146809
rect 61640 146799 61720 146809
rect 62060 146800 62140 146810
rect 60660 146719 60670 146799
rect 60980 146719 60990 146799
rect 61400 146719 61410 146799
rect 61720 146719 61730 146799
rect 62140 146720 62150 146800
rect 62920 146790 63000 146800
rect 63000 146710 63010 146790
rect 63020 146690 63080 146810
rect 60360 146660 60440 146670
rect 62060 146660 62140 146670
rect 50900 146650 50980 146660
rect 50980 146570 50990 146650
rect 60440 146580 60450 146660
rect 60740 146639 60820 146649
rect 61060 146639 61140 146649
rect 61480 146639 61560 146649
rect 61800 146639 61880 146649
rect 60820 146559 60830 146639
rect 61140 146559 61150 146639
rect 61560 146559 61570 146639
rect 61880 146559 61890 146639
rect 62140 146580 62150 146660
rect 62920 146650 63000 146660
rect 63000 146570 63010 146650
rect 60360 146520 60440 146530
rect 62060 146520 62140 146530
rect 49585 146450 49635 146460
rect 50175 146450 50225 146460
rect 50765 146450 50815 146460
rect 60440 146440 60450 146520
rect 60580 146479 60660 146489
rect 60900 146479 60980 146489
rect 61320 146479 61400 146489
rect 61640 146479 61720 146489
rect 60660 146399 60670 146479
rect 60980 146399 60990 146479
rect 61400 146399 61410 146479
rect 61720 146399 61730 146479
rect 62140 146440 62150 146520
rect 63135 146460 63145 147140
rect 63150 146500 63160 147140
rect 63200 147090 63320 147140
rect 63320 146980 63380 147090
rect 63200 146970 63380 146980
rect 63200 146810 63320 146870
rect 63320 146700 63380 146810
rect 63200 146690 63380 146700
rect 63460 146510 63470 147130
rect 63490 147090 63610 147140
rect 63510 147070 63590 147080
rect 63590 146990 63600 147070
rect 63610 146970 63670 147090
rect 63510 146930 63590 146940
rect 63590 146870 63600 146930
rect 63490 146810 63610 146870
rect 63510 146790 63590 146800
rect 63590 146710 63600 146790
rect 63610 146690 63670 146810
rect 63510 146650 63590 146660
rect 63590 146570 63600 146650
rect 63450 146500 63660 146510
rect 63725 146460 63735 147140
rect 63740 146500 63750 147140
rect 63790 147090 63910 147140
rect 63910 146980 63970 147090
rect 63790 146970 63970 146980
rect 63790 146810 63910 146870
rect 63910 146700 63970 146810
rect 63790 146690 63970 146700
rect 64050 146510 64060 147130
rect 64080 147090 64200 147140
rect 64100 147070 64180 147080
rect 64180 146990 64190 147070
rect 64200 146970 64260 147090
rect 64100 146930 64180 146940
rect 64180 146870 64190 146930
rect 64080 146810 64200 146870
rect 64100 146790 64180 146800
rect 64180 146710 64190 146790
rect 64200 146690 64260 146810
rect 64100 146650 64180 146660
rect 64180 146570 64190 146650
rect 64040 146500 64250 146510
rect 64315 146460 64325 147140
rect 64330 146500 64340 147140
rect 64380 147090 64500 147140
rect 74080 147119 74160 147129
rect 74400 147119 74480 147129
rect 74820 147119 74900 147129
rect 75140 147119 75220 147129
rect 64500 146970 64560 147090
rect 73860 147080 73940 147090
rect 73940 147000 73950 147080
rect 74160 147039 74170 147119
rect 74480 147039 74490 147119
rect 74900 147039 74910 147119
rect 75220 147039 75230 147119
rect 76400 147090 76520 147140
rect 75560 147080 75640 147090
rect 75640 147000 75650 147080
rect 76420 147070 76500 147080
rect 76500 146990 76510 147070
rect 76520 146970 76580 147090
rect 74240 146959 74320 146969
rect 74560 146959 74640 146969
rect 74980 146959 75060 146969
rect 75300 146959 75380 146969
rect 73860 146940 73940 146950
rect 64400 146930 64480 146940
rect 64480 146870 64490 146930
rect 64380 146810 64500 146870
rect 73940 146860 73950 146940
rect 74320 146879 74330 146959
rect 74640 146879 74650 146959
rect 75060 146879 75070 146959
rect 75380 146879 75390 146959
rect 75560 146940 75640 146950
rect 75640 146860 75650 146940
rect 76420 146930 76500 146940
rect 76500 146870 76510 146930
rect 76400 146810 76520 146870
rect 64500 146690 64560 146810
rect 73860 146800 73940 146810
rect 73940 146720 73950 146800
rect 74080 146799 74160 146809
rect 74400 146799 74480 146809
rect 74820 146799 74900 146809
rect 75140 146799 75220 146809
rect 75560 146800 75640 146810
rect 74160 146719 74170 146799
rect 74480 146719 74490 146799
rect 74900 146719 74910 146799
rect 75220 146719 75230 146799
rect 75640 146720 75650 146800
rect 76420 146790 76500 146800
rect 76500 146710 76510 146790
rect 76520 146690 76580 146810
rect 73860 146660 73940 146670
rect 75560 146660 75640 146670
rect 64400 146650 64480 146660
rect 64480 146570 64490 146650
rect 73940 146580 73950 146660
rect 74240 146639 74320 146649
rect 74560 146639 74640 146649
rect 74980 146639 75060 146649
rect 75300 146639 75380 146649
rect 74320 146559 74330 146639
rect 74640 146559 74650 146639
rect 75060 146559 75070 146639
rect 75380 146559 75390 146639
rect 75640 146580 75650 146660
rect 76420 146650 76500 146660
rect 76500 146570 76510 146650
rect 73860 146520 73940 146530
rect 75560 146520 75640 146530
rect 63085 146450 63135 146460
rect 63675 146450 63725 146460
rect 64265 146450 64315 146460
rect 73940 146440 73950 146520
rect 74080 146479 74160 146489
rect 74400 146479 74480 146489
rect 74820 146479 74900 146489
rect 75140 146479 75220 146489
rect 74160 146399 74170 146479
rect 74480 146399 74490 146479
rect 74900 146399 74910 146479
rect 75220 146399 75230 146479
rect 75640 146440 75650 146520
rect 76635 146460 76645 147140
rect 76650 146500 76660 147140
rect 76700 147090 76820 147140
rect 76820 146980 76880 147090
rect 76700 146970 76880 146980
rect 76700 146810 76820 146870
rect 76820 146700 76880 146810
rect 76700 146690 76880 146700
rect 76960 146510 76970 147130
rect 76990 147090 77110 147140
rect 77010 147070 77090 147080
rect 77090 146990 77100 147070
rect 77110 146970 77170 147090
rect 77010 146930 77090 146940
rect 77090 146870 77100 146930
rect 76990 146810 77110 146870
rect 77010 146790 77090 146800
rect 77090 146710 77100 146790
rect 77110 146690 77170 146810
rect 77010 146650 77090 146660
rect 77090 146570 77100 146650
rect 76950 146500 77160 146510
rect 77225 146460 77235 147140
rect 77240 146500 77250 147140
rect 77290 147090 77410 147140
rect 77410 146980 77470 147090
rect 77290 146970 77470 146980
rect 77290 146810 77410 146870
rect 77410 146700 77470 146810
rect 77290 146690 77470 146700
rect 77550 146510 77560 147130
rect 77580 147090 77700 147140
rect 77600 147070 77680 147080
rect 77680 146990 77690 147070
rect 77700 146970 77760 147090
rect 77600 146930 77680 146940
rect 77680 146870 77690 146930
rect 77580 146810 77700 146870
rect 77600 146790 77680 146800
rect 77680 146710 77690 146790
rect 77700 146690 77760 146810
rect 77600 146650 77680 146660
rect 77680 146570 77690 146650
rect 77540 146500 77750 146510
rect 77815 146460 77825 147140
rect 77830 146500 77840 147140
rect 77880 147090 78000 147140
rect 87580 147119 87660 147129
rect 87900 147119 87980 147129
rect 88320 147119 88400 147129
rect 88640 147119 88720 147129
rect 78000 146970 78060 147090
rect 87360 147080 87440 147090
rect 87440 147000 87450 147080
rect 87660 147039 87670 147119
rect 87980 147039 87990 147119
rect 88400 147039 88410 147119
rect 88720 147039 88730 147119
rect 89900 147090 90020 147140
rect 89060 147080 89140 147090
rect 89140 147000 89150 147080
rect 89920 147070 90000 147080
rect 90000 146990 90010 147070
rect 90020 146970 90080 147090
rect 87740 146959 87820 146969
rect 88060 146959 88140 146969
rect 88480 146959 88560 146969
rect 88800 146959 88880 146969
rect 87360 146940 87440 146950
rect 77900 146930 77980 146940
rect 77980 146870 77990 146930
rect 77880 146810 78000 146870
rect 87440 146860 87450 146940
rect 87820 146879 87830 146959
rect 88140 146879 88150 146959
rect 88560 146879 88570 146959
rect 88880 146879 88890 146959
rect 89060 146940 89140 146950
rect 89140 146860 89150 146940
rect 89920 146930 90000 146940
rect 90000 146870 90010 146930
rect 89900 146810 90020 146870
rect 78000 146690 78060 146810
rect 87360 146800 87440 146810
rect 87440 146720 87450 146800
rect 87580 146799 87660 146809
rect 87900 146799 87980 146809
rect 88320 146799 88400 146809
rect 88640 146799 88720 146809
rect 89060 146800 89140 146810
rect 87660 146719 87670 146799
rect 87980 146719 87990 146799
rect 88400 146719 88410 146799
rect 88720 146719 88730 146799
rect 89140 146720 89150 146800
rect 89920 146790 90000 146800
rect 90000 146710 90010 146790
rect 90020 146690 90080 146810
rect 87360 146660 87440 146670
rect 89060 146660 89140 146670
rect 77900 146650 77980 146660
rect 77980 146570 77990 146650
rect 87440 146580 87450 146660
rect 87740 146639 87820 146649
rect 88060 146639 88140 146649
rect 88480 146639 88560 146649
rect 88800 146639 88880 146649
rect 87820 146559 87830 146639
rect 88140 146559 88150 146639
rect 88560 146559 88570 146639
rect 88880 146559 88890 146639
rect 89140 146580 89150 146660
rect 89920 146650 90000 146660
rect 90000 146570 90010 146650
rect 87360 146520 87440 146530
rect 89060 146520 89140 146530
rect 76585 146450 76635 146460
rect 77175 146450 77225 146460
rect 77765 146450 77815 146460
rect 87440 146440 87450 146520
rect 87580 146479 87660 146489
rect 87900 146479 87980 146489
rect 88320 146479 88400 146489
rect 88640 146479 88720 146489
rect 87660 146399 87670 146479
rect 87980 146399 87990 146479
rect 88400 146399 88410 146479
rect 88720 146399 88730 146479
rect 89140 146440 89150 146520
rect 90135 146460 90145 147140
rect 90150 146500 90160 147140
rect 90200 147090 90320 147140
rect 90320 146980 90380 147090
rect 90200 146970 90380 146980
rect 90200 146810 90320 146870
rect 90320 146700 90380 146810
rect 90200 146690 90380 146700
rect 90460 146510 90470 147130
rect 90490 147090 90610 147140
rect 90510 147070 90590 147080
rect 90590 146990 90600 147070
rect 90610 146970 90670 147090
rect 90510 146930 90590 146940
rect 90590 146870 90600 146930
rect 90490 146810 90610 146870
rect 90510 146790 90590 146800
rect 90590 146710 90600 146790
rect 90610 146690 90670 146810
rect 90510 146650 90590 146660
rect 90590 146570 90600 146650
rect 90450 146500 90660 146510
rect 90725 146460 90735 147140
rect 90740 146500 90750 147140
rect 90790 147090 90910 147140
rect 90910 146980 90970 147090
rect 90790 146970 90970 146980
rect 90790 146810 90910 146870
rect 90910 146700 90970 146810
rect 90790 146690 90970 146700
rect 91050 146510 91060 147130
rect 91080 147090 91200 147140
rect 91100 147070 91180 147080
rect 91180 146990 91190 147070
rect 91200 146970 91260 147090
rect 91100 146930 91180 146940
rect 91180 146870 91190 146930
rect 91080 146810 91200 146870
rect 91100 146790 91180 146800
rect 91180 146710 91190 146790
rect 91200 146690 91260 146810
rect 91100 146650 91180 146660
rect 91180 146570 91190 146650
rect 91040 146500 91250 146510
rect 91315 146460 91325 147140
rect 91330 146500 91340 147140
rect 91380 147090 91500 147140
rect 101080 147119 101160 147129
rect 101400 147119 101480 147129
rect 101820 147119 101900 147129
rect 102140 147119 102220 147129
rect 114580 147119 114660 147129
rect 114900 147119 114980 147129
rect 115320 147119 115400 147129
rect 115640 147119 115720 147129
rect 91500 146970 91560 147090
rect 100860 147080 100940 147090
rect 100940 147000 100950 147080
rect 101160 147039 101170 147119
rect 101480 147039 101490 147119
rect 101900 147039 101910 147119
rect 102220 147039 102230 147119
rect 103910 147040 103990 147050
rect 104090 147040 104170 147050
rect 104270 147040 104350 147050
rect 104450 147040 104530 147050
rect 104630 147040 104710 147050
rect 104810 147040 104890 147050
rect 104990 147040 105070 147050
rect 105170 147040 105250 147050
rect 105350 147040 105430 147050
rect 105530 147040 105610 147050
rect 105710 147040 105790 147050
rect 105890 147040 105970 147050
rect 106070 147040 106150 147050
rect 106250 147040 106330 147050
rect 106430 147040 106510 147050
rect 106610 147040 106690 147050
rect 106790 147040 106870 147050
rect 106970 147040 107050 147050
rect 107150 147040 107230 147050
rect 107330 147040 107410 147050
rect 107510 147040 107590 147050
rect 107690 147040 107770 147050
rect 107870 147040 107950 147050
rect 108050 147040 108130 147050
rect 108230 147040 108310 147050
rect 108410 147040 108490 147050
rect 108590 147040 108670 147050
rect 108770 147040 108850 147050
rect 108950 147040 109030 147050
rect 109130 147040 109210 147050
rect 109310 147040 109390 147050
rect 109490 147040 109570 147050
rect 109670 147040 109750 147050
rect 109850 147040 109930 147050
rect 110030 147040 110110 147050
rect 110210 147040 110290 147050
rect 110390 147040 110470 147050
rect 110570 147040 110650 147050
rect 110750 147040 110830 147050
rect 110930 147040 111010 147050
rect 111110 147040 111190 147050
rect 111290 147040 111370 147050
rect 111470 147040 111550 147050
rect 111650 147040 111730 147050
rect 111830 147040 111910 147050
rect 112010 147040 112090 147050
rect 112190 147040 112270 147050
rect 112370 147040 112450 147050
rect 112550 147040 112630 147050
rect 112730 147040 112810 147050
rect 112910 147040 112990 147050
rect 101240 146959 101320 146969
rect 101560 146959 101640 146969
rect 101980 146959 102060 146969
rect 102300 146959 102380 146969
rect 103990 146960 104000 147040
rect 104170 146960 104180 147040
rect 104350 146960 104360 147040
rect 104530 146960 104540 147040
rect 104710 146960 104720 147040
rect 104890 146960 104900 147040
rect 105070 146960 105080 147040
rect 105250 146960 105260 147040
rect 105430 146960 105440 147040
rect 105610 146960 105620 147040
rect 105790 146960 105800 147040
rect 105970 146960 105980 147040
rect 106150 146960 106160 147040
rect 106330 146960 106340 147040
rect 106510 146960 106520 147040
rect 106690 146960 106700 147040
rect 106870 146960 106880 147040
rect 107050 146960 107060 147040
rect 107230 146960 107240 147040
rect 107410 146960 107420 147040
rect 107590 146960 107600 147040
rect 107770 146960 107780 147040
rect 107950 146960 107960 147040
rect 108130 146960 108140 147040
rect 108310 146960 108320 147040
rect 108490 146960 108500 147040
rect 108670 146960 108680 147040
rect 108850 146960 108860 147040
rect 109030 146960 109040 147040
rect 109210 146960 109220 147040
rect 109390 146960 109400 147040
rect 109570 146960 109580 147040
rect 109750 146960 109760 147040
rect 109930 146960 109940 147040
rect 110110 146960 110120 147040
rect 110290 146960 110300 147040
rect 110470 146960 110480 147040
rect 110650 146960 110660 147040
rect 110830 146960 110840 147040
rect 111010 146960 111020 147040
rect 111190 146960 111200 147040
rect 111370 146960 111380 147040
rect 111550 146960 111560 147040
rect 111730 146960 111740 147040
rect 111910 146960 111920 147040
rect 112090 146960 112100 147040
rect 112270 146960 112280 147040
rect 112450 146960 112460 147040
rect 112630 146960 112640 147040
rect 112810 146960 112820 147040
rect 112990 146960 113000 147040
rect 114660 147039 114670 147119
rect 114980 147039 114990 147119
rect 115400 147039 115410 147119
rect 115720 147039 115730 147119
rect 116900 147090 117020 147150
rect 116060 147080 116140 147090
rect 116140 147000 116150 147080
rect 116920 147070 117000 147080
rect 117000 146990 117010 147070
rect 117020 146970 117080 147090
rect 114740 146959 114820 146969
rect 115060 146959 115140 146969
rect 115480 146959 115560 146969
rect 115800 146959 115880 146969
rect 100860 146940 100940 146950
rect 91400 146930 91480 146940
rect 91480 146870 91490 146930
rect 91380 146810 91500 146870
rect 100940 146860 100950 146940
rect 101320 146879 101330 146959
rect 101640 146879 101650 146959
rect 102060 146879 102070 146959
rect 102380 146879 102390 146959
rect 114820 146879 114830 146959
rect 115140 146879 115150 146959
rect 115560 146879 115570 146959
rect 115880 146879 115890 146959
rect 116060 146940 116140 146950
rect 103910 146860 103990 146870
rect 104090 146860 104170 146870
rect 104270 146860 104350 146870
rect 104450 146860 104530 146870
rect 104630 146860 104710 146870
rect 104810 146860 104890 146870
rect 104990 146860 105070 146870
rect 105170 146860 105250 146870
rect 105350 146860 105430 146870
rect 105530 146860 105610 146870
rect 105710 146860 105790 146870
rect 105890 146860 105970 146870
rect 106070 146860 106150 146870
rect 106250 146860 106330 146870
rect 106430 146860 106510 146870
rect 106610 146860 106690 146870
rect 106790 146860 106870 146870
rect 106970 146860 107050 146870
rect 107150 146860 107230 146870
rect 107330 146860 107410 146870
rect 107510 146860 107590 146870
rect 107690 146860 107770 146870
rect 107870 146860 107950 146870
rect 108050 146860 108130 146870
rect 108230 146860 108310 146870
rect 108410 146860 108490 146870
rect 108590 146860 108670 146870
rect 108770 146860 108850 146870
rect 108950 146860 109030 146870
rect 109130 146860 109210 146870
rect 109310 146860 109390 146870
rect 109490 146860 109570 146870
rect 109670 146860 109750 146870
rect 109850 146860 109930 146870
rect 110030 146860 110110 146870
rect 110210 146860 110290 146870
rect 110390 146860 110470 146870
rect 110570 146860 110650 146870
rect 110750 146860 110830 146870
rect 110930 146860 111010 146870
rect 111110 146860 111190 146870
rect 111290 146860 111370 146870
rect 111470 146860 111550 146870
rect 111650 146860 111730 146870
rect 111830 146860 111910 146870
rect 112010 146860 112090 146870
rect 112190 146860 112270 146870
rect 112370 146860 112450 146870
rect 112550 146860 112630 146870
rect 112730 146860 112810 146870
rect 112910 146860 112990 146870
rect 116140 146860 116150 146940
rect 116920 146930 117000 146940
rect 117000 146870 117010 146930
rect 91500 146690 91560 146810
rect 100860 146800 100940 146810
rect 100940 146720 100950 146800
rect 101080 146799 101160 146809
rect 101400 146799 101480 146809
rect 101820 146799 101900 146809
rect 102140 146799 102220 146809
rect 101160 146719 101170 146799
rect 101480 146719 101490 146799
rect 101900 146719 101910 146799
rect 102220 146719 102230 146799
rect 103990 146780 104000 146860
rect 104170 146780 104180 146860
rect 104350 146780 104360 146860
rect 104530 146780 104540 146860
rect 104710 146780 104720 146860
rect 104890 146780 104900 146860
rect 105070 146780 105080 146860
rect 105250 146780 105260 146860
rect 105430 146780 105440 146860
rect 105610 146780 105620 146860
rect 105790 146780 105800 146860
rect 105970 146780 105980 146860
rect 106150 146780 106160 146860
rect 106330 146780 106340 146860
rect 106510 146780 106520 146860
rect 106690 146780 106700 146860
rect 106870 146780 106880 146860
rect 107050 146780 107060 146860
rect 107230 146780 107240 146860
rect 107410 146780 107420 146860
rect 107590 146780 107600 146860
rect 107770 146780 107780 146860
rect 107950 146780 107960 146860
rect 108130 146780 108140 146860
rect 108310 146780 108320 146860
rect 108490 146780 108500 146860
rect 108670 146780 108680 146860
rect 108850 146780 108860 146860
rect 109030 146780 109040 146860
rect 109210 146780 109220 146860
rect 109390 146780 109400 146860
rect 109570 146780 109580 146860
rect 109750 146780 109760 146860
rect 109930 146780 109940 146860
rect 110110 146780 110120 146860
rect 110290 146780 110300 146860
rect 110470 146780 110480 146860
rect 110650 146780 110660 146860
rect 110830 146780 110840 146860
rect 111010 146780 111020 146860
rect 111190 146780 111200 146860
rect 111370 146780 111380 146860
rect 111550 146780 111560 146860
rect 111730 146780 111740 146860
rect 111910 146780 111920 146860
rect 112090 146780 112100 146860
rect 112270 146780 112280 146860
rect 112450 146780 112460 146860
rect 112630 146780 112640 146860
rect 112810 146780 112820 146860
rect 112990 146780 113000 146860
rect 116900 146810 117020 146870
rect 114580 146799 114660 146809
rect 114900 146799 114980 146809
rect 115320 146799 115400 146809
rect 115640 146799 115720 146809
rect 116060 146800 116140 146810
rect 114660 146719 114670 146799
rect 114980 146719 114990 146799
rect 115400 146719 115410 146799
rect 115720 146719 115730 146799
rect 116140 146720 116150 146800
rect 116920 146790 117000 146800
rect 117000 146710 117010 146790
rect 117020 146690 117080 146810
rect 103910 146680 103990 146690
rect 104090 146680 104170 146690
rect 104270 146680 104350 146690
rect 104450 146680 104530 146690
rect 104630 146680 104710 146690
rect 104810 146680 104890 146690
rect 104990 146680 105070 146690
rect 105170 146680 105250 146690
rect 105350 146680 105430 146690
rect 105530 146680 105610 146690
rect 105710 146680 105790 146690
rect 105890 146680 105970 146690
rect 106070 146680 106150 146690
rect 106250 146680 106330 146690
rect 106430 146680 106510 146690
rect 106610 146680 106690 146690
rect 106790 146680 106870 146690
rect 106970 146680 107050 146690
rect 107150 146680 107230 146690
rect 107330 146680 107410 146690
rect 107510 146680 107590 146690
rect 107690 146680 107770 146690
rect 107870 146680 107950 146690
rect 108050 146680 108130 146690
rect 108230 146680 108310 146690
rect 108410 146680 108490 146690
rect 108590 146680 108670 146690
rect 108770 146680 108850 146690
rect 108950 146680 109030 146690
rect 109130 146680 109210 146690
rect 109310 146680 109390 146690
rect 109490 146680 109570 146690
rect 109670 146680 109750 146690
rect 109850 146680 109930 146690
rect 110030 146680 110110 146690
rect 110210 146680 110290 146690
rect 110390 146680 110470 146690
rect 110570 146680 110650 146690
rect 110750 146680 110830 146690
rect 110930 146680 111010 146690
rect 111110 146680 111190 146690
rect 111290 146680 111370 146690
rect 111470 146680 111550 146690
rect 111650 146680 111730 146690
rect 111830 146680 111910 146690
rect 112010 146680 112090 146690
rect 112190 146680 112270 146690
rect 112370 146680 112450 146690
rect 112550 146680 112630 146690
rect 112730 146680 112810 146690
rect 112910 146680 112990 146690
rect 100860 146660 100940 146670
rect 91400 146650 91480 146660
rect 91480 146570 91490 146650
rect 100940 146580 100950 146660
rect 101240 146639 101320 146649
rect 101560 146639 101640 146649
rect 101980 146639 102060 146649
rect 102300 146639 102380 146649
rect 101320 146559 101330 146639
rect 101640 146559 101650 146639
rect 102060 146559 102070 146639
rect 102380 146559 102390 146639
rect 103990 146600 104000 146680
rect 104170 146600 104180 146680
rect 104350 146600 104360 146680
rect 104530 146600 104540 146680
rect 104710 146600 104720 146680
rect 104890 146600 104900 146680
rect 105070 146600 105080 146680
rect 105250 146600 105260 146680
rect 105430 146600 105440 146680
rect 105610 146600 105620 146680
rect 105790 146600 105800 146680
rect 105970 146600 105980 146680
rect 106150 146600 106160 146680
rect 106330 146600 106340 146680
rect 106510 146600 106520 146680
rect 106690 146600 106700 146680
rect 106870 146600 106880 146680
rect 107050 146600 107060 146680
rect 107230 146600 107240 146680
rect 107410 146600 107420 146680
rect 107590 146600 107600 146680
rect 107770 146600 107780 146680
rect 107950 146600 107960 146680
rect 108130 146600 108140 146680
rect 108310 146600 108320 146680
rect 108490 146600 108500 146680
rect 108670 146600 108680 146680
rect 108850 146600 108860 146680
rect 109030 146600 109040 146680
rect 109210 146600 109220 146680
rect 109390 146600 109400 146680
rect 109570 146600 109580 146680
rect 109750 146600 109760 146680
rect 109930 146600 109940 146680
rect 110110 146600 110120 146680
rect 110290 146600 110300 146680
rect 110470 146600 110480 146680
rect 110650 146600 110660 146680
rect 110830 146600 110840 146680
rect 111010 146600 111020 146680
rect 111190 146600 111200 146680
rect 111370 146600 111380 146680
rect 111550 146600 111560 146680
rect 111730 146600 111740 146680
rect 111910 146600 111920 146680
rect 112090 146600 112100 146680
rect 112270 146600 112280 146680
rect 112450 146600 112460 146680
rect 112630 146600 112640 146680
rect 112810 146600 112820 146680
rect 112990 146600 113000 146680
rect 116060 146660 116140 146670
rect 114740 146639 114820 146649
rect 115060 146639 115140 146649
rect 115480 146639 115560 146649
rect 115800 146639 115880 146649
rect 114820 146559 114830 146639
rect 115140 146559 115150 146639
rect 115560 146559 115570 146639
rect 115880 146559 115890 146639
rect 116140 146580 116150 146660
rect 116920 146650 117000 146660
rect 117000 146570 117010 146650
rect 100860 146520 100940 146530
rect 116060 146520 116140 146530
rect 90085 146450 90135 146460
rect 90675 146450 90725 146460
rect 91265 146450 91315 146460
rect 100940 146440 100950 146520
rect 103910 146500 103990 146510
rect 104090 146500 104170 146510
rect 104270 146500 104350 146510
rect 104450 146500 104530 146510
rect 104630 146500 104710 146510
rect 104810 146500 104890 146510
rect 104990 146500 105070 146510
rect 105170 146500 105250 146510
rect 105350 146500 105430 146510
rect 105530 146500 105610 146510
rect 105710 146500 105790 146510
rect 105890 146500 105970 146510
rect 106070 146500 106150 146510
rect 106250 146500 106330 146510
rect 106430 146500 106510 146510
rect 106610 146500 106690 146510
rect 106790 146500 106870 146510
rect 106970 146500 107050 146510
rect 107150 146500 107230 146510
rect 107330 146500 107410 146510
rect 107510 146500 107590 146510
rect 107690 146500 107770 146510
rect 107870 146500 107950 146510
rect 108050 146500 108130 146510
rect 108230 146500 108310 146510
rect 108410 146500 108490 146510
rect 108590 146500 108670 146510
rect 108770 146500 108850 146510
rect 108950 146500 109030 146510
rect 109130 146500 109210 146510
rect 109310 146500 109390 146510
rect 109490 146500 109570 146510
rect 109670 146500 109750 146510
rect 109850 146500 109930 146510
rect 110030 146500 110110 146510
rect 110210 146500 110290 146510
rect 110390 146500 110470 146510
rect 110570 146500 110650 146510
rect 110750 146500 110830 146510
rect 110930 146500 111010 146510
rect 111110 146500 111190 146510
rect 111290 146500 111370 146510
rect 111470 146500 111550 146510
rect 111650 146500 111730 146510
rect 111830 146500 111910 146510
rect 112010 146500 112090 146510
rect 112190 146500 112270 146510
rect 112370 146500 112450 146510
rect 112550 146500 112630 146510
rect 112730 146500 112810 146510
rect 112910 146500 112990 146510
rect 101080 146479 101160 146489
rect 101400 146479 101480 146489
rect 101820 146479 101900 146489
rect 102140 146479 102220 146489
rect 101160 146399 101170 146479
rect 101480 146399 101490 146479
rect 101900 146399 101910 146479
rect 102220 146399 102230 146479
rect 103990 146420 104000 146500
rect 104170 146420 104180 146500
rect 104350 146420 104360 146500
rect 104530 146420 104540 146500
rect 104710 146420 104720 146500
rect 104890 146420 104900 146500
rect 105070 146420 105080 146500
rect 105250 146420 105260 146500
rect 105430 146420 105440 146500
rect 105610 146420 105620 146500
rect 105790 146420 105800 146500
rect 105970 146420 105980 146500
rect 106150 146420 106160 146500
rect 106330 146420 106340 146500
rect 106510 146420 106520 146500
rect 106690 146420 106700 146500
rect 106870 146420 106880 146500
rect 107050 146420 107060 146500
rect 107230 146420 107240 146500
rect 107410 146420 107420 146500
rect 107590 146420 107600 146500
rect 107770 146420 107780 146500
rect 107950 146420 107960 146500
rect 108130 146420 108140 146500
rect 108310 146420 108320 146500
rect 108490 146420 108500 146500
rect 108670 146420 108680 146500
rect 108850 146420 108860 146500
rect 109030 146420 109040 146500
rect 109210 146420 109220 146500
rect 109390 146420 109400 146500
rect 109570 146420 109580 146500
rect 109750 146420 109760 146500
rect 109930 146420 109940 146500
rect 110110 146420 110120 146500
rect 110290 146420 110300 146500
rect 110470 146420 110480 146500
rect 110650 146420 110660 146500
rect 110830 146420 110840 146500
rect 111010 146420 111020 146500
rect 111190 146420 111200 146500
rect 111370 146420 111380 146500
rect 111550 146420 111560 146500
rect 111730 146420 111740 146500
rect 111910 146420 111920 146500
rect 112090 146420 112100 146500
rect 112270 146420 112280 146500
rect 112450 146420 112460 146500
rect 112630 146420 112640 146500
rect 112810 146420 112820 146500
rect 112990 146420 113000 146500
rect 114580 146479 114660 146489
rect 114900 146479 114980 146489
rect 115320 146479 115400 146489
rect 115640 146479 115720 146489
rect 114660 146399 114670 146479
rect 114980 146399 114990 146479
rect 115400 146399 115410 146479
rect 115720 146399 115730 146479
rect 116140 146440 116150 146520
rect 117135 146460 117145 147200
rect 117150 146500 117160 147140
rect 117200 147090 117320 147150
rect 127940 147140 127950 147220
rect 128320 147199 128330 147279
rect 128640 147199 128650 147279
rect 129060 147199 129070 147279
rect 129380 147199 129390 147279
rect 129560 147220 129640 147230
rect 141360 147220 141440 147230
rect 129640 147140 129650 147220
rect 141440 147140 141450 147220
rect 141785 147200 141795 147280
rect 142105 147200 142115 147280
rect 145305 147200 145315 147280
rect 145625 147200 145635 147280
rect 145945 147200 145955 147280
rect 146220 147260 146300 147270
rect 146540 147260 146620 147270
rect 146860 147260 146940 147270
rect 147180 147260 147260 147270
rect 148780 147260 148860 147270
rect 149100 147260 149180 147270
rect 149420 147260 149500 147270
rect 149740 147260 149820 147270
rect 152300 147260 152380 147270
rect 152620 147260 152700 147270
rect 152940 147260 153020 147270
rect 153260 147260 153340 147270
rect 153580 147260 153660 147270
rect 153900 147260 153980 147270
rect 154220 147260 154300 147270
rect 154540 147260 154620 147270
rect 154860 147260 154940 147270
rect 155180 147260 155260 147270
rect 155500 147260 155580 147270
rect 155820 147260 155900 147270
rect 146300 147180 146310 147260
rect 146620 147180 146630 147260
rect 146940 147180 146950 147260
rect 147260 147180 147270 147260
rect 148860 147180 148870 147260
rect 149180 147180 149190 147260
rect 149500 147180 149510 147260
rect 149820 147180 149830 147260
rect 152380 147180 152390 147260
rect 152700 147180 152710 147260
rect 153020 147180 153030 147260
rect 153340 147180 153350 147260
rect 153660 147180 153670 147260
rect 153980 147180 153990 147260
rect 154300 147180 154310 147260
rect 154620 147180 154630 147260
rect 154940 147180 154950 147260
rect 155260 147180 155270 147260
rect 155580 147180 155590 147260
rect 155900 147180 155910 147260
rect 128080 147119 128160 147129
rect 128400 147119 128480 147129
rect 128820 147119 128900 147129
rect 129140 147119 129220 147129
rect 117320 146980 117380 147090
rect 127860 147080 127940 147090
rect 127940 147000 127950 147080
rect 128160 147039 128170 147119
rect 128480 147039 128490 147119
rect 128900 147039 128910 147119
rect 129220 147039 129230 147119
rect 130400 147090 130520 147140
rect 129560 147080 129640 147090
rect 129640 147000 129650 147080
rect 130420 147070 130500 147080
rect 130500 146990 130510 147070
rect 117200 146970 117380 146980
rect 130520 146970 130580 147090
rect 128240 146959 128320 146969
rect 128560 146959 128640 146969
rect 128980 146959 129060 146969
rect 129300 146959 129380 146969
rect 127860 146940 127940 146950
rect 117200 146810 117320 146870
rect 127940 146860 127950 146940
rect 128320 146879 128330 146959
rect 128640 146879 128650 146959
rect 129060 146879 129070 146959
rect 129380 146879 129390 146959
rect 129560 146940 129640 146950
rect 129640 146860 129650 146940
rect 130420 146930 130500 146940
rect 130500 146870 130510 146930
rect 130400 146810 130520 146870
rect 117320 146700 117380 146810
rect 127860 146800 127940 146810
rect 127940 146720 127950 146800
rect 128080 146799 128160 146809
rect 128400 146799 128480 146809
rect 128820 146799 128900 146809
rect 129140 146799 129220 146809
rect 129560 146800 129640 146810
rect 128160 146719 128170 146799
rect 128480 146719 128490 146799
rect 128900 146719 128910 146799
rect 129220 146719 129230 146799
rect 129640 146720 129650 146800
rect 130420 146790 130500 146800
rect 130500 146710 130510 146790
rect 117200 146690 117380 146700
rect 130520 146690 130580 146810
rect 127860 146660 127940 146670
rect 129560 146660 129640 146670
rect 127940 146580 127950 146660
rect 128240 146639 128320 146649
rect 128560 146639 128640 146649
rect 128980 146639 129060 146649
rect 129300 146639 129380 146649
rect 128320 146559 128330 146639
rect 128640 146559 128650 146639
rect 129060 146559 129070 146639
rect 129380 146559 129390 146639
rect 129640 146580 129650 146660
rect 130420 146650 130500 146660
rect 130500 146570 130510 146650
rect 127860 146520 127940 146530
rect 129560 146520 129640 146530
rect 117085 146450 117135 146460
rect 127940 146440 127950 146520
rect 128080 146479 128160 146489
rect 128400 146479 128480 146489
rect 128820 146479 128900 146489
rect 129140 146479 129220 146489
rect 128160 146399 128170 146479
rect 128480 146399 128490 146479
rect 128900 146399 128910 146479
rect 129220 146399 129230 146479
rect 129640 146440 129650 146520
rect 130635 146460 130645 147140
rect 130650 146500 130660 147140
rect 130700 147090 130820 147140
rect 141545 147120 141625 147130
rect 141865 147120 141945 147130
rect 142185 147120 142200 147130
rect 145385 147120 145465 147130
rect 145705 147120 145785 147130
rect 146025 147120 146105 147130
rect 130820 146980 130880 147090
rect 141360 147080 141440 147090
rect 141440 147000 141450 147080
rect 141625 147040 141635 147120
rect 141945 147040 141955 147120
rect 145465 147040 145475 147120
rect 145785 147040 145795 147120
rect 146105 147040 146115 147120
rect 146380 147100 146460 147110
rect 146700 147100 146780 147110
rect 147020 147100 147100 147110
rect 147340 147100 147420 147110
rect 148940 147100 149020 147110
rect 149260 147100 149340 147110
rect 149580 147100 149660 147110
rect 152460 147100 152540 147110
rect 152780 147100 152860 147110
rect 153100 147100 153180 147110
rect 153420 147100 153500 147110
rect 153740 147100 153820 147110
rect 154060 147100 154140 147110
rect 154380 147100 154460 147110
rect 154700 147100 154780 147110
rect 155020 147100 155100 147110
rect 155340 147100 155420 147110
rect 155660 147100 155740 147110
rect 155980 147100 156000 147110
rect 146460 147020 146470 147100
rect 146780 147020 146790 147100
rect 147100 147020 147110 147100
rect 147420 147020 147430 147100
rect 149020 147020 149030 147100
rect 149340 147020 149350 147100
rect 149660 147020 149670 147100
rect 152540 147020 152550 147100
rect 152860 147020 152870 147100
rect 153180 147020 153190 147100
rect 153500 147020 153510 147100
rect 153820 147020 153830 147100
rect 154140 147020 154150 147100
rect 154460 147020 154470 147100
rect 154780 147020 154790 147100
rect 155100 147020 155110 147100
rect 155420 147020 155430 147100
rect 155740 147020 155750 147100
rect 156060 147020 156070 147050
rect 156380 147020 156390 147050
rect 156700 147020 156710 147050
rect 157020 147020 157030 147050
rect 157340 147020 157350 147050
rect 157660 147020 157670 147050
rect 157980 147020 157990 147050
rect 158300 147020 158310 147050
rect 158620 147020 158630 147050
rect 158940 147020 158950 147050
rect 159260 147020 159270 147050
rect 159580 147020 159590 147050
rect 163740 147020 163750 147050
rect 164060 147020 164070 147050
rect 164380 147020 164390 147050
rect 164700 147020 164710 147050
rect 165020 147020 165030 147050
rect 165340 147020 165350 147050
rect 165660 147020 165670 147050
rect 165980 147020 165990 147050
rect 166300 147020 166310 147050
rect 166620 147020 166630 147050
rect 166940 147020 166950 147050
rect 167260 147020 167270 147050
rect 167580 147020 167590 147050
rect 167900 147020 167910 147050
rect 168220 147020 168230 147050
rect 168540 147020 168550 147050
rect 168860 147020 168870 147050
rect 169180 147020 169190 147050
rect 169500 147020 169510 147050
rect 169820 147020 169830 147050
rect 170140 147020 170150 147050
rect 170460 147020 170470 147050
rect 170780 147020 170790 147050
rect 130700 146970 130880 146980
rect 141705 146960 141785 146970
rect 142025 146960 142105 146970
rect 145225 146960 145305 146970
rect 145545 146960 145625 146970
rect 145865 146960 145945 146970
rect 141360 146940 141440 146950
rect 130700 146810 130820 146870
rect 141440 146860 141450 146940
rect 141785 146880 141795 146960
rect 142105 146880 142115 146960
rect 145305 146880 145315 146960
rect 145625 146880 145635 146960
rect 145945 146880 145955 146960
rect 146220 146940 146300 146950
rect 146540 146940 146620 146950
rect 146860 146940 146940 146950
rect 147180 146940 147260 146950
rect 147500 146940 147580 146950
rect 148780 146940 148860 146950
rect 149100 146940 149180 146950
rect 149420 146940 149500 146950
rect 149740 146940 149820 146950
rect 152300 146940 152380 146950
rect 152620 146940 152700 146950
rect 152940 146940 153020 146950
rect 153260 146940 153340 146950
rect 153580 146940 153660 146950
rect 153900 146940 153980 146950
rect 154220 146940 154300 146950
rect 154540 146940 154620 146950
rect 154860 146940 154940 146950
rect 155180 146940 155260 146950
rect 155500 146940 155580 146950
rect 155820 146940 155900 146950
rect 156140 146940 156220 146950
rect 156460 146940 156540 146950
rect 156780 146940 156860 146950
rect 157100 146940 157180 146950
rect 157420 146940 157500 146950
rect 157740 146940 157820 146950
rect 158060 146940 158140 146950
rect 158380 146940 158460 146950
rect 158700 146940 158780 146950
rect 159020 146940 159100 146950
rect 159340 146940 159420 146950
rect 163500 146940 163580 146950
rect 163820 146940 163900 146950
rect 164140 146940 164220 146950
rect 164460 146940 164540 146950
rect 164780 146940 164860 146950
rect 165100 146940 165180 146950
rect 165420 146940 165500 146950
rect 165740 146940 165820 146950
rect 166060 146940 166140 146950
rect 166380 146940 166460 146950
rect 166700 146940 166780 146950
rect 167020 146940 167100 146950
rect 167340 146940 167420 146950
rect 167660 146940 167740 146950
rect 167980 146940 168060 146950
rect 168300 146940 168380 146950
rect 168620 146940 168700 146950
rect 168940 146940 169020 146950
rect 169260 146940 169340 146950
rect 169580 146940 169660 146950
rect 169900 146940 169980 146950
rect 170220 146940 170300 146950
rect 170540 146940 170620 146950
rect 170860 146940 170940 146950
rect 146300 146860 146310 146940
rect 146620 146860 146630 146940
rect 146940 146860 146950 146940
rect 147260 146860 147270 146940
rect 147580 146860 147590 146940
rect 148860 146860 148870 146940
rect 149180 146860 149190 146940
rect 149500 146860 149510 146940
rect 149820 146860 149830 146940
rect 152380 146860 152390 146940
rect 152700 146860 152710 146940
rect 153020 146860 153030 146940
rect 153340 146860 153350 146940
rect 153660 146860 153670 146940
rect 153980 146860 153990 146940
rect 154300 146860 154310 146940
rect 154620 146860 154630 146940
rect 154940 146860 154950 146940
rect 155260 146860 155270 146940
rect 155580 146860 155590 146940
rect 155900 146860 155910 146940
rect 156220 146860 156230 146940
rect 156540 146860 156550 146940
rect 156860 146860 156870 146940
rect 157180 146860 157190 146940
rect 157500 146860 157510 146940
rect 157820 146860 157830 146940
rect 158140 146860 158150 146940
rect 158460 146860 158470 146940
rect 158780 146860 158790 146940
rect 159100 146860 159110 146940
rect 159420 146860 159430 146940
rect 163580 146860 163590 146940
rect 163900 146860 163910 146940
rect 164220 146860 164230 146940
rect 164540 146860 164550 146940
rect 164860 146860 164870 146940
rect 165180 146860 165190 146940
rect 165500 146860 165510 146940
rect 165820 146860 165830 146940
rect 166140 146860 166150 146940
rect 166460 146860 166470 146940
rect 166780 146860 166790 146940
rect 167100 146860 167110 146940
rect 167420 146860 167430 146940
rect 167740 146860 167750 146940
rect 168060 146860 168070 146940
rect 168380 146860 168390 146940
rect 168700 146860 168710 146940
rect 169020 146860 169030 146940
rect 169340 146860 169350 146940
rect 169660 146860 169670 146940
rect 169980 146860 169990 146940
rect 170300 146860 170310 146940
rect 170620 146860 170630 146940
rect 170940 146860 170950 146940
rect 130820 146700 130880 146810
rect 141360 146800 141440 146810
rect 141545 146800 141625 146810
rect 141865 146800 141945 146810
rect 142185 146800 142200 146810
rect 145385 146800 145465 146810
rect 145705 146800 145785 146810
rect 146025 146800 146105 146810
rect 141440 146720 141450 146800
rect 141625 146720 141635 146800
rect 141945 146720 141955 146800
rect 145465 146720 145475 146800
rect 145785 146720 145795 146800
rect 146105 146720 146115 146800
rect 146380 146780 146460 146790
rect 146700 146780 146780 146790
rect 147020 146780 147100 146790
rect 147340 146780 147420 146790
rect 148940 146780 149020 146790
rect 149260 146780 149340 146790
rect 149580 146780 149660 146790
rect 152460 146780 152540 146790
rect 152780 146780 152860 146790
rect 153100 146780 153180 146790
rect 153420 146780 153500 146790
rect 153740 146780 153820 146790
rect 154060 146780 154140 146790
rect 154380 146780 154460 146790
rect 154700 146780 154780 146790
rect 155020 146780 155100 146790
rect 155340 146780 155420 146790
rect 155660 146780 155740 146790
rect 155980 146780 156060 146790
rect 156300 146780 156380 146790
rect 156620 146780 156700 146790
rect 156940 146780 157020 146790
rect 157260 146780 157340 146790
rect 157580 146780 157660 146790
rect 157900 146780 157980 146790
rect 158220 146780 158300 146790
rect 158540 146780 158620 146790
rect 158860 146780 158940 146790
rect 159180 146780 159260 146790
rect 159500 146780 159580 146790
rect 163660 146780 163740 146790
rect 163980 146780 164060 146790
rect 164300 146780 164380 146790
rect 164620 146780 164700 146790
rect 164940 146780 165020 146790
rect 165260 146780 165340 146790
rect 165580 146780 165660 146790
rect 165900 146780 165980 146790
rect 166220 146780 166300 146790
rect 166540 146780 166620 146790
rect 166860 146780 166940 146790
rect 167180 146780 167260 146790
rect 167500 146780 167580 146790
rect 167820 146780 167900 146790
rect 168140 146780 168220 146790
rect 168460 146780 168540 146790
rect 168780 146780 168860 146790
rect 169100 146780 169180 146790
rect 169420 146780 169500 146790
rect 169740 146780 169820 146790
rect 170060 146780 170140 146790
rect 170380 146780 170460 146790
rect 170700 146780 170780 146790
rect 146460 146700 146470 146780
rect 146780 146700 146790 146780
rect 147100 146700 147110 146780
rect 147420 146700 147430 146780
rect 149020 146700 149030 146780
rect 149340 146700 149350 146780
rect 149660 146700 149670 146780
rect 152540 146700 152550 146780
rect 152860 146700 152870 146780
rect 153180 146700 153190 146780
rect 153500 146700 153510 146780
rect 153820 146700 153830 146780
rect 154140 146700 154150 146780
rect 154460 146700 154470 146780
rect 154780 146700 154790 146780
rect 155100 146700 155110 146780
rect 155420 146700 155430 146780
rect 155740 146700 155750 146780
rect 156060 146700 156070 146780
rect 156380 146700 156390 146780
rect 156700 146700 156710 146780
rect 157020 146700 157030 146780
rect 157340 146700 157350 146780
rect 157660 146700 157670 146780
rect 157980 146700 157990 146780
rect 158300 146700 158310 146780
rect 158620 146700 158630 146780
rect 158940 146700 158950 146780
rect 159260 146700 159270 146780
rect 159580 146700 159590 146780
rect 163740 146700 163750 146780
rect 164060 146700 164070 146780
rect 164380 146700 164390 146780
rect 164700 146700 164710 146780
rect 165020 146700 165030 146780
rect 165340 146700 165350 146780
rect 165660 146700 165670 146780
rect 165980 146700 165990 146780
rect 166300 146700 166310 146780
rect 166620 146700 166630 146780
rect 166940 146700 166950 146780
rect 167260 146700 167270 146780
rect 167580 146700 167590 146780
rect 167900 146700 167910 146780
rect 168220 146700 168230 146780
rect 168540 146700 168550 146780
rect 168860 146700 168870 146780
rect 169180 146700 169190 146780
rect 169500 146700 169510 146780
rect 169820 146700 169830 146780
rect 170140 146700 170150 146780
rect 170460 146700 170470 146780
rect 170780 146700 170790 146780
rect 130700 146690 130880 146700
rect 141360 146660 141440 146670
rect 141440 146580 141450 146660
rect 141705 146640 141785 146650
rect 142025 146640 142105 146650
rect 145225 146640 145305 146650
rect 145545 146640 145625 146650
rect 145865 146640 145945 146650
rect 141785 146560 141795 146640
rect 142105 146560 142115 146640
rect 145305 146560 145315 146640
rect 145625 146560 145635 146640
rect 145945 146560 145955 146640
rect 146220 146620 146300 146630
rect 146540 146620 146620 146630
rect 146860 146620 146940 146630
rect 147180 146620 147260 146630
rect 147500 146620 147580 146630
rect 148780 146620 148860 146630
rect 149100 146620 149180 146630
rect 149420 146620 149500 146630
rect 149740 146620 149820 146630
rect 152300 146620 152380 146630
rect 152620 146620 152700 146630
rect 152940 146620 153020 146630
rect 153260 146620 153340 146630
rect 153580 146620 153660 146630
rect 153900 146620 153980 146630
rect 154220 146620 154300 146630
rect 154540 146620 154620 146630
rect 154860 146620 154940 146630
rect 155180 146620 155260 146630
rect 155500 146620 155580 146630
rect 155820 146620 155900 146630
rect 156140 146620 156220 146630
rect 156460 146620 156540 146630
rect 156780 146620 156860 146630
rect 157100 146620 157180 146630
rect 157420 146620 157500 146630
rect 157740 146620 157820 146630
rect 158060 146620 158140 146630
rect 158380 146620 158460 146630
rect 158700 146620 158780 146630
rect 159020 146620 159100 146630
rect 159340 146620 159420 146630
rect 163500 146620 163580 146630
rect 163820 146620 163900 146630
rect 164140 146620 164220 146630
rect 164460 146620 164540 146630
rect 164780 146620 164860 146630
rect 165100 146620 165180 146630
rect 165420 146620 165500 146630
rect 165740 146620 165820 146630
rect 166060 146620 166140 146630
rect 166380 146620 166460 146630
rect 166700 146620 166780 146630
rect 167020 146620 167100 146630
rect 167340 146620 167420 146630
rect 167660 146620 167740 146630
rect 167980 146620 168060 146630
rect 168300 146620 168380 146630
rect 168620 146620 168700 146630
rect 168940 146620 169020 146630
rect 169260 146620 169340 146630
rect 169580 146620 169660 146630
rect 169900 146620 169980 146630
rect 170220 146620 170300 146630
rect 170540 146620 170620 146630
rect 170860 146620 170940 146630
rect 146300 146540 146310 146620
rect 146620 146540 146630 146620
rect 146940 146540 146950 146620
rect 147260 146540 147270 146620
rect 147580 146540 147590 146620
rect 148860 146540 148870 146620
rect 149180 146540 149190 146620
rect 149500 146540 149510 146620
rect 149820 146540 149830 146620
rect 152380 146540 152390 146620
rect 152700 146540 152710 146620
rect 153020 146540 153030 146620
rect 153340 146540 153350 146620
rect 153660 146540 153670 146620
rect 153980 146540 153990 146620
rect 154300 146540 154310 146620
rect 154620 146540 154630 146620
rect 154940 146540 154950 146620
rect 155260 146540 155270 146620
rect 155580 146540 155590 146620
rect 155900 146540 155910 146620
rect 156220 146540 156230 146620
rect 156540 146540 156550 146620
rect 156860 146540 156870 146620
rect 157180 146540 157190 146620
rect 157500 146540 157510 146620
rect 157820 146540 157830 146620
rect 158140 146540 158150 146620
rect 158460 146540 158470 146620
rect 158780 146540 158790 146620
rect 159100 146540 159110 146620
rect 159420 146540 159430 146620
rect 163580 146540 163590 146620
rect 163900 146540 163910 146620
rect 164220 146540 164230 146620
rect 164540 146540 164550 146620
rect 164860 146540 164870 146620
rect 165180 146540 165190 146620
rect 165500 146540 165510 146620
rect 165820 146540 165830 146620
rect 166140 146540 166150 146620
rect 166460 146540 166470 146620
rect 166780 146540 166790 146620
rect 167100 146540 167110 146620
rect 167420 146540 167430 146620
rect 167740 146540 167750 146620
rect 168060 146540 168070 146620
rect 168380 146540 168390 146620
rect 168700 146540 168710 146620
rect 169020 146540 169030 146620
rect 169340 146540 169350 146620
rect 169660 146540 169670 146620
rect 169980 146540 169990 146620
rect 170300 146540 170310 146620
rect 170620 146540 170630 146620
rect 170940 146540 170950 146620
rect 141360 146520 141440 146530
rect 130585 146450 130635 146460
rect 141440 146440 141450 146520
rect 141545 146480 141625 146490
rect 141865 146480 141945 146490
rect 142185 146480 142200 146490
rect 145385 146480 145465 146490
rect 145705 146480 145785 146490
rect 146025 146480 146105 146490
rect 141625 146400 141635 146480
rect 141945 146400 141955 146480
rect 145465 146400 145475 146480
rect 145785 146400 145795 146480
rect 146105 146400 146115 146480
rect 146380 146460 146460 146470
rect 146700 146460 146780 146470
rect 147020 146460 147100 146470
rect 147340 146460 147420 146470
rect 48500 146380 48640 146390
rect 60360 146380 60440 146390
rect 62060 146380 62140 146390
rect 73860 146380 73940 146390
rect 75560 146380 75640 146390
rect 87360 146380 87440 146390
rect 89060 146380 89140 146390
rect 100860 146380 100940 146390
rect 116060 146380 116140 146390
rect 127860 146380 127940 146390
rect 129560 146380 129640 146390
rect 141360 146380 141440 146390
rect 146460 146380 146470 146460
rect 146780 146380 146790 146460
rect 147100 146380 147110 146460
rect 147420 146380 147430 146460
rect 42420 146300 42500 146310
rect 42740 146300 42820 146310
rect 43060 146300 43140 146310
rect 43380 146300 43460 146310
rect 43700 146300 43780 146310
rect 30360 146215 30440 146225
rect 30680 146215 30760 146225
rect 31000 146215 31080 146225
rect 31320 146215 31400 146225
rect 31640 146215 31720 146225
rect 31960 146215 32040 146225
rect 32280 146215 32360 146225
rect 32600 146215 32680 146225
rect 32920 146215 33000 146225
rect 33240 146215 33320 146225
rect 33560 146215 33640 146225
rect 33880 146215 33960 146225
rect 34200 146215 34280 146225
rect 34520 146215 34600 146225
rect 34840 146215 34920 146225
rect 35160 146215 35240 146225
rect 35480 146215 35560 146225
rect 35800 146215 35880 146225
rect 36120 146215 36200 146225
rect 36440 146215 36520 146225
rect 36760 146215 36840 146225
rect 37080 146215 37160 146225
rect 37400 146215 37480 146225
rect 37720 146215 37800 146225
rect 40180 146215 40260 146225
rect 40500 146215 40580 146225
rect 40820 146215 40900 146225
rect 41140 146215 41220 146225
rect 42470 146220 42510 146300
rect 42560 146215 42640 146225
rect 42790 146220 42830 146300
rect 42880 146215 42960 146225
rect 43110 146220 43150 146300
rect 43200 146215 43280 146225
rect 43430 146220 43470 146300
rect 43520 146215 43600 146225
rect 43780 146220 43790 146300
rect 30440 146135 30450 146215
rect 30760 146135 30770 146215
rect 31080 146135 31090 146215
rect 31400 146135 31410 146215
rect 31720 146135 31730 146215
rect 32040 146135 32050 146215
rect 32360 146135 32370 146215
rect 32680 146135 32690 146215
rect 33000 146135 33010 146215
rect 33320 146135 33330 146215
rect 33640 146135 33650 146215
rect 33960 146135 33970 146215
rect 34280 146135 34290 146215
rect 34600 146135 34610 146215
rect 34920 146135 34930 146215
rect 35240 146135 35250 146215
rect 35560 146135 35570 146215
rect 35880 146135 35890 146215
rect 36200 146135 36210 146215
rect 36520 146135 36530 146215
rect 36840 146135 36850 146215
rect 37160 146135 37170 146215
rect 37480 146135 37490 146215
rect 37800 146135 37810 146215
rect 40260 146135 40270 146215
rect 40580 146135 40590 146215
rect 40900 146135 40910 146215
rect 41220 146135 41230 146215
rect 42640 146135 42650 146215
rect 42960 146135 42970 146215
rect 43280 146135 43290 146215
rect 43600 146135 43610 146215
rect 19130 146095 19210 146105
rect 19450 146095 19530 146105
rect 19770 146095 19850 146105
rect 20090 146095 20170 146105
rect 20410 146095 20490 146105
rect 20730 146095 20810 146105
rect 21050 146095 21130 146105
rect 21370 146095 21450 146105
rect 21690 146095 21770 146105
rect 22010 146095 22090 146105
rect 22330 146095 22410 146105
rect 22650 146095 22730 146105
rect 22970 146095 23050 146105
rect 23290 146095 23370 146105
rect 23610 146095 23690 146105
rect 23930 146095 24010 146105
rect 24250 146095 24330 146105
rect 24570 146095 24650 146105
rect 24890 146095 24970 146105
rect 25210 146095 25290 146105
rect 25530 146095 25610 146105
rect 25850 146095 25930 146105
rect 26170 146095 26250 146105
rect 19210 146015 19220 146095
rect 19530 146015 19540 146095
rect 19850 146015 19860 146095
rect 20170 146015 20180 146095
rect 20490 146015 20500 146095
rect 20810 146015 20820 146095
rect 21130 146015 21140 146095
rect 21450 146015 21460 146095
rect 21770 146015 21780 146095
rect 22090 146015 22100 146095
rect 22410 146015 22420 146095
rect 22730 146015 22740 146095
rect 23050 146015 23060 146095
rect 23370 146015 23380 146095
rect 23690 146015 23700 146095
rect 24010 146015 24020 146095
rect 24330 146015 24340 146095
rect 24650 146015 24660 146095
rect 24970 146015 24980 146095
rect 25290 146015 25300 146095
rect 25610 146015 25620 146095
rect 25930 146015 25940 146095
rect 26250 146015 26260 146095
rect 30520 146055 30600 146065
rect 30840 146055 30920 146065
rect 31160 146055 31240 146065
rect 31480 146055 31560 146065
rect 31800 146055 31880 146065
rect 32120 146055 32200 146065
rect 32440 146055 32520 146065
rect 32760 146055 32840 146065
rect 33080 146055 33160 146065
rect 33400 146055 33480 146065
rect 33720 146055 33800 146065
rect 34040 146055 34120 146065
rect 34360 146055 34440 146065
rect 34680 146055 34760 146065
rect 35000 146055 35080 146065
rect 35320 146055 35400 146065
rect 35640 146055 35720 146065
rect 35960 146055 36040 146065
rect 36280 146055 36360 146065
rect 36600 146055 36680 146065
rect 36920 146055 37000 146065
rect 37240 146055 37320 146065
rect 37560 146055 37640 146065
rect 40340 146055 40420 146065
rect 40660 146055 40740 146065
rect 40980 146055 41060 146065
rect 42720 146055 42800 146065
rect 43040 146055 43120 146065
rect 43360 146055 43440 146065
rect 30600 145975 30610 146055
rect 30920 145975 30930 146055
rect 31240 145975 31250 146055
rect 31560 145975 31570 146055
rect 31880 145975 31890 146055
rect 32200 145975 32210 146055
rect 32520 145975 32530 146055
rect 32840 145975 32850 146055
rect 33160 145975 33170 146055
rect 33480 145975 33490 146055
rect 33800 145975 33810 146055
rect 34120 145975 34130 146055
rect 34440 145975 34450 146055
rect 34760 145975 34770 146055
rect 35080 145975 35090 146055
rect 35400 145975 35410 146055
rect 35720 145975 35730 146055
rect 36040 145975 36050 146055
rect 36360 145975 36370 146055
rect 36680 145975 36690 146055
rect 37000 145975 37010 146055
rect 37320 145975 37330 146055
rect 37640 145975 37650 146055
rect 40420 145975 40430 146055
rect 40740 145975 40750 146055
rect 41060 145975 41070 146055
rect 42800 145975 42810 146055
rect 43120 145975 43130 146055
rect 43440 145975 43450 146055
rect 48500 146040 48605 146380
rect 48640 146300 48650 146380
rect 49650 146300 51040 146310
rect 60440 146300 60450 146380
rect 62140 146300 62150 146380
rect 63150 146300 64540 146310
rect 73940 146300 73950 146380
rect 75640 146300 75650 146380
rect 76650 146300 78040 146310
rect 87440 146300 87450 146380
rect 89140 146300 89150 146380
rect 90150 146300 91540 146310
rect 100940 146300 100950 146380
rect 103910 146320 103990 146330
rect 104090 146320 104170 146330
rect 104270 146320 104350 146330
rect 104450 146320 104530 146330
rect 104630 146320 104710 146330
rect 104810 146320 104890 146330
rect 104990 146320 105070 146330
rect 105170 146320 105250 146330
rect 105350 146320 105430 146330
rect 105530 146320 105610 146330
rect 105710 146320 105790 146330
rect 105890 146320 105970 146330
rect 106070 146320 106150 146330
rect 106250 146320 106330 146330
rect 106430 146320 106510 146330
rect 106610 146320 106690 146330
rect 106790 146320 106870 146330
rect 106970 146320 107050 146330
rect 107150 146320 107230 146330
rect 107330 146320 107410 146330
rect 107510 146320 107590 146330
rect 107690 146320 107770 146330
rect 107870 146320 107950 146330
rect 108050 146320 108130 146330
rect 108230 146320 108310 146330
rect 108410 146320 108490 146330
rect 108590 146320 108670 146330
rect 108770 146320 108850 146330
rect 108950 146320 109030 146330
rect 109130 146320 109210 146330
rect 109310 146320 109390 146330
rect 109490 146320 109570 146330
rect 109670 146320 109750 146330
rect 109850 146320 109930 146330
rect 110030 146320 110110 146330
rect 110210 146320 110290 146330
rect 110390 146320 110470 146330
rect 110570 146320 110650 146330
rect 110750 146320 110830 146330
rect 110930 146320 111010 146330
rect 111110 146320 111190 146330
rect 111290 146320 111370 146330
rect 111470 146320 111550 146330
rect 111650 146320 111730 146330
rect 111830 146320 111910 146330
rect 112010 146320 112090 146330
rect 112190 146320 112270 146330
rect 112370 146320 112450 146330
rect 112550 146320 112630 146330
rect 112730 146320 112810 146330
rect 112910 146320 112990 146330
rect 103990 146240 104000 146320
rect 104170 146240 104180 146320
rect 104350 146240 104360 146320
rect 104530 146240 104540 146320
rect 104710 146240 104720 146320
rect 104890 146240 104900 146320
rect 105070 146240 105080 146320
rect 105250 146240 105260 146320
rect 105430 146240 105440 146320
rect 105610 146240 105620 146320
rect 105790 146240 105800 146320
rect 105970 146240 105980 146320
rect 106150 146240 106160 146320
rect 106330 146240 106340 146320
rect 106510 146240 106520 146320
rect 106690 146240 106700 146320
rect 106870 146240 106880 146320
rect 107050 146240 107060 146320
rect 107230 146240 107240 146320
rect 107410 146240 107420 146320
rect 107590 146240 107600 146320
rect 107770 146240 107780 146320
rect 107950 146240 107960 146320
rect 108130 146240 108140 146320
rect 108310 146240 108320 146320
rect 108490 146240 108500 146320
rect 108670 146240 108680 146320
rect 108850 146240 108860 146320
rect 109030 146240 109040 146320
rect 109210 146240 109220 146320
rect 109390 146240 109400 146320
rect 109570 146240 109580 146320
rect 109750 146240 109760 146320
rect 109930 146240 109940 146320
rect 110110 146240 110120 146320
rect 110290 146240 110300 146320
rect 110470 146240 110480 146320
rect 110650 146240 110660 146320
rect 110830 146240 110840 146320
rect 111010 146240 111020 146320
rect 111190 146240 111200 146320
rect 111370 146240 111380 146320
rect 111550 146240 111560 146320
rect 111730 146240 111740 146320
rect 111910 146240 111920 146320
rect 112090 146240 112100 146320
rect 112270 146240 112280 146320
rect 112450 146240 112460 146320
rect 112630 146240 112640 146320
rect 112810 146240 112820 146320
rect 112990 146240 113000 146320
rect 116140 146300 116150 146380
rect 117150 146300 117420 146310
rect 127940 146300 127950 146380
rect 129640 146300 129650 146380
rect 130650 146300 130920 146310
rect 141440 146300 141450 146380
rect 146220 146300 146300 146310
rect 146540 146300 146620 146310
rect 146860 146300 146940 146310
rect 147180 146300 147260 146310
rect 147500 146300 147580 146310
rect 146300 146220 146310 146300
rect 146400 146215 146480 146225
rect 146540 146220 146570 146300
rect 146620 146220 146630 146300
rect 146720 146215 146800 146225
rect 146860 146220 146890 146300
rect 146940 146220 146950 146300
rect 147040 146215 147120 146225
rect 147180 146220 147210 146300
rect 147260 146220 147270 146300
rect 147360 146215 147440 146225
rect 147500 146220 147530 146300
rect 147580 146220 147590 146300
rect 148780 146215 148860 146225
rect 149100 146215 149180 146225
rect 149420 146215 149500 146225
rect 149740 146215 149820 146225
rect 152200 146215 152280 146225
rect 152520 146215 152600 146225
rect 152840 146215 152920 146225
rect 153160 146215 153240 146225
rect 153480 146215 153560 146225
rect 153800 146215 153880 146225
rect 154120 146215 154200 146225
rect 154440 146215 154520 146225
rect 154760 146215 154840 146225
rect 155080 146215 155160 146225
rect 155400 146215 155480 146225
rect 155720 146215 155800 146225
rect 156040 146215 156120 146225
rect 156360 146215 156440 146225
rect 156680 146215 156760 146225
rect 157000 146215 157080 146225
rect 157320 146215 157400 146225
rect 157640 146215 157720 146225
rect 157960 146215 158040 146225
rect 158280 146215 158360 146225
rect 158600 146215 158680 146225
rect 158920 146215 159000 146225
rect 159240 146215 159320 146225
rect 159560 146215 159640 146225
rect 48870 146100 48900 146160
rect 48990 146100 49020 146160
rect 49110 146100 49140 146160
rect 49230 146100 49260 146160
rect 49350 146100 49380 146160
rect 49470 146100 49500 146160
rect 49590 146100 49620 146160
rect 49710 146100 49740 146160
rect 49830 146100 49860 146160
rect 49950 146100 49980 146160
rect 50070 146100 50100 146160
rect 50190 146100 50220 146160
rect 50310 146100 50340 146160
rect 50430 146100 50460 146160
rect 50550 146100 50580 146160
rect 50670 146100 50700 146160
rect 50790 146100 50820 146160
rect 50910 146100 50940 146160
rect 51030 146100 51060 146160
rect 51150 146100 51180 146160
rect 51270 146100 51300 146160
rect 51390 146100 51420 146160
rect 51510 146100 51540 146160
rect 51630 146100 51660 146160
rect 51750 146100 51780 146160
rect 51870 146100 51900 146160
rect 51990 146100 52020 146160
rect 52110 146100 52140 146160
rect 52230 146100 52260 146160
rect 52350 146100 52380 146160
rect 52470 146100 52500 146160
rect 52590 146100 52620 146160
rect 52710 146100 52740 146160
rect 52830 146100 52860 146160
rect 52950 146100 52980 146160
rect 53070 146100 53100 146160
rect 53190 146100 53220 146160
rect 53310 146100 53340 146160
rect 53430 146100 53460 146160
rect 53550 146100 53580 146160
rect 53670 146100 53700 146160
rect 53790 146100 53820 146160
rect 53910 146100 53940 146160
rect 54030 146100 54060 146160
rect 54150 146100 54180 146160
rect 54270 146100 54300 146160
rect 54390 146100 54420 146160
rect 54510 146100 54540 146160
rect 54630 146100 54660 146160
rect 54750 146100 54780 146160
rect 54870 146100 54900 146160
rect 54990 146100 55020 146160
rect 55110 146100 55140 146160
rect 55230 146100 55260 146160
rect 55350 146100 55380 146160
rect 55470 146100 55500 146160
rect 55590 146100 55620 146160
rect 55710 146100 55740 146160
rect 55830 146100 55860 146160
rect 55950 146100 55980 146160
rect 56070 146100 56100 146160
rect 56190 146100 56220 146160
rect 56310 146100 56340 146160
rect 56430 146100 56460 146160
rect 56550 146100 56580 146160
rect 56670 146100 56700 146160
rect 56790 146100 56820 146160
rect 56910 146100 56940 146160
rect 57030 146100 57060 146160
rect 57150 146100 57180 146160
rect 57270 146100 57300 146160
rect 57390 146100 57420 146160
rect 57510 146100 57540 146160
rect 57630 146100 57660 146160
rect 57750 146100 57780 146160
rect 57870 146100 57900 146160
rect 57990 146100 58020 146160
rect 58110 146100 58140 146160
rect 58230 146100 58260 146160
rect 58350 146100 58380 146160
rect 58470 146100 58500 146160
rect 58590 146100 58620 146160
rect 58710 146100 58740 146160
rect 58830 146100 58860 146160
rect 58950 146100 58980 146160
rect 59070 146100 59100 146160
rect 59190 146100 59220 146160
rect 59310 146100 59340 146160
rect 59430 146100 59460 146160
rect 59550 146100 59580 146160
rect 59670 146100 59700 146160
rect 59790 146100 59820 146160
rect 59910 146100 59940 146160
rect 60030 146100 60060 146160
rect 60150 146100 60180 146160
rect 62370 146100 62400 146160
rect 62490 146100 62520 146160
rect 62610 146100 62640 146160
rect 62730 146100 62760 146160
rect 62850 146100 62880 146160
rect 62970 146100 63000 146160
rect 63090 146100 63120 146160
rect 63210 146100 63240 146160
rect 63330 146100 63360 146160
rect 63450 146100 63480 146160
rect 63570 146100 63600 146160
rect 63690 146100 63720 146160
rect 63810 146100 63840 146160
rect 63930 146100 63960 146160
rect 64050 146100 64080 146160
rect 64170 146100 64200 146160
rect 64290 146100 64320 146160
rect 64410 146100 64440 146160
rect 64530 146100 64560 146160
rect 64650 146100 64680 146160
rect 64770 146100 64800 146160
rect 64890 146100 64920 146160
rect 65010 146100 65040 146160
rect 65130 146100 65160 146160
rect 65250 146100 65280 146160
rect 65370 146100 65400 146160
rect 65490 146100 65520 146160
rect 65610 146100 65640 146160
rect 65730 146100 65760 146160
rect 65850 146100 65880 146160
rect 65970 146100 66000 146160
rect 66090 146100 66120 146160
rect 66210 146100 66240 146160
rect 66330 146100 66360 146160
rect 66450 146100 66480 146160
rect 66570 146100 66600 146160
rect 66690 146100 66720 146160
rect 66810 146100 66840 146160
rect 66930 146100 66960 146160
rect 67050 146100 67080 146160
rect 67170 146100 67200 146160
rect 67290 146100 67320 146160
rect 67410 146100 67440 146160
rect 67530 146100 67560 146160
rect 67650 146100 67680 146160
rect 67770 146100 67800 146160
rect 67890 146100 67920 146160
rect 68010 146100 68040 146160
rect 68130 146100 68160 146160
rect 68250 146100 68280 146160
rect 68370 146100 68400 146160
rect 68490 146100 68520 146160
rect 68610 146100 68640 146160
rect 68730 146100 68760 146160
rect 68850 146100 68880 146160
rect 68970 146100 69000 146160
rect 69090 146100 69120 146160
rect 69210 146100 69240 146160
rect 69330 146100 69360 146160
rect 69450 146100 69480 146160
rect 69570 146100 69600 146160
rect 69690 146100 69720 146160
rect 69810 146100 69840 146160
rect 69930 146100 69960 146160
rect 70050 146100 70080 146160
rect 70170 146100 70200 146160
rect 70290 146100 70320 146160
rect 70410 146100 70440 146160
rect 70530 146100 70560 146160
rect 70650 146100 70680 146160
rect 70770 146100 70800 146160
rect 70890 146100 70920 146160
rect 71010 146100 71040 146160
rect 71130 146100 71160 146160
rect 71250 146100 71280 146160
rect 71370 146100 71400 146160
rect 71490 146100 71520 146160
rect 71610 146100 71640 146160
rect 71730 146100 71760 146160
rect 71850 146100 71880 146160
rect 71970 146100 72000 146160
rect 72090 146100 72120 146160
rect 72210 146100 72240 146160
rect 72330 146100 72360 146160
rect 72450 146100 72480 146160
rect 72570 146100 72600 146160
rect 72690 146100 72720 146160
rect 72810 146100 72840 146160
rect 72930 146100 72960 146160
rect 73050 146100 73080 146160
rect 73170 146100 73200 146160
rect 73290 146100 73320 146160
rect 73410 146100 73440 146160
rect 73530 146100 73560 146160
rect 73650 146100 73680 146160
rect 75870 146100 75900 146160
rect 75990 146100 76020 146160
rect 76110 146100 76140 146160
rect 76230 146100 76260 146160
rect 76350 146100 76380 146160
rect 76470 146100 76500 146160
rect 76590 146100 76620 146160
rect 76710 146100 76740 146160
rect 76830 146100 76860 146160
rect 76950 146100 76980 146160
rect 77070 146100 77100 146160
rect 77190 146100 77220 146160
rect 77310 146100 77340 146160
rect 77430 146100 77460 146160
rect 77550 146100 77580 146160
rect 77670 146100 77700 146160
rect 77790 146100 77820 146160
rect 77910 146100 77940 146160
rect 78030 146100 78060 146160
rect 78150 146100 78180 146160
rect 78270 146100 78300 146160
rect 78390 146100 78420 146160
rect 78510 146100 78540 146160
rect 78630 146100 78660 146160
rect 78750 146100 78780 146160
rect 78870 146100 78900 146160
rect 78990 146100 79020 146160
rect 79110 146100 79140 146160
rect 79230 146100 79260 146160
rect 79350 146100 79380 146160
rect 79470 146100 79500 146160
rect 79590 146100 79620 146160
rect 79710 146100 79740 146160
rect 79830 146100 79860 146160
rect 79950 146100 79980 146160
rect 80070 146100 80100 146160
rect 80190 146100 80220 146160
rect 80310 146100 80340 146160
rect 80430 146100 80460 146160
rect 80550 146100 80580 146160
rect 80670 146100 80700 146160
rect 80790 146100 80820 146160
rect 80910 146100 80940 146160
rect 81030 146100 81060 146160
rect 81150 146100 81180 146160
rect 81270 146100 81300 146160
rect 81390 146100 81420 146160
rect 81510 146100 81540 146160
rect 81630 146100 81660 146160
rect 81750 146100 81780 146160
rect 81870 146100 81900 146160
rect 81990 146100 82020 146160
rect 82110 146100 82140 146160
rect 82230 146100 82260 146160
rect 82350 146100 82380 146160
rect 82470 146100 82500 146160
rect 82590 146100 82620 146160
rect 82710 146100 82740 146160
rect 82830 146100 82860 146160
rect 82950 146100 82980 146160
rect 83070 146100 83100 146160
rect 83190 146100 83220 146160
rect 83310 146100 83340 146160
rect 83430 146100 83460 146160
rect 83550 146100 83580 146160
rect 83670 146100 83700 146160
rect 83790 146100 83820 146160
rect 83910 146100 83940 146160
rect 84030 146100 84060 146160
rect 84150 146100 84180 146160
rect 84270 146100 84300 146160
rect 84390 146100 84420 146160
rect 84510 146100 84540 146160
rect 84630 146100 84660 146160
rect 84750 146100 84780 146160
rect 84870 146100 84900 146160
rect 84990 146100 85020 146160
rect 85110 146100 85140 146160
rect 85230 146100 85260 146160
rect 85350 146100 85380 146160
rect 85470 146100 85500 146160
rect 85590 146100 85620 146160
rect 85710 146100 85740 146160
rect 85830 146100 85860 146160
rect 85950 146100 85980 146160
rect 86070 146100 86100 146160
rect 86190 146100 86220 146160
rect 86310 146100 86340 146160
rect 86430 146100 86460 146160
rect 86550 146100 86580 146160
rect 86670 146100 86700 146160
rect 86790 146100 86820 146160
rect 86910 146100 86940 146160
rect 87030 146100 87060 146160
rect 87150 146100 87180 146160
rect 89370 146100 89400 146160
rect 89490 146100 89520 146160
rect 89610 146100 89640 146160
rect 89730 146100 89760 146160
rect 89850 146100 89880 146160
rect 89970 146100 90000 146160
rect 90090 146100 90120 146160
rect 90210 146100 90240 146160
rect 90330 146100 90360 146160
rect 90450 146100 90480 146160
rect 90570 146100 90600 146160
rect 90690 146100 90720 146160
rect 90810 146100 90840 146160
rect 90930 146100 90960 146160
rect 91050 146100 91080 146160
rect 91170 146100 91200 146160
rect 91290 146100 91320 146160
rect 91410 146100 91440 146160
rect 91530 146100 91560 146160
rect 91650 146100 91680 146160
rect 91770 146100 91800 146160
rect 91890 146100 91920 146160
rect 92010 146100 92040 146160
rect 92130 146100 92160 146160
rect 92250 146100 92280 146160
rect 92370 146100 92400 146160
rect 92490 146100 92520 146160
rect 92610 146100 92640 146160
rect 92730 146100 92760 146160
rect 92850 146100 92880 146160
rect 92970 146100 93000 146160
rect 93090 146100 93120 146160
rect 93210 146100 93240 146160
rect 93330 146100 93360 146160
rect 93450 146100 93480 146160
rect 93570 146100 93600 146160
rect 93690 146100 93720 146160
rect 93810 146100 93840 146160
rect 93930 146100 93960 146160
rect 94050 146100 94080 146160
rect 94170 146100 94200 146160
rect 94290 146100 94320 146160
rect 94410 146100 94440 146160
rect 94530 146100 94560 146160
rect 94650 146100 94680 146160
rect 94770 146100 94800 146160
rect 94890 146100 94920 146160
rect 95010 146100 95040 146160
rect 95130 146100 95160 146160
rect 95250 146100 95280 146160
rect 95370 146100 95400 146160
rect 95490 146100 95520 146160
rect 95610 146100 95640 146160
rect 95730 146100 95760 146160
rect 95850 146100 95880 146160
rect 95970 146100 96000 146160
rect 96090 146100 96120 146160
rect 96210 146100 96240 146160
rect 96330 146100 96360 146160
rect 96450 146100 96480 146160
rect 96570 146100 96600 146160
rect 96690 146100 96720 146160
rect 96810 146100 96840 146160
rect 96930 146100 96960 146160
rect 97050 146100 97080 146160
rect 97170 146100 97200 146160
rect 97290 146100 97320 146160
rect 97410 146100 97440 146160
rect 97530 146100 97560 146160
rect 97650 146100 97680 146160
rect 97770 146100 97800 146160
rect 97890 146100 97920 146160
rect 98010 146100 98040 146160
rect 98130 146100 98160 146160
rect 98250 146100 98280 146160
rect 98370 146100 98400 146160
rect 98490 146100 98520 146160
rect 98610 146100 98640 146160
rect 98730 146100 98760 146160
rect 98850 146100 98880 146160
rect 98970 146100 99000 146160
rect 99090 146100 99120 146160
rect 99210 146100 99240 146160
rect 99330 146100 99360 146160
rect 99450 146100 99480 146160
rect 99570 146100 99600 146160
rect 99690 146100 99720 146160
rect 99810 146100 99840 146160
rect 99930 146100 99960 146160
rect 100050 146100 100080 146160
rect 100170 146100 100200 146160
rect 100290 146100 100320 146160
rect 100410 146100 100440 146160
rect 100530 146100 100560 146160
rect 100650 146100 100680 146160
rect 116370 146100 116400 146160
rect 116490 146100 116520 146160
rect 116610 146100 116640 146160
rect 116730 146100 116760 146160
rect 116850 146100 116880 146160
rect 116970 146100 117000 146160
rect 117090 146100 117120 146160
rect 117210 146100 117240 146160
rect 117330 146100 117360 146160
rect 127290 146100 127320 146160
rect 127410 146100 127440 146160
rect 127530 146100 127560 146160
rect 127650 146100 127680 146160
rect 129870 146100 129900 146160
rect 129990 146100 130020 146160
rect 130110 146100 130140 146160
rect 130230 146100 130260 146160
rect 130350 146100 130380 146160
rect 130470 146100 130500 146160
rect 130590 146100 130620 146160
rect 130710 146100 130740 146160
rect 130830 146100 130860 146160
rect 140790 146100 140820 146160
rect 140910 146100 140940 146160
rect 141030 146100 141060 146160
rect 141150 146100 141180 146160
rect 146480 146135 146490 146215
rect 146800 146135 146810 146215
rect 147120 146135 147130 146215
rect 147440 146135 147450 146215
rect 148860 146135 148870 146215
rect 149180 146135 149190 146215
rect 149500 146135 149510 146215
rect 149820 146135 149830 146215
rect 152280 146135 152290 146215
rect 152600 146135 152610 146215
rect 152920 146135 152930 146215
rect 153240 146135 153250 146215
rect 153560 146135 153570 146215
rect 153880 146135 153890 146215
rect 154200 146135 154210 146215
rect 154520 146135 154530 146215
rect 154840 146135 154850 146215
rect 155160 146135 155170 146215
rect 155480 146135 155490 146215
rect 155800 146135 155810 146215
rect 156120 146135 156130 146215
rect 156440 146135 156450 146215
rect 156760 146135 156770 146215
rect 157080 146135 157090 146215
rect 157400 146135 157410 146215
rect 157720 146135 157730 146215
rect 158040 146135 158050 146215
rect 158360 146135 158370 146215
rect 158680 146135 158690 146215
rect 159000 146135 159010 146215
rect 159320 146135 159330 146215
rect 159640 146135 159650 146215
rect 163750 146095 163830 146105
rect 164070 146095 164150 146105
rect 164390 146095 164470 146105
rect 164710 146095 164790 146105
rect 165030 146095 165110 146105
rect 165350 146095 165430 146105
rect 165670 146095 165750 146105
rect 165990 146095 166070 146105
rect 166310 146095 166390 146105
rect 166630 146095 166710 146105
rect 166950 146095 167030 146105
rect 167270 146095 167350 146105
rect 167590 146095 167670 146105
rect 167910 146095 167990 146105
rect 168230 146095 168310 146105
rect 168550 146095 168630 146105
rect 168870 146095 168950 146105
rect 169190 146095 169270 146105
rect 169510 146095 169590 146105
rect 169830 146095 169910 146105
rect 170150 146095 170230 146105
rect 170470 146095 170550 146105
rect 170790 146095 170870 146105
rect 146560 146055 146640 146065
rect 146880 146055 146960 146065
rect 147200 146055 147280 146065
rect 148940 146055 149020 146065
rect 149260 146055 149340 146065
rect 149580 146055 149660 146065
rect 152360 146055 152440 146065
rect 152680 146055 152760 146065
rect 153000 146055 153080 146065
rect 153320 146055 153400 146065
rect 153640 146055 153720 146065
rect 153960 146055 154040 146065
rect 154280 146055 154360 146065
rect 154600 146055 154680 146065
rect 154920 146055 155000 146065
rect 155240 146055 155320 146065
rect 155560 146055 155640 146065
rect 155880 146055 155960 146065
rect 156200 146055 156280 146065
rect 156520 146055 156600 146065
rect 156840 146055 156920 146065
rect 157160 146055 157240 146065
rect 157480 146055 157560 146065
rect 157800 146055 157880 146065
rect 158120 146055 158200 146065
rect 158440 146055 158520 146065
rect 158760 146055 158840 146065
rect 159080 146055 159160 146065
rect 159400 146055 159480 146065
rect 146640 145975 146650 146055
rect 146960 145975 146970 146055
rect 147280 145975 147290 146055
rect 149020 145975 149030 146055
rect 149340 145975 149350 146055
rect 149660 145975 149670 146055
rect 152440 145975 152450 146055
rect 152760 145975 152770 146055
rect 153080 145975 153090 146055
rect 153400 145975 153410 146055
rect 153720 145975 153730 146055
rect 154040 145975 154050 146055
rect 154360 145975 154370 146055
rect 154680 145975 154690 146055
rect 155000 145975 155010 146055
rect 155320 145975 155330 146055
rect 155640 145975 155650 146055
rect 155960 145975 155970 146055
rect 156280 145975 156290 146055
rect 156600 145975 156610 146055
rect 156920 145975 156930 146055
rect 157240 145975 157250 146055
rect 157560 145975 157570 146055
rect 157880 145975 157890 146055
rect 158200 145975 158210 146055
rect 158520 145975 158530 146055
rect 158840 145975 158850 146055
rect 159160 145975 159170 146055
rect 159480 145975 159490 146055
rect 163830 146015 163840 146095
rect 164150 146015 164160 146095
rect 164470 146015 164480 146095
rect 164790 146015 164800 146095
rect 165110 146015 165120 146095
rect 165430 146015 165440 146095
rect 165750 146015 165760 146095
rect 166070 146015 166080 146095
rect 166390 146015 166400 146095
rect 166710 146015 166720 146095
rect 167030 146015 167040 146095
rect 167350 146015 167360 146095
rect 167670 146015 167680 146095
rect 167990 146015 168000 146095
rect 168310 146015 168320 146095
rect 168630 146015 168640 146095
rect 168950 146015 168960 146095
rect 169270 146015 169280 146095
rect 169590 146015 169600 146095
rect 169910 146015 169920 146095
rect 170230 146015 170240 146095
rect 170550 146015 170560 146095
rect 170870 146015 170880 146095
rect 18970 145935 19050 145945
rect 19290 145935 19370 145945
rect 19610 145935 19690 145945
rect 19930 145935 20010 145945
rect 20250 145935 20330 145945
rect 20570 145935 20650 145945
rect 20890 145935 20970 145945
rect 21210 145935 21290 145945
rect 21530 145935 21610 145945
rect 21850 145935 21930 145945
rect 22170 145935 22250 145945
rect 22490 145935 22570 145945
rect 22810 145935 22890 145945
rect 23130 145935 23210 145945
rect 23450 145935 23530 145945
rect 23770 145935 23850 145945
rect 24090 145935 24170 145945
rect 24410 145935 24490 145945
rect 24730 145935 24810 145945
rect 25050 145935 25130 145945
rect 25370 145935 25450 145945
rect 25690 145935 25770 145945
rect 26010 145935 26090 145945
rect 26330 145935 26410 145945
rect 163590 145935 163670 145945
rect 163910 145935 163990 145945
rect 164230 145935 164310 145945
rect 164550 145935 164630 145945
rect 164870 145935 164950 145945
rect 165190 145935 165270 145945
rect 165510 145935 165590 145945
rect 165830 145935 165910 145945
rect 166150 145935 166230 145945
rect 166470 145935 166550 145945
rect 166790 145935 166870 145945
rect 167110 145935 167190 145945
rect 167430 145935 167510 145945
rect 167750 145935 167830 145945
rect 168070 145935 168150 145945
rect 168390 145935 168470 145945
rect 168710 145935 168790 145945
rect 169030 145935 169110 145945
rect 169350 145935 169430 145945
rect 169670 145935 169750 145945
rect 169990 145935 170070 145945
rect 170310 145935 170390 145945
rect 170630 145935 170710 145945
rect 170950 145935 171030 145945
rect 19050 145855 19060 145935
rect 19370 145855 19380 145935
rect 19690 145855 19700 145935
rect 20010 145855 20020 145935
rect 20330 145855 20340 145935
rect 20650 145855 20660 145935
rect 20970 145855 20980 145935
rect 21290 145855 21300 145935
rect 21610 145855 21620 145935
rect 21930 145855 21940 145935
rect 22250 145855 22260 145935
rect 22570 145855 22580 145935
rect 22890 145855 22900 145935
rect 23210 145855 23220 145935
rect 23530 145855 23540 145935
rect 23850 145855 23860 145935
rect 24170 145855 24180 145935
rect 24490 145855 24500 145935
rect 24810 145855 24820 145935
rect 25130 145855 25140 145935
rect 25450 145855 25460 145935
rect 25770 145855 25780 145935
rect 26090 145855 26100 145935
rect 26410 145855 26420 145935
rect 30360 145895 30440 145905
rect 30680 145895 30760 145905
rect 31000 145895 31080 145905
rect 31320 145895 31400 145905
rect 31640 145895 31720 145905
rect 31960 145895 32040 145905
rect 32280 145895 32360 145905
rect 32600 145895 32680 145905
rect 32920 145895 33000 145905
rect 33240 145895 33320 145905
rect 33560 145895 33640 145905
rect 33880 145895 33960 145905
rect 34200 145895 34280 145905
rect 34520 145895 34600 145905
rect 34840 145895 34920 145905
rect 35160 145895 35240 145905
rect 35480 145895 35560 145905
rect 35800 145895 35880 145905
rect 36120 145895 36200 145905
rect 36440 145895 36520 145905
rect 36760 145895 36840 145905
rect 37080 145895 37160 145905
rect 37400 145895 37480 145905
rect 37720 145895 37800 145905
rect 40180 145895 40260 145905
rect 40500 145895 40580 145905
rect 40820 145895 40900 145905
rect 41140 145895 41220 145905
rect 42560 145895 42640 145905
rect 42880 145895 42960 145905
rect 43200 145895 43280 145905
rect 43520 145895 43600 145905
rect 146400 145895 146480 145905
rect 146720 145895 146800 145905
rect 147040 145895 147120 145905
rect 147360 145895 147440 145905
rect 148780 145895 148860 145905
rect 149100 145895 149180 145905
rect 149420 145895 149500 145905
rect 149740 145895 149820 145905
rect 152200 145895 152280 145905
rect 152520 145895 152600 145905
rect 152840 145895 152920 145905
rect 153160 145895 153240 145905
rect 153480 145895 153560 145905
rect 153800 145895 153880 145905
rect 154120 145895 154200 145905
rect 154440 145895 154520 145905
rect 154760 145895 154840 145905
rect 155080 145895 155160 145905
rect 155400 145895 155480 145905
rect 155720 145895 155800 145905
rect 156040 145895 156120 145905
rect 156360 145895 156440 145905
rect 156680 145895 156760 145905
rect 157000 145895 157080 145905
rect 157320 145895 157400 145905
rect 157640 145895 157720 145905
rect 157960 145895 158040 145905
rect 158280 145895 158360 145905
rect 158600 145895 158680 145905
rect 158920 145895 159000 145905
rect 159240 145895 159320 145905
rect 159560 145895 159640 145905
rect 30440 145815 30450 145895
rect 30760 145815 30770 145895
rect 31080 145815 31090 145895
rect 31400 145815 31410 145895
rect 31720 145815 31730 145895
rect 32040 145815 32050 145895
rect 32360 145815 32370 145895
rect 32680 145815 32690 145895
rect 33000 145815 33010 145895
rect 33320 145815 33330 145895
rect 33640 145815 33650 145895
rect 33960 145815 33970 145895
rect 34280 145815 34290 145895
rect 34600 145815 34610 145895
rect 34920 145815 34930 145895
rect 35240 145815 35250 145895
rect 35560 145815 35570 145895
rect 35880 145815 35890 145895
rect 36200 145815 36210 145895
rect 36520 145815 36530 145895
rect 36840 145815 36850 145895
rect 37160 145815 37170 145895
rect 37480 145815 37490 145895
rect 37800 145815 37810 145895
rect 40260 145815 40270 145895
rect 40580 145815 40590 145895
rect 40900 145815 40910 145895
rect 41220 145815 41230 145895
rect 42640 145815 42650 145895
rect 42960 145815 42970 145895
rect 43280 145815 43290 145895
rect 43600 145815 43610 145895
rect 146480 145815 146490 145895
rect 146800 145815 146810 145895
rect 147120 145815 147130 145895
rect 147440 145815 147450 145895
rect 148860 145815 148870 145895
rect 149180 145815 149190 145895
rect 149500 145815 149510 145895
rect 149820 145815 149830 145895
rect 152280 145815 152290 145895
rect 152600 145815 152610 145895
rect 152920 145815 152930 145895
rect 153240 145815 153250 145895
rect 153560 145815 153570 145895
rect 153880 145815 153890 145895
rect 154200 145815 154210 145895
rect 154520 145815 154530 145895
rect 154840 145815 154850 145895
rect 155160 145815 155170 145895
rect 155480 145815 155490 145895
rect 155800 145815 155810 145895
rect 156120 145815 156130 145895
rect 156440 145815 156450 145895
rect 156760 145815 156770 145895
rect 157080 145815 157090 145895
rect 157400 145815 157410 145895
rect 157720 145815 157730 145895
rect 158040 145815 158050 145895
rect 158360 145815 158370 145895
rect 158680 145815 158690 145895
rect 159000 145815 159010 145895
rect 159320 145815 159330 145895
rect 159640 145815 159650 145895
rect 163670 145855 163680 145935
rect 163990 145855 164000 145935
rect 164310 145855 164320 145935
rect 164630 145855 164640 145935
rect 164950 145855 164960 145935
rect 165270 145855 165280 145935
rect 165590 145855 165600 145935
rect 165910 145855 165920 145935
rect 166230 145855 166240 145935
rect 166550 145855 166560 145935
rect 166870 145855 166880 145935
rect 167190 145855 167200 145935
rect 167510 145855 167520 145935
rect 167830 145855 167840 145935
rect 168150 145855 168160 145935
rect 168470 145855 168480 145935
rect 168790 145855 168800 145935
rect 169110 145855 169120 145935
rect 169430 145855 169440 145935
rect 169750 145855 169760 145935
rect 170070 145855 170080 145935
rect 170390 145855 170400 145935
rect 170710 145855 170720 145935
rect 171030 145855 171040 145935
rect 19130 145775 19210 145785
rect 19450 145775 19530 145785
rect 19770 145775 19850 145785
rect 20090 145775 20170 145785
rect 20410 145775 20490 145785
rect 20730 145775 20810 145785
rect 21050 145775 21130 145785
rect 21370 145775 21450 145785
rect 21690 145775 21770 145785
rect 22010 145775 22090 145785
rect 22330 145775 22410 145785
rect 22650 145775 22730 145785
rect 22970 145775 23050 145785
rect 23290 145775 23370 145785
rect 23610 145775 23690 145785
rect 23930 145775 24010 145785
rect 24250 145775 24330 145785
rect 24570 145775 24650 145785
rect 24890 145775 24970 145785
rect 25210 145775 25290 145785
rect 25530 145775 25610 145785
rect 25850 145775 25930 145785
rect 26170 145775 26250 145785
rect 163750 145775 163830 145785
rect 164070 145775 164150 145785
rect 164390 145775 164470 145785
rect 164710 145775 164790 145785
rect 165030 145775 165110 145785
rect 165350 145775 165430 145785
rect 165670 145775 165750 145785
rect 165990 145775 166070 145785
rect 166310 145775 166390 145785
rect 166630 145775 166710 145785
rect 166950 145775 167030 145785
rect 167270 145775 167350 145785
rect 167590 145775 167670 145785
rect 167910 145775 167990 145785
rect 168230 145775 168310 145785
rect 168550 145775 168630 145785
rect 168870 145775 168950 145785
rect 169190 145775 169270 145785
rect 169510 145775 169590 145785
rect 169830 145775 169910 145785
rect 170150 145775 170230 145785
rect 170470 145775 170550 145785
rect 170790 145775 170870 145785
rect 19210 145695 19220 145775
rect 19530 145695 19540 145775
rect 19850 145695 19860 145775
rect 20170 145695 20180 145775
rect 20490 145695 20500 145775
rect 20810 145695 20820 145775
rect 21130 145695 21140 145775
rect 21450 145695 21460 145775
rect 21770 145695 21780 145775
rect 22090 145695 22100 145775
rect 22410 145695 22420 145775
rect 22730 145695 22740 145775
rect 23050 145695 23060 145775
rect 23370 145695 23380 145775
rect 23690 145695 23700 145775
rect 24010 145695 24020 145775
rect 24330 145695 24340 145775
rect 24650 145695 24660 145775
rect 24970 145695 24980 145775
rect 25290 145695 25300 145775
rect 25610 145695 25620 145775
rect 25930 145695 25940 145775
rect 26250 145695 26260 145775
rect 30520 145735 30600 145745
rect 30840 145735 30920 145745
rect 31160 145735 31240 145745
rect 31480 145735 31560 145745
rect 31800 145735 31880 145745
rect 32120 145735 32200 145745
rect 32440 145735 32520 145745
rect 32760 145735 32840 145745
rect 33080 145735 33160 145745
rect 33400 145735 33480 145745
rect 33720 145735 33800 145745
rect 34040 145735 34120 145745
rect 34360 145735 34440 145745
rect 34680 145735 34760 145745
rect 35000 145735 35080 145745
rect 35320 145735 35400 145745
rect 35640 145735 35720 145745
rect 35960 145735 36040 145745
rect 36280 145735 36360 145745
rect 36600 145735 36680 145745
rect 36920 145735 37000 145745
rect 37240 145735 37320 145745
rect 37560 145735 37640 145745
rect 40340 145735 40420 145745
rect 40660 145735 40740 145745
rect 40980 145735 41060 145745
rect 42720 145735 42800 145745
rect 43040 145735 43120 145745
rect 43360 145735 43440 145745
rect 146560 145735 146640 145745
rect 146880 145735 146960 145745
rect 147200 145735 147280 145745
rect 148940 145735 149020 145745
rect 149260 145735 149340 145745
rect 149580 145735 149660 145745
rect 152360 145735 152440 145745
rect 152680 145735 152760 145745
rect 153000 145735 153080 145745
rect 153320 145735 153400 145745
rect 153640 145735 153720 145745
rect 153960 145735 154040 145745
rect 154280 145735 154360 145745
rect 154600 145735 154680 145745
rect 154920 145735 155000 145745
rect 155240 145735 155320 145745
rect 155560 145735 155640 145745
rect 155880 145735 155960 145745
rect 156200 145735 156280 145745
rect 156520 145735 156600 145745
rect 156840 145735 156920 145745
rect 157160 145735 157240 145745
rect 157480 145735 157560 145745
rect 157800 145735 157880 145745
rect 158120 145735 158200 145745
rect 158440 145735 158520 145745
rect 158760 145735 158840 145745
rect 159080 145735 159160 145745
rect 159400 145735 159480 145745
rect 30600 145655 30610 145735
rect 30920 145655 30930 145735
rect 31240 145655 31250 145735
rect 31560 145655 31570 145735
rect 31880 145655 31890 145735
rect 32200 145655 32210 145735
rect 32520 145655 32530 145735
rect 32840 145655 32850 145735
rect 33160 145655 33170 145735
rect 33480 145655 33490 145735
rect 33800 145655 33810 145735
rect 34120 145655 34130 145735
rect 34440 145655 34450 145735
rect 34760 145655 34770 145735
rect 35080 145655 35090 145735
rect 35400 145655 35410 145735
rect 35720 145655 35730 145735
rect 36040 145655 36050 145735
rect 36360 145655 36370 145735
rect 36680 145655 36690 145735
rect 37000 145655 37010 145735
rect 37320 145655 37330 145735
rect 37640 145655 37650 145735
rect 40420 145655 40430 145735
rect 40740 145655 40750 145735
rect 41060 145655 41070 145735
rect 42800 145655 42810 145735
rect 43120 145655 43130 145735
rect 43440 145655 43450 145735
rect 146640 145655 146650 145735
rect 146960 145655 146970 145735
rect 147280 145655 147290 145735
rect 149020 145655 149030 145735
rect 149340 145655 149350 145735
rect 149660 145655 149670 145735
rect 152440 145655 152450 145735
rect 152760 145655 152770 145735
rect 153080 145655 153090 145735
rect 153400 145655 153410 145735
rect 153720 145655 153730 145735
rect 154040 145655 154050 145735
rect 154360 145655 154370 145735
rect 154680 145655 154690 145735
rect 155000 145655 155010 145735
rect 155320 145655 155330 145735
rect 155640 145655 155650 145735
rect 155960 145655 155970 145735
rect 156280 145655 156290 145735
rect 156600 145655 156610 145735
rect 156920 145655 156930 145735
rect 157240 145655 157250 145735
rect 157560 145655 157570 145735
rect 157880 145655 157890 145735
rect 158200 145655 158210 145735
rect 158520 145655 158530 145735
rect 158840 145655 158850 145735
rect 159160 145655 159170 145735
rect 159480 145655 159490 145735
rect 163830 145695 163840 145775
rect 164150 145695 164160 145775
rect 164470 145695 164480 145775
rect 164790 145695 164800 145775
rect 165110 145695 165120 145775
rect 165430 145695 165440 145775
rect 165750 145695 165760 145775
rect 166070 145695 166080 145775
rect 166390 145695 166400 145775
rect 166710 145695 166720 145775
rect 167030 145695 167040 145775
rect 167350 145695 167360 145775
rect 167670 145695 167680 145775
rect 167990 145695 168000 145775
rect 168310 145695 168320 145775
rect 168630 145695 168640 145775
rect 168950 145695 168960 145775
rect 169270 145695 169280 145775
rect 169590 145695 169600 145775
rect 169910 145695 169920 145775
rect 170230 145695 170240 145775
rect 170550 145695 170560 145775
rect 170870 145695 170880 145775
rect 18970 145615 19050 145625
rect 19290 145615 19370 145625
rect 19610 145615 19690 145625
rect 19930 145615 20010 145625
rect 20250 145615 20330 145625
rect 20570 145615 20650 145625
rect 20890 145615 20970 145625
rect 21210 145615 21290 145625
rect 21530 145615 21610 145625
rect 21850 145615 21930 145625
rect 22170 145615 22250 145625
rect 22490 145615 22570 145625
rect 22810 145615 22890 145625
rect 23130 145615 23210 145625
rect 23450 145615 23530 145625
rect 23770 145615 23850 145625
rect 24090 145615 24170 145625
rect 24410 145615 24490 145625
rect 24730 145615 24810 145625
rect 25050 145615 25130 145625
rect 25370 145615 25450 145625
rect 25690 145615 25770 145625
rect 26010 145615 26090 145625
rect 26330 145615 26410 145625
rect 163590 145615 163670 145625
rect 163910 145615 163990 145625
rect 164230 145615 164310 145625
rect 164550 145615 164630 145625
rect 164870 145615 164950 145625
rect 165190 145615 165270 145625
rect 165510 145615 165590 145625
rect 165830 145615 165910 145625
rect 166150 145615 166230 145625
rect 166470 145615 166550 145625
rect 166790 145615 166870 145625
rect 167110 145615 167190 145625
rect 167430 145615 167510 145625
rect 167750 145615 167830 145625
rect 168070 145615 168150 145625
rect 168390 145615 168470 145625
rect 168710 145615 168790 145625
rect 169030 145615 169110 145625
rect 169350 145615 169430 145625
rect 169670 145615 169750 145625
rect 169990 145615 170070 145625
rect 170310 145615 170390 145625
rect 170630 145615 170710 145625
rect 170950 145615 171030 145625
rect 19050 145535 19060 145615
rect 19370 145535 19380 145615
rect 19690 145535 19700 145615
rect 20010 145535 20020 145615
rect 20330 145535 20340 145615
rect 20650 145535 20660 145615
rect 20970 145535 20980 145615
rect 21290 145535 21300 145615
rect 21610 145535 21620 145615
rect 21930 145535 21940 145615
rect 22250 145535 22260 145615
rect 22570 145535 22580 145615
rect 22890 145535 22900 145615
rect 23210 145535 23220 145615
rect 23530 145535 23540 145615
rect 23850 145535 23860 145615
rect 24170 145535 24180 145615
rect 24490 145535 24500 145615
rect 24810 145535 24820 145615
rect 25130 145535 25140 145615
rect 25450 145535 25460 145615
rect 25770 145535 25780 145615
rect 26090 145535 26100 145615
rect 26410 145535 26420 145615
rect 30360 145575 30440 145585
rect 30680 145575 30760 145585
rect 31000 145575 31080 145585
rect 31320 145575 31400 145585
rect 31640 145575 31720 145585
rect 31960 145575 32040 145585
rect 32280 145575 32360 145585
rect 32600 145575 32680 145585
rect 32920 145575 33000 145585
rect 33240 145575 33320 145585
rect 33560 145575 33640 145585
rect 33880 145575 33960 145585
rect 34200 145575 34280 145585
rect 34520 145575 34600 145585
rect 34840 145575 34920 145585
rect 35160 145575 35240 145585
rect 35480 145575 35560 145585
rect 35800 145575 35880 145585
rect 36120 145575 36200 145585
rect 36440 145575 36520 145585
rect 36760 145575 36840 145585
rect 37080 145575 37160 145585
rect 37400 145575 37480 145585
rect 37720 145575 37800 145585
rect 40180 145575 40260 145585
rect 40500 145575 40580 145585
rect 40820 145575 40900 145585
rect 41140 145575 41220 145585
rect 42560 145575 42640 145585
rect 42880 145575 42960 145585
rect 43200 145575 43280 145585
rect 43520 145575 43600 145585
rect 146400 145575 146480 145585
rect 146720 145575 146800 145585
rect 147040 145575 147120 145585
rect 147360 145575 147440 145585
rect 148780 145575 148860 145585
rect 149100 145575 149180 145585
rect 149420 145575 149500 145585
rect 149740 145575 149820 145585
rect 152200 145575 152280 145585
rect 152520 145575 152600 145585
rect 152840 145575 152920 145585
rect 153160 145575 153240 145585
rect 153480 145575 153560 145585
rect 153800 145575 153880 145585
rect 154120 145575 154200 145585
rect 154440 145575 154520 145585
rect 154760 145575 154840 145585
rect 155080 145575 155160 145585
rect 155400 145575 155480 145585
rect 155720 145575 155800 145585
rect 156040 145575 156120 145585
rect 156360 145575 156440 145585
rect 156680 145575 156760 145585
rect 157000 145575 157080 145585
rect 157320 145575 157400 145585
rect 157640 145575 157720 145585
rect 157960 145575 158040 145585
rect 158280 145575 158360 145585
rect 158600 145575 158680 145585
rect 158920 145575 159000 145585
rect 159240 145575 159320 145585
rect 159560 145575 159640 145585
rect 30440 145495 30450 145575
rect 30760 145495 30770 145575
rect 31080 145495 31090 145575
rect 31400 145495 31410 145575
rect 31720 145495 31730 145575
rect 32040 145495 32050 145575
rect 32360 145495 32370 145575
rect 32680 145495 32690 145575
rect 33000 145495 33010 145575
rect 33320 145495 33330 145575
rect 33640 145495 33650 145575
rect 33960 145495 33970 145575
rect 34280 145495 34290 145575
rect 34600 145495 34610 145575
rect 34920 145495 34930 145575
rect 35240 145495 35250 145575
rect 35560 145495 35570 145575
rect 35880 145495 35890 145575
rect 36200 145495 36210 145575
rect 36520 145495 36530 145575
rect 36840 145495 36850 145575
rect 37160 145495 37170 145575
rect 37480 145495 37490 145575
rect 37800 145495 37810 145575
rect 40260 145495 40270 145575
rect 40580 145495 40590 145575
rect 40900 145495 40910 145575
rect 41220 145495 41230 145575
rect 42640 145495 42650 145575
rect 42960 145495 42970 145575
rect 43280 145495 43290 145575
rect 43600 145495 43610 145575
rect 146480 145495 146490 145575
rect 146800 145495 146810 145575
rect 147120 145495 147130 145575
rect 147440 145495 147450 145575
rect 148860 145495 148870 145575
rect 149180 145495 149190 145575
rect 149500 145495 149510 145575
rect 149820 145495 149830 145575
rect 152280 145495 152290 145575
rect 152600 145495 152610 145575
rect 152920 145495 152930 145575
rect 153240 145495 153250 145575
rect 153560 145495 153570 145575
rect 153880 145495 153890 145575
rect 154200 145495 154210 145575
rect 154520 145495 154530 145575
rect 154840 145495 154850 145575
rect 155160 145495 155170 145575
rect 155480 145495 155490 145575
rect 155800 145495 155810 145575
rect 156120 145495 156130 145575
rect 156440 145495 156450 145575
rect 156760 145495 156770 145575
rect 157080 145495 157090 145575
rect 157400 145495 157410 145575
rect 157720 145495 157730 145575
rect 158040 145495 158050 145575
rect 158360 145495 158370 145575
rect 158680 145495 158690 145575
rect 159000 145495 159010 145575
rect 159320 145495 159330 145575
rect 159640 145495 159650 145575
rect 163670 145535 163680 145615
rect 163990 145535 164000 145615
rect 164310 145535 164320 145615
rect 164630 145535 164640 145615
rect 164950 145535 164960 145615
rect 165270 145535 165280 145615
rect 165590 145535 165600 145615
rect 165910 145535 165920 145615
rect 166230 145535 166240 145615
rect 166550 145535 166560 145615
rect 166870 145535 166880 145615
rect 167190 145535 167200 145615
rect 167510 145535 167520 145615
rect 167830 145535 167840 145615
rect 168150 145535 168160 145615
rect 168470 145535 168480 145615
rect 168790 145535 168800 145615
rect 169110 145535 169120 145615
rect 169430 145535 169440 145615
rect 169750 145535 169760 145615
rect 170070 145535 170080 145615
rect 170390 145535 170400 145615
rect 170710 145535 170720 145615
rect 171030 145535 171040 145615
rect 19130 145455 19210 145465
rect 19450 145455 19530 145465
rect 19770 145455 19850 145465
rect 20090 145455 20170 145465
rect 20410 145455 20490 145465
rect 20730 145455 20810 145465
rect 21050 145455 21130 145465
rect 21370 145455 21450 145465
rect 21690 145455 21770 145465
rect 22010 145455 22090 145465
rect 22330 145455 22410 145465
rect 22650 145455 22730 145465
rect 22970 145455 23050 145465
rect 23290 145455 23370 145465
rect 23610 145455 23690 145465
rect 23930 145455 24010 145465
rect 24250 145455 24330 145465
rect 24570 145455 24650 145465
rect 24890 145455 24970 145465
rect 25210 145455 25290 145465
rect 25530 145455 25610 145465
rect 25850 145455 25930 145465
rect 26170 145455 26250 145465
rect 163750 145455 163830 145465
rect 164070 145455 164150 145465
rect 164390 145455 164470 145465
rect 164710 145455 164790 145465
rect 165030 145455 165110 145465
rect 165350 145455 165430 145465
rect 165670 145455 165750 145465
rect 165990 145455 166070 145465
rect 166310 145455 166390 145465
rect 166630 145455 166710 145465
rect 166950 145455 167030 145465
rect 167270 145455 167350 145465
rect 167590 145455 167670 145465
rect 167910 145455 167990 145465
rect 168230 145455 168310 145465
rect 168550 145455 168630 145465
rect 168870 145455 168950 145465
rect 169190 145455 169270 145465
rect 169510 145455 169590 145465
rect 169830 145455 169910 145465
rect 170150 145455 170230 145465
rect 170470 145455 170550 145465
rect 170790 145455 170870 145465
rect 19210 145375 19220 145455
rect 19530 145375 19540 145455
rect 19850 145375 19860 145455
rect 20170 145375 20180 145455
rect 20490 145375 20500 145455
rect 20810 145375 20820 145455
rect 21130 145375 21140 145455
rect 21450 145375 21460 145455
rect 21770 145375 21780 145455
rect 22090 145375 22100 145455
rect 22410 145375 22420 145455
rect 22730 145375 22740 145455
rect 23050 145375 23060 145455
rect 23370 145375 23380 145455
rect 23690 145375 23700 145455
rect 24010 145375 24020 145455
rect 24330 145375 24340 145455
rect 24650 145375 24660 145455
rect 24970 145375 24980 145455
rect 25290 145375 25300 145455
rect 25610 145375 25620 145455
rect 25930 145375 25940 145455
rect 26250 145375 26260 145455
rect 30520 145415 30600 145425
rect 30840 145415 30920 145425
rect 31160 145415 31240 145425
rect 31480 145415 31560 145425
rect 31800 145415 31880 145425
rect 32120 145415 32200 145425
rect 32440 145415 32520 145425
rect 32760 145415 32840 145425
rect 33080 145415 33160 145425
rect 33400 145415 33480 145425
rect 33720 145415 33800 145425
rect 34040 145415 34120 145425
rect 34360 145415 34440 145425
rect 34680 145415 34760 145425
rect 35000 145415 35080 145425
rect 35320 145415 35400 145425
rect 35640 145415 35720 145425
rect 35960 145415 36040 145425
rect 36280 145415 36360 145425
rect 36600 145415 36680 145425
rect 36920 145415 37000 145425
rect 37240 145415 37320 145425
rect 37560 145415 37640 145425
rect 40340 145415 40420 145425
rect 40660 145415 40740 145425
rect 40980 145415 41060 145425
rect 42720 145415 42800 145425
rect 43040 145415 43120 145425
rect 43360 145415 43440 145425
rect 146560 145415 146640 145425
rect 146880 145415 146960 145425
rect 147200 145415 147280 145425
rect 148940 145415 149020 145425
rect 149260 145415 149340 145425
rect 149580 145415 149660 145425
rect 152360 145415 152440 145425
rect 152680 145415 152760 145425
rect 153000 145415 153080 145425
rect 153320 145415 153400 145425
rect 153640 145415 153720 145425
rect 153960 145415 154040 145425
rect 154280 145415 154360 145425
rect 154600 145415 154680 145425
rect 154920 145415 155000 145425
rect 155240 145415 155320 145425
rect 155560 145415 155640 145425
rect 155880 145415 155960 145425
rect 156200 145415 156280 145425
rect 156520 145415 156600 145425
rect 156840 145415 156920 145425
rect 157160 145415 157240 145425
rect 157480 145415 157560 145425
rect 157800 145415 157880 145425
rect 158120 145415 158200 145425
rect 158440 145415 158520 145425
rect 158760 145415 158840 145425
rect 159080 145415 159160 145425
rect 159400 145415 159480 145425
rect 30600 145335 30610 145415
rect 30920 145335 30930 145415
rect 31240 145335 31250 145415
rect 31560 145335 31570 145415
rect 31880 145335 31890 145415
rect 32200 145335 32210 145415
rect 32520 145335 32530 145415
rect 32840 145335 32850 145415
rect 33160 145335 33170 145415
rect 33480 145335 33490 145415
rect 33800 145335 33810 145415
rect 34120 145335 34130 145415
rect 34440 145335 34450 145415
rect 34760 145335 34770 145415
rect 35080 145335 35090 145415
rect 35400 145335 35410 145415
rect 35720 145335 35730 145415
rect 36040 145335 36050 145415
rect 36360 145335 36370 145415
rect 36680 145335 36690 145415
rect 37000 145335 37010 145415
rect 37320 145335 37330 145415
rect 37640 145335 37650 145415
rect 40420 145335 40430 145415
rect 40740 145335 40750 145415
rect 41060 145335 41070 145415
rect 42800 145335 42810 145415
rect 43120 145335 43130 145415
rect 43440 145335 43450 145415
rect 146640 145335 146650 145415
rect 146960 145335 146970 145415
rect 147280 145335 147290 145415
rect 149020 145335 149030 145415
rect 149340 145335 149350 145415
rect 149660 145335 149670 145415
rect 152440 145335 152450 145415
rect 152760 145335 152770 145415
rect 153080 145335 153090 145415
rect 153400 145335 153410 145415
rect 153720 145335 153730 145415
rect 154040 145335 154050 145415
rect 154360 145335 154370 145415
rect 154680 145335 154690 145415
rect 155000 145335 155010 145415
rect 155320 145335 155330 145415
rect 155640 145335 155650 145415
rect 155960 145335 155970 145415
rect 156280 145335 156290 145415
rect 156600 145335 156610 145415
rect 156920 145335 156930 145415
rect 157240 145335 157250 145415
rect 157560 145335 157570 145415
rect 157880 145335 157890 145415
rect 158200 145335 158210 145415
rect 158520 145335 158530 145415
rect 158840 145335 158850 145415
rect 159160 145335 159170 145415
rect 159480 145335 159490 145415
rect 163830 145375 163840 145455
rect 164150 145375 164160 145455
rect 164470 145375 164480 145455
rect 164790 145375 164800 145455
rect 165110 145375 165120 145455
rect 165430 145375 165440 145455
rect 165750 145375 165760 145455
rect 166070 145375 166080 145455
rect 166390 145375 166400 145455
rect 166710 145375 166720 145455
rect 167030 145375 167040 145455
rect 167350 145375 167360 145455
rect 167670 145375 167680 145455
rect 167990 145375 168000 145455
rect 168310 145375 168320 145455
rect 168630 145375 168640 145455
rect 168950 145375 168960 145455
rect 169270 145375 169280 145455
rect 169590 145375 169600 145455
rect 169910 145375 169920 145455
rect 170230 145375 170240 145455
rect 170550 145375 170560 145455
rect 170870 145375 170880 145455
rect 18970 145295 19050 145305
rect 19290 145295 19370 145305
rect 19610 145295 19690 145305
rect 19930 145295 20010 145305
rect 20250 145295 20330 145305
rect 20570 145295 20650 145305
rect 20890 145295 20970 145305
rect 21210 145295 21290 145305
rect 21530 145295 21610 145305
rect 21850 145295 21930 145305
rect 22170 145295 22250 145305
rect 22490 145295 22570 145305
rect 22810 145295 22890 145305
rect 23130 145295 23210 145305
rect 23450 145295 23530 145305
rect 23770 145295 23850 145305
rect 24090 145295 24170 145305
rect 24410 145295 24490 145305
rect 24730 145295 24810 145305
rect 25050 145295 25130 145305
rect 25370 145295 25450 145305
rect 25690 145295 25770 145305
rect 26010 145295 26090 145305
rect 26330 145295 26410 145305
rect 163590 145295 163670 145305
rect 163910 145295 163990 145305
rect 164230 145295 164310 145305
rect 164550 145295 164630 145305
rect 164870 145295 164950 145305
rect 165190 145295 165270 145305
rect 165510 145295 165590 145305
rect 165830 145295 165910 145305
rect 166150 145295 166230 145305
rect 166470 145295 166550 145305
rect 166790 145295 166870 145305
rect 167110 145295 167190 145305
rect 167430 145295 167510 145305
rect 167750 145295 167830 145305
rect 168070 145295 168150 145305
rect 168390 145295 168470 145305
rect 168710 145295 168790 145305
rect 169030 145295 169110 145305
rect 169350 145295 169430 145305
rect 169670 145295 169750 145305
rect 169990 145295 170070 145305
rect 170310 145295 170390 145305
rect 170630 145295 170710 145305
rect 170950 145295 171030 145305
rect 19050 145215 19060 145295
rect 19370 145215 19380 145295
rect 19690 145215 19700 145295
rect 20010 145215 20020 145295
rect 20330 145215 20340 145295
rect 20650 145215 20660 145295
rect 20970 145215 20980 145295
rect 21290 145215 21300 145295
rect 21610 145215 21620 145295
rect 21930 145215 21940 145295
rect 22250 145215 22260 145295
rect 22570 145215 22580 145295
rect 22890 145215 22900 145295
rect 23210 145215 23220 145295
rect 23530 145215 23540 145295
rect 23850 145215 23860 145295
rect 24170 145215 24180 145295
rect 24490 145215 24500 145295
rect 24810 145215 24820 145295
rect 25130 145215 25140 145295
rect 25450 145215 25460 145295
rect 25770 145215 25780 145295
rect 26090 145215 26100 145295
rect 26410 145215 26420 145295
rect 30360 145255 30440 145265
rect 30680 145255 30760 145265
rect 31000 145255 31080 145265
rect 31320 145255 31400 145265
rect 31640 145255 31720 145265
rect 31960 145255 32040 145265
rect 32280 145255 32360 145265
rect 32600 145255 32680 145265
rect 32920 145255 33000 145265
rect 33240 145255 33320 145265
rect 33560 145255 33640 145265
rect 33880 145255 33960 145265
rect 34200 145255 34280 145265
rect 34520 145255 34600 145265
rect 34840 145255 34920 145265
rect 35160 145255 35240 145265
rect 35480 145255 35560 145265
rect 35800 145255 35880 145265
rect 36120 145255 36200 145265
rect 36440 145255 36520 145265
rect 36760 145255 36840 145265
rect 37080 145255 37160 145265
rect 37400 145255 37480 145265
rect 37720 145255 37800 145265
rect 40180 145255 40260 145265
rect 40500 145255 40580 145265
rect 40820 145255 40900 145265
rect 41140 145255 41220 145265
rect 42560 145255 42640 145265
rect 42880 145255 42960 145265
rect 43200 145255 43280 145265
rect 43520 145255 43600 145265
rect 146400 145255 146480 145265
rect 146720 145255 146800 145265
rect 147040 145255 147120 145265
rect 147360 145255 147440 145265
rect 148780 145255 148860 145265
rect 149100 145255 149180 145265
rect 149420 145255 149500 145265
rect 149740 145255 149820 145265
rect 152200 145255 152280 145265
rect 152520 145255 152600 145265
rect 152840 145255 152920 145265
rect 153160 145255 153240 145265
rect 153480 145255 153560 145265
rect 153800 145255 153880 145265
rect 154120 145255 154200 145265
rect 154440 145255 154520 145265
rect 154760 145255 154840 145265
rect 155080 145255 155160 145265
rect 155400 145255 155480 145265
rect 155720 145255 155800 145265
rect 156040 145255 156120 145265
rect 156360 145255 156440 145265
rect 156680 145255 156760 145265
rect 157000 145255 157080 145265
rect 157320 145255 157400 145265
rect 157640 145255 157720 145265
rect 157960 145255 158040 145265
rect 158280 145255 158360 145265
rect 158600 145255 158680 145265
rect 158920 145255 159000 145265
rect 159240 145255 159320 145265
rect 159560 145255 159640 145265
rect 30440 145200 30450 145255
rect 30760 145200 30770 145255
rect 31080 145200 31090 145255
rect 31400 145200 31410 145255
rect 31720 145200 31730 145255
rect 32040 145200 32050 145255
rect 32360 145200 32370 145255
rect 32680 145200 32690 145255
rect 33000 145200 33010 145255
rect 33320 145200 33330 145255
rect 33640 145200 33650 145255
rect 33960 145200 33970 145255
rect 34280 145200 34290 145255
rect 34600 145200 34610 145255
rect 34920 145200 34930 145255
rect 35240 145200 35250 145255
rect 35560 145200 35570 145255
rect 35880 145200 35890 145255
rect 36200 145200 36210 145255
rect 36520 145200 36530 145255
rect 36840 145200 36850 145255
rect 37160 145200 37170 145255
rect 37480 145200 37490 145255
rect 37800 145200 37810 145255
rect 40260 145200 40270 145255
rect 40580 145200 40590 145255
rect 40900 145200 40910 145255
rect 41220 145200 41230 145255
rect 42640 145200 42650 145255
rect 42960 145200 42970 145255
rect 43280 145200 43290 145255
rect 43600 145200 43610 145255
rect 146480 145200 146490 145255
rect 146800 145200 146810 145255
rect 147120 145200 147130 145255
rect 147440 145200 147450 145255
rect 148860 145200 148870 145255
rect 149180 145200 149190 145255
rect 149500 145200 149510 145255
rect 149820 145200 149830 145255
rect 152280 145200 152290 145255
rect 152600 145200 152610 145255
rect 152920 145200 152930 145255
rect 153240 145200 153250 145255
rect 153560 145200 153570 145255
rect 153880 145200 153890 145255
rect 154200 145200 154210 145255
rect 154520 145200 154530 145255
rect 154840 145200 154850 145255
rect 155160 145200 155170 145255
rect 155480 145200 155490 145255
rect 155800 145200 155810 145255
rect 156120 145200 156130 145255
rect 156440 145200 156450 145255
rect 156760 145200 156770 145255
rect 157080 145200 157090 145255
rect 157400 145200 157410 145255
rect 157720 145200 157730 145255
rect 158040 145200 158050 145255
rect 158360 145200 158370 145255
rect 158680 145200 158690 145255
rect 159000 145200 159010 145255
rect 159320 145200 159330 145255
rect 159640 145200 159650 145255
rect 163670 145215 163680 145295
rect 163990 145215 164000 145295
rect 164310 145215 164320 145295
rect 164630 145215 164640 145295
rect 164950 145215 164960 145295
rect 165270 145215 165280 145295
rect 165590 145215 165600 145295
rect 165910 145215 165920 145295
rect 166230 145215 166240 145295
rect 166550 145215 166560 145295
rect 166870 145215 166880 145295
rect 167190 145215 167200 145295
rect 167510 145215 167520 145295
rect 167830 145215 167840 145295
rect 168150 145215 168160 145295
rect 168470 145215 168480 145295
rect 168790 145215 168800 145295
rect 169110 145215 169120 145295
rect 169430 145215 169440 145295
rect 169750 145215 169760 145295
rect 170070 145215 170080 145295
rect 170390 145215 170400 145295
rect 170710 145215 170720 145295
rect 171030 145215 171040 145295
rect 19210 142175 19220 142200
rect 19530 142175 19540 142200
rect 19850 142175 19860 142200
rect 20170 142175 20180 142200
rect 20490 142175 20500 142200
rect 20810 142175 20820 142200
rect 21130 142175 21140 142200
rect 21450 142175 21460 142200
rect 21770 142175 21780 142200
rect 22090 142175 22100 142200
rect 22410 142175 22420 142200
rect 22730 142175 22740 142200
rect 23050 142175 23060 142200
rect 23370 142175 23380 142200
rect 23690 142175 23700 142200
rect 24010 142175 24020 142200
rect 24330 142175 24340 142200
rect 24650 142175 24660 142200
rect 24970 142175 24980 142200
rect 25290 142175 25300 142200
rect 25610 142175 25620 142200
rect 25930 142175 25940 142200
rect 26250 142175 26260 142200
rect 30600 142135 30610 142200
rect 30920 142135 30930 142200
rect 31240 142135 31250 142200
rect 31560 142135 31570 142200
rect 31880 142135 31890 142200
rect 32200 142135 32210 142200
rect 32520 142135 32530 142200
rect 32840 142135 32850 142200
rect 33160 142135 33170 142200
rect 33480 142135 33490 142200
rect 33800 142135 33810 142200
rect 34120 142135 34130 142200
rect 34440 142135 34450 142200
rect 34760 142135 34770 142200
rect 35080 142135 35090 142200
rect 35400 142135 35410 142200
rect 35720 142135 35730 142200
rect 36040 142135 36050 142200
rect 36360 142135 36370 142200
rect 36680 142135 36690 142200
rect 37000 142135 37010 142200
rect 37320 142135 37330 142200
rect 37640 142135 37650 142200
rect 40420 142135 40430 142200
rect 40740 142135 40750 142200
rect 41060 142135 41070 142200
rect 42800 142135 42810 142200
rect 43120 142135 43130 142200
rect 43440 142135 43450 142200
rect 146640 142135 146650 142200
rect 146960 142135 146970 142200
rect 147280 142135 147290 142200
rect 149020 142135 149030 142200
rect 149340 142135 149350 142200
rect 149660 142135 149670 142200
rect 152440 142135 152450 142200
rect 152760 142135 152770 142200
rect 153080 142135 153090 142200
rect 153400 142135 153410 142200
rect 153720 142135 153730 142200
rect 154040 142135 154050 142200
rect 154360 142135 154370 142200
rect 154680 142135 154690 142200
rect 155000 142135 155010 142200
rect 155320 142135 155330 142200
rect 155640 142135 155650 142200
rect 155960 142135 155970 142200
rect 156280 142135 156290 142200
rect 156600 142135 156610 142200
rect 156920 142135 156930 142200
rect 157240 142135 157250 142200
rect 157560 142135 157570 142200
rect 157880 142135 157890 142200
rect 158200 142135 158210 142200
rect 158520 142135 158530 142200
rect 158840 142135 158850 142200
rect 159160 142135 159170 142200
rect 159480 142135 159490 142200
rect 163830 142175 163840 142200
rect 164150 142175 164160 142200
rect 164470 142175 164480 142200
rect 164790 142175 164800 142200
rect 165110 142175 165120 142200
rect 165430 142175 165440 142200
rect 165750 142175 165760 142200
rect 166070 142175 166080 142200
rect 166390 142175 166400 142200
rect 166710 142175 166720 142200
rect 167030 142175 167040 142200
rect 167350 142175 167360 142200
rect 167670 142175 167680 142200
rect 167990 142175 168000 142200
rect 168310 142175 168320 142200
rect 168630 142175 168640 142200
rect 168950 142175 168960 142200
rect 169270 142175 169280 142200
rect 169590 142175 169600 142200
rect 169910 142175 169920 142200
rect 170230 142175 170240 142200
rect 170550 142175 170560 142200
rect 170870 142175 170880 142200
rect 18970 142095 19050 142105
rect 19290 142095 19370 142105
rect 19610 142095 19690 142105
rect 19930 142095 20010 142105
rect 20250 142095 20330 142105
rect 20570 142095 20650 142105
rect 20890 142095 20970 142105
rect 21210 142095 21290 142105
rect 21530 142095 21610 142105
rect 21850 142095 21930 142105
rect 22170 142095 22250 142105
rect 22490 142095 22570 142105
rect 22810 142095 22890 142105
rect 23130 142095 23210 142105
rect 23450 142095 23530 142105
rect 23770 142095 23850 142105
rect 24090 142095 24170 142105
rect 24410 142095 24490 142105
rect 24730 142095 24810 142105
rect 25050 142095 25130 142105
rect 25370 142095 25450 142105
rect 25690 142095 25770 142105
rect 26010 142095 26090 142105
rect 26330 142095 26410 142105
rect 163590 142095 163670 142105
rect 163910 142095 163990 142105
rect 164230 142095 164310 142105
rect 164550 142095 164630 142105
rect 164870 142095 164950 142105
rect 165190 142095 165270 142105
rect 165510 142095 165590 142105
rect 165830 142095 165910 142105
rect 166150 142095 166230 142105
rect 166470 142095 166550 142105
rect 166790 142095 166870 142105
rect 167110 142095 167190 142105
rect 167430 142095 167510 142105
rect 167750 142095 167830 142105
rect 168070 142095 168150 142105
rect 168390 142095 168470 142105
rect 168710 142095 168790 142105
rect 169030 142095 169110 142105
rect 169350 142095 169430 142105
rect 169670 142095 169750 142105
rect 169990 142095 170070 142105
rect 170310 142095 170390 142105
rect 170630 142095 170710 142105
rect 170950 142095 171030 142105
rect 19050 142015 19060 142095
rect 19370 142015 19380 142095
rect 19690 142015 19700 142095
rect 20010 142015 20020 142095
rect 20330 142015 20340 142095
rect 20650 142015 20660 142095
rect 20970 142015 20980 142095
rect 21290 142015 21300 142095
rect 21610 142015 21620 142095
rect 21930 142015 21940 142095
rect 22250 142015 22260 142095
rect 22570 142015 22580 142095
rect 22890 142015 22900 142095
rect 23210 142015 23220 142095
rect 23530 142015 23540 142095
rect 23850 142015 23860 142095
rect 24170 142015 24180 142095
rect 24490 142015 24500 142095
rect 24810 142015 24820 142095
rect 25130 142015 25140 142095
rect 25450 142015 25460 142095
rect 25770 142015 25780 142095
rect 26090 142015 26100 142095
rect 26410 142015 26420 142095
rect 30360 142055 30440 142065
rect 30680 142055 30760 142065
rect 31000 142055 31080 142065
rect 31320 142055 31400 142065
rect 31640 142055 31720 142065
rect 31960 142055 32040 142065
rect 32280 142055 32360 142065
rect 32600 142055 32680 142065
rect 32920 142055 33000 142065
rect 33240 142055 33320 142065
rect 33560 142055 33640 142065
rect 33880 142055 33960 142065
rect 34200 142055 34280 142065
rect 34520 142055 34600 142065
rect 34840 142055 34920 142065
rect 35160 142055 35240 142065
rect 35480 142055 35560 142065
rect 35800 142055 35880 142065
rect 36120 142055 36200 142065
rect 36440 142055 36520 142065
rect 36760 142055 36840 142065
rect 37080 142055 37160 142065
rect 37400 142055 37480 142065
rect 37720 142055 37800 142065
rect 40180 142055 40260 142065
rect 40500 142055 40580 142065
rect 40820 142055 40900 142065
rect 41140 142055 41220 142065
rect 42560 142055 42640 142065
rect 42880 142055 42960 142065
rect 43200 142055 43280 142065
rect 43520 142055 43600 142065
rect 146400 142055 146480 142065
rect 146720 142055 146800 142065
rect 147040 142055 147120 142065
rect 147360 142055 147440 142065
rect 148780 142055 148860 142065
rect 149100 142055 149180 142065
rect 149420 142055 149500 142065
rect 149740 142055 149820 142065
rect 152200 142055 152280 142065
rect 152520 142055 152600 142065
rect 152840 142055 152920 142065
rect 153160 142055 153240 142065
rect 153480 142055 153560 142065
rect 153800 142055 153880 142065
rect 154120 142055 154200 142065
rect 154440 142055 154520 142065
rect 154760 142055 154840 142065
rect 155080 142055 155160 142065
rect 155400 142055 155480 142065
rect 155720 142055 155800 142065
rect 156040 142055 156120 142065
rect 156360 142055 156440 142065
rect 156680 142055 156760 142065
rect 157000 142055 157080 142065
rect 157320 142055 157400 142065
rect 157640 142055 157720 142065
rect 157960 142055 158040 142065
rect 158280 142055 158360 142065
rect 158600 142055 158680 142065
rect 158920 142055 159000 142065
rect 159240 142055 159320 142065
rect 159560 142055 159640 142065
rect 30440 141975 30450 142055
rect 30760 141975 30770 142055
rect 31080 141975 31090 142055
rect 31400 141975 31410 142055
rect 31720 141975 31730 142055
rect 32040 141975 32050 142055
rect 32360 141975 32370 142055
rect 32680 141975 32690 142055
rect 33000 141975 33010 142055
rect 33320 141975 33330 142055
rect 33640 141975 33650 142055
rect 33960 141975 33970 142055
rect 34280 141975 34290 142055
rect 34600 141975 34610 142055
rect 34920 141975 34930 142055
rect 35240 141975 35250 142055
rect 35560 141975 35570 142055
rect 35880 141975 35890 142055
rect 36200 141975 36210 142055
rect 36520 141975 36530 142055
rect 36840 141975 36850 142055
rect 37160 141975 37170 142055
rect 37480 141975 37490 142055
rect 37800 141975 37810 142055
rect 40260 141975 40270 142055
rect 40580 141975 40590 142055
rect 40900 141975 40910 142055
rect 41220 141975 41230 142055
rect 42640 141975 42650 142055
rect 42960 141975 42970 142055
rect 43280 141975 43290 142055
rect 43600 141975 43610 142055
rect 146480 141975 146490 142055
rect 146800 141975 146810 142055
rect 147120 141975 147130 142055
rect 147440 141975 147450 142055
rect 148860 141975 148870 142055
rect 149180 141975 149190 142055
rect 149500 141975 149510 142055
rect 149820 141975 149830 142055
rect 152280 141975 152290 142055
rect 152600 141975 152610 142055
rect 152920 141975 152930 142055
rect 153240 141975 153250 142055
rect 153560 141975 153570 142055
rect 153880 141975 153890 142055
rect 154200 141975 154210 142055
rect 154520 141975 154530 142055
rect 154840 141975 154850 142055
rect 155160 141975 155170 142055
rect 155480 141975 155490 142055
rect 155800 141975 155810 142055
rect 156120 141975 156130 142055
rect 156440 141975 156450 142055
rect 156760 141975 156770 142055
rect 157080 141975 157090 142055
rect 157400 141975 157410 142055
rect 157720 141975 157730 142055
rect 158040 141975 158050 142055
rect 158360 141975 158370 142055
rect 158680 141975 158690 142055
rect 159000 141975 159010 142055
rect 159320 141975 159330 142055
rect 159640 141975 159650 142055
rect 163670 142015 163680 142095
rect 163990 142015 164000 142095
rect 164310 142015 164320 142095
rect 164630 142015 164640 142095
rect 164950 142015 164960 142095
rect 165270 142015 165280 142095
rect 165590 142015 165600 142095
rect 165910 142015 165920 142095
rect 166230 142015 166240 142095
rect 166550 142015 166560 142095
rect 166870 142015 166880 142095
rect 167190 142015 167200 142095
rect 167510 142015 167520 142095
rect 167830 142015 167840 142095
rect 168150 142015 168160 142095
rect 168470 142015 168480 142095
rect 168790 142015 168800 142095
rect 169110 142015 169120 142095
rect 169430 142015 169440 142095
rect 169750 142015 169760 142095
rect 170070 142015 170080 142095
rect 170390 142015 170400 142095
rect 170710 142015 170720 142095
rect 171030 142015 171040 142095
rect 19130 141935 19210 141945
rect 19450 141935 19530 141945
rect 19770 141935 19850 141945
rect 20090 141935 20170 141945
rect 20410 141935 20490 141945
rect 20730 141935 20810 141945
rect 21050 141935 21130 141945
rect 21370 141935 21450 141945
rect 21690 141935 21770 141945
rect 22010 141935 22090 141945
rect 22330 141935 22410 141945
rect 22650 141935 22730 141945
rect 22970 141935 23050 141945
rect 23290 141935 23370 141945
rect 23610 141935 23690 141945
rect 23930 141935 24010 141945
rect 24250 141935 24330 141945
rect 24570 141935 24650 141945
rect 24890 141935 24970 141945
rect 25210 141935 25290 141945
rect 25530 141935 25610 141945
rect 25850 141935 25930 141945
rect 26170 141935 26250 141945
rect 163750 141935 163830 141945
rect 164070 141935 164150 141945
rect 164390 141935 164470 141945
rect 164710 141935 164790 141945
rect 165030 141935 165110 141945
rect 165350 141935 165430 141945
rect 165670 141935 165750 141945
rect 165990 141935 166070 141945
rect 166310 141935 166390 141945
rect 166630 141935 166710 141945
rect 166950 141935 167030 141945
rect 167270 141935 167350 141945
rect 167590 141935 167670 141945
rect 167910 141935 167990 141945
rect 168230 141935 168310 141945
rect 168550 141935 168630 141945
rect 168870 141935 168950 141945
rect 169190 141935 169270 141945
rect 169510 141935 169590 141945
rect 169830 141935 169910 141945
rect 170150 141935 170230 141945
rect 170470 141935 170550 141945
rect 170790 141935 170870 141945
rect 19210 141855 19220 141935
rect 19530 141855 19540 141935
rect 19850 141855 19860 141935
rect 20170 141855 20180 141935
rect 20490 141855 20500 141935
rect 20810 141855 20820 141935
rect 21130 141855 21140 141935
rect 21450 141855 21460 141935
rect 21770 141855 21780 141935
rect 22090 141855 22100 141935
rect 22410 141855 22420 141935
rect 22730 141855 22740 141935
rect 23050 141855 23060 141935
rect 23370 141855 23380 141935
rect 23690 141855 23700 141935
rect 24010 141855 24020 141935
rect 24330 141855 24340 141935
rect 24650 141855 24660 141935
rect 24970 141855 24980 141935
rect 25290 141855 25300 141935
rect 25610 141855 25620 141935
rect 25930 141855 25940 141935
rect 26250 141855 26260 141935
rect 30520 141895 30600 141905
rect 30840 141895 30920 141905
rect 31160 141895 31240 141905
rect 31480 141895 31560 141905
rect 31800 141895 31880 141905
rect 32120 141895 32200 141905
rect 32440 141895 32520 141905
rect 32760 141895 32840 141905
rect 33080 141895 33160 141905
rect 33400 141895 33480 141905
rect 33720 141895 33800 141905
rect 34040 141895 34120 141905
rect 34360 141895 34440 141905
rect 34680 141895 34760 141905
rect 35000 141895 35080 141905
rect 35320 141895 35400 141905
rect 35640 141895 35720 141905
rect 35960 141895 36040 141905
rect 36280 141895 36360 141905
rect 36600 141895 36680 141905
rect 36920 141895 37000 141905
rect 37240 141895 37320 141905
rect 37560 141895 37640 141905
rect 40340 141895 40420 141905
rect 40660 141895 40740 141905
rect 40980 141895 41060 141905
rect 42720 141895 42800 141905
rect 43040 141895 43120 141905
rect 43360 141895 43440 141905
rect 146560 141895 146640 141905
rect 146880 141895 146960 141905
rect 147200 141895 147280 141905
rect 148940 141895 149020 141905
rect 149260 141895 149340 141905
rect 149580 141895 149660 141905
rect 152360 141895 152440 141905
rect 152680 141895 152760 141905
rect 153000 141895 153080 141905
rect 153320 141895 153400 141905
rect 153640 141895 153720 141905
rect 153960 141895 154040 141905
rect 154280 141895 154360 141905
rect 154600 141895 154680 141905
rect 154920 141895 155000 141905
rect 155240 141895 155320 141905
rect 155560 141895 155640 141905
rect 155880 141895 155960 141905
rect 156200 141895 156280 141905
rect 156520 141895 156600 141905
rect 156840 141895 156920 141905
rect 157160 141895 157240 141905
rect 157480 141895 157560 141905
rect 157800 141895 157880 141905
rect 158120 141895 158200 141905
rect 158440 141895 158520 141905
rect 158760 141895 158840 141905
rect 159080 141895 159160 141905
rect 159400 141895 159480 141905
rect 30600 141815 30610 141895
rect 30920 141815 30930 141895
rect 31240 141815 31250 141895
rect 31560 141815 31570 141895
rect 31880 141815 31890 141895
rect 32200 141815 32210 141895
rect 32520 141815 32530 141895
rect 32840 141815 32850 141895
rect 33160 141815 33170 141895
rect 33480 141815 33490 141895
rect 33800 141815 33810 141895
rect 34120 141815 34130 141895
rect 34440 141815 34450 141895
rect 34760 141815 34770 141895
rect 35080 141815 35090 141895
rect 35400 141815 35410 141895
rect 35720 141815 35730 141895
rect 36040 141815 36050 141895
rect 36360 141815 36370 141895
rect 36680 141815 36690 141895
rect 37000 141815 37010 141895
rect 37320 141815 37330 141895
rect 37640 141815 37650 141895
rect 40420 141815 40430 141895
rect 40740 141815 40750 141895
rect 41060 141815 41070 141895
rect 42800 141815 42810 141895
rect 43120 141815 43130 141895
rect 43440 141815 43450 141895
rect 146640 141815 146650 141895
rect 146960 141815 146970 141895
rect 147280 141815 147290 141895
rect 149020 141815 149030 141895
rect 149340 141815 149350 141895
rect 149660 141815 149670 141895
rect 152440 141815 152450 141895
rect 152760 141815 152770 141895
rect 153080 141815 153090 141895
rect 153400 141815 153410 141895
rect 153720 141815 153730 141895
rect 154040 141815 154050 141895
rect 154360 141815 154370 141895
rect 154680 141815 154690 141895
rect 155000 141815 155010 141895
rect 155320 141815 155330 141895
rect 155640 141815 155650 141895
rect 155960 141815 155970 141895
rect 156280 141815 156290 141895
rect 156600 141815 156610 141895
rect 156920 141815 156930 141895
rect 157240 141815 157250 141895
rect 157560 141815 157570 141895
rect 157880 141815 157890 141895
rect 158200 141815 158210 141895
rect 158520 141815 158530 141895
rect 158840 141815 158850 141895
rect 159160 141815 159170 141895
rect 159480 141815 159490 141895
rect 163830 141855 163840 141935
rect 164150 141855 164160 141935
rect 164470 141855 164480 141935
rect 164790 141855 164800 141935
rect 165110 141855 165120 141935
rect 165430 141855 165440 141935
rect 165750 141855 165760 141935
rect 166070 141855 166080 141935
rect 166390 141855 166400 141935
rect 166710 141855 166720 141935
rect 167030 141855 167040 141935
rect 167350 141855 167360 141935
rect 167670 141855 167680 141935
rect 167990 141855 168000 141935
rect 168310 141855 168320 141935
rect 168630 141855 168640 141935
rect 168950 141855 168960 141935
rect 169270 141855 169280 141935
rect 169590 141855 169600 141935
rect 169910 141855 169920 141935
rect 170230 141855 170240 141935
rect 170550 141855 170560 141935
rect 170870 141855 170880 141935
rect 18970 141775 19050 141785
rect 19290 141775 19370 141785
rect 19610 141775 19690 141785
rect 19930 141775 20010 141785
rect 20250 141775 20330 141785
rect 20570 141775 20650 141785
rect 20890 141775 20970 141785
rect 21210 141775 21290 141785
rect 21530 141775 21610 141785
rect 21850 141775 21930 141785
rect 22170 141775 22250 141785
rect 22490 141775 22570 141785
rect 22810 141775 22890 141785
rect 23130 141775 23210 141785
rect 23450 141775 23530 141785
rect 23770 141775 23850 141785
rect 24090 141775 24170 141785
rect 24410 141775 24490 141785
rect 24730 141775 24810 141785
rect 25050 141775 25130 141785
rect 25370 141775 25450 141785
rect 25690 141775 25770 141785
rect 26010 141775 26090 141785
rect 26330 141775 26410 141785
rect 163590 141775 163670 141785
rect 163910 141775 163990 141785
rect 164230 141775 164310 141785
rect 164550 141775 164630 141785
rect 164870 141775 164950 141785
rect 165190 141775 165270 141785
rect 165510 141775 165590 141785
rect 165830 141775 165910 141785
rect 166150 141775 166230 141785
rect 166470 141775 166550 141785
rect 166790 141775 166870 141785
rect 167110 141775 167190 141785
rect 167430 141775 167510 141785
rect 167750 141775 167830 141785
rect 168070 141775 168150 141785
rect 168390 141775 168470 141785
rect 168710 141775 168790 141785
rect 169030 141775 169110 141785
rect 169350 141775 169430 141785
rect 169670 141775 169750 141785
rect 169990 141775 170070 141785
rect 170310 141775 170390 141785
rect 170630 141775 170710 141785
rect 170950 141775 171030 141785
rect 19050 141695 19060 141775
rect 19370 141695 19380 141775
rect 19690 141695 19700 141775
rect 20010 141695 20020 141775
rect 20330 141695 20340 141775
rect 20650 141695 20660 141775
rect 20970 141695 20980 141775
rect 21290 141695 21300 141775
rect 21610 141695 21620 141775
rect 21930 141695 21940 141775
rect 22250 141695 22260 141775
rect 22570 141695 22580 141775
rect 22890 141695 22900 141775
rect 23210 141695 23220 141775
rect 23530 141695 23540 141775
rect 23850 141695 23860 141775
rect 24170 141695 24180 141775
rect 24490 141695 24500 141775
rect 24810 141695 24820 141775
rect 25130 141695 25140 141775
rect 25450 141695 25460 141775
rect 25770 141695 25780 141775
rect 26090 141695 26100 141775
rect 26410 141695 26420 141775
rect 30360 141735 30440 141745
rect 30680 141735 30760 141745
rect 31000 141735 31080 141745
rect 31320 141735 31400 141745
rect 31640 141735 31720 141745
rect 31960 141735 32040 141745
rect 32280 141735 32360 141745
rect 32600 141735 32680 141745
rect 32920 141735 33000 141745
rect 33240 141735 33320 141745
rect 33560 141735 33640 141745
rect 33880 141735 33960 141745
rect 34200 141735 34280 141745
rect 34520 141735 34600 141745
rect 34840 141735 34920 141745
rect 35160 141735 35240 141745
rect 35480 141735 35560 141745
rect 35800 141735 35880 141745
rect 36120 141735 36200 141745
rect 36440 141735 36520 141745
rect 36760 141735 36840 141745
rect 37080 141735 37160 141745
rect 37400 141735 37480 141745
rect 37720 141735 37800 141745
rect 40180 141735 40260 141745
rect 40500 141735 40580 141745
rect 40820 141735 40900 141745
rect 41140 141735 41220 141745
rect 42560 141735 42640 141745
rect 42880 141735 42960 141745
rect 43200 141735 43280 141745
rect 43520 141735 43600 141745
rect 146400 141735 146480 141745
rect 146720 141735 146800 141745
rect 147040 141735 147120 141745
rect 147360 141735 147440 141745
rect 148780 141735 148860 141745
rect 149100 141735 149180 141745
rect 149420 141735 149500 141745
rect 149740 141735 149820 141745
rect 152200 141735 152280 141745
rect 152520 141735 152600 141745
rect 152840 141735 152920 141745
rect 153160 141735 153240 141745
rect 153480 141735 153560 141745
rect 153800 141735 153880 141745
rect 154120 141735 154200 141745
rect 154440 141735 154520 141745
rect 154760 141735 154840 141745
rect 155080 141735 155160 141745
rect 155400 141735 155480 141745
rect 155720 141735 155800 141745
rect 156040 141735 156120 141745
rect 156360 141735 156440 141745
rect 156680 141735 156760 141745
rect 157000 141735 157080 141745
rect 157320 141735 157400 141745
rect 157640 141735 157720 141745
rect 157960 141735 158040 141745
rect 158280 141735 158360 141745
rect 158600 141735 158680 141745
rect 158920 141735 159000 141745
rect 159240 141735 159320 141745
rect 159560 141735 159640 141745
rect 30440 141655 30450 141735
rect 30760 141655 30770 141735
rect 31080 141655 31090 141735
rect 31400 141655 31410 141735
rect 31720 141655 31730 141735
rect 32040 141655 32050 141735
rect 32360 141655 32370 141735
rect 32680 141655 32690 141735
rect 33000 141655 33010 141735
rect 33320 141655 33330 141735
rect 33640 141655 33650 141735
rect 33960 141655 33970 141735
rect 34280 141655 34290 141735
rect 34600 141655 34610 141735
rect 34920 141655 34930 141735
rect 35240 141655 35250 141735
rect 35560 141655 35570 141735
rect 35880 141655 35890 141735
rect 36200 141655 36210 141735
rect 36520 141655 36530 141735
rect 36840 141655 36850 141735
rect 37160 141655 37170 141735
rect 37480 141655 37490 141735
rect 37800 141655 37810 141735
rect 40260 141655 40270 141735
rect 40580 141655 40590 141735
rect 40900 141655 40910 141735
rect 41220 141655 41230 141735
rect 42640 141655 42650 141735
rect 42960 141655 42970 141735
rect 43280 141655 43290 141735
rect 43600 141655 43610 141735
rect 146480 141655 146490 141735
rect 146800 141655 146810 141735
rect 147120 141655 147130 141735
rect 147440 141655 147450 141735
rect 148860 141655 148870 141735
rect 149180 141655 149190 141735
rect 149500 141655 149510 141735
rect 149820 141655 149830 141735
rect 152280 141655 152290 141735
rect 152600 141655 152610 141735
rect 152920 141655 152930 141735
rect 153240 141655 153250 141735
rect 153560 141655 153570 141735
rect 153880 141655 153890 141735
rect 154200 141655 154210 141735
rect 154520 141655 154530 141735
rect 154840 141655 154850 141735
rect 155160 141655 155170 141735
rect 155480 141655 155490 141735
rect 155800 141655 155810 141735
rect 156120 141655 156130 141735
rect 156440 141655 156450 141735
rect 156760 141655 156770 141735
rect 157080 141655 157090 141735
rect 157400 141655 157410 141735
rect 157720 141655 157730 141735
rect 158040 141655 158050 141735
rect 158360 141655 158370 141735
rect 158680 141655 158690 141735
rect 159000 141655 159010 141735
rect 159320 141655 159330 141735
rect 159640 141655 159650 141735
rect 163670 141695 163680 141775
rect 163990 141695 164000 141775
rect 164310 141695 164320 141775
rect 164630 141695 164640 141775
rect 164950 141695 164960 141775
rect 165270 141695 165280 141775
rect 165590 141695 165600 141775
rect 165910 141695 165920 141775
rect 166230 141695 166240 141775
rect 166550 141695 166560 141775
rect 166870 141695 166880 141775
rect 167190 141695 167200 141775
rect 167510 141695 167520 141775
rect 167830 141695 167840 141775
rect 168150 141695 168160 141775
rect 168470 141695 168480 141775
rect 168790 141695 168800 141775
rect 169110 141695 169120 141775
rect 169430 141695 169440 141775
rect 169750 141695 169760 141775
rect 170070 141695 170080 141775
rect 170390 141695 170400 141775
rect 170710 141695 170720 141775
rect 171030 141695 171040 141775
rect 18900 141515 26700 141620
rect 30200 141515 38000 141620
rect 40000 141515 41660 141620
rect 42300 141515 43960 141620
rect 146040 141515 147700 141620
rect 148340 141515 150000 141620
rect 152000 141515 159800 141620
rect 163300 141515 171100 141620
rect 18980 141440 19060 141450
rect 19160 141440 19240 141450
rect 19340 141440 19420 141450
rect 19520 141440 19600 141450
rect 19700 141440 19780 141450
rect 19880 141440 19960 141450
rect 20060 141440 20140 141450
rect 20240 141440 20320 141450
rect 20420 141440 20500 141450
rect 20600 141440 20680 141450
rect 20780 141440 20860 141450
rect 20960 141440 21040 141450
rect 21140 141440 21220 141450
rect 21320 141440 21400 141450
rect 21500 141440 21580 141450
rect 21680 141440 21760 141450
rect 21860 141440 21940 141450
rect 22040 141440 22120 141450
rect 22220 141440 22300 141450
rect 22400 141440 22480 141450
rect 22580 141440 22660 141450
rect 22760 141440 22840 141450
rect 22940 141440 23020 141450
rect 23120 141440 23200 141450
rect 23300 141440 23380 141450
rect 23480 141440 23560 141450
rect 23660 141440 23740 141450
rect 23840 141440 23920 141450
rect 24020 141440 24100 141450
rect 24200 141440 24280 141450
rect 24380 141440 24460 141450
rect 24560 141440 24640 141450
rect 24740 141440 24820 141450
rect 24920 141440 25000 141450
rect 25100 141440 25180 141450
rect 25280 141440 25360 141450
rect 25460 141440 25540 141450
rect 25640 141440 25720 141450
rect 25820 141440 25900 141450
rect 26000 141440 26080 141450
rect 26180 141440 26260 141450
rect 26360 141440 26440 141450
rect 26540 141440 26620 141450
rect 30280 141440 30360 141450
rect 30460 141440 30540 141450
rect 30640 141440 30720 141450
rect 30820 141440 30900 141450
rect 31000 141440 31080 141450
rect 31180 141440 31260 141450
rect 31360 141440 31440 141450
rect 31540 141440 31620 141450
rect 31720 141440 31800 141450
rect 31900 141440 31980 141450
rect 32080 141440 32160 141450
rect 32260 141440 32340 141450
rect 32440 141440 32520 141450
rect 32620 141440 32700 141450
rect 32800 141440 32880 141450
rect 32980 141440 33060 141450
rect 33160 141440 33240 141450
rect 33340 141440 33420 141450
rect 33520 141440 33600 141450
rect 33700 141440 33780 141450
rect 33880 141440 33960 141450
rect 34060 141440 34140 141450
rect 34240 141440 34320 141450
rect 34420 141440 34500 141450
rect 34600 141440 34680 141450
rect 34780 141440 34860 141450
rect 34960 141440 35040 141450
rect 35140 141440 35220 141450
rect 35320 141440 35400 141450
rect 35500 141440 35580 141450
rect 35680 141440 35760 141450
rect 35860 141440 35940 141450
rect 36040 141440 36120 141450
rect 36220 141440 36300 141450
rect 36400 141440 36480 141450
rect 36580 141440 36660 141450
rect 36760 141440 36840 141450
rect 36940 141440 37020 141450
rect 37120 141440 37200 141450
rect 37300 141440 37380 141450
rect 37480 141440 37560 141450
rect 37660 141440 37740 141450
rect 37840 141440 37920 141450
rect 40060 141440 40140 141450
rect 40200 141440 40280 141450
rect 40340 141440 40420 141450
rect 40480 141440 40560 141450
rect 40620 141440 40700 141450
rect 40760 141440 40840 141450
rect 40900 141440 40980 141450
rect 41040 141440 41120 141450
rect 41180 141440 41260 141450
rect 41320 141440 41400 141450
rect 42360 141440 42440 141450
rect 42500 141440 42580 141450
rect 42640 141440 42720 141450
rect 42780 141440 42860 141450
rect 42920 141440 43000 141450
rect 43060 141440 43140 141450
rect 43200 141440 43280 141450
rect 43340 141440 43420 141450
rect 43480 141440 43560 141450
rect 43620 141440 43700 141450
rect 146300 141440 146380 141450
rect 146440 141440 146520 141450
rect 146580 141440 146660 141450
rect 146720 141440 146800 141450
rect 146860 141440 146940 141450
rect 147000 141440 147080 141450
rect 147140 141440 147220 141450
rect 147280 141440 147360 141450
rect 147420 141440 147500 141450
rect 147560 141440 147640 141450
rect 19060 141360 19070 141440
rect 19240 141360 19250 141440
rect 19420 141360 19430 141440
rect 19600 141360 19610 141440
rect 19780 141360 19790 141440
rect 19960 141360 19970 141440
rect 20140 141360 20150 141440
rect 20320 141360 20330 141440
rect 20500 141360 20510 141440
rect 20680 141360 20690 141440
rect 20860 141360 20870 141440
rect 21040 141360 21050 141440
rect 21220 141360 21230 141440
rect 21400 141360 21410 141440
rect 21580 141360 21590 141440
rect 21760 141360 21770 141440
rect 21940 141360 21950 141440
rect 22120 141360 22130 141440
rect 22300 141360 22310 141440
rect 22480 141360 22490 141440
rect 22660 141360 22670 141440
rect 22840 141360 22850 141440
rect 23020 141360 23030 141440
rect 23200 141360 23210 141440
rect 23380 141360 23390 141440
rect 23560 141360 23570 141440
rect 23740 141360 23750 141440
rect 23920 141360 23930 141440
rect 24100 141360 24110 141440
rect 24280 141360 24290 141440
rect 24460 141360 24470 141440
rect 24640 141360 24650 141440
rect 24820 141360 24830 141440
rect 25000 141360 25010 141440
rect 25180 141360 25190 141440
rect 25360 141360 25370 141440
rect 25540 141360 25550 141440
rect 25720 141360 25730 141440
rect 25900 141360 25910 141440
rect 26080 141360 26090 141440
rect 26260 141360 26270 141440
rect 26440 141360 26450 141440
rect 26620 141360 26630 141440
rect 30360 141360 30370 141440
rect 30540 141360 30550 141440
rect 30720 141360 30730 141440
rect 30900 141360 30910 141440
rect 31080 141360 31090 141440
rect 31260 141360 31270 141440
rect 31440 141360 31450 141440
rect 31620 141360 31630 141440
rect 31800 141360 31810 141440
rect 31980 141360 31990 141440
rect 32160 141360 32170 141440
rect 32340 141360 32350 141440
rect 32520 141360 32530 141440
rect 32700 141360 32710 141440
rect 32880 141360 32890 141440
rect 33060 141360 33070 141440
rect 33240 141360 33250 141440
rect 33420 141360 33430 141440
rect 33600 141360 33610 141440
rect 33780 141360 33790 141440
rect 33960 141360 33970 141440
rect 34140 141360 34150 141440
rect 34320 141360 34330 141440
rect 34500 141360 34510 141440
rect 34680 141360 34690 141440
rect 34860 141360 34870 141440
rect 35040 141360 35050 141440
rect 35220 141360 35230 141440
rect 35400 141360 35410 141440
rect 35580 141360 35590 141440
rect 35760 141360 35770 141440
rect 35940 141360 35950 141440
rect 36120 141360 36130 141440
rect 36300 141360 36310 141440
rect 36480 141360 36490 141440
rect 36660 141360 36670 141440
rect 36840 141360 36850 141440
rect 37020 141360 37030 141440
rect 37200 141360 37210 141440
rect 37380 141360 37390 141440
rect 37560 141360 37570 141440
rect 37740 141360 37750 141440
rect 37920 141360 37930 141440
rect 40140 141360 40150 141440
rect 40280 141360 40290 141440
rect 40420 141360 40430 141440
rect 40560 141360 40570 141440
rect 40700 141360 40710 141440
rect 40840 141360 40850 141440
rect 40980 141360 40990 141440
rect 41120 141360 41130 141440
rect 41260 141360 41270 141440
rect 41400 141360 41410 141440
rect 42440 141360 42450 141440
rect 42580 141360 42590 141440
rect 42720 141360 42730 141440
rect 42860 141360 42870 141440
rect 43000 141360 43010 141440
rect 43140 141360 43150 141440
rect 43280 141360 43290 141440
rect 43420 141360 43430 141440
rect 43560 141360 43570 141440
rect 43700 141360 43710 141440
rect 146380 141360 146390 141440
rect 146520 141360 146530 141440
rect 146660 141360 146670 141440
rect 146800 141360 146810 141440
rect 146940 141360 146950 141440
rect 147080 141360 147090 141440
rect 147220 141360 147230 141440
rect 147360 141360 147370 141440
rect 147500 141360 147510 141440
rect 147640 141360 147650 141440
rect 28850 141315 28930 141325
rect 29010 141315 29090 141325
rect 29170 141315 29250 141325
rect 29330 141315 29410 141325
rect 29490 141315 29570 141325
rect 18980 141290 19060 141300
rect 19160 141290 19240 141300
rect 19340 141290 19420 141300
rect 19520 141290 19600 141300
rect 19700 141290 19780 141300
rect 19880 141290 19960 141300
rect 20060 141290 20140 141300
rect 20240 141290 20320 141300
rect 20420 141290 20500 141300
rect 20600 141290 20680 141300
rect 20780 141290 20860 141300
rect 20960 141290 21040 141300
rect 21140 141290 21220 141300
rect 21320 141290 21400 141300
rect 21500 141290 21580 141300
rect 21680 141290 21760 141300
rect 21860 141290 21940 141300
rect 22040 141290 22120 141300
rect 22220 141290 22300 141300
rect 22400 141290 22480 141300
rect 22580 141290 22660 141300
rect 22760 141290 22840 141300
rect 22940 141290 23020 141300
rect 23120 141290 23200 141300
rect 23300 141290 23380 141300
rect 23480 141290 23560 141300
rect 23660 141290 23740 141300
rect 23840 141290 23920 141300
rect 24020 141290 24100 141300
rect 24200 141290 24280 141300
rect 24380 141290 24460 141300
rect 24560 141290 24640 141300
rect 24740 141290 24820 141300
rect 24920 141290 25000 141300
rect 25100 141290 25180 141300
rect 25280 141290 25360 141300
rect 25460 141290 25540 141300
rect 25640 141290 25720 141300
rect 25820 141290 25900 141300
rect 26000 141290 26080 141300
rect 26180 141290 26260 141300
rect 26360 141290 26440 141300
rect 26540 141290 26620 141300
rect 19060 141210 19070 141290
rect 19240 141210 19250 141290
rect 19420 141210 19430 141290
rect 19600 141210 19610 141290
rect 19780 141210 19790 141290
rect 19960 141210 19970 141290
rect 20140 141210 20150 141290
rect 20320 141210 20330 141290
rect 20500 141210 20510 141290
rect 20680 141210 20690 141290
rect 20860 141210 20870 141290
rect 21040 141210 21050 141290
rect 21220 141210 21230 141290
rect 21400 141210 21410 141290
rect 21580 141210 21590 141290
rect 21760 141210 21770 141290
rect 21940 141210 21950 141290
rect 22120 141210 22130 141290
rect 22300 141210 22310 141290
rect 22480 141210 22490 141290
rect 22660 141210 22670 141290
rect 22840 141210 22850 141290
rect 23020 141210 23030 141290
rect 23200 141210 23210 141290
rect 23380 141210 23390 141290
rect 23560 141210 23570 141290
rect 23740 141210 23750 141290
rect 23920 141210 23930 141290
rect 24100 141210 24110 141290
rect 24280 141210 24290 141290
rect 24460 141210 24470 141290
rect 24640 141210 24650 141290
rect 24820 141210 24830 141290
rect 25000 141210 25010 141290
rect 25180 141210 25190 141290
rect 25360 141210 25370 141290
rect 25540 141210 25550 141290
rect 25720 141210 25730 141290
rect 25900 141210 25910 141290
rect 26080 141210 26090 141290
rect 26260 141210 26270 141290
rect 26440 141210 26450 141290
rect 26620 141210 26630 141290
rect 28930 141235 28940 141315
rect 29010 141235 29020 141315
rect 29090 141235 29100 141315
rect 29170 141235 29180 141315
rect 29250 141235 29260 141315
rect 29330 141235 29340 141315
rect 29410 141235 29420 141315
rect 29490 141235 29500 141315
rect 29570 141235 29580 141315
rect 148340 141300 150000 141500
rect 152080 141440 152160 141450
rect 152260 141440 152340 141450
rect 152440 141440 152520 141450
rect 152620 141440 152700 141450
rect 152800 141440 152880 141450
rect 152980 141440 153060 141450
rect 153160 141440 153240 141450
rect 153340 141440 153420 141450
rect 153520 141440 153600 141450
rect 153700 141440 153780 141450
rect 153880 141440 153960 141450
rect 154060 141440 154140 141450
rect 154240 141440 154320 141450
rect 154420 141440 154500 141450
rect 154600 141440 154680 141450
rect 154780 141440 154860 141450
rect 154960 141440 155040 141450
rect 155140 141440 155220 141450
rect 155320 141440 155400 141450
rect 155500 141440 155580 141450
rect 155680 141440 155760 141450
rect 155860 141440 155940 141450
rect 156040 141440 156120 141450
rect 156220 141440 156300 141450
rect 156400 141440 156480 141450
rect 156580 141440 156660 141450
rect 156760 141440 156840 141450
rect 156940 141440 157020 141450
rect 157120 141440 157200 141450
rect 157300 141440 157380 141450
rect 157480 141440 157560 141450
rect 157660 141440 157740 141450
rect 157840 141440 157920 141450
rect 158020 141440 158100 141450
rect 158200 141440 158280 141450
rect 158380 141440 158460 141450
rect 158560 141440 158640 141450
rect 158740 141440 158820 141450
rect 158920 141440 159000 141450
rect 159100 141440 159180 141450
rect 159280 141440 159360 141450
rect 159460 141440 159540 141450
rect 159640 141440 159720 141450
rect 163380 141440 163460 141450
rect 163560 141440 163640 141450
rect 163740 141440 163820 141450
rect 163920 141440 164000 141450
rect 164100 141440 164180 141450
rect 164280 141440 164360 141450
rect 164460 141440 164540 141450
rect 164640 141440 164720 141450
rect 164820 141440 164900 141450
rect 165000 141440 165080 141450
rect 165180 141440 165260 141450
rect 165360 141440 165440 141450
rect 165540 141440 165620 141450
rect 165720 141440 165800 141450
rect 165900 141440 165980 141450
rect 166080 141440 166160 141450
rect 166260 141440 166340 141450
rect 166440 141440 166520 141450
rect 166620 141440 166700 141450
rect 166800 141440 166880 141450
rect 166980 141440 167060 141450
rect 167160 141440 167240 141450
rect 167340 141440 167420 141450
rect 167520 141440 167600 141450
rect 167700 141440 167780 141450
rect 167880 141440 167960 141450
rect 168060 141440 168140 141450
rect 168240 141440 168320 141450
rect 168420 141440 168500 141450
rect 168600 141440 168680 141450
rect 168780 141440 168860 141450
rect 168960 141440 169040 141450
rect 169140 141440 169220 141450
rect 169320 141440 169400 141450
rect 169500 141440 169580 141450
rect 169680 141440 169760 141450
rect 169860 141440 169940 141450
rect 170040 141440 170120 141450
rect 170220 141440 170300 141450
rect 170400 141440 170480 141450
rect 170580 141440 170660 141450
rect 170760 141440 170840 141450
rect 170940 141440 171020 141450
rect 152160 141360 152170 141440
rect 152340 141360 152350 141440
rect 152520 141360 152530 141440
rect 152700 141360 152710 141440
rect 152880 141360 152890 141440
rect 153060 141360 153070 141440
rect 153240 141360 153250 141440
rect 153420 141360 153430 141440
rect 153600 141360 153610 141440
rect 153780 141360 153790 141440
rect 153960 141360 153970 141440
rect 154140 141360 154150 141440
rect 154320 141360 154330 141440
rect 154500 141360 154510 141440
rect 154680 141360 154690 141440
rect 154860 141360 154870 141440
rect 155040 141360 155050 141440
rect 155220 141360 155230 141440
rect 155400 141360 155410 141440
rect 155580 141360 155590 141440
rect 155760 141360 155770 141440
rect 155940 141360 155950 141440
rect 156120 141360 156130 141440
rect 156300 141360 156310 141440
rect 156480 141360 156490 141440
rect 156660 141360 156670 141440
rect 156840 141360 156850 141440
rect 157020 141360 157030 141440
rect 157200 141360 157210 141440
rect 157380 141360 157390 141440
rect 157560 141360 157570 141440
rect 157740 141360 157750 141440
rect 157920 141360 157930 141440
rect 158100 141360 158110 141440
rect 158280 141360 158290 141440
rect 158460 141360 158470 141440
rect 158640 141360 158650 141440
rect 158820 141360 158830 141440
rect 159000 141360 159010 141440
rect 159180 141360 159190 141440
rect 159360 141360 159370 141440
rect 159540 141360 159550 141440
rect 159720 141360 159730 141440
rect 163460 141360 163470 141440
rect 163640 141360 163650 141440
rect 163820 141360 163830 141440
rect 164000 141360 164010 141440
rect 164180 141360 164190 141440
rect 164360 141360 164370 141440
rect 164540 141360 164550 141440
rect 164720 141360 164730 141440
rect 164900 141360 164910 141440
rect 165080 141360 165090 141440
rect 165260 141360 165270 141440
rect 165440 141360 165450 141440
rect 165620 141360 165630 141440
rect 165800 141360 165810 141440
rect 165980 141360 165990 141440
rect 166160 141360 166170 141440
rect 166340 141360 166350 141440
rect 166520 141360 166530 141440
rect 166700 141360 166710 141440
rect 166880 141360 166890 141440
rect 167060 141360 167070 141440
rect 167240 141360 167250 141440
rect 167420 141360 167430 141440
rect 167600 141360 167610 141440
rect 167780 141360 167790 141440
rect 167960 141360 167970 141440
rect 168140 141360 168150 141440
rect 168320 141360 168330 141440
rect 168500 141360 168510 141440
rect 168680 141360 168690 141440
rect 168860 141360 168870 141440
rect 169040 141360 169050 141440
rect 169220 141360 169230 141440
rect 169400 141360 169410 141440
rect 169580 141360 169590 141440
rect 169760 141360 169770 141440
rect 169940 141360 169950 141440
rect 170120 141360 170130 141440
rect 170300 141360 170310 141440
rect 170480 141360 170490 141440
rect 170660 141360 170670 141440
rect 170840 141360 170850 141440
rect 171020 141360 171030 141440
rect 161885 141345 161965 141355
rect 162065 141345 162145 141355
rect 162245 141345 162325 141355
rect 162425 141345 162505 141355
rect 162605 141345 162685 141355
rect 30280 141290 30360 141300
rect 30460 141290 30540 141300
rect 30640 141290 30720 141300
rect 30820 141290 30900 141300
rect 31000 141290 31080 141300
rect 31180 141290 31260 141300
rect 31360 141290 31440 141300
rect 31540 141290 31620 141300
rect 31720 141290 31800 141300
rect 31900 141290 31980 141300
rect 32080 141290 32160 141300
rect 32260 141290 32340 141300
rect 32440 141290 32520 141300
rect 32620 141290 32700 141300
rect 32800 141290 32880 141300
rect 32980 141290 33060 141300
rect 33160 141290 33240 141300
rect 33340 141290 33420 141300
rect 33520 141290 33600 141300
rect 33700 141290 33780 141300
rect 33880 141290 33960 141300
rect 34060 141290 34140 141300
rect 34240 141290 34320 141300
rect 34420 141290 34500 141300
rect 34600 141290 34680 141300
rect 34780 141290 34860 141300
rect 34960 141290 35040 141300
rect 35140 141290 35220 141300
rect 35320 141290 35400 141300
rect 35500 141290 35580 141300
rect 35680 141290 35760 141300
rect 35860 141290 35940 141300
rect 36040 141290 36120 141300
rect 36220 141290 36300 141300
rect 36400 141290 36480 141300
rect 36580 141290 36660 141300
rect 36760 141290 36840 141300
rect 36940 141290 37020 141300
rect 37120 141290 37200 141300
rect 37300 141290 37380 141300
rect 37480 141290 37560 141300
rect 37660 141290 37740 141300
rect 37840 141290 37920 141300
rect 30360 141210 30370 141290
rect 30540 141210 30550 141290
rect 30720 141210 30730 141290
rect 30900 141210 30910 141290
rect 31080 141210 31090 141290
rect 31260 141210 31270 141290
rect 31440 141210 31450 141290
rect 31620 141210 31630 141290
rect 31800 141210 31810 141290
rect 31980 141210 31990 141290
rect 32160 141210 32170 141290
rect 32340 141210 32350 141290
rect 32520 141210 32530 141290
rect 32700 141210 32710 141290
rect 32880 141210 32890 141290
rect 33060 141210 33070 141290
rect 33240 141210 33250 141290
rect 33420 141210 33430 141290
rect 33600 141210 33610 141290
rect 33780 141210 33790 141290
rect 33960 141210 33970 141290
rect 34140 141210 34150 141290
rect 34320 141210 34330 141290
rect 34500 141210 34510 141290
rect 34680 141210 34690 141290
rect 34860 141210 34870 141290
rect 35040 141210 35050 141290
rect 35220 141210 35230 141290
rect 35400 141210 35410 141290
rect 35580 141210 35590 141290
rect 35760 141210 35770 141290
rect 35940 141210 35950 141290
rect 36120 141210 36130 141290
rect 36300 141210 36310 141290
rect 36480 141210 36490 141290
rect 36660 141210 36670 141290
rect 36840 141210 36850 141290
rect 37020 141210 37030 141290
rect 37200 141210 37210 141290
rect 37380 141210 37390 141290
rect 37560 141210 37570 141290
rect 37740 141210 37750 141290
rect 37920 141210 37930 141290
rect 40060 141190 40120 141220
rect 41540 141190 41600 141220
rect 42360 141190 42420 141220
rect 43840 141190 43900 141220
rect 146100 141150 146160 141180
rect 147580 141150 147640 141180
rect 148400 141150 148460 141180
rect 40060 141070 40120 141100
rect 41540 141070 41600 141100
rect 42360 141070 42420 141100
rect 43840 141070 43900 141100
rect 146100 141030 146160 141060
rect 147580 141030 147640 141060
rect 148400 141030 148460 141060
rect 40060 140950 40120 140980
rect 41540 140950 41600 140980
rect 42360 140950 42420 140980
rect 43840 140950 43900 140980
rect 19130 140910 19160 140940
rect 19250 140910 19280 140940
rect 26420 140910 26450 140940
rect 26540 140910 26570 140940
rect 30420 140910 30450 140940
rect 30540 140910 30570 140940
rect 37720 140910 37750 140940
rect 37840 140910 37870 140940
rect 146100 140910 146160 140940
rect 147580 140910 147640 140940
rect 148400 140910 148460 140940
rect 19010 140880 19070 140910
rect 19130 140880 19190 140910
rect 19250 140880 19310 140910
rect 26300 140880 26360 140910
rect 26420 140880 26480 140910
rect 26540 140880 26600 140910
rect 30300 140880 30360 140910
rect 30420 140880 30480 140910
rect 30540 140880 30600 140910
rect 37600 140880 37660 140910
rect 37720 140880 37780 140910
rect 37840 140880 37900 140910
rect 40060 140830 40120 140860
rect 41540 140830 41600 140860
rect 42360 140830 42420 140860
rect 43840 140830 43900 140860
rect 19130 140790 19160 140820
rect 19250 140790 19280 140820
rect 26420 140790 26450 140820
rect 26540 140790 26570 140820
rect 30420 140790 30450 140820
rect 30540 140790 30570 140820
rect 37720 140790 37750 140820
rect 37840 140790 37870 140820
rect 146100 140790 146160 140820
rect 147580 140790 147640 140820
rect 148400 140790 148460 140820
rect 19010 140780 19070 140790
rect 19130 140780 19190 140790
rect 19250 140780 19310 140790
rect 26300 140780 26360 140790
rect 26420 140780 26480 140790
rect 26540 140780 26600 140790
rect 30300 140780 30360 140790
rect 30420 140780 30480 140790
rect 30540 140780 30600 140790
rect 37600 140780 37660 140790
rect 37720 140780 37780 140790
rect 37840 140780 37900 140790
rect 148520 140780 148790 141300
rect 149820 140780 150000 141300
rect 152080 141290 152160 141300
rect 152260 141290 152340 141300
rect 152440 141290 152520 141300
rect 152620 141290 152700 141300
rect 152800 141290 152880 141300
rect 152980 141290 153060 141300
rect 153160 141290 153240 141300
rect 153340 141290 153420 141300
rect 153520 141290 153600 141300
rect 153700 141290 153780 141300
rect 153880 141290 153960 141300
rect 154060 141290 154140 141300
rect 154240 141290 154320 141300
rect 154420 141290 154500 141300
rect 154600 141290 154680 141300
rect 154780 141290 154860 141300
rect 154960 141290 155040 141300
rect 155140 141290 155220 141300
rect 155320 141290 155400 141300
rect 155500 141290 155580 141300
rect 155680 141290 155760 141300
rect 155860 141290 155940 141300
rect 156040 141290 156120 141300
rect 156220 141290 156300 141300
rect 156400 141290 156480 141300
rect 156580 141290 156660 141300
rect 156760 141290 156840 141300
rect 156940 141290 157020 141300
rect 157120 141290 157200 141300
rect 157300 141290 157380 141300
rect 157480 141290 157560 141300
rect 157660 141290 157740 141300
rect 157840 141290 157920 141300
rect 158020 141290 158100 141300
rect 158200 141290 158280 141300
rect 158380 141290 158460 141300
rect 158560 141290 158640 141300
rect 158740 141290 158820 141300
rect 158920 141290 159000 141300
rect 159100 141290 159180 141300
rect 159280 141290 159360 141300
rect 159460 141290 159540 141300
rect 159640 141290 159720 141300
rect 152160 141210 152170 141290
rect 152340 141210 152350 141290
rect 152520 141210 152530 141290
rect 152700 141210 152710 141290
rect 152880 141210 152890 141290
rect 153060 141210 153070 141290
rect 153240 141210 153250 141290
rect 153420 141210 153430 141290
rect 153600 141210 153610 141290
rect 153780 141210 153790 141290
rect 153960 141210 153970 141290
rect 154140 141210 154150 141290
rect 154320 141210 154330 141290
rect 154500 141210 154510 141290
rect 154680 141210 154690 141290
rect 154860 141210 154870 141290
rect 155040 141210 155050 141290
rect 155220 141210 155230 141290
rect 155400 141210 155410 141290
rect 155580 141210 155590 141290
rect 155760 141210 155770 141290
rect 155940 141210 155950 141290
rect 156120 141210 156130 141290
rect 156300 141210 156310 141290
rect 156480 141210 156490 141290
rect 156660 141210 156670 141290
rect 156840 141210 156850 141290
rect 157020 141210 157030 141290
rect 157200 141210 157210 141290
rect 157380 141210 157390 141290
rect 157560 141210 157570 141290
rect 157740 141210 157750 141290
rect 157920 141210 157930 141290
rect 158100 141210 158110 141290
rect 158280 141210 158290 141290
rect 158460 141210 158470 141290
rect 158640 141210 158650 141290
rect 158820 141210 158830 141290
rect 159000 141210 159010 141290
rect 159180 141210 159190 141290
rect 159360 141210 159370 141290
rect 159540 141210 159550 141290
rect 159720 141210 159730 141290
rect 161965 141265 161975 141345
rect 162145 141265 162155 141345
rect 162325 141265 162335 141345
rect 162505 141265 162515 141345
rect 162685 141265 162695 141345
rect 163380 141290 163460 141300
rect 163560 141290 163640 141300
rect 163740 141290 163820 141300
rect 163920 141290 164000 141300
rect 164100 141290 164180 141300
rect 164280 141290 164360 141300
rect 164460 141290 164540 141300
rect 164640 141290 164720 141300
rect 164820 141290 164900 141300
rect 165000 141290 165080 141300
rect 165180 141290 165260 141300
rect 165360 141290 165440 141300
rect 165540 141290 165620 141300
rect 165720 141290 165800 141300
rect 165900 141290 165980 141300
rect 166080 141290 166160 141300
rect 166260 141290 166340 141300
rect 166440 141290 166520 141300
rect 166620 141290 166700 141300
rect 166800 141290 166880 141300
rect 166980 141290 167060 141300
rect 167160 141290 167240 141300
rect 167340 141290 167420 141300
rect 167520 141290 167600 141300
rect 167700 141290 167780 141300
rect 167880 141290 167960 141300
rect 168060 141290 168140 141300
rect 168240 141290 168320 141300
rect 168420 141290 168500 141300
rect 168600 141290 168680 141300
rect 168780 141290 168860 141300
rect 168960 141290 169040 141300
rect 169140 141290 169220 141300
rect 169320 141290 169400 141300
rect 169500 141290 169580 141300
rect 169680 141290 169760 141300
rect 169860 141290 169940 141300
rect 170040 141290 170120 141300
rect 170220 141290 170300 141300
rect 170400 141290 170480 141300
rect 170580 141290 170660 141300
rect 170760 141290 170840 141300
rect 170940 141290 171020 141300
rect 163460 141210 163470 141290
rect 163640 141210 163650 141290
rect 163820 141210 163830 141290
rect 164000 141210 164010 141290
rect 164180 141210 164190 141290
rect 164360 141210 164370 141290
rect 164540 141210 164550 141290
rect 164720 141210 164730 141290
rect 164900 141210 164910 141290
rect 165080 141210 165090 141290
rect 165260 141210 165270 141290
rect 165440 141210 165450 141290
rect 165620 141210 165630 141290
rect 165800 141210 165810 141290
rect 165980 141210 165990 141290
rect 166160 141210 166170 141290
rect 166340 141210 166350 141290
rect 166520 141210 166530 141290
rect 166700 141210 166710 141290
rect 166880 141210 166890 141290
rect 167060 141210 167070 141290
rect 167240 141210 167250 141290
rect 167420 141210 167430 141290
rect 167600 141210 167610 141290
rect 167780 141210 167790 141290
rect 167960 141210 167970 141290
rect 168140 141210 168150 141290
rect 168320 141210 168330 141290
rect 168500 141210 168510 141290
rect 168680 141210 168690 141290
rect 168860 141210 168870 141290
rect 169040 141210 169050 141290
rect 169220 141210 169230 141290
rect 169400 141210 169410 141290
rect 169580 141210 169590 141290
rect 169760 141210 169770 141290
rect 169940 141210 169950 141290
rect 170120 141210 170130 141290
rect 170300 141210 170310 141290
rect 170480 141210 170490 141290
rect 170660 141210 170670 141290
rect 170840 141210 170850 141290
rect 171020 141210 171030 141290
rect 161885 141165 161965 141175
rect 162065 141165 162145 141175
rect 162245 141165 162325 141175
rect 162425 141165 162505 141175
rect 162605 141165 162685 141175
rect 152080 141140 152160 141150
rect 152260 141140 152340 141150
rect 152440 141140 152520 141150
rect 152620 141140 152700 141150
rect 152800 141140 152880 141150
rect 152980 141140 153060 141150
rect 153160 141140 153240 141150
rect 153340 141140 153420 141150
rect 153520 141140 153600 141150
rect 153700 141140 153780 141150
rect 153880 141140 153960 141150
rect 154060 141140 154140 141150
rect 154240 141140 154320 141150
rect 154420 141140 154500 141150
rect 154600 141140 154680 141150
rect 154780 141140 154860 141150
rect 154960 141140 155040 141150
rect 155140 141140 155220 141150
rect 155320 141140 155400 141150
rect 155500 141140 155580 141150
rect 155680 141140 155760 141150
rect 155860 141140 155940 141150
rect 156040 141140 156120 141150
rect 156220 141140 156300 141150
rect 156400 141140 156480 141150
rect 156580 141140 156660 141150
rect 156760 141140 156840 141150
rect 156940 141140 157020 141150
rect 157120 141140 157200 141150
rect 157300 141140 157380 141150
rect 157480 141140 157560 141150
rect 157660 141140 157740 141150
rect 157840 141140 157920 141150
rect 158020 141140 158100 141150
rect 158200 141140 158280 141150
rect 158380 141140 158460 141150
rect 158560 141140 158640 141150
rect 158740 141140 158820 141150
rect 158920 141140 159000 141150
rect 159100 141140 159180 141150
rect 159280 141140 159360 141150
rect 159460 141140 159540 141150
rect 159640 141140 159720 141150
rect 152160 141060 152170 141140
rect 152340 141060 152350 141140
rect 152520 141060 152530 141140
rect 152700 141060 152710 141140
rect 152880 141060 152890 141140
rect 153060 141060 153070 141140
rect 153240 141060 153250 141140
rect 153420 141060 153430 141140
rect 153600 141060 153610 141140
rect 153780 141060 153790 141140
rect 153960 141060 153970 141140
rect 154140 141060 154150 141140
rect 154320 141060 154330 141140
rect 154500 141060 154510 141140
rect 154680 141060 154690 141140
rect 154860 141060 154870 141140
rect 155040 141060 155050 141140
rect 155220 141060 155230 141140
rect 155400 141060 155410 141140
rect 155580 141060 155590 141140
rect 155760 141060 155770 141140
rect 155940 141060 155950 141140
rect 156120 141060 156130 141140
rect 156300 141060 156310 141140
rect 156480 141060 156490 141140
rect 156660 141060 156670 141140
rect 156840 141060 156850 141140
rect 157020 141060 157030 141140
rect 157200 141060 157210 141140
rect 157380 141060 157390 141140
rect 157560 141060 157570 141140
rect 157740 141060 157750 141140
rect 157920 141060 157930 141140
rect 158100 141060 158110 141140
rect 158280 141060 158290 141140
rect 158460 141060 158470 141140
rect 158640 141060 158650 141140
rect 158820 141060 158830 141140
rect 159000 141060 159010 141140
rect 159180 141060 159190 141140
rect 159360 141060 159370 141140
rect 159540 141060 159550 141140
rect 159720 141060 159730 141140
rect 161965 141085 161975 141165
rect 162145 141085 162155 141165
rect 162325 141085 162335 141165
rect 162505 141085 162515 141165
rect 162685 141085 162695 141165
rect 163380 141140 163460 141150
rect 163560 141140 163640 141150
rect 163740 141140 163820 141150
rect 163920 141140 164000 141150
rect 164100 141140 164180 141150
rect 164280 141140 164360 141150
rect 164460 141140 164540 141150
rect 164640 141140 164720 141150
rect 164820 141140 164900 141150
rect 165000 141140 165080 141150
rect 165180 141140 165260 141150
rect 165360 141140 165440 141150
rect 165540 141140 165620 141150
rect 165720 141140 165800 141150
rect 165900 141140 165980 141150
rect 166080 141140 166160 141150
rect 166260 141140 166340 141150
rect 166440 141140 166520 141150
rect 166620 141140 166700 141150
rect 166800 141140 166880 141150
rect 166980 141140 167060 141150
rect 167160 141140 167240 141150
rect 167340 141140 167420 141150
rect 167520 141140 167600 141150
rect 167700 141140 167780 141150
rect 167880 141140 167960 141150
rect 168060 141140 168140 141150
rect 168240 141140 168320 141150
rect 168420 141140 168500 141150
rect 168600 141140 168680 141150
rect 168780 141140 168860 141150
rect 168960 141140 169040 141150
rect 169140 141140 169220 141150
rect 169320 141140 169400 141150
rect 169500 141140 169580 141150
rect 169680 141140 169760 141150
rect 169860 141140 169940 141150
rect 170040 141140 170120 141150
rect 170220 141140 170300 141150
rect 170400 141140 170480 141150
rect 170580 141140 170660 141150
rect 170760 141140 170840 141150
rect 170940 141140 171020 141150
rect 163460 141060 163470 141140
rect 163640 141060 163650 141140
rect 163820 141060 163830 141140
rect 164000 141060 164010 141140
rect 164180 141060 164190 141140
rect 164360 141060 164370 141140
rect 164540 141060 164550 141140
rect 164720 141060 164730 141140
rect 164900 141060 164910 141140
rect 165080 141060 165090 141140
rect 165260 141060 165270 141140
rect 165440 141060 165450 141140
rect 165620 141060 165630 141140
rect 165800 141060 165810 141140
rect 165980 141060 165990 141140
rect 166160 141060 166170 141140
rect 166340 141060 166350 141140
rect 166520 141060 166530 141140
rect 166700 141060 166710 141140
rect 166880 141060 166890 141140
rect 167060 141060 167070 141140
rect 167240 141060 167250 141140
rect 167420 141060 167430 141140
rect 167600 141060 167610 141140
rect 167780 141060 167790 141140
rect 167960 141060 167970 141140
rect 168140 141060 168150 141140
rect 168320 141060 168330 141140
rect 168500 141060 168510 141140
rect 168680 141060 168690 141140
rect 168860 141060 168870 141140
rect 169040 141060 169050 141140
rect 169220 141060 169230 141140
rect 169400 141060 169410 141140
rect 169580 141060 169590 141140
rect 169760 141060 169770 141140
rect 169940 141060 169950 141140
rect 170120 141060 170130 141140
rect 170300 141060 170310 141140
rect 170480 141060 170490 141140
rect 170660 141060 170670 141140
rect 170840 141060 170850 141140
rect 171020 141060 171030 141140
rect 152220 140890 152250 140920
rect 152340 140890 152370 140920
rect 159520 140890 159550 140920
rect 159640 140890 159670 140920
rect 152100 140860 152160 140890
rect 152220 140860 152280 140890
rect 152340 140860 152400 140890
rect 159400 140860 159460 140890
rect 159520 140860 159580 140890
rect 159640 140860 159700 140890
rect 152220 140780 152250 140800
rect 152340 140780 152370 140800
rect 159520 140780 159550 140800
rect 159640 140780 159670 140800
rect 163520 140780 163550 140800
rect 163640 140780 163670 140800
rect 170810 140780 170840 140800
rect 170930 140780 170960 140800
rect 77250 140300 90420 140440
rect 101100 140260 105100 140440
rect 132000 140260 143140 140440
rect 146100 130830 146160 130860
rect 36000 130790 37190 130800
rect 37100 130690 37190 130790
rect 40060 130750 40120 130780
rect 37720 130710 37750 130740
rect 37840 130710 37870 130740
rect 36000 130660 37190 130690
rect 37600 130680 37660 130710
rect 37720 130680 37780 130710
rect 37840 130680 37900 130710
rect 36040 130650 36120 130660
rect 36220 130650 36300 130660
rect 36400 130650 36480 130660
rect 36580 130650 36660 130660
rect 36760 130650 36840 130660
rect 36940 130650 37020 130660
rect 36120 130590 36130 130650
rect 36300 130590 36310 130650
rect 36480 130590 36490 130650
rect 36660 130590 36670 130650
rect 36840 130590 36850 130650
rect 37020 130590 37030 130650
rect 37100 130590 37190 130660
rect 40060 130630 40120 130660
rect 37720 130590 37750 130620
rect 37840 130590 37870 130620
rect 36000 130560 37190 130590
rect 37600 130560 37660 130590
rect 37720 130560 37780 130590
rect 37840 130560 37900 130590
rect 36040 130500 36120 130510
rect 36220 130500 36300 130510
rect 36400 130500 36480 130510
rect 36580 130500 36660 130510
rect 36760 130500 36840 130510
rect 36940 130500 37020 130510
rect 36120 130420 36130 130500
rect 36300 130420 36310 130500
rect 36480 130420 36490 130500
rect 36660 130420 36670 130500
rect 36840 130420 36850 130500
rect 37020 130420 37030 130500
rect 36040 130350 36120 130360
rect 36220 130350 36300 130360
rect 36400 130350 36480 130360
rect 36580 130350 36660 130360
rect 36760 130350 36840 130360
rect 36940 130350 37020 130360
rect 36120 130270 36130 130350
rect 36300 130270 36310 130350
rect 36480 130270 36490 130350
rect 36660 130270 36670 130350
rect 36840 130270 36850 130350
rect 37020 130270 37030 130350
rect 37100 130330 37190 130560
rect 40060 130510 40120 130540
rect 37720 130470 37750 130500
rect 37840 130470 37870 130500
rect 37600 130440 37660 130470
rect 37720 130440 37780 130470
rect 37840 130440 37900 130470
rect 40060 130390 40120 130420
rect 37720 130350 37750 130380
rect 37840 130350 37870 130380
rect 37600 130320 37660 130350
rect 37720 130320 37780 130350
rect 37840 130320 37900 130350
rect 40060 130270 40120 130300
rect 19130 130200 19160 130255
rect 19250 130200 19280 130255
rect 26420 130200 26450 130255
rect 26540 130200 26570 130255
rect 30420 130230 30450 130255
rect 30540 130230 30570 130255
rect 37720 130230 37750 130260
rect 37840 130230 37870 130260
rect 30300 130200 30360 130230
rect 30420 130200 30480 130230
rect 30540 130200 30600 130230
rect 37600 130200 37660 130230
rect 37720 130200 37780 130230
rect 37840 130200 37900 130230
rect 40060 130150 40120 130180
rect 30420 130080 30450 130140
rect 30540 130080 30570 130140
rect 37720 130080 37750 130140
rect 37840 130080 37870 130140
rect 40060 130030 40120 130060
rect 18980 129940 19060 129950
rect 19160 129940 19240 129950
rect 19340 129940 19420 129950
rect 19520 129940 19600 129950
rect 19700 129940 19780 129950
rect 19880 129940 19960 129950
rect 20060 129940 20140 129950
rect 20240 129940 20320 129950
rect 20420 129940 20500 129950
rect 20600 129940 20680 129950
rect 20780 129940 20860 129950
rect 20960 129940 21040 129950
rect 21140 129940 21220 129950
rect 21320 129940 21400 129950
rect 21500 129940 21580 129950
rect 21680 129940 21760 129950
rect 21860 129940 21940 129950
rect 22040 129940 22120 129950
rect 22220 129940 22300 129950
rect 22400 129940 22480 129950
rect 22580 129940 22660 129950
rect 22760 129940 22840 129950
rect 22940 129940 23020 129950
rect 23120 129940 23200 129950
rect 23300 129940 23380 129950
rect 23480 129940 23560 129950
rect 23660 129940 23740 129950
rect 23840 129940 23920 129950
rect 24020 129940 24100 129950
rect 24200 129940 24280 129950
rect 24380 129940 24460 129950
rect 24560 129940 24640 129950
rect 24740 129940 24820 129950
rect 24920 129940 25000 129950
rect 25100 129940 25180 129950
rect 25280 129940 25360 129950
rect 25460 129940 25540 129950
rect 25640 129940 25720 129950
rect 25820 129940 25900 129950
rect 26000 129940 26080 129950
rect 26180 129940 26260 129950
rect 26360 129940 26440 129950
rect 26540 129940 26620 129950
rect 30280 129940 30360 129950
rect 30460 129940 30540 129950
rect 30640 129940 30720 129950
rect 30820 129940 30900 129950
rect 31000 129940 31080 129950
rect 31180 129940 31260 129950
rect 31360 129940 31440 129950
rect 31540 129940 31620 129950
rect 31720 129940 31800 129950
rect 31900 129940 31980 129950
rect 32080 129940 32160 129950
rect 32260 129940 32340 129950
rect 32440 129940 32520 129950
rect 32620 129940 32700 129950
rect 32800 129940 32880 129950
rect 32980 129940 33060 129950
rect 33160 129940 33240 129950
rect 33340 129940 33420 129950
rect 33520 129940 33600 129950
rect 33700 129940 33780 129950
rect 33880 129940 33960 129950
rect 34060 129940 34140 129950
rect 34240 129940 34320 129950
rect 34420 129940 34500 129950
rect 34600 129940 34680 129950
rect 34780 129940 34860 129950
rect 34960 129940 35040 129950
rect 35140 129940 35220 129950
rect 35320 129940 35400 129950
rect 35500 129940 35580 129950
rect 35680 129940 35760 129950
rect 35860 129940 35940 129950
rect 36040 129940 36120 129950
rect 36220 129940 36300 129950
rect 36400 129940 36480 129950
rect 36580 129940 36660 129950
rect 36760 129940 36840 129950
rect 36940 129940 37020 129950
rect 37120 129940 37200 129950
rect 37300 129940 37380 129950
rect 37480 129940 37560 129950
rect 37660 129940 37740 129950
rect 37840 129940 37920 129950
rect 40260 129940 40270 130800
rect 41090 130765 41180 130800
rect 40470 130735 41180 130765
rect 40650 130700 40770 130735
rect 40930 130700 41050 130735
rect 41090 130700 41180 130735
rect 41350 130730 41410 130800
rect 40650 130610 40660 130700
rect 40760 130670 40830 130700
rect 40770 130580 40830 130670
rect 40930 130610 40940 130700
rect 41050 130580 41180 130700
rect 41260 130680 41340 130690
rect 41340 130610 41350 130680
rect 41090 130545 41180 130580
rect 41230 130550 41350 130610
rect 40370 130530 40460 130540
rect 40370 130450 40380 130530
rect 40470 130525 41180 130545
rect 40420 130515 41210 130525
rect 41090 130465 41180 130515
rect 40470 130450 41180 130465
rect 40460 130435 41180 130450
rect 40460 130245 40470 130435
rect 40650 130400 40770 130435
rect 40930 130400 41050 130435
rect 41090 130400 41180 130435
rect 41350 130430 41410 130550
rect 40770 130390 40830 130400
rect 40530 130380 40610 130390
rect 40670 130380 40750 130390
rect 40770 130380 40890 130390
rect 40950 130380 41030 130390
rect 40610 130300 40620 130380
rect 40750 130300 40760 130380
rect 40770 130280 40830 130380
rect 40890 130300 40900 130380
rect 41030 130300 41040 130380
rect 41050 130280 41180 130400
rect 41260 130370 41340 130380
rect 41340 130310 41350 130370
rect 41090 130245 41180 130280
rect 41230 130250 41350 130310
rect 40460 130230 41180 130245
rect 40470 130225 41180 130230
rect 40420 130215 41210 130225
rect 41090 130165 41180 130215
rect 40470 130135 41180 130165
rect 40650 130100 40770 130135
rect 40930 130100 41050 130135
rect 41090 130100 41180 130135
rect 41350 130130 41410 130250
rect 41480 130100 41490 130800
rect 41540 130750 41600 130780
rect 42360 130750 42420 130780
rect 41540 130630 41600 130660
rect 42360 130630 42420 130660
rect 41540 130510 41600 130540
rect 42360 130510 42420 130540
rect 41540 130390 41600 130420
rect 42360 130390 42420 130420
rect 41540 130270 41600 130300
rect 42360 130270 42420 130300
rect 41540 130150 41600 130180
rect 42360 130150 42420 130180
rect 42560 130120 42570 130800
rect 42730 130740 42790 130800
rect 43540 130775 43550 130800
rect 42620 130640 42700 130650
rect 42700 130560 42710 130640
rect 42860 130570 42870 130760
rect 42910 130710 43030 130770
rect 43190 130710 43310 130770
rect 43020 130680 43090 130710
rect 43030 130590 43090 130680
rect 43190 130620 43200 130710
rect 43300 130680 43370 130710
rect 43310 130590 43370 130680
rect 42860 130560 43490 130570
rect 42860 130550 42870 130560
rect 42620 130460 42700 130470
rect 42770 130460 42780 130550
rect 42700 130380 42710 130460
rect 42610 130270 42730 130330
rect 42730 130245 42790 130270
rect 42860 130260 42870 130460
rect 42910 130420 43030 130480
rect 43190 130420 43310 130480
rect 43030 130410 43090 130420
rect 43310 130410 43370 130420
rect 42930 130400 43010 130410
rect 43030 130400 43150 130410
rect 43210 130400 43290 130410
rect 43310 130400 43430 130410
rect 43010 130320 43020 130400
rect 43030 130300 43090 130400
rect 43150 130320 43160 130400
rect 43290 130320 43300 130400
rect 43310 130300 43370 130400
rect 43430 130320 43440 130400
rect 42860 130250 43500 130260
rect 43580 130250 43590 130550
rect 42730 130235 43540 130245
rect 42730 130150 42790 130235
rect 43540 130185 43550 130235
rect 42860 130120 42870 130170
rect 42910 130120 43030 130180
rect 43190 130120 43310 130180
rect 43030 130110 43090 130120
rect 43310 130110 43370 130120
rect 43030 130100 43150 130110
rect 43310 130100 43430 130110
rect 40770 130090 40830 130100
rect 40530 130080 40610 130090
rect 40770 130080 40890 130090
rect 40610 130000 40620 130080
rect 40770 129980 40830 130080
rect 40890 130000 40900 130080
rect 41050 129980 41180 130100
rect 41540 130030 41600 130060
rect 42360 130030 42420 130060
rect 43030 130000 43090 130100
rect 43150 130020 43160 130100
rect 43310 130000 43370 130100
rect 43430 130020 43440 130100
rect 41090 129950 41180 129980
rect 43780 129960 43790 130800
rect 43840 130750 43900 130780
rect 146100 130710 146160 130740
rect 43840 130630 43900 130660
rect 146300 130650 146310 130920
rect 146690 130820 146810 130880
rect 146970 130820 147090 130880
rect 146690 130730 146700 130820
rect 146800 130790 146870 130820
rect 146810 130700 146870 130790
rect 146970 130730 146980 130820
rect 147090 130700 147140 130820
rect 146410 130650 147140 130660
rect 146460 130635 147140 130645
rect 146100 130590 146160 130620
rect 146450 130585 146460 130635
rect 43840 130510 43900 130540
rect 146690 130520 146810 130580
rect 146970 130520 147090 130580
rect 146810 130510 146870 130520
rect 146570 130500 146650 130510
rect 146710 130500 146790 130510
rect 146810 130500 146930 130510
rect 146990 130500 147070 130510
rect 146100 130470 146160 130500
rect 146650 130420 146660 130500
rect 146790 130420 146800 130500
rect 43840 130390 43900 130420
rect 146810 130400 146870 130500
rect 146930 130420 146940 130500
rect 147070 130420 147080 130500
rect 147090 130400 147140 130520
rect 146100 130350 146160 130380
rect 43840 130270 43900 130300
rect 146100 130230 146160 130260
rect 147580 130230 147640 130246
rect 148400 130230 148460 130246
rect 148600 130220 148610 130246
rect 148950 130220 149070 130246
rect 149230 130220 149350 130246
rect 149060 130190 149130 130220
rect 43840 130150 43900 130180
rect 146100 130110 146160 130140
rect 147580 130110 147640 130140
rect 148400 130110 148460 130140
rect 149070 130100 149130 130190
rect 149230 130130 149240 130220
rect 149340 130190 149410 130220
rect 149350 130100 149410 130190
rect 149530 130070 149620 130246
rect 149820 130060 149830 130246
rect 149880 130230 149940 130246
rect 152220 130210 152250 130240
rect 152340 130210 152370 130240
rect 159520 130210 159550 130240
rect 159640 130210 159670 130240
rect 163520 130210 163550 130240
rect 163640 130210 163670 130240
rect 163960 130235 164040 130245
rect 152100 130180 152160 130210
rect 152220 130180 152280 130210
rect 152340 130180 152400 130210
rect 159400 130180 159460 130210
rect 159520 130180 159580 130210
rect 159640 130180 159700 130210
rect 163400 130180 163460 130210
rect 163520 130180 163580 130210
rect 163640 130180 163700 130210
rect 164040 130155 164050 130235
rect 170810 130210 170840 130240
rect 170930 130210 170960 130240
rect 170690 130180 170750 130210
rect 170810 130180 170870 130210
rect 170930 130180 170990 130210
rect 149880 130110 149940 130140
rect 152220 130060 152250 130120
rect 152340 130060 152370 130120
rect 159520 130060 159550 130120
rect 159640 130060 159670 130120
rect 163520 130060 163550 130120
rect 163640 130060 163670 130120
rect 170810 130060 170840 130120
rect 170930 130060 170960 130120
rect 43840 130030 43900 130060
rect 146100 129990 146160 130020
rect 147580 129990 147640 130020
rect 148400 129990 148460 130020
rect 149880 129990 149940 130020
rect 19060 129860 19070 129940
rect 19240 129860 19250 129940
rect 19420 129860 19430 129940
rect 19600 129860 19610 129940
rect 19780 129860 19790 129940
rect 19960 129860 19970 129940
rect 20140 129860 20150 129940
rect 20320 129860 20330 129940
rect 20500 129860 20510 129940
rect 20680 129860 20690 129940
rect 20860 129860 20870 129940
rect 21040 129860 21050 129940
rect 21220 129860 21230 129940
rect 21400 129860 21410 129940
rect 21580 129860 21590 129940
rect 21760 129860 21770 129940
rect 21940 129860 21950 129940
rect 22120 129860 22130 129940
rect 22300 129860 22310 129940
rect 22480 129860 22490 129940
rect 22660 129860 22670 129940
rect 22840 129860 22850 129940
rect 23020 129860 23030 129940
rect 23200 129860 23210 129940
rect 23380 129860 23390 129940
rect 23560 129860 23570 129940
rect 23740 129860 23750 129940
rect 23920 129860 23930 129940
rect 24100 129860 24110 129940
rect 24280 129860 24290 129940
rect 24460 129860 24470 129940
rect 24640 129860 24650 129940
rect 24820 129860 24830 129940
rect 25000 129860 25010 129940
rect 25180 129860 25190 129940
rect 25360 129860 25370 129940
rect 25540 129860 25550 129940
rect 25720 129860 25730 129940
rect 25900 129860 25910 129940
rect 26080 129860 26090 129940
rect 26260 129860 26270 129940
rect 26440 129860 26450 129940
rect 26620 129860 26630 129940
rect 27315 129915 27395 129925
rect 27495 129915 27575 129925
rect 27675 129915 27755 129925
rect 27855 129915 27935 129925
rect 28035 129915 28115 129925
rect 27395 129835 27405 129915
rect 27575 129835 27585 129915
rect 27755 129835 27765 129915
rect 27935 129835 27945 129915
rect 28115 129835 28125 129915
rect 30360 129860 30370 129940
rect 30540 129860 30550 129940
rect 30720 129860 30730 129940
rect 30900 129860 30910 129940
rect 31080 129860 31090 129940
rect 31260 129860 31270 129940
rect 31440 129860 31450 129940
rect 31620 129860 31630 129940
rect 31800 129860 31810 129940
rect 31980 129860 31990 129940
rect 32160 129860 32170 129940
rect 32340 129860 32350 129940
rect 32520 129860 32530 129940
rect 32700 129860 32710 129940
rect 32880 129860 32890 129940
rect 33060 129860 33070 129940
rect 33240 129860 33250 129940
rect 33420 129860 33430 129940
rect 33600 129860 33610 129940
rect 33780 129860 33790 129940
rect 33960 129860 33970 129940
rect 34140 129860 34150 129940
rect 34320 129860 34330 129940
rect 34500 129860 34510 129940
rect 34680 129860 34690 129940
rect 34860 129860 34870 129940
rect 35040 129860 35050 129940
rect 35220 129860 35230 129940
rect 35400 129860 35410 129940
rect 35580 129860 35590 129940
rect 35760 129860 35770 129940
rect 35940 129860 35950 129940
rect 36120 129860 36130 129940
rect 36300 129860 36310 129940
rect 36480 129860 36490 129940
rect 36660 129860 36670 129940
rect 36840 129860 36850 129940
rect 37020 129860 37030 129940
rect 37200 129860 37210 129940
rect 37380 129860 37390 129940
rect 37560 129860 37570 129940
rect 37740 129860 37750 129940
rect 37920 129860 37930 129940
rect 40060 129910 40120 129940
rect 41540 129910 41600 129940
rect 42360 129910 42420 129940
rect 43840 129910 43900 129940
rect 146100 129870 146160 129900
rect 147580 129870 147640 129900
rect 148400 129870 148460 129900
rect 149880 129870 149940 129900
rect 18980 129790 19060 129800
rect 19160 129790 19240 129800
rect 19340 129790 19420 129800
rect 19520 129790 19600 129800
rect 19700 129790 19780 129800
rect 19880 129790 19960 129800
rect 20060 129790 20140 129800
rect 20240 129790 20320 129800
rect 20420 129790 20500 129800
rect 20600 129790 20680 129800
rect 20780 129790 20860 129800
rect 20960 129790 21040 129800
rect 21140 129790 21220 129800
rect 21320 129790 21400 129800
rect 21500 129790 21580 129800
rect 21680 129790 21760 129800
rect 21860 129790 21940 129800
rect 22040 129790 22120 129800
rect 22220 129790 22300 129800
rect 22400 129790 22480 129800
rect 22580 129790 22660 129800
rect 22760 129790 22840 129800
rect 22940 129790 23020 129800
rect 23120 129790 23200 129800
rect 23300 129790 23380 129800
rect 23480 129790 23560 129800
rect 23660 129790 23740 129800
rect 23840 129790 23920 129800
rect 24020 129790 24100 129800
rect 24200 129790 24280 129800
rect 24380 129790 24460 129800
rect 24560 129790 24640 129800
rect 24740 129790 24820 129800
rect 24920 129790 25000 129800
rect 25100 129790 25180 129800
rect 25280 129790 25360 129800
rect 25460 129790 25540 129800
rect 25640 129790 25720 129800
rect 25820 129790 25900 129800
rect 26000 129790 26080 129800
rect 26180 129790 26260 129800
rect 26360 129790 26440 129800
rect 26540 129790 26620 129800
rect 30280 129790 30360 129800
rect 30460 129790 30540 129800
rect 30640 129790 30720 129800
rect 30820 129790 30900 129800
rect 31000 129790 31080 129800
rect 31180 129790 31260 129800
rect 31360 129790 31440 129800
rect 31540 129790 31620 129800
rect 31720 129790 31800 129800
rect 31900 129790 31980 129800
rect 32080 129790 32160 129800
rect 32260 129790 32340 129800
rect 32440 129790 32520 129800
rect 32620 129790 32700 129800
rect 32800 129790 32880 129800
rect 32980 129790 33060 129800
rect 33160 129790 33240 129800
rect 33340 129790 33420 129800
rect 33520 129790 33600 129800
rect 33700 129790 33780 129800
rect 33880 129790 33960 129800
rect 34060 129790 34140 129800
rect 34240 129790 34320 129800
rect 34420 129790 34500 129800
rect 34600 129790 34680 129800
rect 34780 129790 34860 129800
rect 34960 129790 35040 129800
rect 35140 129790 35220 129800
rect 35320 129790 35400 129800
rect 35500 129790 35580 129800
rect 35680 129790 35760 129800
rect 35860 129790 35940 129800
rect 36040 129790 36120 129800
rect 36220 129790 36300 129800
rect 36400 129790 36480 129800
rect 36580 129790 36660 129800
rect 36760 129790 36840 129800
rect 36940 129790 37020 129800
rect 37120 129790 37200 129800
rect 37300 129790 37380 129800
rect 37480 129790 37560 129800
rect 37660 129790 37740 129800
rect 37840 129790 37920 129800
rect 152080 129790 152160 129800
rect 152260 129790 152340 129800
rect 152440 129790 152520 129800
rect 152620 129790 152700 129800
rect 152800 129790 152880 129800
rect 152980 129790 153060 129800
rect 153160 129790 153240 129800
rect 153340 129790 153420 129800
rect 153520 129790 153600 129800
rect 153700 129790 153780 129800
rect 153880 129790 153960 129800
rect 154060 129790 154140 129800
rect 154240 129790 154320 129800
rect 154420 129790 154500 129800
rect 154600 129790 154680 129800
rect 154780 129790 154860 129800
rect 154960 129790 155040 129800
rect 155140 129790 155220 129800
rect 155320 129790 155400 129800
rect 155500 129790 155580 129800
rect 155680 129790 155760 129800
rect 155860 129790 155940 129800
rect 156040 129790 156120 129800
rect 156220 129790 156300 129800
rect 156400 129790 156480 129800
rect 156580 129790 156660 129800
rect 156760 129790 156840 129800
rect 156940 129790 157020 129800
rect 157120 129790 157200 129800
rect 157300 129790 157380 129800
rect 157480 129790 157560 129800
rect 157660 129790 157740 129800
rect 157840 129790 157920 129800
rect 158020 129790 158100 129800
rect 158200 129790 158280 129800
rect 158380 129790 158460 129800
rect 158560 129790 158640 129800
rect 158740 129790 158820 129800
rect 158920 129790 159000 129800
rect 159100 129790 159180 129800
rect 159280 129790 159360 129800
rect 159460 129790 159540 129800
rect 159640 129790 159720 129800
rect 163380 129790 163460 129800
rect 163560 129790 163640 129800
rect 163740 129790 163820 129800
rect 163920 129790 164000 129800
rect 164100 129790 164180 129800
rect 164280 129790 164360 129800
rect 164460 129790 164540 129800
rect 164640 129790 164720 129800
rect 164820 129790 164900 129800
rect 165000 129790 165080 129800
rect 165180 129790 165260 129800
rect 165360 129790 165440 129800
rect 165540 129790 165620 129800
rect 165720 129790 165800 129800
rect 165900 129790 165980 129800
rect 166080 129790 166160 129800
rect 166260 129790 166340 129800
rect 166440 129790 166520 129800
rect 166620 129790 166700 129800
rect 166800 129790 166880 129800
rect 166980 129790 167060 129800
rect 167160 129790 167240 129800
rect 167340 129790 167420 129800
rect 167520 129790 167600 129800
rect 167700 129790 167780 129800
rect 167880 129790 167960 129800
rect 168060 129790 168140 129800
rect 168240 129790 168320 129800
rect 168420 129790 168500 129800
rect 168600 129790 168680 129800
rect 168780 129790 168860 129800
rect 168960 129790 169040 129800
rect 169140 129790 169220 129800
rect 169320 129790 169400 129800
rect 169500 129790 169580 129800
rect 169680 129790 169760 129800
rect 169860 129790 169940 129800
rect 170040 129790 170120 129800
rect 170220 129790 170300 129800
rect 170400 129790 170480 129800
rect 170580 129790 170660 129800
rect 170760 129790 170840 129800
rect 170940 129790 171020 129800
rect 19060 129710 19070 129790
rect 19240 129710 19250 129790
rect 19420 129710 19430 129790
rect 19600 129710 19610 129790
rect 19780 129710 19790 129790
rect 19960 129710 19970 129790
rect 20140 129710 20150 129790
rect 20320 129710 20330 129790
rect 20500 129710 20510 129790
rect 20680 129710 20690 129790
rect 20860 129710 20870 129790
rect 21040 129710 21050 129790
rect 21220 129710 21230 129790
rect 21400 129710 21410 129790
rect 21580 129710 21590 129790
rect 21760 129710 21770 129790
rect 21940 129710 21950 129790
rect 22120 129710 22130 129790
rect 22300 129710 22310 129790
rect 22480 129710 22490 129790
rect 22660 129710 22670 129790
rect 22840 129710 22850 129790
rect 23020 129710 23030 129790
rect 23200 129710 23210 129790
rect 23380 129710 23390 129790
rect 23560 129710 23570 129790
rect 23740 129710 23750 129790
rect 23920 129710 23930 129790
rect 24100 129710 24110 129790
rect 24280 129710 24290 129790
rect 24460 129710 24470 129790
rect 24640 129710 24650 129790
rect 24820 129710 24830 129790
rect 25000 129710 25010 129790
rect 25180 129710 25190 129790
rect 25360 129710 25370 129790
rect 25540 129710 25550 129790
rect 25720 129710 25730 129790
rect 25900 129710 25910 129790
rect 26080 129710 26090 129790
rect 26260 129710 26270 129790
rect 26440 129710 26450 129790
rect 26620 129710 26630 129790
rect 27315 129735 27395 129745
rect 27495 129735 27575 129745
rect 27675 129735 27755 129745
rect 27855 129735 27935 129745
rect 28035 129735 28115 129745
rect 27395 129655 27405 129735
rect 27575 129655 27585 129735
rect 27755 129655 27765 129735
rect 27935 129655 27945 129735
rect 28115 129655 28125 129735
rect 30360 129710 30370 129790
rect 30540 129710 30550 129790
rect 30720 129710 30730 129790
rect 30900 129710 30910 129790
rect 31080 129710 31090 129790
rect 31260 129710 31270 129790
rect 31440 129710 31450 129790
rect 31620 129710 31630 129790
rect 31800 129710 31810 129790
rect 31980 129710 31990 129790
rect 32160 129710 32170 129790
rect 32340 129710 32350 129790
rect 32520 129710 32530 129790
rect 32700 129710 32710 129790
rect 32880 129710 32890 129790
rect 33060 129710 33070 129790
rect 33240 129710 33250 129790
rect 33420 129710 33430 129790
rect 33600 129710 33610 129790
rect 33780 129710 33790 129790
rect 33960 129710 33970 129790
rect 34140 129710 34150 129790
rect 34320 129710 34330 129790
rect 34500 129710 34510 129790
rect 34680 129710 34690 129790
rect 34860 129710 34870 129790
rect 35040 129710 35050 129790
rect 35220 129710 35230 129790
rect 35400 129710 35410 129790
rect 35580 129710 35590 129790
rect 35760 129710 35770 129790
rect 35940 129710 35950 129790
rect 36120 129710 36130 129790
rect 36300 129710 36310 129790
rect 36480 129710 36490 129790
rect 36660 129710 36670 129790
rect 36840 129710 36850 129790
rect 37020 129710 37030 129790
rect 37200 129710 37210 129790
rect 37380 129710 37390 129790
rect 37560 129710 37570 129790
rect 37740 129710 37750 129790
rect 37920 129710 37930 129790
rect 152160 129710 152170 129790
rect 152340 129710 152350 129790
rect 152520 129710 152530 129790
rect 152700 129710 152710 129790
rect 152880 129710 152890 129790
rect 153060 129710 153070 129790
rect 153240 129710 153250 129790
rect 153420 129710 153430 129790
rect 153600 129710 153610 129790
rect 153780 129710 153790 129790
rect 153960 129710 153970 129790
rect 154140 129710 154150 129790
rect 154320 129710 154330 129790
rect 154500 129710 154510 129790
rect 154680 129710 154690 129790
rect 154860 129710 154870 129790
rect 155040 129710 155050 129790
rect 155220 129710 155230 129790
rect 155400 129710 155410 129790
rect 155580 129710 155590 129790
rect 155760 129710 155770 129790
rect 155940 129710 155950 129790
rect 156120 129710 156130 129790
rect 156300 129710 156310 129790
rect 156480 129710 156490 129790
rect 156660 129710 156670 129790
rect 156840 129710 156850 129790
rect 157020 129710 157030 129790
rect 157200 129710 157210 129790
rect 157380 129710 157390 129790
rect 157560 129710 157570 129790
rect 157740 129710 157750 129790
rect 157920 129710 157930 129790
rect 158100 129710 158110 129790
rect 158280 129710 158290 129790
rect 158460 129710 158470 129790
rect 158640 129710 158650 129790
rect 158820 129710 158830 129790
rect 159000 129710 159010 129790
rect 159180 129710 159190 129790
rect 159360 129710 159370 129790
rect 159540 129710 159550 129790
rect 159720 129710 159730 129790
rect 160430 129765 160510 129775
rect 160590 129765 160670 129775
rect 160750 129765 160830 129775
rect 160910 129765 160990 129775
rect 161070 129765 161150 129775
rect 160510 129685 160520 129765
rect 160590 129685 160600 129765
rect 160670 129685 160680 129765
rect 160750 129685 160760 129765
rect 160830 129685 160840 129765
rect 160910 129685 160920 129765
rect 160990 129685 161000 129765
rect 161070 129685 161080 129765
rect 161150 129685 161160 129765
rect 163460 129710 163470 129790
rect 163640 129710 163650 129790
rect 163820 129710 163830 129790
rect 164000 129710 164010 129790
rect 164180 129710 164190 129790
rect 164360 129710 164370 129790
rect 164540 129710 164550 129790
rect 164720 129710 164730 129790
rect 164900 129710 164910 129790
rect 165080 129710 165090 129790
rect 165260 129710 165270 129790
rect 165440 129710 165450 129790
rect 165620 129710 165630 129790
rect 165800 129710 165810 129790
rect 165980 129710 165990 129790
rect 166160 129710 166170 129790
rect 166340 129710 166350 129790
rect 166520 129710 166530 129790
rect 166700 129710 166710 129790
rect 166880 129710 166890 129790
rect 167060 129710 167070 129790
rect 167240 129710 167250 129790
rect 167420 129710 167430 129790
rect 167600 129710 167610 129790
rect 167780 129710 167790 129790
rect 167960 129710 167970 129790
rect 168140 129710 168150 129790
rect 168320 129710 168330 129790
rect 168500 129710 168510 129790
rect 168680 129710 168690 129790
rect 168860 129710 168870 129790
rect 169040 129710 169050 129790
rect 169220 129710 169230 129790
rect 169400 129710 169410 129790
rect 169580 129710 169590 129790
rect 169760 129710 169770 129790
rect 169940 129710 169950 129790
rect 170120 129710 170130 129790
rect 170300 129710 170310 129790
rect 170480 129710 170490 129790
rect 170660 129710 170670 129790
rect 170840 129710 170850 129790
rect 171020 129710 171030 129790
rect 18980 129640 19060 129650
rect 19160 129640 19240 129650
rect 19340 129640 19420 129650
rect 19520 129640 19600 129650
rect 19700 129640 19780 129650
rect 19880 129640 19960 129650
rect 20060 129640 20140 129650
rect 20240 129640 20320 129650
rect 20420 129640 20500 129650
rect 20600 129640 20680 129650
rect 20780 129640 20860 129650
rect 20960 129640 21040 129650
rect 21140 129640 21220 129650
rect 21320 129640 21400 129650
rect 21500 129640 21580 129650
rect 21680 129640 21760 129650
rect 21860 129640 21940 129650
rect 22040 129640 22120 129650
rect 22220 129640 22300 129650
rect 22400 129640 22480 129650
rect 22580 129640 22660 129650
rect 22760 129640 22840 129650
rect 22940 129640 23020 129650
rect 23120 129640 23200 129650
rect 23300 129640 23380 129650
rect 23480 129640 23560 129650
rect 23660 129640 23740 129650
rect 23840 129640 23920 129650
rect 24020 129640 24100 129650
rect 24200 129640 24280 129650
rect 24380 129640 24460 129650
rect 24560 129640 24640 129650
rect 24740 129640 24820 129650
rect 24920 129640 25000 129650
rect 25100 129640 25180 129650
rect 25280 129640 25360 129650
rect 25460 129640 25540 129650
rect 25640 129640 25720 129650
rect 25820 129640 25900 129650
rect 26000 129640 26080 129650
rect 26180 129640 26260 129650
rect 26360 129640 26440 129650
rect 26540 129640 26620 129650
rect 30280 129640 30360 129650
rect 30460 129640 30540 129650
rect 30640 129640 30720 129650
rect 30820 129640 30900 129650
rect 31000 129640 31080 129650
rect 31180 129640 31260 129650
rect 31360 129640 31440 129650
rect 31540 129640 31620 129650
rect 31720 129640 31800 129650
rect 31900 129640 31980 129650
rect 32080 129640 32160 129650
rect 32260 129640 32340 129650
rect 32440 129640 32520 129650
rect 32620 129640 32700 129650
rect 32800 129640 32880 129650
rect 32980 129640 33060 129650
rect 33160 129640 33240 129650
rect 33340 129640 33420 129650
rect 33520 129640 33600 129650
rect 33700 129640 33780 129650
rect 33880 129640 33960 129650
rect 34060 129640 34140 129650
rect 34240 129640 34320 129650
rect 34420 129640 34500 129650
rect 34600 129640 34680 129650
rect 34780 129640 34860 129650
rect 34960 129640 35040 129650
rect 35140 129640 35220 129650
rect 35320 129640 35400 129650
rect 35500 129640 35580 129650
rect 35680 129640 35760 129650
rect 35860 129640 35940 129650
rect 36040 129640 36120 129650
rect 36220 129640 36300 129650
rect 36400 129640 36480 129650
rect 36580 129640 36660 129650
rect 36760 129640 36840 129650
rect 36940 129640 37020 129650
rect 37120 129640 37200 129650
rect 37300 129640 37380 129650
rect 37480 129640 37560 129650
rect 37660 129640 37740 129650
rect 37840 129640 37920 129650
rect 40060 129640 40140 129650
rect 40200 129640 40280 129650
rect 40340 129640 40420 129650
rect 40480 129640 40560 129650
rect 40620 129640 40700 129650
rect 40760 129640 40840 129650
rect 40900 129640 40980 129650
rect 41040 129640 41120 129650
rect 41180 129640 41260 129650
rect 41320 129640 41400 129650
rect 42360 129640 42440 129650
rect 42500 129640 42580 129650
rect 42640 129640 42720 129650
rect 42780 129640 42860 129650
rect 42920 129640 43000 129650
rect 43060 129640 43140 129650
rect 43200 129640 43280 129650
rect 43340 129640 43420 129650
rect 43480 129640 43560 129650
rect 43620 129640 43700 129650
rect 146300 129640 146380 129650
rect 146440 129640 146520 129650
rect 146580 129640 146660 129650
rect 146720 129640 146800 129650
rect 146860 129640 146940 129650
rect 147000 129640 147080 129650
rect 147140 129640 147220 129650
rect 147280 129640 147360 129650
rect 147420 129640 147500 129650
rect 147560 129640 147640 129650
rect 148600 129640 148680 129650
rect 148740 129640 148820 129650
rect 148880 129640 148960 129650
rect 149020 129640 149100 129650
rect 149160 129640 149240 129650
rect 149300 129640 149380 129650
rect 149440 129640 149520 129650
rect 149580 129640 149660 129650
rect 149720 129640 149800 129650
rect 149860 129640 149940 129650
rect 152080 129640 152160 129650
rect 152260 129640 152340 129650
rect 152440 129640 152520 129650
rect 152620 129640 152700 129650
rect 152800 129640 152880 129650
rect 152980 129640 153060 129650
rect 153160 129640 153240 129650
rect 153340 129640 153420 129650
rect 153520 129640 153600 129650
rect 153700 129640 153780 129650
rect 153880 129640 153960 129650
rect 154060 129640 154140 129650
rect 154240 129640 154320 129650
rect 154420 129640 154500 129650
rect 154600 129640 154680 129650
rect 154780 129640 154860 129650
rect 154960 129640 155040 129650
rect 155140 129640 155220 129650
rect 155320 129640 155400 129650
rect 155500 129640 155580 129650
rect 155680 129640 155760 129650
rect 155860 129640 155940 129650
rect 156040 129640 156120 129650
rect 156220 129640 156300 129650
rect 156400 129640 156480 129650
rect 156580 129640 156660 129650
rect 156760 129640 156840 129650
rect 156940 129640 157020 129650
rect 157120 129640 157200 129650
rect 157300 129640 157380 129650
rect 157480 129640 157560 129650
rect 157660 129640 157740 129650
rect 157840 129640 157920 129650
rect 158020 129640 158100 129650
rect 158200 129640 158280 129650
rect 158380 129640 158460 129650
rect 158560 129640 158640 129650
rect 158740 129640 158820 129650
rect 158920 129640 159000 129650
rect 159100 129640 159180 129650
rect 159280 129640 159360 129650
rect 159460 129640 159540 129650
rect 159640 129640 159720 129650
rect 163380 129640 163460 129650
rect 163560 129640 163640 129650
rect 163740 129640 163820 129650
rect 163920 129640 164000 129650
rect 164100 129640 164180 129650
rect 164280 129640 164360 129650
rect 164460 129640 164540 129650
rect 164640 129640 164720 129650
rect 164820 129640 164900 129650
rect 165000 129640 165080 129650
rect 165180 129640 165260 129650
rect 165360 129640 165440 129650
rect 165540 129640 165620 129650
rect 165720 129640 165800 129650
rect 165900 129640 165980 129650
rect 166080 129640 166160 129650
rect 166260 129640 166340 129650
rect 166440 129640 166520 129650
rect 166620 129640 166700 129650
rect 166800 129640 166880 129650
rect 166980 129640 167060 129650
rect 167160 129640 167240 129650
rect 167340 129640 167420 129650
rect 167520 129640 167600 129650
rect 167700 129640 167780 129650
rect 167880 129640 167960 129650
rect 168060 129640 168140 129650
rect 168240 129640 168320 129650
rect 168420 129640 168500 129650
rect 168600 129640 168680 129650
rect 168780 129640 168860 129650
rect 168960 129640 169040 129650
rect 169140 129640 169220 129650
rect 169320 129640 169400 129650
rect 169500 129640 169580 129650
rect 169680 129640 169760 129650
rect 169860 129640 169940 129650
rect 170040 129640 170120 129650
rect 170220 129640 170300 129650
rect 170400 129640 170480 129650
rect 170580 129640 170660 129650
rect 170760 129640 170840 129650
rect 170940 129640 171020 129650
rect 19060 129560 19070 129640
rect 19240 129560 19250 129640
rect 19420 129560 19430 129640
rect 19600 129560 19610 129640
rect 19780 129560 19790 129640
rect 19960 129560 19970 129640
rect 20140 129560 20150 129640
rect 20320 129560 20330 129640
rect 20500 129560 20510 129640
rect 20680 129560 20690 129640
rect 20860 129560 20870 129640
rect 21040 129560 21050 129640
rect 21220 129560 21230 129640
rect 21400 129560 21410 129640
rect 21580 129560 21590 129640
rect 21760 129560 21770 129640
rect 21940 129560 21950 129640
rect 22120 129560 22130 129640
rect 22300 129560 22310 129640
rect 22480 129560 22490 129640
rect 22660 129560 22670 129640
rect 22840 129560 22850 129640
rect 23020 129560 23030 129640
rect 23200 129560 23210 129640
rect 23380 129560 23390 129640
rect 23560 129560 23570 129640
rect 23740 129560 23750 129640
rect 23920 129560 23930 129640
rect 24100 129560 24110 129640
rect 24280 129560 24290 129640
rect 24460 129560 24470 129640
rect 24640 129560 24650 129640
rect 24820 129560 24830 129640
rect 25000 129560 25010 129640
rect 25180 129560 25190 129640
rect 25360 129560 25370 129640
rect 25540 129560 25550 129640
rect 25720 129560 25730 129640
rect 25900 129560 25910 129640
rect 26080 129560 26090 129640
rect 26260 129560 26270 129640
rect 26440 129560 26450 129640
rect 26620 129560 26630 129640
rect 30360 129560 30370 129640
rect 30540 129560 30550 129640
rect 30720 129560 30730 129640
rect 30900 129560 30910 129640
rect 31080 129560 31090 129640
rect 31260 129560 31270 129640
rect 31440 129560 31450 129640
rect 31620 129560 31630 129640
rect 31800 129560 31810 129640
rect 31980 129560 31990 129640
rect 32160 129560 32170 129640
rect 32340 129560 32350 129640
rect 32520 129560 32530 129640
rect 32700 129560 32710 129640
rect 32880 129560 32890 129640
rect 33060 129560 33070 129640
rect 33240 129560 33250 129640
rect 33420 129560 33430 129640
rect 33600 129560 33610 129640
rect 33780 129560 33790 129640
rect 33960 129560 33970 129640
rect 34140 129560 34150 129640
rect 34320 129560 34330 129640
rect 34500 129560 34510 129640
rect 34680 129560 34690 129640
rect 34860 129560 34870 129640
rect 35040 129560 35050 129640
rect 35220 129560 35230 129640
rect 35400 129560 35410 129640
rect 35580 129560 35590 129640
rect 35760 129560 35770 129640
rect 35940 129560 35950 129640
rect 36120 129560 36130 129640
rect 36300 129560 36310 129640
rect 36480 129560 36490 129640
rect 36660 129560 36670 129640
rect 36840 129560 36850 129640
rect 37020 129560 37030 129640
rect 37200 129560 37210 129640
rect 37380 129560 37390 129640
rect 37560 129560 37570 129640
rect 37740 129560 37750 129640
rect 37920 129560 37930 129640
rect 40140 129560 40150 129640
rect 40280 129560 40290 129640
rect 40420 129560 40430 129640
rect 40560 129560 40570 129640
rect 40700 129560 40710 129640
rect 40840 129560 40850 129640
rect 40980 129560 40990 129640
rect 41120 129560 41130 129640
rect 41260 129560 41270 129640
rect 41400 129560 41410 129640
rect 42440 129560 42450 129640
rect 42580 129560 42590 129640
rect 42720 129560 42730 129640
rect 42860 129560 42870 129640
rect 43000 129560 43010 129640
rect 43140 129560 43150 129640
rect 43280 129560 43290 129640
rect 43420 129560 43430 129640
rect 43560 129560 43570 129640
rect 43700 129560 43710 129640
rect 146380 129581 146390 129640
rect 146520 129581 146530 129640
rect 146660 129581 146670 129640
rect 146800 129581 146810 129640
rect 146940 129581 146950 129640
rect 147080 129581 147090 129640
rect 147220 129581 147230 129640
rect 147360 129581 147370 129640
rect 147500 129581 147510 129640
rect 147640 129581 147650 129640
rect 148680 129581 148690 129640
rect 148820 129581 148830 129640
rect 148960 129581 148970 129640
rect 149100 129581 149110 129640
rect 149240 129581 149250 129640
rect 149380 129581 149390 129640
rect 149520 129581 149530 129640
rect 149660 129581 149670 129640
rect 149800 129581 149810 129640
rect 149940 129581 149950 129640
rect 152160 129581 152170 129640
rect 152340 129581 152350 129640
rect 152520 129581 152530 129640
rect 152700 129581 152710 129640
rect 152880 129581 152890 129640
rect 153060 129581 153070 129640
rect 153240 129581 153250 129640
rect 153420 129581 153430 129640
rect 153600 129581 153610 129640
rect 153780 129581 153790 129640
rect 153960 129581 153970 129640
rect 154140 129581 154150 129640
rect 154320 129581 154330 129640
rect 154500 129581 154510 129640
rect 154680 129581 154690 129640
rect 154860 129581 154870 129640
rect 155040 129581 155050 129640
rect 155220 129581 155230 129640
rect 155400 129581 155410 129640
rect 155580 129581 155590 129640
rect 155760 129581 155770 129640
rect 155940 129581 155950 129640
rect 156120 129581 156130 129640
rect 156300 129581 156310 129640
rect 156480 129581 156490 129640
rect 156660 129581 156670 129640
rect 156840 129581 156850 129640
rect 157020 129581 157030 129640
rect 157200 129581 157210 129640
rect 157380 129581 157390 129640
rect 157560 129581 157570 129640
rect 157740 129581 157750 129640
rect 157920 129581 157930 129640
rect 158100 129581 158110 129640
rect 158280 129581 158290 129640
rect 158460 129581 158470 129640
rect 158640 129581 158650 129640
rect 158820 129581 158830 129640
rect 159000 129581 159010 129640
rect 159180 129581 159190 129640
rect 159360 129581 159370 129640
rect 159540 129581 159550 129640
rect 159720 129581 159730 129640
rect 163460 129581 163470 129640
rect 163640 129581 163650 129640
rect 163820 129581 163830 129640
rect 164000 129581 164010 129640
rect 164180 129581 164190 129640
rect 164360 129581 164370 129640
rect 164540 129581 164550 129640
rect 164720 129581 164730 129640
rect 164900 129581 164910 129640
rect 165080 129581 165090 129640
rect 165260 129581 165270 129640
rect 165440 129581 165450 129640
rect 165620 129581 165630 129640
rect 165800 129581 165810 129640
rect 165980 129581 165990 129640
rect 166160 129581 166170 129640
rect 166340 129581 166350 129640
rect 166520 129581 166530 129640
rect 166700 129581 166710 129640
rect 166880 129581 166890 129640
rect 167060 129581 167070 129640
rect 167240 129581 167250 129640
rect 167420 129581 167430 129640
rect 167600 129581 167610 129640
rect 167780 129581 167790 129640
rect 167960 129581 167970 129640
rect 168140 129581 168150 129640
rect 168320 129581 168330 129640
rect 168500 129581 168510 129640
rect 168680 129581 168690 129640
rect 168860 129581 168870 129640
rect 169040 129581 169050 129640
rect 169220 129581 169230 129640
rect 169400 129581 169410 129640
rect 169580 129581 169590 129640
rect 169760 129581 169770 129640
rect 169940 129581 169950 129640
rect 170120 129581 170130 129640
rect 170300 129581 170310 129640
rect 170480 129581 170490 129640
rect 170660 129581 170670 129640
rect 170840 129581 170850 129640
rect 171020 129581 171030 129640
rect 146040 129500 147700 129581
rect 148340 129500 150000 129581
rect 152000 129500 159800 129581
rect 163210 129560 171100 129581
rect 163300 129500 171100 129560
rect 30360 129420 30440 129430
rect 30680 129420 30760 129430
rect 31000 129420 31080 129430
rect 31320 129420 31400 129430
rect 31640 129420 31720 129430
rect 31960 129420 32040 129430
rect 32280 129420 32360 129430
rect 32600 129420 32680 129430
rect 32920 129420 33000 129430
rect 33240 129420 33320 129430
rect 33560 129420 33640 129430
rect 33880 129420 33960 129430
rect 34200 129420 34280 129430
rect 34520 129420 34600 129430
rect 34840 129420 34920 129430
rect 35160 129420 35240 129430
rect 35480 129420 35560 129430
rect 35800 129420 35880 129430
rect 36120 129420 36200 129430
rect 36440 129420 36520 129430
rect 36760 129420 36840 129430
rect 37080 129420 37160 129430
rect 37400 129420 37480 129430
rect 37720 129420 37800 129430
rect 40180 129420 40260 129430
rect 40500 129420 40580 129430
rect 40820 129420 40900 129430
rect 41140 129420 41220 129430
rect 42560 129420 42640 129430
rect 42880 129420 42960 129430
rect 43200 129420 43280 129430
rect 43520 129420 43600 129430
rect 18970 129390 19050 129400
rect 19290 129390 19370 129400
rect 19610 129390 19690 129400
rect 19930 129390 20010 129400
rect 20250 129390 20330 129400
rect 20570 129390 20650 129400
rect 20890 129390 20970 129400
rect 21210 129390 21290 129400
rect 21530 129390 21610 129400
rect 21850 129390 21930 129400
rect 22170 129390 22250 129400
rect 22490 129390 22570 129400
rect 22810 129390 22890 129400
rect 23130 129390 23210 129400
rect 23450 129390 23530 129400
rect 23770 129390 23850 129400
rect 24090 129390 24170 129400
rect 24410 129390 24490 129400
rect 24730 129390 24810 129400
rect 25050 129390 25130 129400
rect 25370 129390 25450 129400
rect 25690 129390 25770 129400
rect 26010 129390 26090 129400
rect 26330 129390 26410 129400
rect 19050 129310 19060 129390
rect 19370 129310 19380 129390
rect 19690 129310 19700 129390
rect 20010 129310 20020 129390
rect 20330 129310 20340 129390
rect 20650 129310 20660 129390
rect 20970 129310 20980 129390
rect 21290 129310 21300 129390
rect 21610 129310 21620 129390
rect 21930 129310 21940 129390
rect 22250 129310 22260 129390
rect 22570 129310 22580 129390
rect 22890 129310 22900 129390
rect 23210 129310 23220 129390
rect 23530 129310 23540 129390
rect 23850 129310 23860 129390
rect 24170 129310 24180 129390
rect 24490 129310 24500 129390
rect 24810 129310 24820 129390
rect 25130 129310 25140 129390
rect 25450 129310 25460 129390
rect 25770 129310 25780 129390
rect 26090 129310 26100 129390
rect 26410 129310 26420 129390
rect 30440 129340 30450 129420
rect 30760 129340 30770 129420
rect 31080 129340 31090 129420
rect 31400 129340 31410 129420
rect 31720 129340 31730 129420
rect 32040 129340 32050 129420
rect 32360 129340 32370 129420
rect 32680 129340 32690 129420
rect 33000 129340 33010 129420
rect 33320 129340 33330 129420
rect 33640 129340 33650 129420
rect 33960 129340 33970 129420
rect 34280 129340 34290 129420
rect 34600 129340 34610 129420
rect 34920 129340 34930 129420
rect 35240 129340 35250 129420
rect 35560 129340 35570 129420
rect 35880 129340 35890 129420
rect 36200 129340 36210 129420
rect 36520 129340 36530 129420
rect 36840 129340 36850 129420
rect 37160 129340 37170 129420
rect 37480 129340 37490 129420
rect 37800 129340 37810 129420
rect 40260 129340 40270 129420
rect 40580 129340 40590 129420
rect 40900 129340 40910 129420
rect 41220 129340 41230 129420
rect 42640 129340 42650 129420
rect 42960 129340 42970 129420
rect 43280 129340 43290 129420
rect 43600 129340 43610 129420
rect 146400 129411 146480 129421
rect 146720 129411 146800 129421
rect 147040 129411 147120 129421
rect 147360 129411 147440 129421
rect 148780 129411 148860 129421
rect 149100 129411 149180 129421
rect 149420 129411 149500 129421
rect 149740 129411 149820 129421
rect 152200 129411 152280 129421
rect 152520 129411 152600 129421
rect 152840 129411 152920 129421
rect 153160 129411 153240 129421
rect 153480 129411 153560 129421
rect 153800 129411 153880 129421
rect 154120 129411 154200 129421
rect 154440 129411 154520 129421
rect 154760 129411 154840 129421
rect 155080 129411 155160 129421
rect 155400 129411 155480 129421
rect 155720 129411 155800 129421
rect 156040 129411 156120 129421
rect 156360 129411 156440 129421
rect 156680 129411 156760 129421
rect 157000 129411 157080 129421
rect 157320 129411 157400 129421
rect 157640 129411 157720 129421
rect 157960 129411 158040 129421
rect 158280 129411 158360 129421
rect 158600 129411 158680 129421
rect 158920 129411 159000 129421
rect 159240 129411 159320 129421
rect 159560 129411 159640 129421
rect 146480 129331 146490 129411
rect 146800 129331 146810 129411
rect 147120 129331 147130 129411
rect 147440 129331 147450 129411
rect 148860 129331 148870 129411
rect 149180 129331 149190 129411
rect 149500 129331 149510 129411
rect 149820 129331 149830 129411
rect 152280 129331 152290 129411
rect 152600 129331 152610 129411
rect 152920 129331 152930 129411
rect 153240 129331 153250 129411
rect 153560 129331 153570 129411
rect 153880 129331 153890 129411
rect 154200 129331 154210 129411
rect 154520 129331 154530 129411
rect 154840 129331 154850 129411
rect 155160 129331 155170 129411
rect 155480 129331 155490 129411
rect 155800 129331 155810 129411
rect 156120 129331 156130 129411
rect 156440 129331 156450 129411
rect 156760 129331 156770 129411
rect 157080 129331 157090 129411
rect 157400 129331 157410 129411
rect 157720 129331 157730 129411
rect 158040 129331 158050 129411
rect 158360 129331 158370 129411
rect 158680 129331 158690 129411
rect 159000 129331 159010 129411
rect 159320 129331 159330 129411
rect 159640 129331 159650 129411
rect 163590 129381 163670 129391
rect 163910 129381 163990 129391
rect 164230 129381 164310 129391
rect 164550 129381 164630 129391
rect 164870 129381 164950 129391
rect 165190 129381 165270 129391
rect 165510 129381 165590 129391
rect 165830 129381 165910 129391
rect 166150 129381 166230 129391
rect 166470 129381 166550 129391
rect 166790 129381 166870 129391
rect 167110 129381 167190 129391
rect 167430 129381 167510 129391
rect 167750 129381 167830 129391
rect 168070 129381 168150 129391
rect 168390 129381 168470 129391
rect 168710 129381 168790 129391
rect 169030 129381 169110 129391
rect 169350 129381 169430 129391
rect 169670 129381 169750 129391
rect 169990 129381 170070 129391
rect 170310 129381 170390 129391
rect 170630 129381 170710 129391
rect 170950 129381 171030 129391
rect 163670 129301 163680 129381
rect 163990 129301 164000 129381
rect 164310 129301 164320 129381
rect 164630 129301 164640 129381
rect 164950 129301 164960 129381
rect 165270 129301 165280 129381
rect 165590 129301 165600 129381
rect 165910 129301 165920 129381
rect 166230 129301 166240 129381
rect 166550 129301 166560 129381
rect 166870 129301 166880 129381
rect 167190 129301 167200 129381
rect 167510 129301 167520 129381
rect 167830 129301 167840 129381
rect 168150 129301 168160 129381
rect 168470 129301 168480 129381
rect 168790 129301 168800 129381
rect 169110 129301 169120 129381
rect 169430 129301 169440 129381
rect 169750 129301 169760 129381
rect 170070 129301 170080 129381
rect 170390 129301 170400 129381
rect 170710 129301 170720 129381
rect 171030 129301 171040 129381
rect 30520 129260 30600 129270
rect 30840 129260 30920 129270
rect 31160 129260 31240 129270
rect 31480 129260 31560 129270
rect 31800 129260 31880 129270
rect 32120 129260 32200 129270
rect 32440 129260 32520 129270
rect 32760 129260 32840 129270
rect 33080 129260 33160 129270
rect 33400 129260 33480 129270
rect 33720 129260 33800 129270
rect 34040 129260 34120 129270
rect 34360 129260 34440 129270
rect 34680 129260 34760 129270
rect 35000 129260 35080 129270
rect 35320 129260 35400 129270
rect 35640 129260 35720 129270
rect 35960 129260 36040 129270
rect 36280 129260 36360 129270
rect 36600 129260 36680 129270
rect 36920 129260 37000 129270
rect 37240 129260 37320 129270
rect 37560 129260 37640 129270
rect 40340 129260 40420 129270
rect 40660 129260 40740 129270
rect 40980 129260 41060 129270
rect 42720 129260 42800 129270
rect 43040 129260 43120 129270
rect 43360 129260 43440 129270
rect 19130 129230 19210 129240
rect 19450 129230 19530 129240
rect 19770 129230 19850 129240
rect 20090 129230 20170 129240
rect 20410 129230 20490 129240
rect 20730 129230 20810 129240
rect 21050 129230 21130 129240
rect 21370 129230 21450 129240
rect 21690 129230 21770 129240
rect 22010 129230 22090 129240
rect 22330 129230 22410 129240
rect 22650 129230 22730 129240
rect 22970 129230 23050 129240
rect 23290 129230 23370 129240
rect 23610 129230 23690 129240
rect 23930 129230 24010 129240
rect 24250 129230 24330 129240
rect 24570 129230 24650 129240
rect 24890 129230 24970 129240
rect 25210 129230 25290 129240
rect 25530 129230 25610 129240
rect 25850 129230 25930 129240
rect 26170 129230 26250 129240
rect 19210 129150 19220 129230
rect 19530 129150 19540 129230
rect 19850 129150 19860 129230
rect 20170 129150 20180 129230
rect 20490 129150 20500 129230
rect 20810 129150 20820 129230
rect 21130 129150 21140 129230
rect 21450 129150 21460 129230
rect 21770 129150 21780 129230
rect 22090 129150 22100 129230
rect 22410 129150 22420 129230
rect 22730 129150 22740 129230
rect 23050 129150 23060 129230
rect 23370 129150 23380 129230
rect 23690 129150 23700 129230
rect 24010 129150 24020 129230
rect 24330 129150 24340 129230
rect 24650 129150 24660 129230
rect 24970 129150 24980 129230
rect 25290 129150 25300 129230
rect 25610 129150 25620 129230
rect 25930 129150 25940 129230
rect 26250 129150 26260 129230
rect 30600 129180 30610 129260
rect 30920 129180 30930 129260
rect 31240 129180 31250 129260
rect 31560 129180 31570 129260
rect 31880 129180 31890 129260
rect 32200 129180 32210 129260
rect 32520 129180 32530 129260
rect 32840 129180 32850 129260
rect 33160 129180 33170 129260
rect 33480 129180 33490 129260
rect 33800 129180 33810 129260
rect 34120 129180 34130 129260
rect 34440 129180 34450 129260
rect 34760 129180 34770 129260
rect 35080 129180 35090 129260
rect 35400 129180 35410 129260
rect 35720 129180 35730 129260
rect 36040 129180 36050 129260
rect 36360 129180 36370 129260
rect 36680 129180 36690 129260
rect 37000 129180 37010 129260
rect 37320 129180 37330 129260
rect 37640 129180 37650 129260
rect 40420 129180 40430 129260
rect 40740 129180 40750 129260
rect 41060 129180 41070 129260
rect 42800 129180 42810 129260
rect 43120 129180 43130 129260
rect 43440 129180 43450 129260
rect 146560 129251 146640 129261
rect 146880 129251 146960 129261
rect 147200 129251 147280 129261
rect 148940 129251 149020 129261
rect 149260 129251 149340 129261
rect 149580 129251 149660 129261
rect 152360 129251 152440 129261
rect 152680 129251 152760 129261
rect 153000 129251 153080 129261
rect 153320 129251 153400 129261
rect 153640 129251 153720 129261
rect 153960 129251 154040 129261
rect 154280 129251 154360 129261
rect 154600 129251 154680 129261
rect 154920 129251 155000 129261
rect 155240 129251 155320 129261
rect 155560 129251 155640 129261
rect 155880 129251 155960 129261
rect 156200 129251 156280 129261
rect 156520 129251 156600 129261
rect 156840 129251 156920 129261
rect 157160 129251 157240 129261
rect 157480 129251 157560 129261
rect 157800 129251 157880 129261
rect 158120 129251 158200 129261
rect 158440 129251 158520 129261
rect 158760 129251 158840 129261
rect 159080 129251 159160 129261
rect 159400 129251 159480 129261
rect 146640 129171 146650 129251
rect 146960 129171 146970 129251
rect 147280 129171 147290 129251
rect 149020 129171 149030 129251
rect 149340 129171 149350 129251
rect 149660 129171 149670 129251
rect 152440 129171 152450 129251
rect 152760 129171 152770 129251
rect 153080 129171 153090 129251
rect 153400 129171 153410 129251
rect 153720 129171 153730 129251
rect 154040 129171 154050 129251
rect 154360 129171 154370 129251
rect 154680 129171 154690 129251
rect 155000 129171 155010 129251
rect 155320 129171 155330 129251
rect 155640 129171 155650 129251
rect 155960 129171 155970 129251
rect 156280 129171 156290 129251
rect 156600 129171 156610 129251
rect 156920 129171 156930 129251
rect 157240 129171 157250 129251
rect 157560 129171 157570 129251
rect 157880 129171 157890 129251
rect 158200 129171 158210 129251
rect 158520 129171 158530 129251
rect 158840 129171 158850 129251
rect 159160 129171 159170 129251
rect 159480 129171 159490 129251
rect 163750 129221 163830 129231
rect 164070 129221 164150 129231
rect 164390 129221 164470 129231
rect 164710 129221 164790 129231
rect 165030 129221 165110 129231
rect 165350 129221 165430 129231
rect 165670 129221 165750 129231
rect 165990 129221 166070 129231
rect 166310 129221 166390 129231
rect 166630 129221 166710 129231
rect 166950 129221 167030 129231
rect 167270 129221 167350 129231
rect 167590 129221 167670 129231
rect 167910 129221 167990 129231
rect 168230 129221 168310 129231
rect 168550 129221 168630 129231
rect 168870 129221 168950 129231
rect 169190 129221 169270 129231
rect 169510 129221 169590 129231
rect 169830 129221 169910 129231
rect 170150 129221 170230 129231
rect 170470 129221 170550 129231
rect 170790 129221 170870 129231
rect 163830 129141 163840 129221
rect 164150 129141 164160 129221
rect 164470 129141 164480 129221
rect 164790 129141 164800 129221
rect 165110 129141 165120 129221
rect 165430 129141 165440 129221
rect 165750 129141 165760 129221
rect 166070 129141 166080 129221
rect 166390 129141 166400 129221
rect 166710 129141 166720 129221
rect 167030 129141 167040 129221
rect 167350 129141 167360 129221
rect 167670 129141 167680 129221
rect 167990 129141 168000 129221
rect 168310 129141 168320 129221
rect 168630 129141 168640 129221
rect 168950 129141 168960 129221
rect 169270 129141 169280 129221
rect 169590 129141 169600 129221
rect 169910 129141 169920 129221
rect 170230 129141 170240 129221
rect 170550 129141 170560 129221
rect 170870 129141 170880 129221
rect 30360 129100 30440 129110
rect 30680 129100 30760 129110
rect 31000 129100 31080 129110
rect 31320 129100 31400 129110
rect 31640 129100 31720 129110
rect 31960 129100 32040 129110
rect 32280 129100 32360 129110
rect 32600 129100 32680 129110
rect 32920 129100 33000 129110
rect 33240 129100 33320 129110
rect 33560 129100 33640 129110
rect 33880 129100 33960 129110
rect 34200 129100 34280 129110
rect 34520 129100 34600 129110
rect 34840 129100 34920 129110
rect 35160 129100 35240 129110
rect 35480 129100 35560 129110
rect 35800 129100 35880 129110
rect 36120 129100 36200 129110
rect 36440 129100 36520 129110
rect 36760 129100 36840 129110
rect 37080 129100 37160 129110
rect 37400 129100 37480 129110
rect 37720 129100 37800 129110
rect 40180 129100 40260 129110
rect 40500 129100 40580 129110
rect 40820 129100 40900 129110
rect 41140 129100 41220 129110
rect 42560 129100 42640 129110
rect 42880 129100 42960 129110
rect 43200 129100 43280 129110
rect 43520 129100 43600 129110
rect 18970 129070 19050 129080
rect 19290 129070 19370 129080
rect 19610 129070 19690 129080
rect 19930 129070 20010 129080
rect 20250 129070 20330 129080
rect 20570 129070 20650 129080
rect 20890 129070 20970 129080
rect 21210 129070 21290 129080
rect 21530 129070 21610 129080
rect 21850 129070 21930 129080
rect 22170 129070 22250 129080
rect 22490 129070 22570 129080
rect 22810 129070 22890 129080
rect 23130 129070 23210 129080
rect 23450 129070 23530 129080
rect 23770 129070 23850 129080
rect 24090 129070 24170 129080
rect 24410 129070 24490 129080
rect 24730 129070 24810 129080
rect 25050 129070 25130 129080
rect 25370 129070 25450 129080
rect 25690 129070 25770 129080
rect 26010 129070 26090 129080
rect 26330 129070 26410 129080
rect 19050 128990 19060 129070
rect 19370 128990 19380 129070
rect 19690 128990 19700 129070
rect 20010 128990 20020 129070
rect 20330 128990 20340 129070
rect 20650 128990 20660 129070
rect 20970 128990 20980 129070
rect 21290 128990 21300 129070
rect 21610 128990 21620 129070
rect 21930 128990 21940 129070
rect 22250 128990 22260 129070
rect 22570 128990 22580 129070
rect 22890 128990 22900 129070
rect 23210 128990 23220 129070
rect 23530 128990 23540 129070
rect 23850 128990 23860 129070
rect 24170 128990 24180 129070
rect 24490 128990 24500 129070
rect 24810 128990 24820 129070
rect 25130 128990 25140 129070
rect 25450 128990 25460 129070
rect 25770 128990 25780 129070
rect 26090 128990 26100 129070
rect 26410 128990 26420 129070
rect 30440 129020 30450 129100
rect 30760 129020 30770 129100
rect 31080 129020 31090 129100
rect 31400 129020 31410 129100
rect 31720 129020 31730 129100
rect 32040 129020 32050 129100
rect 32360 129020 32370 129100
rect 32680 129020 32690 129100
rect 33000 129020 33010 129100
rect 33320 129020 33330 129100
rect 33640 129020 33650 129100
rect 33960 129020 33970 129100
rect 34280 129020 34290 129100
rect 34600 129020 34610 129100
rect 34920 129020 34930 129100
rect 35240 129020 35250 129100
rect 35560 129020 35570 129100
rect 35880 129020 35890 129100
rect 36200 129020 36210 129100
rect 36520 129020 36530 129100
rect 36840 129020 36850 129100
rect 37160 129020 37170 129100
rect 37480 129020 37490 129100
rect 37800 129020 37810 129100
rect 40260 129020 40270 129100
rect 40580 129020 40590 129100
rect 40900 129020 40910 129100
rect 41220 129020 41230 129100
rect 42640 129020 42650 129100
rect 42960 129020 42970 129100
rect 43280 129020 43290 129100
rect 43600 129020 43610 129100
rect 146400 129091 146480 129101
rect 146720 129091 146800 129101
rect 147040 129091 147120 129101
rect 147360 129091 147440 129101
rect 148780 129091 148860 129101
rect 149100 129091 149180 129101
rect 149420 129091 149500 129101
rect 149740 129091 149820 129101
rect 152200 129091 152280 129101
rect 152520 129091 152600 129101
rect 152840 129091 152920 129101
rect 153160 129091 153240 129101
rect 153480 129091 153560 129101
rect 153800 129091 153880 129101
rect 154120 129091 154200 129101
rect 154440 129091 154520 129101
rect 154760 129091 154840 129101
rect 155080 129091 155160 129101
rect 155400 129091 155480 129101
rect 155720 129091 155800 129101
rect 156040 129091 156120 129101
rect 156360 129091 156440 129101
rect 156680 129091 156760 129101
rect 157000 129091 157080 129101
rect 157320 129091 157400 129101
rect 157640 129091 157720 129101
rect 157960 129091 158040 129101
rect 158280 129091 158360 129101
rect 158600 129091 158680 129101
rect 158920 129091 159000 129101
rect 159240 129091 159320 129101
rect 159560 129091 159640 129101
rect 146480 129011 146490 129091
rect 146800 129011 146810 129091
rect 147120 129011 147130 129091
rect 147440 129011 147450 129091
rect 148860 129011 148870 129091
rect 149180 129011 149190 129091
rect 149500 129011 149510 129091
rect 149820 129011 149830 129091
rect 152280 129011 152290 129091
rect 152600 129011 152610 129091
rect 152920 129011 152930 129091
rect 153240 129011 153250 129091
rect 153560 129011 153570 129091
rect 153880 129011 153890 129091
rect 154200 129011 154210 129091
rect 154520 129011 154530 129091
rect 154840 129011 154850 129091
rect 155160 129011 155170 129091
rect 155480 129011 155490 129091
rect 155800 129011 155810 129091
rect 156120 129011 156130 129091
rect 156440 129011 156450 129091
rect 156760 129011 156770 129091
rect 157080 129011 157090 129091
rect 157400 129011 157410 129091
rect 157720 129011 157730 129091
rect 158040 129011 158050 129091
rect 158360 129011 158370 129091
rect 158680 129011 158690 129091
rect 159000 129011 159010 129091
rect 159320 129011 159330 129091
rect 159640 129011 159650 129091
rect 163590 129061 163670 129071
rect 163910 129061 163990 129071
rect 164230 129061 164310 129071
rect 164550 129061 164630 129071
rect 164870 129061 164950 129071
rect 165190 129061 165270 129071
rect 165510 129061 165590 129071
rect 165830 129061 165910 129071
rect 166150 129061 166230 129071
rect 166470 129061 166550 129071
rect 166790 129061 166870 129071
rect 167110 129061 167190 129071
rect 167430 129061 167510 129071
rect 167750 129061 167830 129071
rect 168070 129061 168150 129071
rect 168390 129061 168470 129071
rect 168710 129061 168790 129071
rect 169030 129061 169110 129071
rect 169350 129061 169430 129071
rect 169670 129061 169750 129071
rect 169990 129061 170070 129071
rect 170310 129061 170390 129071
rect 170630 129061 170710 129071
rect 170950 129061 171030 129071
rect 163670 128981 163680 129061
rect 163990 128981 164000 129061
rect 164310 128981 164320 129061
rect 164630 128981 164640 129061
rect 164950 128981 164960 129061
rect 165270 128981 165280 129061
rect 165590 128981 165600 129061
rect 165910 128981 165920 129061
rect 166230 128981 166240 129061
rect 166550 128981 166560 129061
rect 166870 128981 166880 129061
rect 167190 128981 167200 129061
rect 167510 128981 167520 129061
rect 167830 128981 167840 129061
rect 168150 128981 168160 129061
rect 168470 128981 168480 129061
rect 168790 128981 168800 129061
rect 169110 128981 169120 129061
rect 169430 128981 169440 129061
rect 169750 128981 169760 129061
rect 170070 128981 170080 129061
rect 170390 128981 170400 129061
rect 170710 128981 170720 129061
rect 171030 128981 171040 129061
rect 30520 128940 30600 128950
rect 30840 128940 30920 128950
rect 31160 128940 31240 128950
rect 31480 128940 31560 128950
rect 31800 128940 31880 128950
rect 32120 128940 32200 128950
rect 32440 128940 32520 128950
rect 32760 128940 32840 128950
rect 33080 128940 33160 128950
rect 33400 128940 33480 128950
rect 33720 128940 33800 128950
rect 34040 128940 34120 128950
rect 34360 128940 34440 128950
rect 34680 128940 34760 128950
rect 35000 128940 35080 128950
rect 35320 128940 35400 128950
rect 35640 128940 35720 128950
rect 35960 128940 36040 128950
rect 36280 128940 36360 128950
rect 36600 128940 36680 128950
rect 36920 128940 37000 128950
rect 37240 128940 37320 128950
rect 37560 128940 37640 128950
rect 40340 128940 40420 128950
rect 40660 128940 40740 128950
rect 40980 128940 41060 128950
rect 42720 128940 42800 128950
rect 43040 128940 43120 128950
rect 43360 128940 43440 128950
rect 19130 128910 19210 128920
rect 19450 128910 19530 128920
rect 19770 128910 19850 128920
rect 20090 128910 20170 128920
rect 20410 128910 20490 128920
rect 20730 128910 20810 128920
rect 21050 128910 21130 128920
rect 21370 128910 21450 128920
rect 21690 128910 21770 128920
rect 22010 128910 22090 128920
rect 22330 128910 22410 128920
rect 22650 128910 22730 128920
rect 22970 128910 23050 128920
rect 23290 128910 23370 128920
rect 23610 128910 23690 128920
rect 23930 128910 24010 128920
rect 24250 128910 24330 128920
rect 24570 128910 24650 128920
rect 24890 128910 24970 128920
rect 25210 128910 25290 128920
rect 25530 128910 25610 128920
rect 25850 128910 25930 128920
rect 26170 128910 26250 128920
rect 19210 128830 19220 128910
rect 19530 128830 19540 128910
rect 19850 128830 19860 128910
rect 20170 128830 20180 128910
rect 20490 128830 20500 128910
rect 20810 128830 20820 128910
rect 21130 128830 21140 128910
rect 21450 128830 21460 128910
rect 21770 128830 21780 128910
rect 22090 128830 22100 128910
rect 22410 128830 22420 128910
rect 22730 128830 22740 128910
rect 23050 128830 23060 128910
rect 23370 128830 23380 128910
rect 23690 128830 23700 128910
rect 24010 128830 24020 128910
rect 24330 128830 24340 128910
rect 24650 128830 24660 128910
rect 24970 128830 24980 128910
rect 25290 128830 25300 128910
rect 25610 128830 25620 128910
rect 25930 128830 25940 128910
rect 26250 128830 26260 128910
rect 30600 128860 30610 128940
rect 30920 128860 30930 128940
rect 31240 128860 31250 128940
rect 31560 128860 31570 128940
rect 31880 128860 31890 128940
rect 32200 128860 32210 128940
rect 32520 128860 32530 128940
rect 32840 128860 32850 128940
rect 33160 128860 33170 128940
rect 33480 128860 33490 128940
rect 33800 128860 33810 128940
rect 34120 128860 34130 128940
rect 34440 128860 34450 128940
rect 34760 128860 34770 128940
rect 35080 128860 35090 128940
rect 35400 128860 35410 128940
rect 35720 128860 35730 128940
rect 36040 128860 36050 128940
rect 36360 128860 36370 128940
rect 36680 128860 36690 128940
rect 37000 128860 37010 128940
rect 37320 128860 37330 128940
rect 37640 128860 37650 128940
rect 40420 128860 40430 128940
rect 40740 128860 40750 128940
rect 41060 128860 41070 128940
rect 42800 128860 42810 128940
rect 43120 128860 43130 128940
rect 43440 128860 43450 128940
rect 146560 128931 146640 128941
rect 146880 128931 146960 128941
rect 147200 128931 147280 128941
rect 148940 128931 149020 128941
rect 149260 128931 149340 128941
rect 149580 128931 149660 128941
rect 152360 128931 152440 128941
rect 152680 128931 152760 128941
rect 153000 128931 153080 128941
rect 153320 128931 153400 128941
rect 153640 128931 153720 128941
rect 153960 128931 154040 128941
rect 154280 128931 154360 128941
rect 154600 128931 154680 128941
rect 154920 128931 155000 128941
rect 155240 128931 155320 128941
rect 155560 128931 155640 128941
rect 155880 128931 155960 128941
rect 156200 128931 156280 128941
rect 156520 128931 156600 128941
rect 156840 128931 156920 128941
rect 157160 128931 157240 128941
rect 157480 128931 157560 128941
rect 157800 128931 157880 128941
rect 158120 128931 158200 128941
rect 158440 128931 158520 128941
rect 158760 128931 158840 128941
rect 159080 128931 159160 128941
rect 159400 128931 159480 128941
rect 146640 128851 146650 128931
rect 146960 128851 146970 128931
rect 147280 128851 147290 128931
rect 149020 128851 149030 128931
rect 149340 128851 149350 128931
rect 149660 128851 149670 128931
rect 152440 128851 152450 128931
rect 152760 128851 152770 128931
rect 153080 128851 153090 128931
rect 153400 128851 153410 128931
rect 153720 128851 153730 128931
rect 154040 128851 154050 128931
rect 154360 128851 154370 128931
rect 154680 128851 154690 128931
rect 155000 128851 155010 128931
rect 155320 128851 155330 128931
rect 155640 128851 155650 128931
rect 155960 128851 155970 128931
rect 156280 128851 156290 128931
rect 156600 128851 156610 128931
rect 156920 128851 156930 128931
rect 157240 128851 157250 128931
rect 157560 128851 157570 128931
rect 157880 128851 157890 128931
rect 158200 128851 158210 128931
rect 158520 128851 158530 128931
rect 158840 128851 158850 128931
rect 159160 128851 159170 128931
rect 159480 128851 159490 128931
rect 163750 128901 163830 128911
rect 164070 128901 164150 128911
rect 164390 128901 164470 128911
rect 164710 128901 164790 128911
rect 165030 128901 165110 128911
rect 165350 128901 165430 128911
rect 165670 128901 165750 128911
rect 165990 128901 166070 128911
rect 166310 128901 166390 128911
rect 166630 128901 166710 128911
rect 166950 128901 167030 128911
rect 167270 128901 167350 128911
rect 167590 128901 167670 128911
rect 167910 128901 167990 128911
rect 168230 128901 168310 128911
rect 168550 128901 168630 128911
rect 168870 128901 168950 128911
rect 169190 128901 169270 128911
rect 169510 128901 169590 128911
rect 169830 128901 169910 128911
rect 170150 128901 170230 128911
rect 170470 128901 170550 128911
rect 170790 128901 170870 128911
rect 163830 128821 163840 128901
rect 164150 128821 164160 128901
rect 164470 128821 164480 128901
rect 164790 128821 164800 128901
rect 165110 128821 165120 128901
rect 165430 128821 165440 128901
rect 165750 128821 165760 128901
rect 166070 128821 166080 128901
rect 166390 128821 166400 128901
rect 166710 128821 166720 128901
rect 167030 128821 167040 128901
rect 167350 128821 167360 128901
rect 167670 128821 167680 128901
rect 167990 128821 168000 128901
rect 168310 128821 168320 128901
rect 168630 128821 168640 128901
rect 168950 128821 168960 128901
rect 169270 128821 169280 128901
rect 169590 128821 169600 128901
rect 169910 128821 169920 128901
rect 170230 128821 170240 128901
rect 170550 128821 170560 128901
rect 170870 128821 170880 128901
rect 30360 128680 30440 128690
rect 30680 128680 30760 128690
rect 31000 128680 31080 128690
rect 31320 128680 31400 128690
rect 31640 128680 31720 128690
rect 31960 128680 32040 128690
rect 32280 128680 32360 128690
rect 32600 128680 32680 128690
rect 32920 128680 33000 128690
rect 33240 128680 33320 128690
rect 33560 128680 33640 128690
rect 33880 128680 33960 128690
rect 34200 128680 34280 128690
rect 34520 128680 34600 128690
rect 34840 128680 34920 128690
rect 35160 128680 35240 128690
rect 35480 128680 35560 128690
rect 35800 128680 35880 128690
rect 36120 128680 36200 128690
rect 36440 128680 36520 128690
rect 36760 128680 36840 128690
rect 37080 128680 37160 128690
rect 37400 128680 37480 128690
rect 37720 128680 37800 128690
rect 40180 128680 40260 128690
rect 40500 128680 40580 128690
rect 40820 128680 40900 128690
rect 41140 128680 41220 128690
rect 42560 128680 42640 128690
rect 42880 128680 42960 128690
rect 43200 128680 43280 128690
rect 43520 128680 43600 128690
rect 18970 128650 19050 128660
rect 19290 128650 19370 128660
rect 19610 128650 19690 128660
rect 19930 128650 20010 128660
rect 20250 128650 20330 128660
rect 20570 128650 20650 128660
rect 20890 128650 20970 128660
rect 21210 128650 21290 128660
rect 21530 128650 21610 128660
rect 21850 128650 21930 128660
rect 22170 128650 22250 128660
rect 22490 128650 22570 128660
rect 22810 128650 22890 128660
rect 23130 128650 23210 128660
rect 23450 128650 23530 128660
rect 23770 128650 23850 128660
rect 24090 128650 24170 128660
rect 24410 128650 24490 128660
rect 24730 128650 24810 128660
rect 25050 128650 25130 128660
rect 25370 128650 25450 128660
rect 25690 128650 25770 128660
rect 26010 128650 26090 128660
rect 26330 128650 26410 128660
rect 19050 128570 19060 128650
rect 19370 128570 19380 128650
rect 19690 128570 19700 128650
rect 20010 128570 20020 128650
rect 20330 128570 20340 128650
rect 20650 128570 20660 128650
rect 20970 128570 20980 128650
rect 21290 128570 21300 128650
rect 21610 128570 21620 128650
rect 21930 128570 21940 128650
rect 22250 128570 22260 128650
rect 22570 128570 22580 128650
rect 22890 128570 22900 128650
rect 23210 128570 23220 128650
rect 23530 128570 23540 128650
rect 23850 128570 23860 128650
rect 24170 128570 24180 128650
rect 24490 128570 24500 128650
rect 24810 128570 24820 128650
rect 25130 128570 25140 128650
rect 25450 128570 25460 128650
rect 25770 128570 25780 128650
rect 26090 128570 26100 128650
rect 26410 128570 26420 128650
rect 30440 128600 30450 128680
rect 30760 128600 30770 128680
rect 31080 128600 31090 128680
rect 31400 128600 31410 128680
rect 31720 128600 31730 128680
rect 32040 128600 32050 128680
rect 32360 128600 32370 128680
rect 32680 128600 32690 128680
rect 33000 128600 33010 128680
rect 33320 128600 33330 128680
rect 33640 128600 33650 128680
rect 33960 128600 33970 128680
rect 34280 128600 34290 128680
rect 34600 128600 34610 128680
rect 34920 128600 34930 128680
rect 35240 128600 35250 128680
rect 35560 128600 35570 128680
rect 35880 128600 35890 128680
rect 36200 128600 36210 128680
rect 36520 128600 36530 128680
rect 36840 128600 36850 128680
rect 37160 128600 37170 128680
rect 37480 128600 37490 128680
rect 37800 128600 37810 128680
rect 40260 128600 40270 128680
rect 40580 128600 40590 128680
rect 40900 128600 40910 128680
rect 41220 128600 41230 128680
rect 42640 128600 42650 128680
rect 42960 128600 42970 128680
rect 43280 128600 43290 128680
rect 43600 128600 43610 128680
rect 146400 128671 146480 128681
rect 146720 128671 146800 128681
rect 147040 128671 147120 128681
rect 147360 128671 147440 128681
rect 148780 128671 148860 128681
rect 149100 128671 149180 128681
rect 149420 128671 149500 128681
rect 149740 128671 149820 128681
rect 152200 128671 152280 128681
rect 152520 128671 152600 128681
rect 152840 128671 152920 128681
rect 153160 128671 153240 128681
rect 153480 128671 153560 128681
rect 153800 128671 153880 128681
rect 154120 128671 154200 128681
rect 154440 128671 154520 128681
rect 154760 128671 154840 128681
rect 155080 128671 155160 128681
rect 155400 128671 155480 128681
rect 155720 128671 155800 128681
rect 156040 128671 156120 128681
rect 156360 128671 156440 128681
rect 156680 128671 156760 128681
rect 157000 128671 157080 128681
rect 157320 128671 157400 128681
rect 157640 128671 157720 128681
rect 157960 128671 158040 128681
rect 158280 128671 158360 128681
rect 158600 128671 158680 128681
rect 158920 128671 159000 128681
rect 159240 128671 159320 128681
rect 159560 128671 159640 128681
rect 146480 128591 146490 128671
rect 146800 128591 146810 128671
rect 147120 128591 147130 128671
rect 147440 128591 147450 128671
rect 148860 128591 148870 128671
rect 149180 128591 149190 128671
rect 149500 128591 149510 128671
rect 149820 128591 149830 128671
rect 152280 128591 152290 128671
rect 152600 128591 152610 128671
rect 152920 128591 152930 128671
rect 153240 128591 153250 128671
rect 153560 128591 153570 128671
rect 153880 128591 153890 128671
rect 154200 128591 154210 128671
rect 154520 128591 154530 128671
rect 154840 128591 154850 128671
rect 155160 128591 155170 128671
rect 155480 128591 155490 128671
rect 155800 128591 155810 128671
rect 156120 128591 156130 128671
rect 156440 128591 156450 128671
rect 156760 128591 156770 128671
rect 157080 128591 157090 128671
rect 157400 128591 157410 128671
rect 157720 128591 157730 128671
rect 158040 128591 158050 128671
rect 158360 128591 158370 128671
rect 158680 128591 158690 128671
rect 159000 128591 159010 128671
rect 159320 128591 159330 128671
rect 159640 128591 159650 128671
rect 163590 128641 163670 128651
rect 163910 128641 163990 128651
rect 164230 128641 164310 128651
rect 164550 128641 164630 128651
rect 164870 128641 164950 128651
rect 165190 128641 165270 128651
rect 165510 128641 165590 128651
rect 165830 128641 165910 128651
rect 166150 128641 166230 128651
rect 166470 128641 166550 128651
rect 166790 128641 166870 128651
rect 167110 128641 167190 128651
rect 167430 128641 167510 128651
rect 167750 128641 167830 128651
rect 168070 128641 168150 128651
rect 168390 128641 168470 128651
rect 168710 128641 168790 128651
rect 169030 128641 169110 128651
rect 169350 128641 169430 128651
rect 169670 128641 169750 128651
rect 169990 128641 170070 128651
rect 170310 128641 170390 128651
rect 170630 128641 170710 128651
rect 170950 128641 171030 128651
rect 163670 128561 163680 128641
rect 163990 128561 164000 128641
rect 164310 128561 164320 128641
rect 164630 128561 164640 128641
rect 164950 128561 164960 128641
rect 165270 128561 165280 128641
rect 165590 128561 165600 128641
rect 165910 128561 165920 128641
rect 166230 128561 166240 128641
rect 166550 128561 166560 128641
rect 166870 128561 166880 128641
rect 167190 128561 167200 128641
rect 167510 128561 167520 128641
rect 167830 128561 167840 128641
rect 168150 128561 168160 128641
rect 168470 128561 168480 128641
rect 168790 128561 168800 128641
rect 169110 128561 169120 128641
rect 169430 128561 169440 128641
rect 169750 128561 169760 128641
rect 170070 128561 170080 128641
rect 170390 128561 170400 128641
rect 170710 128561 170720 128641
rect 171030 128561 171040 128641
rect 30520 128520 30600 128530
rect 30840 128520 30920 128530
rect 31160 128520 31240 128530
rect 31480 128520 31560 128530
rect 31800 128520 31880 128530
rect 32120 128520 32200 128530
rect 32440 128520 32520 128530
rect 32760 128520 32840 128530
rect 33080 128520 33160 128530
rect 33400 128520 33480 128530
rect 33720 128520 33800 128530
rect 34040 128520 34120 128530
rect 34360 128520 34440 128530
rect 34680 128520 34760 128530
rect 35000 128520 35080 128530
rect 35320 128520 35400 128530
rect 35640 128520 35720 128530
rect 35960 128520 36040 128530
rect 36280 128520 36360 128530
rect 36600 128520 36680 128530
rect 36920 128520 37000 128530
rect 37240 128520 37320 128530
rect 37560 128520 37640 128530
rect 40340 128520 40420 128530
rect 40660 128520 40740 128530
rect 40980 128520 41060 128530
rect 42720 128520 42800 128530
rect 43040 128520 43120 128530
rect 43360 128520 43440 128530
rect 19130 128490 19210 128500
rect 19450 128490 19530 128500
rect 19770 128490 19850 128500
rect 20090 128490 20170 128500
rect 20410 128490 20490 128500
rect 20730 128490 20810 128500
rect 21050 128490 21130 128500
rect 21370 128490 21450 128500
rect 21690 128490 21770 128500
rect 22010 128490 22090 128500
rect 22330 128490 22410 128500
rect 22650 128490 22730 128500
rect 22970 128490 23050 128500
rect 23290 128490 23370 128500
rect 23610 128490 23690 128500
rect 23930 128490 24010 128500
rect 24250 128490 24330 128500
rect 24570 128490 24650 128500
rect 24890 128490 24970 128500
rect 25210 128490 25290 128500
rect 25530 128490 25610 128500
rect 25850 128490 25930 128500
rect 26170 128490 26250 128500
rect 19210 128410 19220 128490
rect 19530 128410 19540 128490
rect 19850 128410 19860 128490
rect 20170 128410 20180 128490
rect 20490 128410 20500 128490
rect 20810 128410 20820 128490
rect 21130 128410 21140 128490
rect 21450 128410 21460 128490
rect 21770 128410 21780 128490
rect 22090 128410 22100 128490
rect 22410 128410 22420 128490
rect 22730 128410 22740 128490
rect 23050 128410 23060 128490
rect 23370 128410 23380 128490
rect 23690 128410 23700 128490
rect 24010 128410 24020 128490
rect 24330 128410 24340 128490
rect 24650 128410 24660 128490
rect 24970 128410 24980 128490
rect 25290 128410 25300 128490
rect 25610 128410 25620 128490
rect 25930 128410 25940 128490
rect 26250 128410 26260 128490
rect 30600 128440 30610 128520
rect 30920 128440 30930 128520
rect 31240 128440 31250 128520
rect 31560 128440 31570 128520
rect 31880 128440 31890 128520
rect 32200 128440 32210 128520
rect 32520 128440 32530 128520
rect 32840 128440 32850 128520
rect 33160 128440 33170 128520
rect 33480 128440 33490 128520
rect 33800 128440 33810 128520
rect 34120 128440 34130 128520
rect 34440 128440 34450 128520
rect 34760 128440 34770 128520
rect 35080 128440 35090 128520
rect 35400 128440 35410 128520
rect 35720 128440 35730 128520
rect 36040 128440 36050 128520
rect 36360 128440 36370 128520
rect 36680 128440 36690 128520
rect 37000 128440 37010 128520
rect 37320 128440 37330 128520
rect 37640 128440 37650 128520
rect 40420 128440 40430 128520
rect 40740 128440 40750 128520
rect 41060 128440 41070 128520
rect 42800 128440 42810 128520
rect 43120 128440 43130 128520
rect 43440 128440 43450 128520
rect 146560 128511 146640 128521
rect 146880 128511 146960 128521
rect 147200 128511 147280 128521
rect 148940 128511 149020 128521
rect 149260 128511 149340 128521
rect 149580 128511 149660 128521
rect 152360 128511 152440 128521
rect 152680 128511 152760 128521
rect 153000 128511 153080 128521
rect 153320 128511 153400 128521
rect 153640 128511 153720 128521
rect 153960 128511 154040 128521
rect 154280 128511 154360 128521
rect 154600 128511 154680 128521
rect 154920 128511 155000 128521
rect 155240 128511 155320 128521
rect 155560 128511 155640 128521
rect 155880 128511 155960 128521
rect 156200 128511 156280 128521
rect 156520 128511 156600 128521
rect 156840 128511 156920 128521
rect 157160 128511 157240 128521
rect 157480 128511 157560 128521
rect 157800 128511 157880 128521
rect 158120 128511 158200 128521
rect 158440 128511 158520 128521
rect 158760 128511 158840 128521
rect 159080 128511 159160 128521
rect 159400 128511 159480 128521
rect 146640 128431 146650 128511
rect 146960 128431 146970 128511
rect 147280 128431 147290 128511
rect 149020 128431 149030 128511
rect 149340 128431 149350 128511
rect 149660 128431 149670 128511
rect 152440 128431 152450 128511
rect 152760 128431 152770 128511
rect 153080 128431 153090 128511
rect 153400 128431 153410 128511
rect 153720 128431 153730 128511
rect 154040 128431 154050 128511
rect 154360 128431 154370 128511
rect 154680 128431 154690 128511
rect 155000 128431 155010 128511
rect 155320 128431 155330 128511
rect 155640 128431 155650 128511
rect 155960 128431 155970 128511
rect 156280 128431 156290 128511
rect 156600 128431 156610 128511
rect 156920 128431 156930 128511
rect 157240 128431 157250 128511
rect 157560 128431 157570 128511
rect 157880 128431 157890 128511
rect 158200 128431 158210 128511
rect 158520 128431 158530 128511
rect 158840 128431 158850 128511
rect 159160 128431 159170 128511
rect 159480 128431 159490 128511
rect 163750 128481 163830 128491
rect 164070 128481 164150 128491
rect 164390 128481 164470 128491
rect 164710 128481 164790 128491
rect 165030 128481 165110 128491
rect 165350 128481 165430 128491
rect 165670 128481 165750 128491
rect 165990 128481 166070 128491
rect 166310 128481 166390 128491
rect 166630 128481 166710 128491
rect 166950 128481 167030 128491
rect 167270 128481 167350 128491
rect 167590 128481 167670 128491
rect 167910 128481 167990 128491
rect 168230 128481 168310 128491
rect 168550 128481 168630 128491
rect 168870 128481 168950 128491
rect 169190 128481 169270 128491
rect 169510 128481 169590 128491
rect 169830 128481 169910 128491
rect 170150 128481 170230 128491
rect 170470 128481 170550 128491
rect 170790 128481 170870 128491
rect 163830 128401 163840 128481
rect 164150 128401 164160 128481
rect 164470 128401 164480 128481
rect 164790 128401 164800 128481
rect 165110 128401 165120 128481
rect 165430 128401 165440 128481
rect 165750 128401 165760 128481
rect 166070 128401 166080 128481
rect 166390 128401 166400 128481
rect 166710 128401 166720 128481
rect 167030 128401 167040 128481
rect 167350 128401 167360 128481
rect 167670 128401 167680 128481
rect 167990 128401 168000 128481
rect 168310 128401 168320 128481
rect 168630 128401 168640 128481
rect 168950 128401 168960 128481
rect 169270 128401 169280 128481
rect 169590 128401 169600 128481
rect 169910 128401 169920 128481
rect 170230 128401 170240 128481
rect 170550 128401 170560 128481
rect 170870 128401 170880 128481
rect 30360 128360 30440 128370
rect 30680 128360 30760 128370
rect 31000 128360 31080 128370
rect 31320 128360 31400 128370
rect 31640 128360 31720 128370
rect 31960 128360 32040 128370
rect 32280 128360 32360 128370
rect 32600 128360 32680 128370
rect 32920 128360 33000 128370
rect 33240 128360 33320 128370
rect 33560 128360 33640 128370
rect 33880 128360 33960 128370
rect 34200 128360 34280 128370
rect 34520 128360 34600 128370
rect 34840 128360 34920 128370
rect 35160 128360 35240 128370
rect 35480 128360 35560 128370
rect 35800 128360 35880 128370
rect 36120 128360 36200 128370
rect 36440 128360 36520 128370
rect 36760 128360 36840 128370
rect 37080 128360 37160 128370
rect 37400 128360 37480 128370
rect 37720 128360 37800 128370
rect 40180 128360 40260 128370
rect 40500 128360 40580 128370
rect 40820 128360 40900 128370
rect 41140 128360 41220 128370
rect 42560 128360 42640 128370
rect 42880 128360 42960 128370
rect 43200 128360 43280 128370
rect 43520 128360 43600 128370
rect 18970 128330 19050 128340
rect 19290 128330 19370 128340
rect 19610 128330 19690 128340
rect 19930 128330 20010 128340
rect 20250 128330 20330 128340
rect 20570 128330 20650 128340
rect 20890 128330 20970 128340
rect 21210 128330 21290 128340
rect 21530 128330 21610 128340
rect 21850 128330 21930 128340
rect 22170 128330 22250 128340
rect 22490 128330 22570 128340
rect 22810 128330 22890 128340
rect 23130 128330 23210 128340
rect 23450 128330 23530 128340
rect 23770 128330 23850 128340
rect 24090 128330 24170 128340
rect 24410 128330 24490 128340
rect 24730 128330 24810 128340
rect 25050 128330 25130 128340
rect 25370 128330 25450 128340
rect 25690 128330 25770 128340
rect 26010 128330 26090 128340
rect 26330 128330 26410 128340
rect 19050 128250 19060 128330
rect 19370 128250 19380 128330
rect 19690 128250 19700 128330
rect 20010 128250 20020 128330
rect 20330 128250 20340 128330
rect 20650 128250 20660 128330
rect 20970 128250 20980 128330
rect 21290 128250 21300 128330
rect 21610 128250 21620 128330
rect 21930 128250 21940 128330
rect 22250 128250 22260 128330
rect 22570 128250 22580 128330
rect 22890 128250 22900 128330
rect 23210 128250 23220 128330
rect 23530 128250 23540 128330
rect 23850 128250 23860 128330
rect 24170 128250 24180 128330
rect 24490 128250 24500 128330
rect 24810 128250 24820 128330
rect 25130 128250 25140 128330
rect 25450 128250 25460 128330
rect 25770 128250 25780 128330
rect 26090 128250 26100 128330
rect 26410 128250 26420 128330
rect 30440 128280 30450 128360
rect 30760 128280 30770 128360
rect 31080 128280 31090 128360
rect 31400 128280 31410 128360
rect 31720 128280 31730 128360
rect 32040 128280 32050 128360
rect 32360 128280 32370 128360
rect 32680 128280 32690 128360
rect 33000 128280 33010 128360
rect 33320 128280 33330 128360
rect 33640 128280 33650 128360
rect 33960 128280 33970 128360
rect 34280 128280 34290 128360
rect 34600 128280 34610 128360
rect 34920 128280 34930 128360
rect 35240 128280 35250 128360
rect 35560 128280 35570 128360
rect 35880 128280 35890 128360
rect 36200 128280 36210 128360
rect 36520 128280 36530 128360
rect 36840 128280 36850 128360
rect 37160 128280 37170 128360
rect 37480 128280 37490 128360
rect 37800 128280 37810 128360
rect 40260 128280 40270 128360
rect 40580 128280 40590 128360
rect 40900 128280 40910 128360
rect 41220 128280 41230 128360
rect 42640 128280 42650 128360
rect 42960 128280 42970 128360
rect 43280 128280 43290 128360
rect 43600 128280 43610 128360
rect 146400 128351 146480 128361
rect 146720 128351 146800 128361
rect 147040 128351 147120 128361
rect 147360 128351 147440 128361
rect 148780 128351 148860 128361
rect 149100 128351 149180 128361
rect 149420 128351 149500 128361
rect 149740 128351 149820 128361
rect 152200 128351 152280 128361
rect 152520 128351 152600 128361
rect 152840 128351 152920 128361
rect 153160 128351 153240 128361
rect 153480 128351 153560 128361
rect 153800 128351 153880 128361
rect 154120 128351 154200 128361
rect 154440 128351 154520 128361
rect 154760 128351 154840 128361
rect 155080 128351 155160 128361
rect 155400 128351 155480 128361
rect 155720 128351 155800 128361
rect 156040 128351 156120 128361
rect 156360 128351 156440 128361
rect 156680 128351 156760 128361
rect 157000 128351 157080 128361
rect 157320 128351 157400 128361
rect 157640 128351 157720 128361
rect 157960 128351 158040 128361
rect 158280 128351 158360 128361
rect 158600 128351 158680 128361
rect 158920 128351 159000 128361
rect 159240 128351 159320 128361
rect 159560 128351 159640 128361
rect 146480 128271 146490 128351
rect 146800 128271 146810 128351
rect 147120 128271 147130 128351
rect 147440 128271 147450 128351
rect 148860 128271 148870 128351
rect 149180 128271 149190 128351
rect 149500 128271 149510 128351
rect 149820 128271 149830 128351
rect 152280 128271 152290 128351
rect 152600 128271 152610 128351
rect 152920 128271 152930 128351
rect 153240 128271 153250 128351
rect 153560 128271 153570 128351
rect 153880 128271 153890 128351
rect 154200 128271 154210 128351
rect 154520 128271 154530 128351
rect 154840 128271 154850 128351
rect 155160 128271 155170 128351
rect 155480 128271 155490 128351
rect 155800 128271 155810 128351
rect 156120 128271 156130 128351
rect 156440 128271 156450 128351
rect 156760 128271 156770 128351
rect 157080 128271 157090 128351
rect 157400 128271 157410 128351
rect 157720 128271 157730 128351
rect 158040 128271 158050 128351
rect 158360 128271 158370 128351
rect 158680 128271 158690 128351
rect 159000 128271 159010 128351
rect 159320 128271 159330 128351
rect 159640 128271 159650 128351
rect 163590 128321 163670 128331
rect 163910 128321 163990 128331
rect 164230 128321 164310 128331
rect 164550 128321 164630 128331
rect 164870 128321 164950 128331
rect 165190 128321 165270 128331
rect 165510 128321 165590 128331
rect 165830 128321 165910 128331
rect 166150 128321 166230 128331
rect 166470 128321 166550 128331
rect 166790 128321 166870 128331
rect 167110 128321 167190 128331
rect 167430 128321 167510 128331
rect 167750 128321 167830 128331
rect 168070 128321 168150 128331
rect 168390 128321 168470 128331
rect 168710 128321 168790 128331
rect 169030 128321 169110 128331
rect 169350 128321 169430 128331
rect 169670 128321 169750 128331
rect 169990 128321 170070 128331
rect 170310 128321 170390 128331
rect 170630 128321 170710 128331
rect 170950 128321 171030 128331
rect 163670 128241 163680 128321
rect 163990 128241 164000 128321
rect 164310 128241 164320 128321
rect 164630 128241 164640 128321
rect 164950 128241 164960 128321
rect 165270 128241 165280 128321
rect 165590 128241 165600 128321
rect 165910 128241 165920 128321
rect 166230 128241 166240 128321
rect 166550 128241 166560 128321
rect 166870 128241 166880 128321
rect 167190 128241 167200 128321
rect 167510 128241 167520 128321
rect 167830 128241 167840 128321
rect 168150 128241 168160 128321
rect 168470 128241 168480 128321
rect 168790 128241 168800 128321
rect 169110 128241 169120 128321
rect 169430 128241 169440 128321
rect 169750 128241 169760 128321
rect 170070 128241 170080 128321
rect 170390 128241 170400 128321
rect 170710 128241 170720 128321
rect 171030 128241 171040 128321
rect 30520 128200 30600 128210
rect 30840 128200 30920 128210
rect 31160 128200 31240 128210
rect 31480 128200 31560 128210
rect 31800 128200 31880 128210
rect 32120 128200 32200 128210
rect 32440 128200 32520 128210
rect 32760 128200 32840 128210
rect 33080 128200 33160 128210
rect 33400 128200 33480 128210
rect 33720 128200 33800 128210
rect 34040 128200 34120 128210
rect 34360 128200 34440 128210
rect 34680 128200 34760 128210
rect 35000 128200 35080 128210
rect 35320 128200 35400 128210
rect 35640 128200 35720 128210
rect 35960 128200 36040 128210
rect 36280 128200 36360 128210
rect 36600 128200 36680 128210
rect 36920 128200 37000 128210
rect 37240 128200 37320 128210
rect 37560 128200 37640 128210
rect 40340 128200 40420 128210
rect 40660 128200 40740 128210
rect 40980 128200 41060 128210
rect 42720 128200 42800 128210
rect 43040 128200 43120 128210
rect 43360 128200 43440 128210
rect 19130 128170 19210 128180
rect 19450 128170 19530 128180
rect 19770 128170 19850 128180
rect 20090 128170 20170 128180
rect 20410 128170 20490 128180
rect 20730 128170 20810 128180
rect 21050 128170 21130 128180
rect 21370 128170 21450 128180
rect 21690 128170 21770 128180
rect 22010 128170 22090 128180
rect 22330 128170 22410 128180
rect 22650 128170 22730 128180
rect 22970 128170 23050 128180
rect 23290 128170 23370 128180
rect 23610 128170 23690 128180
rect 23930 128170 24010 128180
rect 24250 128170 24330 128180
rect 24570 128170 24650 128180
rect 24890 128170 24970 128180
rect 25210 128170 25290 128180
rect 25530 128170 25610 128180
rect 25850 128170 25930 128180
rect 26170 128170 26250 128180
rect 19210 128090 19220 128170
rect 19530 128090 19540 128170
rect 19850 128090 19860 128170
rect 20170 128090 20180 128170
rect 20490 128090 20500 128170
rect 20810 128090 20820 128170
rect 21130 128090 21140 128170
rect 21450 128090 21460 128170
rect 21770 128090 21780 128170
rect 22090 128090 22100 128170
rect 22410 128090 22420 128170
rect 22730 128090 22740 128170
rect 23050 128090 23060 128170
rect 23370 128090 23380 128170
rect 23690 128090 23700 128170
rect 24010 128090 24020 128170
rect 24330 128090 24340 128170
rect 24650 128090 24660 128170
rect 24970 128090 24980 128170
rect 25290 128090 25300 128170
rect 25610 128090 25620 128170
rect 25930 128090 25940 128170
rect 26250 128090 26260 128170
rect 30600 128120 30610 128200
rect 30920 128120 30930 128200
rect 31240 128120 31250 128200
rect 31560 128120 31570 128200
rect 31880 128120 31890 128200
rect 32200 128120 32210 128200
rect 32520 128120 32530 128200
rect 32840 128120 32850 128200
rect 33160 128120 33170 128200
rect 33480 128120 33490 128200
rect 33800 128120 33810 128200
rect 34120 128120 34130 128200
rect 34440 128120 34450 128200
rect 34760 128120 34770 128200
rect 35080 128120 35090 128200
rect 35400 128120 35410 128200
rect 35720 128120 35730 128200
rect 36040 128120 36050 128200
rect 36360 128120 36370 128200
rect 36680 128120 36690 128200
rect 37000 128120 37010 128200
rect 37320 128120 37330 128200
rect 37640 128120 37650 128200
rect 40420 128120 40430 128200
rect 40740 128120 40750 128200
rect 41060 128120 41070 128200
rect 42800 128120 42810 128200
rect 43120 128120 43130 128200
rect 43440 128120 43450 128200
rect 146560 128191 146640 128201
rect 146880 128191 146960 128201
rect 147200 128191 147280 128201
rect 148940 128191 149020 128201
rect 149260 128191 149340 128201
rect 149580 128191 149660 128201
rect 152360 128191 152440 128201
rect 152680 128191 152760 128201
rect 153000 128191 153080 128201
rect 153320 128191 153400 128201
rect 153640 128191 153720 128201
rect 153960 128191 154040 128201
rect 154280 128191 154360 128201
rect 154600 128191 154680 128201
rect 154920 128191 155000 128201
rect 155240 128191 155320 128201
rect 155560 128191 155640 128201
rect 155880 128191 155960 128201
rect 156200 128191 156280 128201
rect 156520 128191 156600 128201
rect 156840 128191 156920 128201
rect 157160 128191 157240 128201
rect 157480 128191 157560 128201
rect 157800 128191 157880 128201
rect 158120 128191 158200 128201
rect 158440 128191 158520 128201
rect 158760 128191 158840 128201
rect 159080 128191 159160 128201
rect 159400 128191 159480 128201
rect 146640 128111 146650 128191
rect 146960 128111 146970 128191
rect 147280 128111 147290 128191
rect 149020 128111 149030 128191
rect 149340 128111 149350 128191
rect 149660 128111 149670 128191
rect 152440 128111 152450 128191
rect 152760 128111 152770 128191
rect 153080 128111 153090 128191
rect 153400 128111 153410 128191
rect 153720 128111 153730 128191
rect 154040 128111 154050 128191
rect 154360 128111 154370 128191
rect 154680 128111 154690 128191
rect 155000 128111 155010 128191
rect 155320 128111 155330 128191
rect 155640 128111 155650 128191
rect 155960 128111 155970 128191
rect 156280 128111 156290 128191
rect 156600 128111 156610 128191
rect 156920 128111 156930 128191
rect 157240 128111 157250 128191
rect 157560 128111 157570 128191
rect 157880 128111 157890 128191
rect 158200 128111 158210 128191
rect 158520 128111 158530 128191
rect 158840 128111 158850 128191
rect 159160 128111 159170 128191
rect 159480 128111 159490 128191
rect 163750 128161 163830 128171
rect 164070 128161 164150 128171
rect 164390 128161 164470 128171
rect 164710 128161 164790 128171
rect 165030 128161 165110 128171
rect 165350 128161 165430 128171
rect 165670 128161 165750 128171
rect 165990 128161 166070 128171
rect 166310 128161 166390 128171
rect 166630 128161 166710 128171
rect 166950 128161 167030 128171
rect 167270 128161 167350 128171
rect 167590 128161 167670 128171
rect 167910 128161 167990 128171
rect 168230 128161 168310 128171
rect 168550 128161 168630 128171
rect 168870 128161 168950 128171
rect 169190 128161 169270 128171
rect 169510 128161 169590 128171
rect 169830 128161 169910 128171
rect 170150 128161 170230 128171
rect 170470 128161 170550 128171
rect 170790 128161 170870 128171
rect 163830 128081 163840 128161
rect 164150 128081 164160 128161
rect 164470 128081 164480 128161
rect 164790 128081 164800 128161
rect 165110 128081 165120 128161
rect 165430 128081 165440 128161
rect 165750 128081 165760 128161
rect 166070 128081 166080 128161
rect 166390 128081 166400 128161
rect 166710 128081 166720 128161
rect 167030 128081 167040 128161
rect 167350 128081 167360 128161
rect 167670 128081 167680 128161
rect 167990 128081 168000 128161
rect 168310 128081 168320 128161
rect 168630 128081 168640 128161
rect 168950 128081 168960 128161
rect 169270 128081 169280 128161
rect 169590 128081 169600 128161
rect 169910 128081 169920 128161
rect 170230 128081 170240 128161
rect 170550 128081 170560 128161
rect 170870 128081 170880 128161
rect 18980 127940 19060 127950
rect 19160 127940 19240 127950
rect 19340 127940 19420 127950
rect 19520 127940 19600 127950
rect 19700 127940 19780 127950
rect 19880 127940 19960 127950
rect 20060 127940 20140 127950
rect 20240 127940 20320 127950
rect 20420 127940 20500 127950
rect 20600 127940 20680 127950
rect 20780 127940 20860 127950
rect 20960 127940 21040 127950
rect 21140 127940 21220 127950
rect 21320 127940 21400 127950
rect 21500 127940 21580 127950
rect 21680 127940 21760 127950
rect 21860 127940 21940 127950
rect 22040 127940 22120 127950
rect 22220 127940 22300 127950
rect 22400 127940 22480 127950
rect 22580 127940 22660 127950
rect 22760 127940 22840 127950
rect 22940 127940 23020 127950
rect 23120 127940 23200 127950
rect 23300 127940 23380 127950
rect 23480 127940 23560 127950
rect 23660 127940 23740 127950
rect 23840 127940 23920 127950
rect 24020 127940 24100 127950
rect 24200 127940 24280 127950
rect 24380 127940 24460 127950
rect 24560 127940 24640 127950
rect 24740 127940 24820 127950
rect 24920 127940 25000 127950
rect 25100 127940 25180 127950
rect 25280 127940 25360 127950
rect 25460 127940 25540 127950
rect 25640 127940 25720 127950
rect 25820 127940 25900 127950
rect 26000 127940 26080 127950
rect 26180 127940 26260 127950
rect 26360 127940 26440 127950
rect 26540 127940 26620 127950
rect 30280 127940 30360 127950
rect 30460 127940 30540 127950
rect 30640 127940 30720 127950
rect 30820 127940 30900 127950
rect 31000 127940 31080 127950
rect 31180 127940 31260 127950
rect 31360 127940 31440 127950
rect 31540 127940 31620 127950
rect 31720 127940 31800 127950
rect 31900 127940 31980 127950
rect 32080 127940 32160 127950
rect 32260 127940 32340 127950
rect 32440 127940 32520 127950
rect 32620 127940 32700 127950
rect 32800 127940 32880 127950
rect 32980 127940 33060 127950
rect 33160 127940 33240 127950
rect 33340 127940 33420 127950
rect 33520 127940 33600 127950
rect 33700 127940 33780 127950
rect 33880 127940 33960 127950
rect 34060 127940 34140 127950
rect 34240 127940 34320 127950
rect 34420 127940 34500 127950
rect 34600 127940 34680 127950
rect 34780 127940 34860 127950
rect 34960 127940 35040 127950
rect 35140 127940 35220 127950
rect 35320 127940 35400 127950
rect 35500 127940 35580 127950
rect 35680 127940 35760 127950
rect 35860 127940 35940 127950
rect 36040 127940 36120 127950
rect 36220 127940 36300 127950
rect 36400 127940 36480 127950
rect 36580 127940 36660 127950
rect 36760 127940 36840 127950
rect 36940 127940 37020 127950
rect 37120 127940 37200 127950
rect 37300 127940 37380 127950
rect 37480 127940 37560 127950
rect 37660 127940 37740 127950
rect 37840 127940 37920 127950
rect 40060 127940 40140 127950
rect 40200 127940 40280 127950
rect 40340 127940 40420 127950
rect 40480 127940 40560 127950
rect 40620 127940 40700 127950
rect 40760 127940 40840 127950
rect 40900 127940 40980 127950
rect 41040 127940 41120 127950
rect 41180 127940 41260 127950
rect 41320 127940 41400 127950
rect 42360 127940 42440 127950
rect 42500 127940 42580 127950
rect 42640 127940 42720 127950
rect 42780 127940 42860 127950
rect 42920 127940 43000 127950
rect 43060 127940 43140 127950
rect 43200 127940 43280 127950
rect 43340 127940 43420 127950
rect 43480 127940 43560 127950
rect 43620 127940 43700 127950
rect 146300 127940 146380 127950
rect 146440 127940 146520 127950
rect 146580 127940 146660 127950
rect 146720 127940 146800 127950
rect 146860 127940 146940 127950
rect 147000 127940 147080 127950
rect 147140 127940 147220 127950
rect 147280 127940 147360 127950
rect 147420 127940 147500 127950
rect 147560 127940 147640 127950
rect 19060 127860 19070 127940
rect 19240 127860 19250 127940
rect 19420 127860 19430 127940
rect 19600 127860 19610 127940
rect 19780 127860 19790 127940
rect 19960 127860 19970 127940
rect 20140 127860 20150 127940
rect 20320 127860 20330 127940
rect 20500 127860 20510 127940
rect 20680 127860 20690 127940
rect 20860 127860 20870 127940
rect 21040 127860 21050 127940
rect 21220 127860 21230 127940
rect 21400 127860 21410 127940
rect 21580 127860 21590 127940
rect 21760 127860 21770 127940
rect 21940 127860 21950 127940
rect 22120 127860 22130 127940
rect 22300 127860 22310 127940
rect 22480 127860 22490 127940
rect 22660 127860 22670 127940
rect 22840 127860 22850 127940
rect 23020 127860 23030 127940
rect 23200 127860 23210 127940
rect 23380 127860 23390 127940
rect 23560 127860 23570 127940
rect 23740 127860 23750 127940
rect 23920 127860 23930 127940
rect 24100 127860 24110 127940
rect 24280 127860 24290 127940
rect 24460 127860 24470 127940
rect 24640 127860 24650 127940
rect 24820 127860 24830 127940
rect 25000 127860 25010 127940
rect 25180 127860 25190 127940
rect 25360 127860 25370 127940
rect 25540 127860 25550 127940
rect 25720 127860 25730 127940
rect 25900 127860 25910 127940
rect 26080 127860 26090 127940
rect 26260 127860 26270 127940
rect 26440 127860 26450 127940
rect 26620 127860 26630 127940
rect 30360 127860 30370 127940
rect 30540 127860 30550 127940
rect 30720 127860 30730 127940
rect 30900 127860 30910 127940
rect 31080 127860 31090 127940
rect 31260 127860 31270 127940
rect 31440 127860 31450 127940
rect 31620 127860 31630 127940
rect 31800 127860 31810 127940
rect 31980 127860 31990 127940
rect 32160 127860 32170 127940
rect 32340 127860 32350 127940
rect 32520 127860 32530 127940
rect 32700 127860 32710 127940
rect 32880 127860 32890 127940
rect 33060 127860 33070 127940
rect 33240 127860 33250 127940
rect 33420 127860 33430 127940
rect 33600 127860 33610 127940
rect 33780 127860 33790 127940
rect 33960 127860 33970 127940
rect 34140 127860 34150 127940
rect 34320 127860 34330 127940
rect 34500 127860 34510 127940
rect 34680 127860 34690 127940
rect 34860 127860 34870 127940
rect 35040 127860 35050 127940
rect 35220 127860 35230 127940
rect 35400 127860 35410 127940
rect 35580 127860 35590 127940
rect 35760 127860 35770 127940
rect 35940 127860 35950 127940
rect 36120 127860 36130 127940
rect 36300 127860 36310 127940
rect 36480 127860 36490 127940
rect 36660 127860 36670 127940
rect 36840 127860 36850 127940
rect 37020 127860 37030 127940
rect 37200 127860 37210 127940
rect 37380 127860 37390 127940
rect 37560 127860 37570 127940
rect 37740 127860 37750 127940
rect 37920 127860 37930 127940
rect 40140 127860 40150 127940
rect 40280 127860 40290 127940
rect 40420 127860 40430 127940
rect 40560 127860 40570 127940
rect 40700 127860 40710 127940
rect 40840 127860 40850 127940
rect 40980 127860 40990 127940
rect 41120 127860 41130 127940
rect 41260 127860 41270 127940
rect 41400 127860 41410 127940
rect 42440 127860 42450 127940
rect 42580 127860 42590 127940
rect 42720 127860 42730 127940
rect 42860 127860 42870 127940
rect 43000 127860 43010 127940
rect 43140 127860 43150 127940
rect 43280 127860 43290 127940
rect 43420 127860 43430 127940
rect 43560 127860 43570 127940
rect 43700 127860 43710 127940
rect 146380 127860 146390 127940
rect 146520 127860 146530 127940
rect 146660 127860 146670 127940
rect 146800 127860 146810 127940
rect 146940 127860 146950 127940
rect 147080 127860 147090 127940
rect 147220 127860 147230 127940
rect 147360 127860 147370 127940
rect 147500 127860 147510 127940
rect 147640 127860 147650 127940
rect 28850 127815 28930 127825
rect 29010 127815 29090 127825
rect 29170 127815 29250 127825
rect 29330 127815 29410 127825
rect 29490 127815 29570 127825
rect 18980 127790 19060 127800
rect 19160 127790 19240 127800
rect 19340 127790 19420 127800
rect 19520 127790 19600 127800
rect 19700 127790 19780 127800
rect 19880 127790 19960 127800
rect 20060 127790 20140 127800
rect 20240 127790 20320 127800
rect 20420 127790 20500 127800
rect 20600 127790 20680 127800
rect 20780 127790 20860 127800
rect 20960 127790 21040 127800
rect 21140 127790 21220 127800
rect 21320 127790 21400 127800
rect 21500 127790 21580 127800
rect 21680 127790 21760 127800
rect 21860 127790 21940 127800
rect 22040 127790 22120 127800
rect 22220 127790 22300 127800
rect 22400 127790 22480 127800
rect 22580 127790 22660 127800
rect 22760 127790 22840 127800
rect 22940 127790 23020 127800
rect 23120 127790 23200 127800
rect 23300 127790 23380 127800
rect 23480 127790 23560 127800
rect 23660 127790 23740 127800
rect 23840 127790 23920 127800
rect 24020 127790 24100 127800
rect 24200 127790 24280 127800
rect 24380 127790 24460 127800
rect 24560 127790 24640 127800
rect 24740 127790 24820 127800
rect 24920 127790 25000 127800
rect 25100 127790 25180 127800
rect 25280 127790 25360 127800
rect 25460 127790 25540 127800
rect 25640 127790 25720 127800
rect 25820 127790 25900 127800
rect 26000 127790 26080 127800
rect 26180 127790 26260 127800
rect 26360 127790 26440 127800
rect 26540 127790 26620 127800
rect 19060 127710 19070 127790
rect 19240 127710 19250 127790
rect 19420 127710 19430 127790
rect 19600 127710 19610 127790
rect 19780 127710 19790 127790
rect 19960 127710 19970 127790
rect 20140 127710 20150 127790
rect 20320 127710 20330 127790
rect 20500 127710 20510 127790
rect 20680 127710 20690 127790
rect 20860 127710 20870 127790
rect 21040 127710 21050 127790
rect 21220 127710 21230 127790
rect 21400 127710 21410 127790
rect 21580 127710 21590 127790
rect 21760 127710 21770 127790
rect 21940 127710 21950 127790
rect 22120 127710 22130 127790
rect 22300 127710 22310 127790
rect 22480 127710 22490 127790
rect 22660 127710 22670 127790
rect 22840 127710 22850 127790
rect 23020 127710 23030 127790
rect 23200 127710 23210 127790
rect 23380 127710 23390 127790
rect 23560 127710 23570 127790
rect 23740 127710 23750 127790
rect 23920 127710 23930 127790
rect 24100 127710 24110 127790
rect 24280 127710 24290 127790
rect 24460 127710 24470 127790
rect 24640 127710 24650 127790
rect 24820 127710 24830 127790
rect 25000 127710 25010 127790
rect 25180 127710 25190 127790
rect 25360 127710 25370 127790
rect 25540 127710 25550 127790
rect 25720 127710 25730 127790
rect 25900 127710 25910 127790
rect 26080 127710 26090 127790
rect 26260 127710 26270 127790
rect 26440 127710 26450 127790
rect 26620 127710 26630 127790
rect 28930 127735 28940 127815
rect 29010 127735 29020 127815
rect 29090 127735 29100 127815
rect 29170 127735 29180 127815
rect 29250 127735 29260 127815
rect 29330 127735 29340 127815
rect 29410 127735 29420 127815
rect 29490 127735 29500 127815
rect 29570 127735 29580 127815
rect 148340 127800 150000 128070
rect 152080 127940 152160 127950
rect 152260 127940 152340 127950
rect 152440 127940 152520 127950
rect 152620 127940 152700 127950
rect 152800 127940 152880 127950
rect 152980 127940 153060 127950
rect 153160 127940 153240 127950
rect 153340 127940 153420 127950
rect 153520 127940 153600 127950
rect 153700 127940 153780 127950
rect 153880 127940 153960 127950
rect 154060 127940 154140 127950
rect 154240 127940 154320 127950
rect 154420 127940 154500 127950
rect 154600 127940 154680 127950
rect 154780 127940 154860 127950
rect 154960 127940 155040 127950
rect 155140 127940 155220 127950
rect 155320 127940 155400 127950
rect 155500 127940 155580 127950
rect 155680 127940 155760 127950
rect 155860 127940 155940 127950
rect 156040 127940 156120 127950
rect 156220 127940 156300 127950
rect 156400 127940 156480 127950
rect 156580 127940 156660 127950
rect 156760 127940 156840 127950
rect 156940 127940 157020 127950
rect 157120 127940 157200 127950
rect 157300 127940 157380 127950
rect 157480 127940 157560 127950
rect 157660 127940 157740 127950
rect 157840 127940 157920 127950
rect 158020 127940 158100 127950
rect 158200 127940 158280 127950
rect 158380 127940 158460 127950
rect 158560 127940 158640 127950
rect 158740 127940 158820 127950
rect 158920 127940 159000 127950
rect 159100 127940 159180 127950
rect 159280 127940 159360 127950
rect 159460 127940 159540 127950
rect 159640 127940 159720 127950
rect 163380 127940 163460 127950
rect 163560 127940 163640 127950
rect 163740 127940 163820 127950
rect 163920 127940 164000 127950
rect 164100 127940 164180 127950
rect 164280 127940 164360 127950
rect 164460 127940 164540 127950
rect 164640 127940 164720 127950
rect 164820 127940 164900 127950
rect 165000 127940 165080 127950
rect 165180 127940 165260 127950
rect 165360 127940 165440 127950
rect 165540 127940 165620 127950
rect 165720 127940 165800 127950
rect 165900 127940 165980 127950
rect 166080 127940 166160 127950
rect 166260 127940 166340 127950
rect 166440 127940 166520 127950
rect 166620 127940 166700 127950
rect 166800 127940 166880 127950
rect 166980 127940 167060 127950
rect 167160 127940 167240 127950
rect 167340 127940 167420 127950
rect 167520 127940 167600 127950
rect 167700 127940 167780 127950
rect 167880 127940 167960 127950
rect 168060 127940 168140 127950
rect 168240 127940 168320 127950
rect 168420 127940 168500 127950
rect 168600 127940 168680 127950
rect 168780 127940 168860 127950
rect 168960 127940 169040 127950
rect 169140 127940 169220 127950
rect 169320 127940 169400 127950
rect 169500 127940 169580 127950
rect 169680 127940 169760 127950
rect 169860 127940 169940 127950
rect 170040 127940 170120 127950
rect 170220 127940 170300 127950
rect 170400 127940 170480 127950
rect 170580 127940 170660 127950
rect 170760 127940 170840 127950
rect 170940 127940 171020 127950
rect 152160 127860 152170 127940
rect 152340 127860 152350 127940
rect 152520 127860 152530 127940
rect 152700 127860 152710 127940
rect 152880 127860 152890 127940
rect 153060 127860 153070 127940
rect 153240 127860 153250 127940
rect 153420 127860 153430 127940
rect 153600 127860 153610 127940
rect 153780 127860 153790 127940
rect 153960 127860 153970 127940
rect 154140 127860 154150 127940
rect 154320 127860 154330 127940
rect 154500 127860 154510 127940
rect 154680 127860 154690 127940
rect 154860 127860 154870 127940
rect 155040 127860 155050 127940
rect 155220 127860 155230 127940
rect 155400 127860 155410 127940
rect 155580 127860 155590 127940
rect 155760 127860 155770 127940
rect 155940 127860 155950 127940
rect 156120 127860 156130 127940
rect 156300 127860 156310 127940
rect 156480 127860 156490 127940
rect 156660 127860 156670 127940
rect 156840 127860 156850 127940
rect 157020 127860 157030 127940
rect 157200 127860 157210 127940
rect 157380 127860 157390 127940
rect 157560 127860 157570 127940
rect 157740 127860 157750 127940
rect 157920 127860 157930 127940
rect 158100 127860 158110 127940
rect 158280 127860 158290 127940
rect 158460 127860 158470 127940
rect 158640 127860 158650 127940
rect 158820 127860 158830 127940
rect 159000 127860 159010 127940
rect 159180 127860 159190 127940
rect 159360 127860 159370 127940
rect 159540 127860 159550 127940
rect 159720 127860 159730 127940
rect 163460 127860 163470 127940
rect 163640 127860 163650 127940
rect 163820 127860 163830 127940
rect 164000 127860 164010 127940
rect 164180 127860 164190 127940
rect 164360 127860 164370 127940
rect 164540 127860 164550 127940
rect 164720 127860 164730 127940
rect 164900 127860 164910 127940
rect 165080 127860 165090 127940
rect 165260 127860 165270 127940
rect 165440 127860 165450 127940
rect 165620 127860 165630 127940
rect 165800 127860 165810 127940
rect 165980 127860 165990 127940
rect 166160 127860 166170 127940
rect 166340 127860 166350 127940
rect 166520 127860 166530 127940
rect 166700 127860 166710 127940
rect 166880 127860 166890 127940
rect 167060 127860 167070 127940
rect 167240 127860 167250 127940
rect 167420 127860 167430 127940
rect 167600 127860 167610 127940
rect 167780 127860 167790 127940
rect 167960 127860 167970 127940
rect 168140 127860 168150 127940
rect 168320 127860 168330 127940
rect 168500 127860 168510 127940
rect 168680 127860 168690 127940
rect 168860 127860 168870 127940
rect 169040 127860 169050 127940
rect 169220 127860 169230 127940
rect 169400 127860 169410 127940
rect 169580 127860 169590 127940
rect 169760 127860 169770 127940
rect 169940 127860 169950 127940
rect 170120 127860 170130 127940
rect 170300 127860 170310 127940
rect 170480 127860 170490 127940
rect 170660 127860 170670 127940
rect 170840 127860 170850 127940
rect 171020 127860 171030 127940
rect 161885 127845 161965 127855
rect 162065 127845 162145 127855
rect 162245 127845 162325 127855
rect 162425 127845 162505 127855
rect 162605 127845 162685 127855
rect 30280 127790 30360 127800
rect 30460 127790 30540 127800
rect 30640 127790 30720 127800
rect 30820 127790 30900 127800
rect 31000 127790 31080 127800
rect 31180 127790 31260 127800
rect 31360 127790 31440 127800
rect 31540 127790 31620 127800
rect 31720 127790 31800 127800
rect 31900 127790 31980 127800
rect 32080 127790 32160 127800
rect 32260 127790 32340 127800
rect 32440 127790 32520 127800
rect 32620 127790 32700 127800
rect 32800 127790 32880 127800
rect 32980 127790 33060 127800
rect 33160 127790 33240 127800
rect 33340 127790 33420 127800
rect 33520 127790 33600 127800
rect 33700 127790 33780 127800
rect 33880 127790 33960 127800
rect 34060 127790 34140 127800
rect 34240 127790 34320 127800
rect 34420 127790 34500 127800
rect 34600 127790 34680 127800
rect 34780 127790 34860 127800
rect 34960 127790 35040 127800
rect 35140 127790 35220 127800
rect 35320 127790 35400 127800
rect 35500 127790 35580 127800
rect 35680 127790 35760 127800
rect 35860 127790 35940 127800
rect 36040 127790 36120 127800
rect 36220 127790 36300 127800
rect 36400 127790 36480 127800
rect 36580 127790 36660 127800
rect 36760 127790 36840 127800
rect 36940 127790 37020 127800
rect 37120 127790 37200 127800
rect 37300 127790 37380 127800
rect 37480 127790 37560 127800
rect 37660 127790 37740 127800
rect 37840 127790 37920 127800
rect 30360 127710 30370 127790
rect 30540 127710 30550 127790
rect 30720 127710 30730 127790
rect 30900 127710 30910 127790
rect 31080 127710 31090 127790
rect 31260 127710 31270 127790
rect 31440 127710 31450 127790
rect 31620 127710 31630 127790
rect 31800 127710 31810 127790
rect 31980 127710 31990 127790
rect 32160 127710 32170 127790
rect 32340 127710 32350 127790
rect 32520 127710 32530 127790
rect 32700 127710 32710 127790
rect 32880 127710 32890 127790
rect 33060 127710 33070 127790
rect 33240 127710 33250 127790
rect 33420 127710 33430 127790
rect 33600 127710 33610 127790
rect 33780 127710 33790 127790
rect 33960 127710 33970 127790
rect 34140 127710 34150 127790
rect 34320 127710 34330 127790
rect 34500 127710 34510 127790
rect 34680 127710 34690 127790
rect 34860 127710 34870 127790
rect 35040 127710 35050 127790
rect 35220 127710 35230 127790
rect 35400 127710 35410 127790
rect 35580 127710 35590 127790
rect 35760 127710 35770 127790
rect 35940 127710 35950 127790
rect 36120 127710 36130 127790
rect 36300 127710 36310 127790
rect 36480 127710 36490 127790
rect 36660 127710 36670 127790
rect 36840 127710 36850 127790
rect 37020 127710 37030 127790
rect 37200 127710 37210 127790
rect 37380 127710 37390 127790
rect 37560 127710 37570 127790
rect 37740 127710 37750 127790
rect 37920 127710 37930 127790
rect 40060 127690 40120 127720
rect 41540 127690 41600 127720
rect 42360 127690 42420 127720
rect 43840 127690 43900 127720
rect 146100 127650 146160 127680
rect 147580 127650 147640 127680
rect 148400 127650 148460 127680
rect 40060 127570 40120 127600
rect 41540 127570 41600 127600
rect 42360 127570 42420 127600
rect 43840 127570 43900 127600
rect 146100 127530 146160 127560
rect 147580 127530 147640 127560
rect 148400 127530 148460 127560
rect 40060 127450 40120 127480
rect 41540 127450 41600 127480
rect 42360 127450 42420 127480
rect 43840 127450 43900 127480
rect 19130 127410 19160 127440
rect 19250 127410 19280 127440
rect 26420 127410 26450 127440
rect 26540 127410 26570 127440
rect 30420 127410 30450 127440
rect 30540 127410 30570 127440
rect 37720 127410 37750 127440
rect 37840 127410 37870 127440
rect 146100 127410 146160 127440
rect 147580 127410 147640 127440
rect 148400 127410 148460 127440
rect 19010 127380 19070 127410
rect 19130 127380 19190 127410
rect 19250 127380 19310 127410
rect 26300 127380 26360 127410
rect 26420 127380 26480 127410
rect 26540 127380 26600 127410
rect 30300 127380 30360 127410
rect 30420 127380 30480 127410
rect 30540 127380 30600 127410
rect 37600 127380 37660 127410
rect 37720 127380 37780 127410
rect 37840 127380 37900 127410
rect 40060 127330 40120 127360
rect 41540 127330 41600 127360
rect 42360 127330 42420 127360
rect 43840 127330 43900 127360
rect 19130 127290 19160 127320
rect 19250 127290 19280 127320
rect 26420 127290 26450 127320
rect 26540 127290 26570 127320
rect 30420 127290 30450 127320
rect 30540 127290 30570 127320
rect 37720 127290 37750 127320
rect 37840 127290 37870 127320
rect 146100 127290 146160 127320
rect 147580 127290 147640 127320
rect 148400 127290 148460 127320
rect 19010 127260 19070 127290
rect 19130 127260 19190 127290
rect 19250 127260 19310 127290
rect 26300 127260 26360 127290
rect 26420 127260 26480 127290
rect 26540 127260 26600 127290
rect 30300 127260 30360 127290
rect 30420 127260 30480 127290
rect 30540 127260 30600 127290
rect 37600 127260 37660 127290
rect 37720 127260 37780 127290
rect 37840 127260 37900 127290
rect 31010 127245 37190 127260
rect 36000 127170 37190 127245
rect 40060 127210 40120 127240
rect 41540 127210 41600 127240
rect 42360 127210 42420 127240
rect 43840 127210 43900 127240
rect 148520 127236 148790 127800
rect 149820 127236 150000 127800
rect 152080 127790 152160 127800
rect 152260 127790 152340 127800
rect 152440 127790 152520 127800
rect 152620 127790 152700 127800
rect 152800 127790 152880 127800
rect 152980 127790 153060 127800
rect 153160 127790 153240 127800
rect 153340 127790 153420 127800
rect 153520 127790 153600 127800
rect 153700 127790 153780 127800
rect 153880 127790 153960 127800
rect 154060 127790 154140 127800
rect 154240 127790 154320 127800
rect 154420 127790 154500 127800
rect 154600 127790 154680 127800
rect 154780 127790 154860 127800
rect 154960 127790 155040 127800
rect 155140 127790 155220 127800
rect 155320 127790 155400 127800
rect 155500 127790 155580 127800
rect 155680 127790 155760 127800
rect 155860 127790 155940 127800
rect 156040 127790 156120 127800
rect 156220 127790 156300 127800
rect 156400 127790 156480 127800
rect 156580 127790 156660 127800
rect 156760 127790 156840 127800
rect 156940 127790 157020 127800
rect 157120 127790 157200 127800
rect 157300 127790 157380 127800
rect 157480 127790 157560 127800
rect 157660 127790 157740 127800
rect 157840 127790 157920 127800
rect 158020 127790 158100 127800
rect 158200 127790 158280 127800
rect 158380 127790 158460 127800
rect 158560 127790 158640 127800
rect 158740 127790 158820 127800
rect 158920 127790 159000 127800
rect 159100 127790 159180 127800
rect 159280 127790 159360 127800
rect 159460 127790 159540 127800
rect 159640 127790 159720 127800
rect 152160 127710 152170 127790
rect 152340 127710 152350 127790
rect 152520 127710 152530 127790
rect 152700 127710 152710 127790
rect 152880 127710 152890 127790
rect 153060 127710 153070 127790
rect 153240 127710 153250 127790
rect 153420 127710 153430 127790
rect 153600 127710 153610 127790
rect 153780 127710 153790 127790
rect 153960 127710 153970 127790
rect 154140 127710 154150 127790
rect 154320 127710 154330 127790
rect 154500 127710 154510 127790
rect 154680 127710 154690 127790
rect 154860 127710 154870 127790
rect 155040 127710 155050 127790
rect 155220 127710 155230 127790
rect 155400 127710 155410 127790
rect 155580 127710 155590 127790
rect 155760 127710 155770 127790
rect 155940 127710 155950 127790
rect 156120 127710 156130 127790
rect 156300 127710 156310 127790
rect 156480 127710 156490 127790
rect 156660 127710 156670 127790
rect 156840 127710 156850 127790
rect 157020 127710 157030 127790
rect 157200 127710 157210 127790
rect 157380 127710 157390 127790
rect 157560 127710 157570 127790
rect 157740 127710 157750 127790
rect 157920 127710 157930 127790
rect 158100 127710 158110 127790
rect 158280 127710 158290 127790
rect 158460 127710 158470 127790
rect 158640 127710 158650 127790
rect 158820 127710 158830 127790
rect 159000 127710 159010 127790
rect 159180 127710 159190 127790
rect 159360 127710 159370 127790
rect 159540 127710 159550 127790
rect 159720 127710 159730 127790
rect 161965 127765 161975 127845
rect 162145 127765 162155 127845
rect 162325 127765 162335 127845
rect 162505 127765 162515 127845
rect 162685 127765 162695 127845
rect 163380 127790 163460 127800
rect 163560 127790 163640 127800
rect 163740 127790 163820 127800
rect 163920 127790 164000 127800
rect 164100 127790 164180 127800
rect 164280 127790 164360 127800
rect 164460 127790 164540 127800
rect 164640 127790 164720 127800
rect 164820 127790 164900 127800
rect 165000 127790 165080 127800
rect 165180 127790 165260 127800
rect 165360 127790 165440 127800
rect 165540 127790 165620 127800
rect 165720 127790 165800 127800
rect 165900 127790 165980 127800
rect 166080 127790 166160 127800
rect 166260 127790 166340 127800
rect 166440 127790 166520 127800
rect 166620 127790 166700 127800
rect 166800 127790 166880 127800
rect 166980 127790 167060 127800
rect 167160 127790 167240 127800
rect 167340 127790 167420 127800
rect 167520 127790 167600 127800
rect 167700 127790 167780 127800
rect 167880 127790 167960 127800
rect 168060 127790 168140 127800
rect 168240 127790 168320 127800
rect 168420 127790 168500 127800
rect 168600 127790 168680 127800
rect 168780 127790 168860 127800
rect 168960 127790 169040 127800
rect 169140 127790 169220 127800
rect 169320 127790 169400 127800
rect 169500 127790 169580 127800
rect 169680 127790 169760 127800
rect 169860 127790 169940 127800
rect 170040 127790 170120 127800
rect 170220 127790 170300 127800
rect 170400 127790 170480 127800
rect 170580 127790 170660 127800
rect 170760 127790 170840 127800
rect 170940 127790 171020 127800
rect 163460 127710 163470 127790
rect 163640 127710 163650 127790
rect 163820 127710 163830 127790
rect 164000 127710 164010 127790
rect 164180 127710 164190 127790
rect 164360 127710 164370 127790
rect 164540 127710 164550 127790
rect 164720 127710 164730 127790
rect 164900 127710 164910 127790
rect 165080 127710 165090 127790
rect 165260 127710 165270 127790
rect 165440 127710 165450 127790
rect 165620 127710 165630 127790
rect 165800 127710 165810 127790
rect 165980 127710 165990 127790
rect 166160 127710 166170 127790
rect 166340 127710 166350 127790
rect 166520 127710 166530 127790
rect 166700 127710 166710 127790
rect 166880 127710 166890 127790
rect 167060 127710 167070 127790
rect 167240 127710 167250 127790
rect 167420 127710 167430 127790
rect 167600 127710 167610 127790
rect 167780 127710 167790 127790
rect 167960 127710 167970 127790
rect 168140 127710 168150 127790
rect 168320 127710 168330 127790
rect 168500 127710 168510 127790
rect 168680 127710 168690 127790
rect 168860 127710 168870 127790
rect 169040 127710 169050 127790
rect 169220 127710 169230 127790
rect 169400 127710 169410 127790
rect 169580 127710 169590 127790
rect 169760 127710 169770 127790
rect 169940 127710 169950 127790
rect 170120 127710 170130 127790
rect 170300 127710 170310 127790
rect 170480 127710 170490 127790
rect 170660 127710 170670 127790
rect 170840 127710 170850 127790
rect 171020 127710 171030 127790
rect 161885 127665 161965 127675
rect 162065 127665 162145 127675
rect 162245 127665 162325 127675
rect 162425 127665 162505 127675
rect 162605 127665 162685 127675
rect 152080 127640 152160 127650
rect 152260 127640 152340 127650
rect 152440 127640 152520 127650
rect 152620 127640 152700 127650
rect 152800 127640 152880 127650
rect 152980 127640 153060 127650
rect 153160 127640 153240 127650
rect 153340 127640 153420 127650
rect 153520 127640 153600 127650
rect 153700 127640 153780 127650
rect 153880 127640 153960 127650
rect 154060 127640 154140 127650
rect 154240 127640 154320 127650
rect 154420 127640 154500 127650
rect 154600 127640 154680 127650
rect 154780 127640 154860 127650
rect 154960 127640 155040 127650
rect 155140 127640 155220 127650
rect 155320 127640 155400 127650
rect 155500 127640 155580 127650
rect 155680 127640 155760 127650
rect 155860 127640 155940 127650
rect 156040 127640 156120 127650
rect 156220 127640 156300 127650
rect 156400 127640 156480 127650
rect 156580 127640 156660 127650
rect 156760 127640 156840 127650
rect 156940 127640 157020 127650
rect 157120 127640 157200 127650
rect 157300 127640 157380 127650
rect 157480 127640 157560 127650
rect 157660 127640 157740 127650
rect 157840 127640 157920 127650
rect 158020 127640 158100 127650
rect 158200 127640 158280 127650
rect 158380 127640 158460 127650
rect 158560 127640 158640 127650
rect 158740 127640 158820 127650
rect 158920 127640 159000 127650
rect 159100 127640 159180 127650
rect 159280 127640 159360 127650
rect 159460 127640 159540 127650
rect 159640 127640 159720 127650
rect 152160 127560 152170 127640
rect 152340 127560 152350 127640
rect 152520 127560 152530 127640
rect 152700 127560 152710 127640
rect 152880 127560 152890 127640
rect 153060 127560 153070 127640
rect 153240 127560 153250 127640
rect 153420 127560 153430 127640
rect 153600 127560 153610 127640
rect 153780 127560 153790 127640
rect 153960 127560 153970 127640
rect 154140 127560 154150 127640
rect 154320 127560 154330 127640
rect 154500 127560 154510 127640
rect 154680 127560 154690 127640
rect 154860 127560 154870 127640
rect 155040 127560 155050 127640
rect 155220 127560 155230 127640
rect 155400 127560 155410 127640
rect 155580 127560 155590 127640
rect 155760 127560 155770 127640
rect 155940 127560 155950 127640
rect 156120 127560 156130 127640
rect 156300 127560 156310 127640
rect 156480 127560 156490 127640
rect 156660 127560 156670 127640
rect 156840 127560 156850 127640
rect 157020 127560 157030 127640
rect 157200 127560 157210 127640
rect 157380 127560 157390 127640
rect 157560 127560 157570 127640
rect 157740 127560 157750 127640
rect 157920 127560 157930 127640
rect 158100 127560 158110 127640
rect 158280 127560 158290 127640
rect 158460 127560 158470 127640
rect 158640 127560 158650 127640
rect 158820 127560 158830 127640
rect 159000 127560 159010 127640
rect 159180 127560 159190 127640
rect 159360 127560 159370 127640
rect 159540 127560 159550 127640
rect 159720 127560 159730 127640
rect 161965 127585 161975 127665
rect 162145 127585 162155 127665
rect 162325 127585 162335 127665
rect 162505 127585 162515 127665
rect 162685 127585 162695 127665
rect 163380 127640 163460 127650
rect 163560 127640 163640 127650
rect 163740 127640 163820 127650
rect 163920 127640 164000 127650
rect 164100 127640 164180 127650
rect 164280 127640 164360 127650
rect 164460 127640 164540 127650
rect 164640 127640 164720 127650
rect 164820 127640 164900 127650
rect 165000 127640 165080 127650
rect 165180 127640 165260 127650
rect 165360 127640 165440 127650
rect 165540 127640 165620 127650
rect 165720 127640 165800 127650
rect 165900 127640 165980 127650
rect 166080 127640 166160 127650
rect 166260 127640 166340 127650
rect 166440 127640 166520 127650
rect 166620 127640 166700 127650
rect 166800 127640 166880 127650
rect 166980 127640 167060 127650
rect 167160 127640 167240 127650
rect 167340 127640 167420 127650
rect 167520 127640 167600 127650
rect 167700 127640 167780 127650
rect 167880 127640 167960 127650
rect 168060 127640 168140 127650
rect 168240 127640 168320 127650
rect 168420 127640 168500 127650
rect 168600 127640 168680 127650
rect 168780 127640 168860 127650
rect 168960 127640 169040 127650
rect 169140 127640 169220 127650
rect 169320 127640 169400 127650
rect 169500 127640 169580 127650
rect 169680 127640 169760 127650
rect 169860 127640 169940 127650
rect 170040 127640 170120 127650
rect 170220 127640 170300 127650
rect 170400 127640 170480 127650
rect 170580 127640 170660 127650
rect 170760 127640 170840 127650
rect 170940 127640 171020 127650
rect 163460 127560 163470 127640
rect 163640 127560 163650 127640
rect 163820 127560 163830 127640
rect 164000 127560 164010 127640
rect 164180 127560 164190 127640
rect 164360 127560 164370 127640
rect 164540 127560 164550 127640
rect 164720 127560 164730 127640
rect 164900 127560 164910 127640
rect 165080 127560 165090 127640
rect 165260 127560 165270 127640
rect 165440 127560 165450 127640
rect 165620 127560 165630 127640
rect 165800 127560 165810 127640
rect 165980 127560 165990 127640
rect 166160 127560 166170 127640
rect 166340 127560 166350 127640
rect 166520 127560 166530 127640
rect 166700 127560 166710 127640
rect 166880 127560 166890 127640
rect 167060 127560 167070 127640
rect 167240 127560 167250 127640
rect 167420 127560 167430 127640
rect 167600 127560 167610 127640
rect 167780 127560 167790 127640
rect 167960 127560 167970 127640
rect 168140 127560 168150 127640
rect 168320 127560 168330 127640
rect 168500 127560 168510 127640
rect 168680 127560 168690 127640
rect 168860 127560 168870 127640
rect 169040 127560 169050 127640
rect 169220 127560 169230 127640
rect 169400 127560 169410 127640
rect 169580 127560 169590 127640
rect 169760 127560 169770 127640
rect 169940 127560 169950 127640
rect 170120 127560 170130 127640
rect 170300 127560 170310 127640
rect 170480 127560 170490 127640
rect 170660 127560 170670 127640
rect 170840 127560 170850 127640
rect 171020 127560 171030 127640
rect 152220 127390 152250 127420
rect 152340 127390 152370 127420
rect 159520 127390 159550 127420
rect 159640 127390 159670 127420
rect 152100 127360 152160 127390
rect 152220 127360 152280 127390
rect 152340 127360 152400 127390
rect 159400 127360 159460 127390
rect 159520 127360 159580 127390
rect 159640 127360 159700 127390
rect 152220 127270 152250 127300
rect 152340 127270 152370 127300
rect 159520 127270 159550 127300
rect 159640 127270 159670 127300
rect 163520 127270 163550 127300
rect 163640 127270 163670 127300
rect 170810 127270 170840 127300
rect 170930 127270 170960 127300
rect 152100 127240 152160 127270
rect 152220 127240 152280 127270
rect 152340 127240 152400 127270
rect 152810 127236 158990 127260
rect 159400 127240 159460 127270
rect 159520 127240 159580 127270
rect 159640 127240 159700 127270
rect 163400 127240 163460 127270
rect 163520 127240 163580 127270
rect 163640 127240 163700 127270
rect 170690 127240 170750 127270
rect 170810 127240 170870 127270
rect 170930 127240 170990 127270
rect 164280 127236 164360 127240
rect 164460 127236 164540 127240
rect 164640 127236 164720 127240
rect 164820 127236 164900 127240
rect 165000 127236 165080 127240
rect 165180 127236 165260 127240
rect 165360 127236 165440 127240
rect 165540 127236 165620 127240
rect 165720 127236 165800 127240
rect 165900 127236 165980 127240
rect 166080 127236 166160 127240
rect 166260 127236 166340 127240
rect 166440 127236 166520 127240
rect 166620 127236 166700 127240
rect 166800 127236 166880 127240
rect 166980 127236 167060 127240
rect 167160 127236 167240 127240
rect 167340 127236 167420 127240
rect 167520 127236 167600 127240
rect 167700 127236 167780 127240
rect 167880 127236 167960 127240
rect 168060 127236 168140 127240
rect 168240 127236 168320 127240
rect 168420 127236 168500 127240
rect 168600 127236 168680 127240
rect 168780 127236 168860 127240
rect 168960 127236 169040 127240
rect 169140 127236 169220 127240
rect 169320 127236 169400 127240
rect 169500 127236 169580 127240
rect 169680 127236 169760 127240
rect 169860 127236 169940 127240
rect 170040 127236 170120 127240
rect 37720 127170 37750 127200
rect 37840 127170 37870 127200
rect 36120 127150 36130 127170
rect 36300 127150 36310 127170
rect 36480 127150 36490 127170
rect 36660 127150 36670 127170
rect 36840 127150 36850 127170
rect 37020 127150 37030 127170
rect 36040 127080 36120 127090
rect 36220 127080 36300 127090
rect 36400 127080 36480 127090
rect 36580 127080 36660 127090
rect 36760 127080 36840 127090
rect 36940 127080 37020 127090
rect 36120 127000 36130 127080
rect 36300 127000 36310 127080
rect 36480 127000 36490 127080
rect 36660 127000 36670 127080
rect 36840 127000 36850 127080
rect 37020 127000 37030 127080
rect 37100 126940 37190 127170
rect 37600 127140 37660 127170
rect 37720 127140 37780 127170
rect 37840 127140 37900 127170
rect 40060 127090 40120 127120
rect 41540 127090 41600 127120
rect 42360 127090 42420 127120
rect 43840 127090 43900 127120
rect 37720 127050 37750 127080
rect 37840 127050 37870 127080
rect 37600 127020 37660 127050
rect 37720 127020 37780 127050
rect 37840 127020 37900 127050
rect 40060 126970 40120 127000
rect 41540 126970 41600 127000
rect 42360 126970 42420 127000
rect 43840 126970 43900 127000
rect 36000 126910 37190 126940
rect 37720 126930 37750 126960
rect 37840 126930 37870 126960
rect 36120 126850 36130 126910
rect 36300 126850 36310 126910
rect 36480 126850 36490 126910
rect 36660 126850 36670 126910
rect 36840 126850 36850 126910
rect 37020 126850 37030 126910
rect 37100 126840 37190 126910
rect 37600 126900 37660 126930
rect 37720 126900 37780 126930
rect 37840 126900 37900 126930
rect 40060 126850 40120 126880
rect 41540 126850 41600 126880
rect 42360 126850 42420 126880
rect 43840 126850 43900 126880
rect 36000 126810 37190 126840
rect 37720 126810 37750 126840
rect 37840 126810 37870 126840
rect 37100 126800 37190 126810
rect 36000 126790 37190 126800
rect 36040 126610 36120 126620
rect 36220 126610 36300 126620
rect 36400 126610 36480 126620
rect 36580 126610 36660 126620
rect 36760 126610 36840 126620
rect 36940 126610 37020 126620
rect 36120 126530 36130 126610
rect 36300 126530 36310 126610
rect 36480 126530 36490 126610
rect 36660 126530 36670 126610
rect 36840 126530 36850 126610
rect 37020 126530 37030 126610
rect 36040 126290 36120 126300
rect 36220 126290 36300 126300
rect 36400 126290 36480 126300
rect 36580 126290 36660 126300
rect 36760 126290 36840 126300
rect 36940 126290 37020 126300
rect 36120 126210 36130 126290
rect 36300 126210 36310 126290
rect 36480 126210 36490 126290
rect 36660 126210 36670 126290
rect 36840 126210 36850 126290
rect 37020 126210 37030 126290
rect 37100 126120 37190 126790
rect 37600 126780 37660 126810
rect 37720 126780 37780 126810
rect 37840 126780 37900 126810
rect 40060 126730 40120 126760
rect 41540 126730 41600 126760
rect 42360 126730 42420 126760
rect 43840 126730 43900 126760
rect 37720 126690 37750 126720
rect 37840 126690 37870 126720
rect 37600 126660 37660 126690
rect 37720 126660 37780 126690
rect 37840 126660 37900 126690
rect 40060 126610 40120 126640
rect 41540 126610 41600 126640
rect 42360 126610 42420 126640
rect 43840 126610 43900 126640
rect 37720 126570 37750 126600
rect 37840 126570 37870 126600
rect 37600 126540 37660 126570
rect 37720 126540 37780 126570
rect 37840 126540 37900 126570
rect 40060 126490 40120 126520
rect 41540 126490 41600 126520
rect 42360 126490 42420 126520
rect 43840 126490 43900 126520
rect 37720 126450 37750 126480
rect 37840 126450 37870 126480
rect 37600 126420 37660 126450
rect 37720 126420 37780 126450
rect 37840 126420 37900 126450
rect 40060 126370 40120 126400
rect 41540 126370 41600 126400
rect 42360 126370 42420 126400
rect 43840 126370 43900 126400
rect 37720 126330 37750 126360
rect 37840 126330 37870 126360
rect 37600 126300 37660 126330
rect 37720 126300 37780 126330
rect 37840 126300 37900 126330
rect 40060 126250 40120 126280
rect 41540 126250 41600 126280
rect 42360 126250 42420 126280
rect 43840 126250 43900 126280
rect 37720 126210 37750 126240
rect 37840 126210 37870 126240
rect 37600 126180 37660 126210
rect 37720 126180 37780 126210
rect 37840 126180 37900 126210
rect 40060 126130 40120 126160
rect 41540 126130 41600 126160
rect 42360 126130 42420 126160
rect 43840 126130 43900 126160
rect 36000 126110 37190 126120
rect 37100 126010 37190 126110
rect 37720 126090 37750 126120
rect 37840 126090 37870 126120
rect 37600 126060 37660 126090
rect 37720 126060 37780 126090
rect 37840 126060 37900 126090
rect 40060 126010 40120 126040
rect 41540 126010 41600 126040
rect 42360 126010 42420 126040
rect 43840 126010 43900 126040
rect 36000 125980 37190 126010
rect 36040 125970 36120 125980
rect 36220 125970 36300 125980
rect 36400 125970 36480 125980
rect 36580 125970 36660 125980
rect 36760 125970 36840 125980
rect 36940 125970 37020 125980
rect 36120 125910 36130 125970
rect 36300 125910 36310 125970
rect 36480 125910 36490 125970
rect 36660 125910 36670 125970
rect 36840 125910 36850 125970
rect 37020 125910 37030 125970
rect 37100 125910 37190 125980
rect 37720 125970 37750 126000
rect 37840 125970 37870 126000
rect 37600 125940 37660 125970
rect 37720 125940 37780 125970
rect 37840 125940 37900 125970
rect 36000 125880 37190 125910
rect 40060 125890 40120 125920
rect 41540 125890 41600 125920
rect 42360 125890 42420 125920
rect 43840 125890 43900 125920
rect 36040 125820 36120 125830
rect 36220 125820 36300 125830
rect 36400 125820 36480 125830
rect 36580 125820 36660 125830
rect 36760 125820 36840 125830
rect 36940 125820 37020 125830
rect 36120 125740 36130 125820
rect 36300 125740 36310 125820
rect 36480 125740 36490 125820
rect 36660 125740 36670 125820
rect 36840 125740 36850 125820
rect 37020 125740 37030 125820
rect 37100 125680 37190 125880
rect 37720 125850 37750 125880
rect 37840 125850 37870 125880
rect 37600 125820 37660 125850
rect 37720 125820 37780 125850
rect 37840 125820 37900 125850
rect 40060 125770 40120 125800
rect 41540 125770 41600 125800
rect 42360 125770 42420 125800
rect 43840 125770 43900 125800
rect 37720 125730 37750 125760
rect 37840 125730 37870 125760
rect 37600 125700 37660 125730
rect 37720 125700 37780 125730
rect 37840 125700 37900 125730
rect 36000 125650 37190 125680
rect 40060 125650 40120 125680
rect 41540 125650 41600 125680
rect 42360 125650 42420 125680
rect 43840 125650 43900 125680
rect 36120 125590 36130 125650
rect 36300 125590 36310 125650
rect 36480 125590 36490 125650
rect 36660 125590 36670 125650
rect 36840 125590 36850 125650
rect 37020 125590 37030 125650
rect 37100 125580 37190 125650
rect 37720 125610 37750 125640
rect 37840 125610 37870 125640
rect 37600 125580 37660 125610
rect 37720 125580 37780 125610
rect 37840 125580 37900 125610
rect 36000 125550 37190 125580
rect 37100 125540 37190 125550
rect 36000 125530 37190 125540
rect 40060 125530 40120 125560
rect 41540 125530 41600 125560
rect 42360 125530 42420 125560
rect 43840 125530 43900 125560
rect 36040 125350 36120 125360
rect 36220 125350 36300 125360
rect 36400 125350 36480 125360
rect 36580 125350 36660 125360
rect 36760 125350 36840 125360
rect 36940 125350 37020 125360
rect 36120 125270 36130 125350
rect 36300 125270 36310 125350
rect 36480 125270 36490 125350
rect 36660 125270 36670 125350
rect 36840 125270 36850 125350
rect 37020 125270 37030 125350
rect 36040 125030 36120 125040
rect 36220 125030 36300 125040
rect 36400 125030 36480 125040
rect 36580 125030 36660 125040
rect 36760 125030 36840 125040
rect 36940 125030 37020 125040
rect 36120 124950 36130 125030
rect 36300 124950 36310 125030
rect 36480 124950 36490 125030
rect 36660 124950 36670 125030
rect 36840 124950 36850 125030
rect 37020 124950 37030 125030
rect 37100 124860 37190 125530
rect 37720 125490 37750 125520
rect 37840 125490 37870 125520
rect 37600 125460 37660 125490
rect 37720 125460 37780 125490
rect 37840 125460 37900 125490
rect 40060 125410 40120 125440
rect 41540 125410 41600 125440
rect 42360 125410 42420 125440
rect 43840 125410 43900 125440
rect 37720 125370 37750 125400
rect 37840 125370 37870 125400
rect 37600 125340 37660 125370
rect 37720 125340 37780 125370
rect 37840 125340 37900 125370
rect 40060 125290 40120 125320
rect 41540 125290 41600 125320
rect 42360 125290 42420 125320
rect 43840 125290 43900 125320
rect 37720 125250 37750 125280
rect 37840 125250 37870 125280
rect 37600 125220 37660 125250
rect 37720 125220 37780 125250
rect 37840 125220 37900 125250
rect 40060 125170 40120 125200
rect 41540 125170 41600 125200
rect 42360 125170 42420 125200
rect 43840 125170 43900 125200
rect 37720 125130 37750 125160
rect 37840 125130 37870 125160
rect 37600 125100 37660 125130
rect 37720 125100 37780 125130
rect 37840 125100 37900 125130
rect 40060 125050 40120 125080
rect 41540 125050 41600 125080
rect 42360 125050 42420 125080
rect 43840 125050 43900 125080
rect 37720 125010 37750 125040
rect 37840 125010 37870 125040
rect 37600 124980 37660 125010
rect 37720 124980 37780 125010
rect 37840 124980 37900 125010
rect 40060 124930 40120 124960
rect 41540 124930 41600 124960
rect 42360 124930 42420 124960
rect 43840 124930 43900 124960
rect 37720 124890 37750 124920
rect 37840 124890 37870 124920
rect 37600 124860 37660 124890
rect 37720 124860 37780 124890
rect 37840 124860 37900 124890
rect 36000 124850 37190 124860
rect 37100 124750 37190 124850
rect 40060 124810 40120 124840
rect 41540 124810 41600 124840
rect 42360 124810 42420 124840
rect 43840 124810 43900 124840
rect 37720 124770 37750 124800
rect 37840 124770 37870 124800
rect 36000 124720 37190 124750
rect 37600 124740 37660 124770
rect 37720 124740 37780 124770
rect 37840 124740 37900 124770
rect 36040 124710 36120 124720
rect 36220 124710 36300 124720
rect 36400 124710 36480 124720
rect 36580 124710 36660 124720
rect 36760 124710 36840 124720
rect 36940 124710 37020 124720
rect 36120 124650 36130 124710
rect 36300 124650 36310 124710
rect 36480 124650 36490 124710
rect 36660 124650 36670 124710
rect 36840 124650 36850 124710
rect 37020 124650 37030 124710
rect 37100 124650 37190 124720
rect 40060 124690 40120 124720
rect 41540 124690 41600 124720
rect 42360 124690 42420 124720
rect 43840 124690 43900 124720
rect 37720 124650 37750 124680
rect 37840 124650 37870 124680
rect 36000 124620 37190 124650
rect 37600 124620 37660 124650
rect 37720 124620 37780 124650
rect 37840 124620 37900 124650
rect 36040 124560 36120 124570
rect 36220 124560 36300 124570
rect 36400 124560 36480 124570
rect 36580 124560 36660 124570
rect 36760 124560 36840 124570
rect 36940 124560 37020 124570
rect 36120 124480 36130 124560
rect 36300 124480 36310 124560
rect 36480 124480 36490 124560
rect 36660 124480 36670 124560
rect 36840 124480 36850 124560
rect 37020 124480 37030 124560
rect 37100 124420 37190 124620
rect 40060 124570 40120 124600
rect 41540 124570 41600 124600
rect 42360 124570 42420 124600
rect 43840 124570 43900 124600
rect 37720 124530 37750 124560
rect 37840 124530 37870 124560
rect 37600 124500 37660 124530
rect 37720 124500 37780 124530
rect 37840 124500 37900 124530
rect 40060 124450 40120 124480
rect 41540 124450 41600 124480
rect 42360 124450 42420 124480
rect 43840 124450 43900 124480
rect 36000 124390 37190 124420
rect 37720 124410 37750 124440
rect 37840 124410 37870 124440
rect 36120 124330 36130 124390
rect 36300 124330 36310 124390
rect 36480 124330 36490 124390
rect 36660 124330 36670 124390
rect 36840 124330 36850 124390
rect 37020 124330 37030 124390
rect 37100 124320 37190 124390
rect 37600 124380 37660 124410
rect 37720 124380 37780 124410
rect 37840 124380 37900 124410
rect 40060 124330 40120 124360
rect 41540 124330 41600 124360
rect 42360 124330 42420 124360
rect 43840 124330 43900 124360
rect 36000 124290 37190 124320
rect 37720 124290 37750 124320
rect 37840 124290 37870 124320
rect 37100 124280 37190 124290
rect 36000 124270 37190 124280
rect 36040 124090 36120 124100
rect 36220 124090 36300 124100
rect 36400 124090 36480 124100
rect 36580 124090 36660 124100
rect 36760 124090 36840 124100
rect 36940 124090 37020 124100
rect 36120 124010 36130 124090
rect 36300 124010 36310 124090
rect 36480 124010 36490 124090
rect 36660 124010 36670 124090
rect 36840 124010 36850 124090
rect 37020 124010 37030 124090
rect 36040 123770 36120 123780
rect 36220 123770 36300 123780
rect 36400 123770 36480 123780
rect 36580 123770 36660 123780
rect 36760 123770 36840 123780
rect 36940 123770 37020 123780
rect 36120 123690 36130 123770
rect 36300 123690 36310 123770
rect 36480 123690 36490 123770
rect 36660 123690 36670 123770
rect 36840 123690 36850 123770
rect 37020 123690 37030 123770
rect 37100 123600 37190 124270
rect 37600 124260 37660 124290
rect 37720 124260 37780 124290
rect 37840 124260 37900 124290
rect 40060 124210 40120 124240
rect 41540 124210 41600 124240
rect 42360 124210 42420 124240
rect 43840 124210 43900 124240
rect 37720 124170 37750 124200
rect 37840 124170 37870 124200
rect 37600 124140 37660 124170
rect 37720 124140 37780 124170
rect 37840 124140 37900 124170
rect 40060 124090 40120 124120
rect 41540 124090 41600 124120
rect 42360 124090 42420 124120
rect 43840 124090 43900 124120
rect 37720 124050 37750 124080
rect 37840 124050 37870 124080
rect 37600 124020 37660 124050
rect 37720 124020 37780 124050
rect 37840 124020 37900 124050
rect 40060 123970 40120 124000
rect 41540 123970 41600 124000
rect 42360 123970 42420 124000
rect 43840 123970 43900 124000
rect 37720 123930 37750 123960
rect 37840 123930 37870 123960
rect 37600 123900 37660 123930
rect 37720 123900 37780 123930
rect 37840 123900 37900 123930
rect 40060 123850 40120 123880
rect 41540 123850 41600 123880
rect 42360 123850 42420 123880
rect 43840 123850 43900 123880
rect 37720 123810 37750 123840
rect 37840 123810 37870 123840
rect 37600 123780 37660 123810
rect 37720 123780 37780 123810
rect 37840 123780 37900 123810
rect 40060 123730 40120 123760
rect 41540 123730 41600 123760
rect 42360 123730 42420 123760
rect 43840 123730 43900 123760
rect 37720 123690 37750 123720
rect 37840 123690 37870 123720
rect 37600 123660 37660 123690
rect 37720 123660 37780 123690
rect 37840 123660 37900 123690
rect 40060 123610 40120 123640
rect 41540 123610 41600 123640
rect 42360 123610 42420 123640
rect 43840 123610 43900 123640
rect 36000 123590 37190 123600
rect 37100 123490 37190 123590
rect 37720 123570 37750 123600
rect 37840 123570 37870 123600
rect 37600 123540 37660 123570
rect 37720 123540 37780 123570
rect 37840 123540 37900 123570
rect 40060 123490 40120 123520
rect 41540 123490 41600 123520
rect 42360 123490 42420 123520
rect 43840 123490 43900 123520
rect 36000 123460 37190 123490
rect 36040 123450 36120 123460
rect 36220 123450 36300 123460
rect 36400 123450 36480 123460
rect 36580 123450 36660 123460
rect 36760 123450 36840 123460
rect 36940 123450 37020 123460
rect 36120 123390 36130 123450
rect 36300 123390 36310 123450
rect 36480 123390 36490 123450
rect 36660 123390 36670 123450
rect 36840 123390 36850 123450
rect 37020 123390 37030 123450
rect 37100 123390 37190 123460
rect 37720 123450 37750 123480
rect 37840 123450 37870 123480
rect 37600 123420 37660 123450
rect 37720 123420 37780 123450
rect 37840 123420 37900 123450
rect 36000 123360 37190 123390
rect 40060 123370 40120 123400
rect 41540 123370 41600 123400
rect 42360 123370 42420 123400
rect 43840 123370 43900 123400
rect 36040 123300 36120 123310
rect 36220 123300 36300 123310
rect 36400 123300 36480 123310
rect 36580 123300 36660 123310
rect 36760 123300 36840 123310
rect 36940 123300 37020 123310
rect 36120 123220 36130 123300
rect 36300 123220 36310 123300
rect 36480 123220 36490 123300
rect 36660 123220 36670 123300
rect 36840 123220 36850 123300
rect 37020 123220 37030 123300
rect 37100 123160 37190 123360
rect 37720 123330 37750 123360
rect 37840 123330 37870 123360
rect 37600 123300 37660 123330
rect 37720 123300 37780 123330
rect 37840 123300 37900 123330
rect 40060 123250 40120 123280
rect 41540 123250 41600 123280
rect 42360 123250 42420 123280
rect 43840 123250 43900 123280
rect 37720 123210 37750 123240
rect 37840 123210 37870 123240
rect 37600 123180 37660 123210
rect 37720 123180 37780 123210
rect 37840 123180 37900 123210
rect 36000 123130 37190 123160
rect 40060 123130 40120 123160
rect 41540 123130 41600 123160
rect 42360 123130 42420 123160
rect 43840 123130 43900 123160
rect 36120 123070 36130 123130
rect 36300 123070 36310 123130
rect 36480 123070 36490 123130
rect 36660 123070 36670 123130
rect 36840 123070 36850 123130
rect 37020 123070 37030 123130
rect 37100 123060 37190 123130
rect 37720 123090 37750 123120
rect 37840 123090 37870 123120
rect 37600 123060 37660 123090
rect 37720 123060 37780 123090
rect 37840 123060 37900 123090
rect 36000 123030 37190 123060
rect 37100 123020 37190 123030
rect 36000 123010 37190 123020
rect 40060 123010 40120 123040
rect 41540 123010 41600 123040
rect 42360 123010 42420 123040
rect 43840 123010 43900 123040
rect 36040 122830 36120 122840
rect 36220 122830 36300 122840
rect 36400 122830 36480 122840
rect 36580 122830 36660 122840
rect 36760 122830 36840 122840
rect 36940 122830 37020 122840
rect 36120 122750 36130 122830
rect 36300 122750 36310 122830
rect 36480 122750 36490 122830
rect 36660 122750 36670 122830
rect 36840 122750 36850 122830
rect 37020 122750 37030 122830
rect 36040 122510 36120 122520
rect 36220 122510 36300 122520
rect 36400 122510 36480 122520
rect 36580 122510 36660 122520
rect 36760 122510 36840 122520
rect 36940 122510 37020 122520
rect 36120 122430 36130 122510
rect 36300 122430 36310 122510
rect 36480 122430 36490 122510
rect 36660 122430 36670 122510
rect 36840 122430 36850 122510
rect 37020 122430 37030 122510
rect 37100 122340 37190 123010
rect 37720 122970 37750 123000
rect 37840 122970 37870 123000
rect 37600 122940 37660 122970
rect 37720 122940 37780 122970
rect 37840 122940 37900 122970
rect 40060 122890 40120 122920
rect 41540 122890 41600 122920
rect 42360 122890 42420 122920
rect 43840 122890 43900 122920
rect 37720 122850 37750 122880
rect 37840 122850 37870 122880
rect 37600 122820 37660 122850
rect 37720 122820 37780 122850
rect 37840 122820 37900 122850
rect 40060 122770 40120 122800
rect 41540 122770 41600 122800
rect 42360 122770 42420 122800
rect 43840 122770 43900 122800
rect 37720 122730 37750 122760
rect 37840 122730 37870 122760
rect 37600 122700 37660 122730
rect 37720 122700 37780 122730
rect 37840 122700 37900 122730
rect 40060 122650 40120 122680
rect 41540 122650 41600 122680
rect 42360 122650 42420 122680
rect 43840 122650 43900 122680
rect 37720 122610 37750 122640
rect 37840 122610 37870 122640
rect 37600 122580 37660 122610
rect 37720 122580 37780 122610
rect 37840 122580 37900 122610
rect 40060 122530 40120 122560
rect 41540 122530 41600 122560
rect 42360 122530 42420 122560
rect 43840 122530 43900 122560
rect 37720 122490 37750 122520
rect 37840 122490 37870 122520
rect 37600 122460 37660 122490
rect 37720 122460 37780 122490
rect 37840 122460 37900 122490
rect 40060 122410 40120 122440
rect 41540 122410 41600 122440
rect 42360 122410 42420 122440
rect 43840 122410 43900 122440
rect 37720 122370 37750 122400
rect 37840 122370 37870 122400
rect 37600 122340 37660 122370
rect 37720 122340 37780 122370
rect 37840 122340 37900 122370
rect 36000 122330 37190 122340
rect 37100 122230 37190 122330
rect 40060 122290 40120 122320
rect 41540 122290 41600 122320
rect 42360 122290 42420 122320
rect 43840 122290 43900 122320
rect 37720 122250 37750 122280
rect 37840 122250 37870 122280
rect 36000 122200 37190 122230
rect 37600 122220 37660 122250
rect 37720 122220 37780 122250
rect 37840 122220 37900 122250
rect 40685 122210 40925 122240
rect 36040 122190 36120 122200
rect 36220 122190 36300 122200
rect 36400 122190 36480 122200
rect 36580 122190 36660 122200
rect 36760 122190 36840 122200
rect 36940 122190 37020 122200
rect 36120 122130 36130 122190
rect 36300 122130 36310 122190
rect 36480 122130 36490 122190
rect 36660 122130 36670 122190
rect 36840 122130 36850 122190
rect 37020 122130 37030 122190
rect 37100 122130 37190 122200
rect 40060 122170 40120 122200
rect 37720 122130 37750 122160
rect 37840 122130 37870 122160
rect 40685 122150 40715 122210
rect 40775 122150 40865 122210
rect 40895 122150 40925 122210
rect 41540 122170 41600 122200
rect 42360 122170 42420 122200
rect 43840 122170 43900 122200
rect 36000 122100 37190 122130
rect 37600 122100 37660 122130
rect 37720 122100 37780 122130
rect 37840 122100 37900 122130
rect 40685 122120 40925 122150
rect 36040 122040 36120 122050
rect 36220 122040 36300 122050
rect 36400 122040 36480 122050
rect 36580 122040 36660 122050
rect 36760 122040 36840 122050
rect 36940 122040 37020 122050
rect 36120 121960 36130 122040
rect 36300 121960 36310 122040
rect 36480 121960 36490 122040
rect 36660 121960 36670 122040
rect 36840 121960 36850 122040
rect 37020 121960 37030 122040
rect 37100 121900 37190 122100
rect 40060 122050 40120 122080
rect 41540 122050 41600 122080
rect 42360 122050 42420 122080
rect 43840 122050 43900 122080
rect 37720 122010 37750 122040
rect 37840 122010 37870 122040
rect 37600 121980 37660 122010
rect 37720 121980 37780 122010
rect 37840 121980 37900 122010
rect 40060 121930 40120 121960
rect 41540 121930 41600 121960
rect 42360 121930 42420 121960
rect 43840 121930 43900 121960
rect 36000 121870 37190 121900
rect 37720 121890 37750 121920
rect 37840 121890 37870 121920
rect 36120 121810 36130 121870
rect 36300 121810 36310 121870
rect 36480 121810 36490 121870
rect 36660 121810 36670 121870
rect 36840 121810 36850 121870
rect 37020 121810 37030 121870
rect 37100 121800 37190 121870
rect 37600 121860 37660 121890
rect 37720 121860 37780 121890
rect 37840 121860 37900 121890
rect 40060 121810 40120 121840
rect 41540 121810 41600 121840
rect 42360 121810 42420 121840
rect 43840 121810 43900 121840
rect 36000 121770 37190 121800
rect 37720 121770 37750 121800
rect 37840 121770 37870 121800
rect 37100 121760 37190 121770
rect 36000 121750 37190 121760
rect 36040 121570 36120 121580
rect 36220 121570 36300 121580
rect 36400 121570 36480 121580
rect 36580 121570 36660 121580
rect 36760 121570 36840 121580
rect 36940 121570 37020 121580
rect 36120 121490 36130 121570
rect 36300 121490 36310 121570
rect 36480 121490 36490 121570
rect 36660 121490 36670 121570
rect 36840 121490 36850 121570
rect 37020 121490 37030 121570
rect 36040 121250 36120 121260
rect 36220 121250 36300 121260
rect 36400 121250 36480 121260
rect 36580 121250 36660 121260
rect 36760 121250 36840 121260
rect 36940 121250 37020 121260
rect 36120 121170 36130 121250
rect 36300 121170 36310 121250
rect 36480 121170 36490 121250
rect 36660 121170 36670 121250
rect 36840 121170 36850 121250
rect 37020 121170 37030 121250
rect 37100 121080 37190 121750
rect 37600 121740 37660 121770
rect 37720 121740 37780 121770
rect 37840 121740 37900 121770
rect 40060 121690 40120 121720
rect 41540 121690 41600 121720
rect 42360 121690 42420 121720
rect 43840 121690 43900 121720
rect 37720 121650 37750 121680
rect 37840 121650 37870 121680
rect 37600 121620 37660 121650
rect 37720 121620 37780 121650
rect 37840 121620 37900 121650
rect 40060 121570 40120 121600
rect 41540 121570 41600 121600
rect 42360 121570 42420 121600
rect 43840 121570 43900 121600
rect 37720 121530 37750 121560
rect 37840 121530 37870 121560
rect 37600 121500 37660 121530
rect 37720 121500 37780 121530
rect 37840 121500 37900 121530
rect 40678 121504 40758 121514
rect 40838 121504 40918 121514
rect 40060 121450 40120 121480
rect 37720 121410 37750 121440
rect 37840 121410 37870 121440
rect 40758 121434 40768 121504
rect 40678 121424 40768 121434
rect 40838 121434 40848 121504
rect 40918 121434 40928 121504
rect 41540 121450 41600 121480
rect 42360 121450 42420 121480
rect 43840 121450 43900 121480
rect 40838 121424 40928 121434
rect 37600 121380 37660 121410
rect 37720 121380 37780 121410
rect 37840 121380 37900 121410
rect 40060 121330 40120 121360
rect 40678 121344 40758 121354
rect 40838 121344 40918 121354
rect 37720 121290 37750 121320
rect 37840 121290 37870 121320
rect 37600 121260 37660 121290
rect 37720 121260 37780 121290
rect 37840 121260 37900 121290
rect 40758 121264 40768 121344
rect 40838 121264 40848 121344
rect 40918 121264 40928 121344
rect 41540 121330 41600 121360
rect 42360 121330 42420 121360
rect 43840 121330 43900 121360
rect 40060 121210 40120 121240
rect 41540 121210 41600 121240
rect 42360 121210 42420 121240
rect 43840 121210 43900 121240
rect 37720 121170 37750 121200
rect 37840 121170 37870 121200
rect 37600 121140 37660 121170
rect 37720 121140 37780 121170
rect 37840 121140 37900 121170
rect 40060 121090 40120 121120
rect 41540 121090 41600 121120
rect 42360 121090 42420 121120
rect 43840 121090 43900 121120
rect 36000 121070 37190 121080
rect 37100 120970 37190 121070
rect 37720 121050 37750 121080
rect 37840 121050 37870 121080
rect 37600 121020 37660 121050
rect 37720 121020 37780 121050
rect 37840 121020 37900 121050
rect 40060 120970 40120 121000
rect 41540 120970 41600 121000
rect 42360 120970 42420 121000
rect 43840 120970 43900 121000
rect 36000 120940 37190 120970
rect 36040 120930 36120 120940
rect 36220 120930 36300 120940
rect 36400 120930 36480 120940
rect 36580 120930 36660 120940
rect 36760 120930 36840 120940
rect 36940 120930 37020 120940
rect 36120 120870 36130 120930
rect 36300 120870 36310 120930
rect 36480 120870 36490 120930
rect 36660 120870 36670 120930
rect 36840 120870 36850 120930
rect 37020 120870 37030 120930
rect 37100 120870 37190 120940
rect 37720 120930 37750 120960
rect 37840 120930 37870 120960
rect 37600 120900 37660 120930
rect 37720 120900 37780 120930
rect 37840 120900 37900 120930
rect 36000 120840 37190 120870
rect 40060 120850 40120 120880
rect 41540 120850 41600 120880
rect 42360 120850 42420 120880
rect 43840 120850 43900 120880
rect 36040 120780 36120 120790
rect 36220 120780 36300 120790
rect 36400 120780 36480 120790
rect 36580 120780 36660 120790
rect 36760 120780 36840 120790
rect 36940 120780 37020 120790
rect 36120 120700 36130 120780
rect 36300 120700 36310 120780
rect 36480 120700 36490 120780
rect 36660 120700 36670 120780
rect 36840 120700 36850 120780
rect 37020 120700 37030 120780
rect 37100 120640 37190 120840
rect 37720 120810 37750 120840
rect 37840 120810 37870 120840
rect 37600 120780 37660 120810
rect 37720 120780 37780 120810
rect 37840 120780 37900 120810
rect 40060 120730 40120 120760
rect 41540 120730 41600 120760
rect 42360 120730 42420 120760
rect 43840 120730 43900 120760
rect 37720 120690 37750 120720
rect 37840 120690 37870 120720
rect 37600 120660 37660 120690
rect 37720 120660 37780 120690
rect 37840 120660 37900 120690
rect 36000 120610 37190 120640
rect 40060 120610 40120 120640
rect 41540 120610 41600 120640
rect 42360 120610 42420 120640
rect 43840 120610 43900 120640
rect 36120 120550 36130 120610
rect 36300 120550 36310 120610
rect 36480 120550 36490 120610
rect 36660 120550 36670 120610
rect 36840 120550 36850 120610
rect 37020 120550 37030 120610
rect 37100 120540 37190 120610
rect 37720 120570 37750 120600
rect 37840 120570 37870 120600
rect 37600 120540 37660 120570
rect 37720 120540 37780 120570
rect 37840 120540 37900 120570
rect 36000 120510 37190 120540
rect 37100 120500 37190 120510
rect 36000 120490 37190 120500
rect 40060 120490 40120 120520
rect 41540 120490 41600 120520
rect 42360 120490 42420 120520
rect 43840 120490 43900 120520
rect 36040 120310 36120 120320
rect 36220 120310 36300 120320
rect 36400 120310 36480 120320
rect 36580 120310 36660 120320
rect 36760 120310 36840 120320
rect 36940 120310 37020 120320
rect 36120 120230 36130 120310
rect 36300 120230 36310 120310
rect 36480 120230 36490 120310
rect 36660 120230 36670 120310
rect 36840 120230 36850 120310
rect 37020 120230 37030 120310
rect 36040 119990 36120 120000
rect 36220 119990 36300 120000
rect 36400 119990 36480 120000
rect 36580 119990 36660 120000
rect 36760 119990 36840 120000
rect 36940 119990 37020 120000
rect 36120 119910 36130 119990
rect 36300 119910 36310 119990
rect 36480 119910 36490 119990
rect 36660 119910 36670 119990
rect 36840 119910 36850 119990
rect 37020 119910 37030 119990
rect 37100 119820 37190 120490
rect 37720 120450 37750 120480
rect 37840 120450 37870 120480
rect 42595 120475 42675 120485
rect 37600 120420 37660 120450
rect 37720 120420 37780 120450
rect 37840 120420 37900 120450
rect 42675 120405 42685 120475
rect 40060 120370 40120 120400
rect 41540 120370 41600 120400
rect 42360 120370 42420 120400
rect 42595 120395 42685 120405
rect 43840 120370 43900 120400
rect 37720 120330 37750 120360
rect 37840 120330 37870 120360
rect 37600 120300 37660 120330
rect 37720 120300 37780 120330
rect 37840 120300 37900 120330
rect 42595 120315 42675 120325
rect 40060 120250 40120 120280
rect 41540 120250 41600 120280
rect 42360 120250 42420 120280
rect 37720 120210 37750 120240
rect 37840 120210 37870 120240
rect 42675 120235 42685 120315
rect 43030 120300 43390 120360
rect 43840 120250 43900 120280
rect 38595 120215 38675 120225
rect 38775 120215 38855 120225
rect 38955 120215 39035 120225
rect 39135 120215 39215 120225
rect 39315 120215 39395 120225
rect 37600 120180 37660 120210
rect 37720 120180 37780 120210
rect 37840 120180 37900 120210
rect 38675 120135 38685 120215
rect 38855 120135 38865 120215
rect 39035 120135 39045 120215
rect 39215 120135 39225 120215
rect 39395 120135 39405 120215
rect 43580 120170 43700 120230
rect 40060 120130 40120 120160
rect 41540 120130 41600 120160
rect 42360 120130 42420 120160
rect 42950 120150 43560 120160
rect 43550 120145 43560 120150
rect 42910 120135 43560 120145
rect 37720 120090 37750 120120
rect 37840 120090 37870 120120
rect 37600 120060 37660 120090
rect 37720 120060 37780 120090
rect 37840 120060 37900 120090
rect 42900 120085 42910 120135
rect 38595 120035 38675 120045
rect 38775 120035 38855 120045
rect 38955 120035 39035 120045
rect 39135 120035 39215 120045
rect 39315 120035 39395 120045
rect 43030 120040 43390 120100
rect 37720 119970 37750 120000
rect 37840 119970 37870 120000
rect 37600 119940 37660 119970
rect 37720 119940 37780 119970
rect 37840 119940 37900 119970
rect 38675 119955 38685 120035
rect 38855 119955 38865 120035
rect 39035 119955 39045 120035
rect 39215 119955 39225 120035
rect 39395 119955 39405 120035
rect 40060 120010 40120 120040
rect 41540 120010 41600 120040
rect 42360 120010 42420 120040
rect 42682 119960 42822 120030
rect 40060 119890 40120 119920
rect 40678 119899 40758 119909
rect 40838 119899 40918 119909
rect 37720 119850 37750 119880
rect 37840 119850 37870 119880
rect 38595 119855 38675 119865
rect 38775 119855 38855 119865
rect 38955 119855 39035 119865
rect 39135 119855 39215 119865
rect 39315 119855 39395 119865
rect 37600 119820 37660 119850
rect 37720 119820 37780 119850
rect 37840 119820 37900 119850
rect 36000 119810 37190 119820
rect 37100 119710 37190 119810
rect 38675 119775 38685 119855
rect 38855 119775 38865 119855
rect 39035 119775 39045 119855
rect 39215 119775 39225 119855
rect 39395 119775 39405 119855
rect 40758 119819 40768 119899
rect 40838 119819 40848 119899
rect 40918 119819 40928 119899
rect 41540 119890 41600 119920
rect 42360 119890 42420 119920
rect 42822 119900 42892 119960
rect 42822 119890 43470 119900
rect 43550 119890 43560 120135
rect 43700 120050 43760 120170
rect 43840 120130 43900 120160
rect 43840 120010 43900 120040
rect 43580 119910 43700 119970
rect 42822 119820 42892 119890
rect 42910 119875 43560 119885
rect 42900 119825 42910 119875
rect 40060 119770 40120 119800
rect 37720 119730 37750 119760
rect 37840 119730 37870 119760
rect 40685 119750 40925 119780
rect 41540 119770 41600 119800
rect 42360 119770 42420 119800
rect 42682 119760 42822 119820
rect 43030 119780 43390 119840
rect 43700 119790 43760 119910
rect 43840 119890 43900 119920
rect 43840 119770 43900 119800
rect 36000 119680 37190 119710
rect 37600 119700 37660 119730
rect 37720 119700 37780 119730
rect 37840 119700 37900 119730
rect 40685 119690 40715 119750
rect 40775 119690 40865 119750
rect 40895 119690 40925 119750
rect 36040 119670 36120 119680
rect 36220 119670 36300 119680
rect 36400 119670 36480 119680
rect 36580 119670 36660 119680
rect 36760 119670 36840 119680
rect 36940 119670 37020 119680
rect 36120 119610 36130 119670
rect 36300 119610 36310 119670
rect 36480 119610 36490 119670
rect 36660 119610 36670 119670
rect 36840 119610 36850 119670
rect 37020 119610 37030 119670
rect 37100 119610 37190 119680
rect 38595 119675 38675 119685
rect 38775 119675 38855 119685
rect 38955 119675 39035 119685
rect 39135 119675 39215 119685
rect 39315 119675 39395 119685
rect 37720 119610 37750 119640
rect 37840 119610 37870 119640
rect 36000 119580 37190 119610
rect 37600 119580 37660 119610
rect 37720 119580 37780 119610
rect 37840 119580 37900 119610
rect 38675 119595 38685 119675
rect 38855 119595 38865 119675
rect 39035 119595 39045 119675
rect 39215 119595 39225 119675
rect 39395 119595 39405 119675
rect 40060 119650 40120 119680
rect 40685 119660 40925 119690
rect 41540 119650 41600 119680
rect 42360 119650 42420 119680
rect 40678 119629 40758 119639
rect 40838 119629 40918 119639
rect 36040 119520 36120 119530
rect 36220 119520 36300 119530
rect 36400 119520 36480 119530
rect 36580 119520 36660 119530
rect 36760 119520 36840 119530
rect 36940 119520 37020 119530
rect 36120 119440 36130 119520
rect 36300 119440 36310 119520
rect 36480 119440 36490 119520
rect 36660 119440 36670 119520
rect 36840 119440 36850 119520
rect 37020 119440 37030 119520
rect 37100 119380 37190 119580
rect 40060 119530 40120 119560
rect 40758 119549 40768 119629
rect 40838 119549 40848 119629
rect 40918 119549 40928 119629
rect 42822 119620 42892 119760
rect 43580 119650 43700 119710
rect 43840 119650 43900 119680
rect 42950 119630 43560 119640
rect 43550 119625 43560 119630
rect 42682 119560 42822 119620
rect 42910 119615 43560 119625
rect 42900 119565 42910 119615
rect 41540 119530 41600 119560
rect 42360 119530 42420 119560
rect 37720 119490 37750 119520
rect 37840 119490 37870 119520
rect 38595 119495 38675 119505
rect 38775 119495 38855 119505
rect 38955 119495 39035 119505
rect 39135 119495 39215 119505
rect 39315 119495 39395 119505
rect 37600 119460 37660 119490
rect 37720 119460 37780 119490
rect 37840 119460 37900 119490
rect 38675 119415 38685 119495
rect 38855 119415 38865 119495
rect 39035 119415 39045 119495
rect 39215 119415 39225 119495
rect 39395 119415 39405 119495
rect 40060 119410 40120 119440
rect 41540 119410 41600 119440
rect 42360 119410 42420 119440
rect 42822 119420 42892 119560
rect 43030 119520 43390 119580
rect 36000 119350 37190 119380
rect 37720 119370 37750 119400
rect 37840 119370 37870 119400
rect 36120 119290 36130 119350
rect 36300 119290 36310 119350
rect 36480 119290 36490 119350
rect 36660 119290 36670 119350
rect 36840 119290 36850 119350
rect 37020 119290 37030 119350
rect 37100 119280 37190 119350
rect 37600 119340 37660 119370
rect 37720 119340 37780 119370
rect 37840 119340 37900 119370
rect 40170 119320 40180 119410
rect 40060 119290 40120 119320
rect 36000 119250 37190 119280
rect 37720 119250 37750 119280
rect 37840 119250 37870 119280
rect 37100 119240 37190 119250
rect 36000 119230 37190 119240
rect 36040 119050 36120 119060
rect 36220 119050 36300 119060
rect 36400 119050 36480 119060
rect 36580 119050 36660 119060
rect 36760 119050 36840 119060
rect 36940 119050 37020 119060
rect 36120 118970 36130 119050
rect 36300 118970 36310 119050
rect 36480 118970 36490 119050
rect 36660 118970 36670 119050
rect 36840 118970 36850 119050
rect 37020 118970 37030 119050
rect 36040 118730 36120 118740
rect 36220 118730 36300 118740
rect 36400 118730 36480 118740
rect 36580 118730 36660 118740
rect 36760 118730 36840 118740
rect 36940 118730 37020 118740
rect 36120 118650 36130 118730
rect 36300 118650 36310 118730
rect 36480 118650 36490 118730
rect 36660 118650 36670 118730
rect 36840 118650 36850 118730
rect 37020 118650 37030 118730
rect 37100 118560 37190 119230
rect 37600 119220 37660 119250
rect 37720 119220 37780 119250
rect 37840 119220 37900 119250
rect 40060 119170 40120 119200
rect 37720 119130 37750 119160
rect 37840 119130 37870 119160
rect 37600 119100 37660 119130
rect 37720 119100 37780 119130
rect 37840 119100 37900 119130
rect 40060 119050 40120 119080
rect 37720 119010 37750 119040
rect 37840 119010 37870 119040
rect 37600 118980 37660 119010
rect 37720 118980 37780 119010
rect 37840 118980 37900 119010
rect 40060 118930 40120 118960
rect 37720 118890 37750 118920
rect 37840 118890 37870 118920
rect 37600 118860 37660 118890
rect 37720 118860 37780 118890
rect 37840 118860 37900 118890
rect 40060 118810 40120 118840
rect 37720 118770 37750 118800
rect 37840 118770 37870 118800
rect 37600 118740 37660 118770
rect 37720 118740 37780 118770
rect 37840 118740 37900 118770
rect 40060 118690 40120 118720
rect 37720 118650 37750 118680
rect 37840 118650 37870 118680
rect 37600 118620 37660 118650
rect 37720 118620 37780 118650
rect 37840 118620 37900 118650
rect 40060 118570 40120 118600
rect 36000 118550 37190 118560
rect 37100 118450 37190 118550
rect 37720 118530 37750 118560
rect 37840 118530 37870 118560
rect 40260 118530 40270 119320
rect 40380 119310 41180 119400
rect 40650 119280 40770 119310
rect 40930 119280 41050 119310
rect 41090 119280 41180 119310
rect 40650 119190 40660 119280
rect 40760 119250 40830 119280
rect 40770 119160 40830 119250
rect 40930 119190 40940 119280
rect 41050 119160 41180 119280
rect 41260 119240 41340 119250
rect 41340 119190 41350 119240
rect 41090 119125 41180 119160
rect 41230 119130 41350 119190
rect 40470 119120 41180 119125
rect 40370 119110 41180 119120
rect 40370 119030 40380 119110
rect 40470 119105 41180 119110
rect 40420 119095 41210 119105
rect 41090 119045 41180 119095
rect 40470 119030 41180 119045
rect 40460 119015 41180 119030
rect 40460 118825 40470 119015
rect 40650 118980 40770 119015
rect 40930 118980 41050 119015
rect 41090 118980 41180 119015
rect 41350 119010 41410 119130
rect 40770 118970 40830 118980
rect 40530 118960 40610 118970
rect 40670 118960 40750 118970
rect 40770 118960 40890 118970
rect 40950 118960 41030 118970
rect 40610 118880 40620 118960
rect 40750 118880 40760 118960
rect 40770 118860 40830 118960
rect 40890 118880 40900 118960
rect 41030 118880 41040 118960
rect 41050 118860 41180 118980
rect 41260 118960 41340 118970
rect 41340 118890 41350 118960
rect 41090 118825 41180 118860
rect 41230 118830 41350 118890
rect 40460 118810 41180 118825
rect 40470 118805 41180 118810
rect 40420 118795 41210 118805
rect 41090 118745 41180 118795
rect 40470 118715 41180 118745
rect 40650 118680 40770 118715
rect 40930 118680 41050 118715
rect 41090 118680 41180 118715
rect 41350 118710 41410 118830
rect 41480 118680 41490 119390
rect 42860 119370 43470 119380
rect 43550 119370 43560 119615
rect 43700 119530 43760 119650
rect 43840 119530 43900 119560
rect 43580 119390 43700 119450
rect 43840 119410 43900 119440
rect 42910 119355 43560 119365
rect 41540 119290 41600 119320
rect 42360 119290 42420 119320
rect 42900 119305 42910 119355
rect 43030 119260 43390 119320
rect 43700 119270 43760 119390
rect 43840 119290 43900 119320
rect 41540 119170 41600 119200
rect 42360 119170 42420 119200
rect 42470 119160 42480 119250
rect 43840 119170 43900 119200
rect 41540 119050 41600 119080
rect 42360 119050 42420 119080
rect 41540 118930 41600 118960
rect 42360 118930 42420 118960
rect 41540 118810 41600 118840
rect 42360 118810 42420 118840
rect 41540 118690 41600 118720
rect 42360 118690 42420 118720
rect 42560 118680 42570 119160
rect 42960 119120 43460 119130
rect 42620 119100 42700 119110
rect 42700 119030 42710 119100
rect 42620 119020 42710 119030
rect 42770 119020 42780 119110
rect 43840 119050 43900 119080
rect 42620 118940 42700 118950
rect 42700 118890 42710 118940
rect 42610 118830 42730 118890
rect 42730 118805 42790 118830
rect 42860 118820 42870 119020
rect 42910 118980 43030 119040
rect 43190 118980 43310 119040
rect 43030 118970 43090 118980
rect 43310 118970 43370 118980
rect 42930 118960 43010 118970
rect 43030 118960 43150 118970
rect 43210 118960 43290 118970
rect 43310 118960 43430 118970
rect 43010 118880 43020 118960
rect 43030 118860 43090 118960
rect 43150 118880 43160 118960
rect 43290 118880 43300 118960
rect 43310 118860 43370 118960
rect 43430 118880 43440 118960
rect 43840 118930 43900 118960
rect 42860 118810 43500 118820
rect 43840 118810 43900 118840
rect 42730 118795 43540 118805
rect 42730 118710 42790 118795
rect 43540 118745 43550 118795
rect 42860 118680 42870 118730
rect 42910 118680 43030 118740
rect 43190 118680 43310 118740
rect 43840 118690 43900 118720
rect 40770 118670 40830 118680
rect 40530 118660 40610 118670
rect 40770 118660 40890 118670
rect 40610 118580 40620 118660
rect 40770 118560 40830 118660
rect 40890 118580 40900 118660
rect 41050 118560 41180 118680
rect 43030 118670 43090 118680
rect 43310 118670 43370 118680
rect 43030 118660 43150 118670
rect 43310 118660 43430 118670
rect 41540 118570 41600 118600
rect 42360 118570 42420 118600
rect 43030 118560 43090 118660
rect 43150 118580 43160 118660
rect 43310 118560 43370 118660
rect 43430 118580 43440 118660
rect 43840 118570 43900 118600
rect 41090 118550 41180 118560
rect 40470 118530 41180 118550
rect 37600 118500 37660 118530
rect 37720 118500 37780 118530
rect 37840 118500 37900 118530
rect 40060 118450 40120 118480
rect 36000 118420 37190 118450
rect 40170 118440 40180 118530
rect 40260 118520 41100 118530
rect 36040 118410 36120 118420
rect 36220 118410 36300 118420
rect 36400 118410 36480 118420
rect 36580 118410 36660 118420
rect 36760 118410 36840 118420
rect 36940 118410 37020 118420
rect 36120 118350 36130 118410
rect 36300 118350 36310 118410
rect 36480 118350 36490 118410
rect 36660 118350 36670 118410
rect 36840 118350 36850 118410
rect 37020 118350 37030 118410
rect 37100 118350 37190 118420
rect 37720 118410 37750 118440
rect 37840 118410 37870 118440
rect 37600 118380 37660 118410
rect 37720 118380 37780 118410
rect 37840 118380 37900 118410
rect 36000 118320 37190 118350
rect 40060 118330 40120 118360
rect 36040 118260 36120 118270
rect 36220 118260 36300 118270
rect 36400 118260 36480 118270
rect 36580 118260 36660 118270
rect 36760 118260 36840 118270
rect 36940 118260 37020 118270
rect 36120 118180 36130 118260
rect 36300 118180 36310 118260
rect 36480 118180 36490 118260
rect 36660 118180 36670 118260
rect 36840 118180 36850 118260
rect 37020 118180 37030 118260
rect 37100 118120 37190 118320
rect 37720 118290 37750 118320
rect 37840 118290 37870 118320
rect 37600 118260 37660 118290
rect 37720 118260 37780 118290
rect 37840 118260 37900 118290
rect 40060 118210 40120 118240
rect 37720 118170 37750 118200
rect 37840 118170 37870 118200
rect 37600 118140 37660 118170
rect 37720 118140 37780 118170
rect 37840 118140 37900 118170
rect 36000 118090 37190 118120
rect 40060 118090 40120 118120
rect 36120 118030 36130 118090
rect 36300 118030 36310 118090
rect 36480 118030 36490 118090
rect 36660 118030 36670 118090
rect 36840 118030 36850 118090
rect 37020 118030 37030 118090
rect 37100 118020 37190 118090
rect 37720 118050 37750 118080
rect 37840 118050 37870 118080
rect 37600 118020 37660 118050
rect 37720 118020 37780 118050
rect 37840 118020 37900 118050
rect 36000 117990 37190 118020
rect 37100 117980 37190 117990
rect 36000 117970 37190 117980
rect 40060 117970 40120 118000
rect 36040 117790 36120 117800
rect 36220 117790 36300 117800
rect 36400 117790 36480 117800
rect 36580 117790 36660 117800
rect 36760 117790 36840 117800
rect 36940 117790 37020 117800
rect 36120 117710 36130 117790
rect 36300 117710 36310 117790
rect 36480 117710 36490 117790
rect 36660 117710 36670 117790
rect 36840 117710 36850 117790
rect 37020 117710 37030 117790
rect 36040 117470 36120 117480
rect 36220 117470 36300 117480
rect 36400 117470 36480 117480
rect 36580 117470 36660 117480
rect 36760 117470 36840 117480
rect 36940 117470 37020 117480
rect 36120 117390 36130 117470
rect 36300 117390 36310 117470
rect 36480 117390 36490 117470
rect 36660 117390 36670 117470
rect 36840 117390 36850 117470
rect 37020 117390 37030 117470
rect 37100 117300 37190 117970
rect 37720 117930 37750 117960
rect 37840 117930 37870 117960
rect 37600 117900 37660 117930
rect 37720 117900 37780 117930
rect 37840 117900 37900 117930
rect 40060 117850 40120 117880
rect 37720 117810 37750 117840
rect 37840 117810 37870 117840
rect 37600 117780 37660 117810
rect 37720 117780 37780 117810
rect 37840 117780 37900 117810
rect 40060 117730 40120 117760
rect 37720 117690 37750 117720
rect 37840 117690 37870 117720
rect 37600 117660 37660 117690
rect 37720 117660 37780 117690
rect 37840 117660 37900 117690
rect 40060 117610 40120 117640
rect 37720 117570 37750 117600
rect 37840 117570 37870 117600
rect 37600 117540 37660 117570
rect 37720 117540 37780 117570
rect 37840 117540 37900 117570
rect 40060 117490 40120 117520
rect 37720 117450 37750 117480
rect 37840 117450 37870 117480
rect 37600 117420 37660 117450
rect 37720 117420 37780 117450
rect 37840 117420 37900 117450
rect 40060 117370 40120 117400
rect 37720 117330 37750 117360
rect 37840 117330 37870 117360
rect 37600 117300 37660 117330
rect 37720 117300 37780 117330
rect 37840 117300 37900 117330
rect 36000 117290 37190 117300
rect 37100 117190 37190 117290
rect 40060 117250 40120 117280
rect 37720 117210 37750 117240
rect 37840 117210 37870 117240
rect 36000 117160 37190 117190
rect 37600 117180 37660 117210
rect 37720 117180 37780 117210
rect 37840 117180 37900 117210
rect 36040 117150 36120 117160
rect 36220 117150 36300 117160
rect 36400 117150 36480 117160
rect 36580 117150 36660 117160
rect 36760 117150 36840 117160
rect 36940 117150 37020 117160
rect 36120 117090 36130 117150
rect 36300 117090 36310 117150
rect 36480 117090 36490 117150
rect 36660 117090 36670 117150
rect 36840 117090 36850 117150
rect 37020 117090 37030 117150
rect 37100 117090 37190 117160
rect 40060 117130 40120 117160
rect 37720 117090 37750 117120
rect 37840 117090 37870 117120
rect 36000 117060 37190 117090
rect 37600 117060 37660 117090
rect 37720 117060 37780 117090
rect 37840 117060 37900 117090
rect 36040 117000 36120 117010
rect 36220 117000 36300 117010
rect 36400 117000 36480 117010
rect 36580 117000 36660 117010
rect 36760 117000 36840 117010
rect 36940 117000 37020 117010
rect 36120 116920 36130 117000
rect 36300 116920 36310 117000
rect 36480 116920 36490 117000
rect 36660 116920 36670 117000
rect 36840 116920 36850 117000
rect 37020 116920 37030 117000
rect 36040 116850 36120 116860
rect 36220 116850 36300 116860
rect 36400 116850 36480 116860
rect 36580 116850 36660 116860
rect 36760 116850 36840 116860
rect 36940 116850 37020 116860
rect 36120 116770 36130 116850
rect 36300 116770 36310 116850
rect 36480 116770 36490 116850
rect 36660 116770 36670 116850
rect 36840 116770 36850 116850
rect 37020 116770 37030 116850
rect 37100 116830 37190 117060
rect 40060 117010 40120 117040
rect 37720 116970 37750 117000
rect 37840 116970 37870 117000
rect 37600 116940 37660 116970
rect 37720 116940 37780 116970
rect 37840 116940 37900 116970
rect 40060 116890 40120 116920
rect 37720 116850 37750 116880
rect 37840 116850 37870 116880
rect 37600 116820 37660 116850
rect 37720 116820 37780 116850
rect 37840 116820 37900 116850
rect 40060 116770 40120 116800
rect 19130 116700 19160 116755
rect 19250 116700 19280 116755
rect 26420 116700 26450 116755
rect 26540 116700 26570 116755
rect 30420 116730 30450 116755
rect 30540 116730 30570 116755
rect 37720 116730 37750 116760
rect 37840 116730 37870 116760
rect 30300 116700 30360 116730
rect 30420 116700 30480 116730
rect 30540 116700 30600 116730
rect 37600 116700 37660 116730
rect 37720 116700 37780 116730
rect 37840 116700 37900 116730
rect 40060 116650 40120 116680
rect 30420 116580 30450 116640
rect 30540 116580 30570 116640
rect 37720 116580 37750 116640
rect 37840 116580 37870 116640
rect 40060 116530 40120 116560
rect 18980 116440 19060 116450
rect 19160 116440 19240 116450
rect 19340 116440 19420 116450
rect 19520 116440 19600 116450
rect 19700 116440 19780 116450
rect 19880 116440 19960 116450
rect 20060 116440 20140 116450
rect 20240 116440 20320 116450
rect 20420 116440 20500 116450
rect 20600 116440 20680 116450
rect 20780 116440 20860 116450
rect 20960 116440 21040 116450
rect 21140 116440 21220 116450
rect 21320 116440 21400 116450
rect 21500 116440 21580 116450
rect 21680 116440 21760 116450
rect 21860 116440 21940 116450
rect 22040 116440 22120 116450
rect 22220 116440 22300 116450
rect 22400 116440 22480 116450
rect 22580 116440 22660 116450
rect 22760 116440 22840 116450
rect 22940 116440 23020 116450
rect 23120 116440 23200 116450
rect 23300 116440 23380 116450
rect 23480 116440 23560 116450
rect 23660 116440 23740 116450
rect 23840 116440 23920 116450
rect 24020 116440 24100 116450
rect 24200 116440 24280 116450
rect 24380 116440 24460 116450
rect 24560 116440 24640 116450
rect 24740 116440 24820 116450
rect 24920 116440 25000 116450
rect 25100 116440 25180 116450
rect 25280 116440 25360 116450
rect 25460 116440 25540 116450
rect 25640 116440 25720 116450
rect 25820 116440 25900 116450
rect 26000 116440 26080 116450
rect 26180 116440 26260 116450
rect 26360 116440 26440 116450
rect 26540 116440 26620 116450
rect 30280 116440 30360 116450
rect 30460 116440 30540 116450
rect 30640 116440 30720 116450
rect 30820 116440 30900 116450
rect 31000 116440 31080 116450
rect 31180 116440 31260 116450
rect 31360 116440 31440 116450
rect 31540 116440 31620 116450
rect 31720 116440 31800 116450
rect 31900 116440 31980 116450
rect 32080 116440 32160 116450
rect 32260 116440 32340 116450
rect 32440 116440 32520 116450
rect 32620 116440 32700 116450
rect 32800 116440 32880 116450
rect 32980 116440 33060 116450
rect 33160 116440 33240 116450
rect 33340 116440 33420 116450
rect 33520 116440 33600 116450
rect 33700 116440 33780 116450
rect 33880 116440 33960 116450
rect 34060 116440 34140 116450
rect 34240 116440 34320 116450
rect 34420 116440 34500 116450
rect 34600 116440 34680 116450
rect 34780 116440 34860 116450
rect 34960 116440 35040 116450
rect 35140 116440 35220 116450
rect 35320 116440 35400 116450
rect 35500 116440 35580 116450
rect 35680 116440 35760 116450
rect 35860 116440 35940 116450
rect 36040 116440 36120 116450
rect 36220 116440 36300 116450
rect 36400 116440 36480 116450
rect 36580 116440 36660 116450
rect 36760 116440 36840 116450
rect 36940 116440 37020 116450
rect 37120 116440 37200 116450
rect 37300 116440 37380 116450
rect 37480 116440 37560 116450
rect 37660 116440 37740 116450
rect 37840 116440 37920 116450
rect 40260 116440 40270 118440
rect 40380 118430 41180 118520
rect 41540 118450 41600 118480
rect 42360 118450 42420 118480
rect 43840 118450 43900 118480
rect 40650 118400 40770 118430
rect 40930 118400 41050 118430
rect 41090 118400 41180 118430
rect 40650 118310 40660 118400
rect 40760 118370 40830 118400
rect 40770 118280 40830 118370
rect 40930 118310 40940 118400
rect 41050 118280 41180 118400
rect 41090 118245 41180 118280
rect 41230 118250 41350 118310
rect 40470 118240 41180 118245
rect 40370 118230 41180 118240
rect 40370 118150 40380 118230
rect 40470 118225 41180 118230
rect 40420 118215 41210 118225
rect 41090 118165 41180 118215
rect 40470 118150 41180 118165
rect 40460 118135 41180 118150
rect 40460 117945 40470 118135
rect 40650 118100 40770 118135
rect 40930 118100 41050 118135
rect 41090 118100 41180 118135
rect 41350 118130 41410 118250
rect 40770 118090 40830 118100
rect 40530 118080 40610 118090
rect 40670 118080 40750 118090
rect 40770 118080 40890 118090
rect 40950 118080 41030 118090
rect 40610 118000 40620 118080
rect 40750 118000 40760 118080
rect 40770 117980 40830 118080
rect 40890 118000 40900 118080
rect 41030 118000 41040 118080
rect 41050 117980 41180 118100
rect 41260 118080 41340 118090
rect 41340 118010 41350 118080
rect 41090 117945 41180 117980
rect 41230 117950 41350 118010
rect 40460 117930 41180 117945
rect 40470 117925 41180 117930
rect 40420 117915 41210 117925
rect 41090 117865 41180 117915
rect 40470 117835 41180 117865
rect 40650 117800 40770 117835
rect 40930 117800 41050 117835
rect 41090 117800 41180 117835
rect 41350 117830 41410 117950
rect 40650 117710 40660 117800
rect 40760 117770 40830 117800
rect 40770 117680 40830 117770
rect 40930 117710 40940 117800
rect 41050 117680 41180 117800
rect 41260 117780 41340 117790
rect 41340 117710 41350 117780
rect 41090 117645 41180 117680
rect 41230 117650 41350 117710
rect 40370 117630 40460 117640
rect 40370 117550 40380 117630
rect 40470 117625 41180 117645
rect 40420 117615 41210 117625
rect 41090 117565 41180 117615
rect 40470 117550 41180 117565
rect 40460 117535 41180 117550
rect 40460 117345 40470 117535
rect 40650 117500 40770 117535
rect 40930 117500 41050 117535
rect 41090 117500 41180 117535
rect 41350 117530 41410 117650
rect 40770 117490 40830 117500
rect 40530 117480 40610 117490
rect 40670 117480 40750 117490
rect 40770 117480 40890 117490
rect 40950 117480 41030 117490
rect 40610 117400 40620 117480
rect 40750 117400 40760 117480
rect 40770 117380 40830 117480
rect 40890 117400 40900 117480
rect 41030 117400 41040 117480
rect 41050 117380 41180 117500
rect 41260 117480 41340 117490
rect 41340 117410 41350 117480
rect 41090 117345 41180 117380
rect 41230 117350 41350 117410
rect 40460 117330 41180 117345
rect 40470 117325 41180 117330
rect 40420 117315 41210 117325
rect 41090 117265 41180 117315
rect 40470 117235 41180 117265
rect 40650 117200 40770 117235
rect 40930 117200 41050 117235
rect 41090 117200 41180 117235
rect 41350 117230 41410 117350
rect 40650 117110 40660 117200
rect 40760 117170 40830 117200
rect 40770 117080 40830 117170
rect 40930 117110 40940 117200
rect 41050 117080 41180 117200
rect 41260 117180 41340 117190
rect 41340 117110 41350 117180
rect 41090 117045 41180 117080
rect 41230 117050 41350 117110
rect 40370 117030 40460 117040
rect 40370 116950 40380 117030
rect 40470 117025 41180 117045
rect 40420 117015 41210 117025
rect 41090 116965 41180 117015
rect 40470 116950 41180 116965
rect 40460 116935 41180 116950
rect 40460 116745 40470 116935
rect 40650 116900 40770 116935
rect 40930 116900 41050 116935
rect 41090 116900 41180 116935
rect 41350 116930 41410 117050
rect 40770 116890 40830 116900
rect 40530 116880 40610 116890
rect 40670 116880 40750 116890
rect 40770 116880 40890 116890
rect 40950 116880 41030 116890
rect 40610 116800 40620 116880
rect 40750 116800 40760 116880
rect 40770 116780 40830 116880
rect 40890 116800 40900 116880
rect 41030 116800 41040 116880
rect 41050 116780 41180 116900
rect 41260 116870 41340 116880
rect 41340 116810 41350 116870
rect 41090 116745 41180 116780
rect 41230 116750 41350 116810
rect 40460 116730 41180 116745
rect 40470 116725 41180 116730
rect 40420 116715 41210 116725
rect 41090 116665 41180 116715
rect 40470 116635 41180 116665
rect 40650 116600 40770 116635
rect 40930 116600 41050 116635
rect 41090 116600 41180 116635
rect 41350 116630 41410 116750
rect 41480 116600 41490 118370
rect 41540 118330 41600 118360
rect 42360 118330 42420 118360
rect 43840 118330 43900 118360
rect 41540 118210 41600 118240
rect 42360 118210 42420 118240
rect 43840 118210 43900 118240
rect 41540 118090 41600 118120
rect 42360 118090 42420 118120
rect 42910 118100 43030 118160
rect 43190 118100 43310 118160
rect 43030 118090 43090 118100
rect 43310 118090 43370 118100
rect 43840 118090 43900 118120
rect 42930 118080 43010 118090
rect 43030 118080 43150 118090
rect 43210 118080 43290 118090
rect 43310 118080 43430 118090
rect 41540 117970 41600 118000
rect 42360 117970 42420 118000
rect 42470 117980 42480 118070
rect 41540 117850 41600 117880
rect 42360 117850 42420 117880
rect 41540 117730 41600 117760
rect 42360 117730 42420 117760
rect 41540 117610 41600 117640
rect 42360 117610 42420 117640
rect 41540 117490 41600 117520
rect 42360 117490 42420 117520
rect 41540 117370 41600 117400
rect 42360 117370 42420 117400
rect 41540 117250 41600 117280
rect 42360 117250 42420 117280
rect 41540 117130 41600 117160
rect 42360 117130 42420 117160
rect 41540 117010 41600 117040
rect 42360 117010 42420 117040
rect 41540 116890 41600 116920
rect 42360 116890 42420 116920
rect 41540 116770 41600 116800
rect 42360 116770 42420 116800
rect 41540 116650 41600 116680
rect 42360 116650 42420 116680
rect 42560 116620 42570 117980
rect 42610 117950 42730 118010
rect 42730 117925 42790 117950
rect 42860 117940 42870 118070
rect 43010 118000 43020 118080
rect 43030 117980 43090 118080
rect 43150 118000 43160 118080
rect 43290 118000 43300 118080
rect 43310 117980 43370 118080
rect 43430 118000 43440 118080
rect 43840 117970 43900 118000
rect 42860 117930 43500 117940
rect 42730 117915 43540 117925
rect 42730 117830 42790 117915
rect 43540 117865 43550 117915
rect 42620 117740 42700 117750
rect 42700 117660 42710 117740
rect 42860 117660 42870 117850
rect 42910 117800 43030 117860
rect 43190 117800 43310 117860
rect 43020 117770 43090 117800
rect 43030 117680 43090 117770
rect 43190 117710 43200 117800
rect 43300 117770 43370 117800
rect 43310 117680 43370 117770
rect 42860 117650 43490 117660
rect 42860 117640 42870 117650
rect 42620 117560 42700 117570
rect 42700 117480 42710 117560
rect 42770 117550 42780 117640
rect 42610 117360 42730 117420
rect 42730 117335 42790 117360
rect 42860 117350 42870 117550
rect 42910 117510 43030 117570
rect 43190 117510 43310 117570
rect 43030 117500 43090 117510
rect 43310 117500 43370 117510
rect 42930 117490 43010 117500
rect 43030 117490 43150 117500
rect 43210 117490 43290 117500
rect 43310 117490 43430 117500
rect 43010 117410 43020 117490
rect 43030 117390 43090 117490
rect 43150 117410 43160 117490
rect 43290 117410 43300 117490
rect 43310 117390 43370 117490
rect 43430 117410 43440 117490
rect 42860 117340 43500 117350
rect 43580 117340 43590 117640
rect 42730 117325 43540 117335
rect 42730 117240 42790 117325
rect 43540 117275 43550 117325
rect 42620 117140 42700 117150
rect 42700 117060 42710 117140
rect 42860 117070 42870 117260
rect 42910 117210 43030 117270
rect 43190 117210 43310 117270
rect 43020 117180 43090 117210
rect 43030 117090 43090 117180
rect 43190 117120 43200 117210
rect 43300 117180 43370 117210
rect 43310 117090 43370 117180
rect 42860 117060 43490 117070
rect 42860 117050 42870 117060
rect 42620 116960 42700 116970
rect 42770 116960 42780 117050
rect 42700 116880 42710 116960
rect 42610 116770 42730 116830
rect 42730 116745 42790 116770
rect 42860 116760 42870 116960
rect 42910 116920 43030 116980
rect 43190 116920 43310 116980
rect 43030 116910 43090 116920
rect 43310 116910 43370 116920
rect 42930 116900 43010 116910
rect 43030 116900 43150 116910
rect 43210 116900 43290 116910
rect 43310 116900 43430 116910
rect 43010 116820 43020 116900
rect 43030 116800 43090 116900
rect 43150 116820 43160 116900
rect 43290 116820 43300 116900
rect 43310 116800 43370 116900
rect 43430 116820 43440 116900
rect 42860 116750 43500 116760
rect 43580 116750 43590 117050
rect 42730 116735 43540 116745
rect 42730 116650 42790 116735
rect 43540 116685 43550 116735
rect 42860 116620 42870 116670
rect 42910 116620 43030 116680
rect 43190 116620 43310 116680
rect 43030 116610 43090 116620
rect 43310 116610 43370 116620
rect 43030 116600 43150 116610
rect 43310 116600 43430 116610
rect 40770 116590 40830 116600
rect 40530 116580 40610 116590
rect 40770 116580 40890 116590
rect 40610 116500 40620 116580
rect 40770 116480 40830 116580
rect 40890 116500 40900 116580
rect 41050 116480 41180 116600
rect 41540 116530 41600 116560
rect 42360 116530 42420 116560
rect 43030 116500 43090 116600
rect 43150 116520 43160 116600
rect 43310 116500 43370 116600
rect 43430 116520 43440 116600
rect 41090 116450 41180 116480
rect 43780 116460 43790 117940
rect 43840 117850 43900 117880
rect 43840 117730 43900 117760
rect 43840 117610 43900 117640
rect 43840 117490 43900 117520
rect 43840 117370 43900 117400
rect 146100 117330 146160 117360
rect 43840 117250 43900 117280
rect 146100 117210 146160 117240
rect 43840 117130 43900 117160
rect 146300 117150 146310 117420
rect 146690 117320 146810 117380
rect 146970 117320 147090 117380
rect 146690 117230 146700 117320
rect 146800 117290 146870 117320
rect 146810 117200 146870 117290
rect 146970 117230 146980 117320
rect 147090 117200 147150 117320
rect 146410 117150 147140 117160
rect 146460 117135 147150 117145
rect 146100 117090 146160 117120
rect 146450 117085 146460 117135
rect 43840 117010 43900 117040
rect 43840 116890 43900 116920
rect 146690 117020 146810 117080
rect 146970 117020 147090 117080
rect 146810 117010 146870 117020
rect 146570 117000 146650 117010
rect 146710 117000 146790 117010
rect 146810 117000 146930 117010
rect 146990 117000 147070 117010
rect 146100 116970 146160 117000
rect 146650 116920 146660 117000
rect 146790 116920 146800 117000
rect 146810 116900 146870 117000
rect 146930 116920 146940 117000
rect 147070 116920 147080 117000
rect 147090 116900 147150 117020
rect 146100 116850 146160 116880
rect 43840 116770 43900 116800
rect 146100 116730 146160 116760
rect 147580 116730 147640 116746
rect 148400 116730 148460 116746
rect 148600 116720 148610 116746
rect 148950 116720 149070 116746
rect 149230 116720 149350 116746
rect 149060 116690 149130 116720
rect 43840 116650 43900 116680
rect 146100 116610 146160 116640
rect 147580 116610 147640 116640
rect 148400 116610 148460 116640
rect 149070 116600 149130 116690
rect 149230 116630 149240 116720
rect 149340 116690 149410 116720
rect 149350 116600 149410 116690
rect 149530 116570 149620 116746
rect 149820 116560 149830 116746
rect 149880 116730 149940 116746
rect 152220 116710 152250 116740
rect 152340 116710 152370 116740
rect 159520 116710 159550 116740
rect 159640 116710 159670 116740
rect 163520 116710 163550 116740
rect 163640 116710 163670 116740
rect 163960 116735 164040 116745
rect 152100 116680 152160 116710
rect 152220 116680 152280 116710
rect 152340 116680 152400 116710
rect 159400 116680 159460 116710
rect 159520 116680 159580 116710
rect 159640 116680 159700 116710
rect 163400 116680 163460 116710
rect 163520 116680 163580 116710
rect 163640 116680 163700 116710
rect 164040 116655 164050 116735
rect 170810 116710 170840 116740
rect 170930 116710 170960 116740
rect 170690 116680 170750 116710
rect 170810 116680 170870 116710
rect 170930 116680 170990 116710
rect 149880 116610 149940 116640
rect 152220 116560 152250 116620
rect 152340 116560 152370 116620
rect 159520 116560 159550 116620
rect 159640 116560 159670 116620
rect 163520 116560 163550 116620
rect 163640 116560 163670 116620
rect 170810 116560 170840 116620
rect 170930 116560 170960 116620
rect 43840 116530 43900 116560
rect 146100 116490 146160 116520
rect 147580 116490 147640 116520
rect 148400 116490 148460 116520
rect 149880 116490 149940 116520
rect 19060 116360 19070 116440
rect 19240 116360 19250 116440
rect 19420 116360 19430 116440
rect 19600 116360 19610 116440
rect 19780 116360 19790 116440
rect 19960 116360 19970 116440
rect 20140 116360 20150 116440
rect 20320 116360 20330 116440
rect 20500 116360 20510 116440
rect 20680 116360 20690 116440
rect 20860 116360 20870 116440
rect 21040 116360 21050 116440
rect 21220 116360 21230 116440
rect 21400 116360 21410 116440
rect 21580 116360 21590 116440
rect 21760 116360 21770 116440
rect 21940 116360 21950 116440
rect 22120 116360 22130 116440
rect 22300 116360 22310 116440
rect 22480 116360 22490 116440
rect 22660 116360 22670 116440
rect 22840 116360 22850 116440
rect 23020 116360 23030 116440
rect 23200 116360 23210 116440
rect 23380 116360 23390 116440
rect 23560 116360 23570 116440
rect 23740 116360 23750 116440
rect 23920 116360 23930 116440
rect 24100 116360 24110 116440
rect 24280 116360 24290 116440
rect 24460 116360 24470 116440
rect 24640 116360 24650 116440
rect 24820 116360 24830 116440
rect 25000 116360 25010 116440
rect 25180 116360 25190 116440
rect 25360 116360 25370 116440
rect 25540 116360 25550 116440
rect 25720 116360 25730 116440
rect 25900 116360 25910 116440
rect 26080 116360 26090 116440
rect 26260 116360 26270 116440
rect 26440 116360 26450 116440
rect 26620 116360 26630 116440
rect 27315 116415 27395 116425
rect 27495 116415 27575 116425
rect 27675 116415 27755 116425
rect 27855 116415 27935 116425
rect 28035 116415 28115 116425
rect 27395 116335 27405 116415
rect 27575 116335 27585 116415
rect 27755 116335 27765 116415
rect 27935 116335 27945 116415
rect 28115 116335 28125 116415
rect 30360 116360 30370 116440
rect 30540 116360 30550 116440
rect 30720 116360 30730 116440
rect 30900 116360 30910 116440
rect 31080 116360 31090 116440
rect 31260 116360 31270 116440
rect 31440 116360 31450 116440
rect 31620 116360 31630 116440
rect 31800 116360 31810 116440
rect 31980 116360 31990 116440
rect 32160 116360 32170 116440
rect 32340 116360 32350 116440
rect 32520 116360 32530 116440
rect 32700 116360 32710 116440
rect 32880 116360 32890 116440
rect 33060 116360 33070 116440
rect 33240 116360 33250 116440
rect 33420 116360 33430 116440
rect 33600 116360 33610 116440
rect 33780 116360 33790 116440
rect 33960 116360 33970 116440
rect 34140 116360 34150 116440
rect 34320 116360 34330 116440
rect 34500 116360 34510 116440
rect 34680 116360 34690 116440
rect 34860 116360 34870 116440
rect 35040 116360 35050 116440
rect 35220 116360 35230 116440
rect 35400 116360 35410 116440
rect 35580 116360 35590 116440
rect 35760 116360 35770 116440
rect 35940 116360 35950 116440
rect 36120 116360 36130 116440
rect 36300 116360 36310 116440
rect 36480 116360 36490 116440
rect 36660 116360 36670 116440
rect 36840 116360 36850 116440
rect 37020 116360 37030 116440
rect 37200 116360 37210 116440
rect 37380 116360 37390 116440
rect 37560 116360 37570 116440
rect 37740 116360 37750 116440
rect 37920 116360 37930 116440
rect 40060 116410 40120 116440
rect 41540 116410 41600 116440
rect 42360 116410 42420 116440
rect 43840 116410 43900 116440
rect 146100 116370 146160 116400
rect 147580 116370 147640 116400
rect 148400 116370 148460 116400
rect 149880 116370 149940 116400
rect 18980 116290 19060 116300
rect 19160 116290 19240 116300
rect 19340 116290 19420 116300
rect 19520 116290 19600 116300
rect 19700 116290 19780 116300
rect 19880 116290 19960 116300
rect 20060 116290 20140 116300
rect 20240 116290 20320 116300
rect 20420 116290 20500 116300
rect 20600 116290 20680 116300
rect 20780 116290 20860 116300
rect 20960 116290 21040 116300
rect 21140 116290 21220 116300
rect 21320 116290 21400 116300
rect 21500 116290 21580 116300
rect 21680 116290 21760 116300
rect 21860 116290 21940 116300
rect 22040 116290 22120 116300
rect 22220 116290 22300 116300
rect 22400 116290 22480 116300
rect 22580 116290 22660 116300
rect 22760 116290 22840 116300
rect 22940 116290 23020 116300
rect 23120 116290 23200 116300
rect 23300 116290 23380 116300
rect 23480 116290 23560 116300
rect 23660 116290 23740 116300
rect 23840 116290 23920 116300
rect 24020 116290 24100 116300
rect 24200 116290 24280 116300
rect 24380 116290 24460 116300
rect 24560 116290 24640 116300
rect 24740 116290 24820 116300
rect 24920 116290 25000 116300
rect 25100 116290 25180 116300
rect 25280 116290 25360 116300
rect 25460 116290 25540 116300
rect 25640 116290 25720 116300
rect 25820 116290 25900 116300
rect 26000 116290 26080 116300
rect 26180 116290 26260 116300
rect 26360 116290 26440 116300
rect 26540 116290 26620 116300
rect 30280 116290 30360 116300
rect 30460 116290 30540 116300
rect 30640 116290 30720 116300
rect 30820 116290 30900 116300
rect 31000 116290 31080 116300
rect 31180 116290 31260 116300
rect 31360 116290 31440 116300
rect 31540 116290 31620 116300
rect 31720 116290 31800 116300
rect 31900 116290 31980 116300
rect 32080 116290 32160 116300
rect 32260 116290 32340 116300
rect 32440 116290 32520 116300
rect 32620 116290 32700 116300
rect 32800 116290 32880 116300
rect 32980 116290 33060 116300
rect 33160 116290 33240 116300
rect 33340 116290 33420 116300
rect 33520 116290 33600 116300
rect 33700 116290 33780 116300
rect 33880 116290 33960 116300
rect 34060 116290 34140 116300
rect 34240 116290 34320 116300
rect 34420 116290 34500 116300
rect 34600 116290 34680 116300
rect 34780 116290 34860 116300
rect 34960 116290 35040 116300
rect 35140 116290 35220 116300
rect 35320 116290 35400 116300
rect 35500 116290 35580 116300
rect 35680 116290 35760 116300
rect 35860 116290 35940 116300
rect 36040 116290 36120 116300
rect 36220 116290 36300 116300
rect 36400 116290 36480 116300
rect 36580 116290 36660 116300
rect 36760 116290 36840 116300
rect 36940 116290 37020 116300
rect 37120 116290 37200 116300
rect 37300 116290 37380 116300
rect 37480 116290 37560 116300
rect 37660 116290 37740 116300
rect 37840 116290 37920 116300
rect 152080 116290 152160 116300
rect 152260 116290 152340 116300
rect 152440 116290 152520 116300
rect 152620 116290 152700 116300
rect 152800 116290 152880 116300
rect 152980 116290 153060 116300
rect 153160 116290 153240 116300
rect 153340 116290 153420 116300
rect 153520 116290 153600 116300
rect 153700 116290 153780 116300
rect 153880 116290 153960 116300
rect 154060 116290 154140 116300
rect 154240 116290 154320 116300
rect 154420 116290 154500 116300
rect 154600 116290 154680 116300
rect 154780 116290 154860 116300
rect 154960 116290 155040 116300
rect 155140 116290 155220 116300
rect 155320 116290 155400 116300
rect 155500 116290 155580 116300
rect 155680 116290 155760 116300
rect 155860 116290 155940 116300
rect 156040 116290 156120 116300
rect 156220 116290 156300 116300
rect 156400 116290 156480 116300
rect 156580 116290 156660 116300
rect 156760 116290 156840 116300
rect 156940 116290 157020 116300
rect 157120 116290 157200 116300
rect 157300 116290 157380 116300
rect 157480 116290 157560 116300
rect 157660 116290 157740 116300
rect 157840 116290 157920 116300
rect 158020 116290 158100 116300
rect 158200 116290 158280 116300
rect 158380 116290 158460 116300
rect 158560 116290 158640 116300
rect 158740 116290 158820 116300
rect 158920 116290 159000 116300
rect 159100 116290 159180 116300
rect 159280 116290 159360 116300
rect 159460 116290 159540 116300
rect 159640 116290 159720 116300
rect 163380 116290 163460 116300
rect 163560 116290 163640 116300
rect 163740 116290 163820 116300
rect 163920 116290 164000 116300
rect 164100 116290 164180 116300
rect 164280 116290 164360 116300
rect 164460 116290 164540 116300
rect 164640 116290 164720 116300
rect 164820 116290 164900 116300
rect 165000 116290 165080 116300
rect 165180 116290 165260 116300
rect 165360 116290 165440 116300
rect 165540 116290 165620 116300
rect 165720 116290 165800 116300
rect 165900 116290 165980 116300
rect 166080 116290 166160 116300
rect 166260 116290 166340 116300
rect 166440 116290 166520 116300
rect 166620 116290 166700 116300
rect 166800 116290 166880 116300
rect 166980 116290 167060 116300
rect 167160 116290 167240 116300
rect 167340 116290 167420 116300
rect 167520 116290 167600 116300
rect 167700 116290 167780 116300
rect 167880 116290 167960 116300
rect 168060 116290 168140 116300
rect 168240 116290 168320 116300
rect 168420 116290 168500 116300
rect 168600 116290 168680 116300
rect 168780 116290 168860 116300
rect 168960 116290 169040 116300
rect 169140 116290 169220 116300
rect 169320 116290 169400 116300
rect 169500 116290 169580 116300
rect 169680 116290 169760 116300
rect 169860 116290 169940 116300
rect 170040 116290 170120 116300
rect 170220 116290 170300 116300
rect 170400 116290 170480 116300
rect 170580 116290 170660 116300
rect 170760 116290 170840 116300
rect 170940 116290 171020 116300
rect 19060 116210 19070 116290
rect 19240 116210 19250 116290
rect 19420 116210 19430 116290
rect 19600 116210 19610 116290
rect 19780 116210 19790 116290
rect 19960 116210 19970 116290
rect 20140 116210 20150 116290
rect 20320 116210 20330 116290
rect 20500 116210 20510 116290
rect 20680 116210 20690 116290
rect 20860 116210 20870 116290
rect 21040 116210 21050 116290
rect 21220 116210 21230 116290
rect 21400 116210 21410 116290
rect 21580 116210 21590 116290
rect 21760 116210 21770 116290
rect 21940 116210 21950 116290
rect 22120 116210 22130 116290
rect 22300 116210 22310 116290
rect 22480 116210 22490 116290
rect 22660 116210 22670 116290
rect 22840 116210 22850 116290
rect 23020 116210 23030 116290
rect 23200 116210 23210 116290
rect 23380 116210 23390 116290
rect 23560 116210 23570 116290
rect 23740 116210 23750 116290
rect 23920 116210 23930 116290
rect 24100 116210 24110 116290
rect 24280 116210 24290 116290
rect 24460 116210 24470 116290
rect 24640 116210 24650 116290
rect 24820 116210 24830 116290
rect 25000 116210 25010 116290
rect 25180 116210 25190 116290
rect 25360 116210 25370 116290
rect 25540 116210 25550 116290
rect 25720 116210 25730 116290
rect 25900 116210 25910 116290
rect 26080 116210 26090 116290
rect 26260 116210 26270 116290
rect 26440 116210 26450 116290
rect 26620 116210 26630 116290
rect 27315 116235 27395 116245
rect 27495 116235 27575 116245
rect 27675 116235 27755 116245
rect 27855 116235 27935 116245
rect 28035 116235 28115 116245
rect 27395 116155 27405 116235
rect 27575 116155 27585 116235
rect 27755 116155 27765 116235
rect 27935 116155 27945 116235
rect 28115 116155 28125 116235
rect 30360 116210 30370 116290
rect 30540 116210 30550 116290
rect 30720 116210 30730 116290
rect 30900 116210 30910 116290
rect 31080 116210 31090 116290
rect 31260 116210 31270 116290
rect 31440 116210 31450 116290
rect 31620 116210 31630 116290
rect 31800 116210 31810 116290
rect 31980 116210 31990 116290
rect 32160 116210 32170 116290
rect 32340 116210 32350 116290
rect 32520 116210 32530 116290
rect 32700 116210 32710 116290
rect 32880 116210 32890 116290
rect 33060 116210 33070 116290
rect 33240 116210 33250 116290
rect 33420 116210 33430 116290
rect 33600 116210 33610 116290
rect 33780 116210 33790 116290
rect 33960 116210 33970 116290
rect 34140 116210 34150 116290
rect 34320 116210 34330 116290
rect 34500 116210 34510 116290
rect 34680 116210 34690 116290
rect 34860 116210 34870 116290
rect 35040 116210 35050 116290
rect 35220 116210 35230 116290
rect 35400 116210 35410 116290
rect 35580 116210 35590 116290
rect 35760 116210 35770 116290
rect 35940 116210 35950 116290
rect 36120 116210 36130 116290
rect 36300 116210 36310 116290
rect 36480 116210 36490 116290
rect 36660 116210 36670 116290
rect 36840 116210 36850 116290
rect 37020 116210 37030 116290
rect 37200 116210 37210 116290
rect 37380 116210 37390 116290
rect 37560 116210 37570 116290
rect 37740 116210 37750 116290
rect 37920 116210 37930 116290
rect 152160 116210 152170 116290
rect 152340 116210 152350 116290
rect 152520 116210 152530 116290
rect 152700 116210 152710 116290
rect 152880 116210 152890 116290
rect 153060 116210 153070 116290
rect 153240 116210 153250 116290
rect 153420 116210 153430 116290
rect 153600 116210 153610 116290
rect 153780 116210 153790 116290
rect 153960 116210 153970 116290
rect 154140 116210 154150 116290
rect 154320 116210 154330 116290
rect 154500 116210 154510 116290
rect 154680 116210 154690 116290
rect 154860 116210 154870 116290
rect 155040 116210 155050 116290
rect 155220 116210 155230 116290
rect 155400 116210 155410 116290
rect 155580 116210 155590 116290
rect 155760 116210 155770 116290
rect 155940 116210 155950 116290
rect 156120 116210 156130 116290
rect 156300 116210 156310 116290
rect 156480 116210 156490 116290
rect 156660 116210 156670 116290
rect 156840 116210 156850 116290
rect 157020 116210 157030 116290
rect 157200 116210 157210 116290
rect 157380 116210 157390 116290
rect 157560 116210 157570 116290
rect 157740 116210 157750 116290
rect 157920 116210 157930 116290
rect 158100 116210 158110 116290
rect 158280 116210 158290 116290
rect 158460 116210 158470 116290
rect 158640 116210 158650 116290
rect 158820 116210 158830 116290
rect 159000 116210 159010 116290
rect 159180 116210 159190 116290
rect 159360 116210 159370 116290
rect 159540 116210 159550 116290
rect 159720 116210 159730 116290
rect 160430 116265 160510 116275
rect 160590 116265 160670 116275
rect 160750 116265 160830 116275
rect 160910 116265 160990 116275
rect 161070 116265 161150 116275
rect 160510 116185 160520 116265
rect 160590 116185 160600 116265
rect 160670 116185 160680 116265
rect 160750 116185 160760 116265
rect 160830 116185 160840 116265
rect 160910 116185 160920 116265
rect 160990 116185 161000 116265
rect 161070 116185 161080 116265
rect 161150 116185 161160 116265
rect 163460 116210 163470 116290
rect 163640 116210 163650 116290
rect 163820 116210 163830 116290
rect 164000 116210 164010 116290
rect 164180 116210 164190 116290
rect 164360 116210 164370 116290
rect 164540 116210 164550 116290
rect 164720 116210 164730 116290
rect 164900 116210 164910 116290
rect 165080 116210 165090 116290
rect 165260 116210 165270 116290
rect 165440 116210 165450 116290
rect 165620 116210 165630 116290
rect 165800 116210 165810 116290
rect 165980 116210 165990 116290
rect 166160 116210 166170 116290
rect 166340 116210 166350 116290
rect 166520 116210 166530 116290
rect 166700 116210 166710 116290
rect 166880 116210 166890 116290
rect 167060 116210 167070 116290
rect 167240 116210 167250 116290
rect 167420 116210 167430 116290
rect 167600 116210 167610 116290
rect 167780 116210 167790 116290
rect 167960 116210 167970 116290
rect 168140 116210 168150 116290
rect 168320 116210 168330 116290
rect 168500 116210 168510 116290
rect 168680 116210 168690 116290
rect 168860 116210 168870 116290
rect 169040 116210 169050 116290
rect 169220 116210 169230 116290
rect 169400 116210 169410 116290
rect 169580 116210 169590 116290
rect 169760 116210 169770 116290
rect 169940 116210 169950 116290
rect 170120 116210 170130 116290
rect 170300 116210 170310 116290
rect 170480 116210 170490 116290
rect 170660 116210 170670 116290
rect 170840 116210 170850 116290
rect 171020 116210 171030 116290
rect 18980 116140 19060 116150
rect 19160 116140 19240 116150
rect 19340 116140 19420 116150
rect 19520 116140 19600 116150
rect 19700 116140 19780 116150
rect 19880 116140 19960 116150
rect 20060 116140 20140 116150
rect 20240 116140 20320 116150
rect 20420 116140 20500 116150
rect 20600 116140 20680 116150
rect 20780 116140 20860 116150
rect 20960 116140 21040 116150
rect 21140 116140 21220 116150
rect 21320 116140 21400 116150
rect 21500 116140 21580 116150
rect 21680 116140 21760 116150
rect 21860 116140 21940 116150
rect 22040 116140 22120 116150
rect 22220 116140 22300 116150
rect 22400 116140 22480 116150
rect 22580 116140 22660 116150
rect 22760 116140 22840 116150
rect 22940 116140 23020 116150
rect 23120 116140 23200 116150
rect 23300 116140 23380 116150
rect 23480 116140 23560 116150
rect 23660 116140 23740 116150
rect 23840 116140 23920 116150
rect 24020 116140 24100 116150
rect 24200 116140 24280 116150
rect 24380 116140 24460 116150
rect 24560 116140 24640 116150
rect 24740 116140 24820 116150
rect 24920 116140 25000 116150
rect 25100 116140 25180 116150
rect 25280 116140 25360 116150
rect 25460 116140 25540 116150
rect 25640 116140 25720 116150
rect 25820 116140 25900 116150
rect 26000 116140 26080 116150
rect 26180 116140 26260 116150
rect 26360 116140 26440 116150
rect 26540 116140 26620 116150
rect 30280 116140 30360 116150
rect 30460 116140 30540 116150
rect 30640 116140 30720 116150
rect 30820 116140 30900 116150
rect 31000 116140 31080 116150
rect 31180 116140 31260 116150
rect 31360 116140 31440 116150
rect 31540 116140 31620 116150
rect 31720 116140 31800 116150
rect 31900 116140 31980 116150
rect 32080 116140 32160 116150
rect 32260 116140 32340 116150
rect 32440 116140 32520 116150
rect 32620 116140 32700 116150
rect 32800 116140 32880 116150
rect 32980 116140 33060 116150
rect 33160 116140 33240 116150
rect 33340 116140 33420 116150
rect 33520 116140 33600 116150
rect 33700 116140 33780 116150
rect 33880 116140 33960 116150
rect 34060 116140 34140 116150
rect 34240 116140 34320 116150
rect 34420 116140 34500 116150
rect 34600 116140 34680 116150
rect 34780 116140 34860 116150
rect 34960 116140 35040 116150
rect 35140 116140 35220 116150
rect 35320 116140 35400 116150
rect 35500 116140 35580 116150
rect 35680 116140 35760 116150
rect 35860 116140 35940 116150
rect 36040 116140 36120 116150
rect 36220 116140 36300 116150
rect 36400 116140 36480 116150
rect 36580 116140 36660 116150
rect 36760 116140 36840 116150
rect 36940 116140 37020 116150
rect 37120 116140 37200 116150
rect 37300 116140 37380 116150
rect 37480 116140 37560 116150
rect 37660 116140 37740 116150
rect 37840 116140 37920 116150
rect 40060 116140 40140 116150
rect 40200 116140 40280 116150
rect 40340 116140 40420 116150
rect 40480 116140 40560 116150
rect 40620 116140 40700 116150
rect 40760 116140 40840 116150
rect 40900 116140 40980 116150
rect 41040 116140 41120 116150
rect 41180 116140 41260 116150
rect 41320 116140 41400 116150
rect 42360 116140 42440 116150
rect 42500 116140 42580 116150
rect 42640 116140 42720 116150
rect 42780 116140 42860 116150
rect 42920 116140 43000 116150
rect 43060 116140 43140 116150
rect 43200 116140 43280 116150
rect 43340 116140 43420 116150
rect 43480 116140 43560 116150
rect 43620 116140 43700 116150
rect 146300 116140 146380 116150
rect 146440 116140 146520 116150
rect 146580 116140 146660 116150
rect 146720 116140 146800 116150
rect 146860 116140 146940 116150
rect 147000 116140 147080 116150
rect 147140 116140 147220 116150
rect 147280 116140 147360 116150
rect 147420 116140 147500 116150
rect 147560 116140 147640 116150
rect 148600 116140 148680 116150
rect 148740 116140 148820 116150
rect 148880 116140 148960 116150
rect 149020 116140 149100 116150
rect 149160 116140 149240 116150
rect 149300 116140 149380 116150
rect 149440 116140 149520 116150
rect 149580 116140 149660 116150
rect 149720 116140 149800 116150
rect 149860 116140 149940 116150
rect 152080 116140 152160 116150
rect 152260 116140 152340 116150
rect 152440 116140 152520 116150
rect 152620 116140 152700 116150
rect 152800 116140 152880 116150
rect 152980 116140 153060 116150
rect 153160 116140 153240 116150
rect 153340 116140 153420 116150
rect 153520 116140 153600 116150
rect 153700 116140 153780 116150
rect 153880 116140 153960 116150
rect 154060 116140 154140 116150
rect 154240 116140 154320 116150
rect 154420 116140 154500 116150
rect 154600 116140 154680 116150
rect 154780 116140 154860 116150
rect 154960 116140 155040 116150
rect 155140 116140 155220 116150
rect 155320 116140 155400 116150
rect 155500 116140 155580 116150
rect 155680 116140 155760 116150
rect 155860 116140 155940 116150
rect 156040 116140 156120 116150
rect 156220 116140 156300 116150
rect 156400 116140 156480 116150
rect 156580 116140 156660 116150
rect 156760 116140 156840 116150
rect 156940 116140 157020 116150
rect 157120 116140 157200 116150
rect 157300 116140 157380 116150
rect 157480 116140 157560 116150
rect 157660 116140 157740 116150
rect 157840 116140 157920 116150
rect 158020 116140 158100 116150
rect 158200 116140 158280 116150
rect 158380 116140 158460 116150
rect 158560 116140 158640 116150
rect 158740 116140 158820 116150
rect 158920 116140 159000 116150
rect 159100 116140 159180 116150
rect 159280 116140 159360 116150
rect 159460 116140 159540 116150
rect 159640 116140 159720 116150
rect 163380 116140 163460 116150
rect 163560 116140 163640 116150
rect 163740 116140 163820 116150
rect 163920 116140 164000 116150
rect 164100 116140 164180 116150
rect 164280 116140 164360 116150
rect 164460 116140 164540 116150
rect 164640 116140 164720 116150
rect 164820 116140 164900 116150
rect 165000 116140 165080 116150
rect 165180 116140 165260 116150
rect 165360 116140 165440 116150
rect 165540 116140 165620 116150
rect 165720 116140 165800 116150
rect 165900 116140 165980 116150
rect 166080 116140 166160 116150
rect 166260 116140 166340 116150
rect 166440 116140 166520 116150
rect 166620 116140 166700 116150
rect 166800 116140 166880 116150
rect 166980 116140 167060 116150
rect 167160 116140 167240 116150
rect 167340 116140 167420 116150
rect 167520 116140 167600 116150
rect 167700 116140 167780 116150
rect 167880 116140 167960 116150
rect 168060 116140 168140 116150
rect 168240 116140 168320 116150
rect 168420 116140 168500 116150
rect 168600 116140 168680 116150
rect 168780 116140 168860 116150
rect 168960 116140 169040 116150
rect 169140 116140 169220 116150
rect 169320 116140 169400 116150
rect 169500 116140 169580 116150
rect 169680 116140 169760 116150
rect 169860 116140 169940 116150
rect 170040 116140 170120 116150
rect 170220 116140 170300 116150
rect 170400 116140 170480 116150
rect 170580 116140 170660 116150
rect 170760 116140 170840 116150
rect 170940 116140 171020 116150
rect 19060 116060 19070 116140
rect 19240 116060 19250 116140
rect 19420 116060 19430 116140
rect 19600 116060 19610 116140
rect 19780 116060 19790 116140
rect 19960 116060 19970 116140
rect 20140 116060 20150 116140
rect 20320 116060 20330 116140
rect 20500 116060 20510 116140
rect 20680 116060 20690 116140
rect 20860 116060 20870 116140
rect 21040 116060 21050 116140
rect 21220 116060 21230 116140
rect 21400 116060 21410 116140
rect 21580 116060 21590 116140
rect 21760 116060 21770 116140
rect 21940 116060 21950 116140
rect 22120 116060 22130 116140
rect 22300 116060 22310 116140
rect 22480 116060 22490 116140
rect 22660 116060 22670 116140
rect 22840 116060 22850 116140
rect 23020 116060 23030 116140
rect 23200 116060 23210 116140
rect 23380 116060 23390 116140
rect 23560 116060 23570 116140
rect 23740 116060 23750 116140
rect 23920 116060 23930 116140
rect 24100 116060 24110 116140
rect 24280 116060 24290 116140
rect 24460 116060 24470 116140
rect 24640 116060 24650 116140
rect 24820 116060 24830 116140
rect 25000 116060 25010 116140
rect 25180 116060 25190 116140
rect 25360 116060 25370 116140
rect 25540 116060 25550 116140
rect 25720 116060 25730 116140
rect 25900 116060 25910 116140
rect 26080 116060 26090 116140
rect 26260 116060 26270 116140
rect 26440 116060 26450 116140
rect 26620 116060 26630 116140
rect 30360 116060 30370 116140
rect 30540 116060 30550 116140
rect 30720 116060 30730 116140
rect 30900 116060 30910 116140
rect 31080 116060 31090 116140
rect 31260 116060 31270 116140
rect 31440 116060 31450 116140
rect 31620 116060 31630 116140
rect 31800 116060 31810 116140
rect 31980 116060 31990 116140
rect 32160 116060 32170 116140
rect 32340 116060 32350 116140
rect 32520 116060 32530 116140
rect 32700 116060 32710 116140
rect 32880 116060 32890 116140
rect 33060 116060 33070 116140
rect 33240 116060 33250 116140
rect 33420 116060 33430 116140
rect 33600 116060 33610 116140
rect 33780 116060 33790 116140
rect 33960 116060 33970 116140
rect 34140 116060 34150 116140
rect 34320 116060 34330 116140
rect 34500 116060 34510 116140
rect 34680 116060 34690 116140
rect 34860 116060 34870 116140
rect 35040 116060 35050 116140
rect 35220 116060 35230 116140
rect 35400 116060 35410 116140
rect 35580 116060 35590 116140
rect 35760 116060 35770 116140
rect 35940 116060 35950 116140
rect 36120 116060 36130 116140
rect 36300 116060 36310 116140
rect 36480 116060 36490 116140
rect 36660 116060 36670 116140
rect 36840 116060 36850 116140
rect 37020 116060 37030 116140
rect 37200 116060 37210 116140
rect 37380 116060 37390 116140
rect 37560 116060 37570 116140
rect 37740 116060 37750 116140
rect 37920 116060 37930 116140
rect 40140 116060 40150 116140
rect 40280 116060 40290 116140
rect 40420 116060 40430 116140
rect 40560 116060 40570 116140
rect 40700 116060 40710 116140
rect 40840 116060 40850 116140
rect 40980 116060 40990 116140
rect 41120 116060 41130 116140
rect 41260 116060 41270 116140
rect 41400 116060 41410 116140
rect 42440 116060 42450 116140
rect 42580 116060 42590 116140
rect 42720 116060 42730 116140
rect 42860 116060 42870 116140
rect 43000 116060 43010 116140
rect 43140 116060 43150 116140
rect 43280 116060 43290 116140
rect 43420 116060 43430 116140
rect 43560 116060 43570 116140
rect 43700 116060 43710 116140
rect 146380 116081 146390 116140
rect 146520 116081 146530 116140
rect 146660 116081 146670 116140
rect 146800 116081 146810 116140
rect 146940 116081 146950 116140
rect 147080 116081 147090 116140
rect 147220 116081 147230 116140
rect 147360 116081 147370 116140
rect 147500 116081 147510 116140
rect 147640 116081 147650 116140
rect 148680 116081 148690 116140
rect 148820 116081 148830 116140
rect 148960 116081 148970 116140
rect 149100 116081 149110 116140
rect 149240 116081 149250 116140
rect 149380 116081 149390 116140
rect 149520 116081 149530 116140
rect 149660 116081 149670 116140
rect 149800 116081 149810 116140
rect 149940 116081 149950 116140
rect 152160 116081 152170 116140
rect 152340 116081 152350 116140
rect 152520 116081 152530 116140
rect 152700 116081 152710 116140
rect 152880 116081 152890 116140
rect 153060 116081 153070 116140
rect 153240 116081 153250 116140
rect 153420 116081 153430 116140
rect 153600 116081 153610 116140
rect 153780 116081 153790 116140
rect 153960 116081 153970 116140
rect 154140 116081 154150 116140
rect 154320 116081 154330 116140
rect 154500 116081 154510 116140
rect 154680 116081 154690 116140
rect 154860 116081 154870 116140
rect 155040 116081 155050 116140
rect 155220 116081 155230 116140
rect 155400 116081 155410 116140
rect 155580 116081 155590 116140
rect 155760 116081 155770 116140
rect 155940 116081 155950 116140
rect 156120 116081 156130 116140
rect 156300 116081 156310 116140
rect 156480 116081 156490 116140
rect 156660 116081 156670 116140
rect 156840 116081 156850 116140
rect 157020 116081 157030 116140
rect 157200 116081 157210 116140
rect 157380 116081 157390 116140
rect 157560 116081 157570 116140
rect 157740 116081 157750 116140
rect 157920 116081 157930 116140
rect 158100 116081 158110 116140
rect 158280 116081 158290 116140
rect 158460 116081 158470 116140
rect 158640 116081 158650 116140
rect 158820 116081 158830 116140
rect 159000 116081 159010 116140
rect 159180 116081 159190 116140
rect 159360 116081 159370 116140
rect 159540 116081 159550 116140
rect 159720 116081 159730 116140
rect 163460 116081 163470 116140
rect 163640 116081 163650 116140
rect 163820 116081 163830 116140
rect 164000 116081 164010 116140
rect 164180 116081 164190 116140
rect 164360 116081 164370 116140
rect 164540 116081 164550 116140
rect 164720 116081 164730 116140
rect 164900 116081 164910 116140
rect 165080 116081 165090 116140
rect 165260 116081 165270 116140
rect 165440 116081 165450 116140
rect 165620 116081 165630 116140
rect 165800 116081 165810 116140
rect 165980 116081 165990 116140
rect 166160 116081 166170 116140
rect 166340 116081 166350 116140
rect 166520 116081 166530 116140
rect 166700 116081 166710 116140
rect 166880 116081 166890 116140
rect 167060 116081 167070 116140
rect 167240 116081 167250 116140
rect 167420 116081 167430 116140
rect 167600 116081 167610 116140
rect 167780 116081 167790 116140
rect 167960 116081 167970 116140
rect 168140 116081 168150 116140
rect 168320 116081 168330 116140
rect 168500 116081 168510 116140
rect 168680 116081 168690 116140
rect 168860 116081 168870 116140
rect 169040 116081 169050 116140
rect 169220 116081 169230 116140
rect 169400 116081 169410 116140
rect 169580 116081 169590 116140
rect 169760 116081 169770 116140
rect 169940 116081 169950 116140
rect 170120 116081 170130 116140
rect 170300 116081 170310 116140
rect 170480 116081 170490 116140
rect 170660 116081 170670 116140
rect 170840 116081 170850 116140
rect 171020 116081 171030 116140
rect 146040 116000 147700 116081
rect 148340 116000 150000 116081
rect 152000 116000 159800 116081
rect 163210 116060 171100 116081
rect 163300 116000 171100 116060
rect 30360 115920 30440 115930
rect 30680 115920 30760 115930
rect 31000 115920 31080 115930
rect 31320 115920 31400 115930
rect 31640 115920 31720 115930
rect 31960 115920 32040 115930
rect 32280 115920 32360 115930
rect 32600 115920 32680 115930
rect 32920 115920 33000 115930
rect 33240 115920 33320 115930
rect 33560 115920 33640 115930
rect 33880 115920 33960 115930
rect 34200 115920 34280 115930
rect 34520 115920 34600 115930
rect 34840 115920 34920 115930
rect 35160 115920 35240 115930
rect 35480 115920 35560 115930
rect 35800 115920 35880 115930
rect 36120 115920 36200 115930
rect 36440 115920 36520 115930
rect 36760 115920 36840 115930
rect 37080 115920 37160 115930
rect 37400 115920 37480 115930
rect 37720 115920 37800 115930
rect 40180 115920 40260 115930
rect 40500 115920 40580 115930
rect 40820 115920 40900 115930
rect 41140 115920 41220 115930
rect 42560 115920 42640 115930
rect 42880 115920 42960 115930
rect 43200 115920 43280 115930
rect 43520 115920 43600 115930
rect 18970 115890 19050 115900
rect 19290 115890 19370 115900
rect 19610 115890 19690 115900
rect 19930 115890 20010 115900
rect 20250 115890 20330 115900
rect 20570 115890 20650 115900
rect 20890 115890 20970 115900
rect 21210 115890 21290 115900
rect 21530 115890 21610 115900
rect 21850 115890 21930 115900
rect 22170 115890 22250 115900
rect 22490 115890 22570 115900
rect 22810 115890 22890 115900
rect 23130 115890 23210 115900
rect 23450 115890 23530 115900
rect 23770 115890 23850 115900
rect 24090 115890 24170 115900
rect 24410 115890 24490 115900
rect 24730 115890 24810 115900
rect 25050 115890 25130 115900
rect 25370 115890 25450 115900
rect 25690 115890 25770 115900
rect 26010 115890 26090 115900
rect 26330 115890 26410 115900
rect 19050 115810 19060 115890
rect 19370 115810 19380 115890
rect 19690 115810 19700 115890
rect 20010 115810 20020 115890
rect 20330 115810 20340 115890
rect 20650 115810 20660 115890
rect 20970 115810 20980 115890
rect 21290 115810 21300 115890
rect 21610 115810 21620 115890
rect 21930 115810 21940 115890
rect 22250 115810 22260 115890
rect 22570 115810 22580 115890
rect 22890 115810 22900 115890
rect 23210 115810 23220 115890
rect 23530 115810 23540 115890
rect 23850 115810 23860 115890
rect 24170 115810 24180 115890
rect 24490 115810 24500 115890
rect 24810 115810 24820 115890
rect 25130 115810 25140 115890
rect 25450 115810 25460 115890
rect 25770 115810 25780 115890
rect 26090 115810 26100 115890
rect 26410 115810 26420 115890
rect 30440 115840 30450 115920
rect 30760 115840 30770 115920
rect 31080 115840 31090 115920
rect 31400 115840 31410 115920
rect 31720 115840 31730 115920
rect 32040 115840 32050 115920
rect 32360 115840 32370 115920
rect 32680 115840 32690 115920
rect 33000 115840 33010 115920
rect 33320 115840 33330 115920
rect 33640 115840 33650 115920
rect 33960 115840 33970 115920
rect 34280 115840 34290 115920
rect 34600 115840 34610 115920
rect 34920 115840 34930 115920
rect 35240 115840 35250 115920
rect 35560 115840 35570 115920
rect 35880 115840 35890 115920
rect 36200 115840 36210 115920
rect 36520 115840 36530 115920
rect 36840 115840 36850 115920
rect 37160 115840 37170 115920
rect 37480 115840 37490 115920
rect 37800 115840 37810 115920
rect 40260 115840 40270 115920
rect 40580 115840 40590 115920
rect 40900 115840 40910 115920
rect 41220 115840 41230 115920
rect 42640 115840 42650 115920
rect 42960 115840 42970 115920
rect 43280 115840 43290 115920
rect 43600 115840 43610 115920
rect 146400 115911 146480 115921
rect 146720 115911 146800 115921
rect 147040 115911 147120 115921
rect 147360 115911 147440 115921
rect 148780 115911 148860 115921
rect 149100 115911 149180 115921
rect 149420 115911 149500 115921
rect 149740 115911 149820 115921
rect 152200 115911 152280 115921
rect 152520 115911 152600 115921
rect 152840 115911 152920 115921
rect 153160 115911 153240 115921
rect 153480 115911 153560 115921
rect 153800 115911 153880 115921
rect 154120 115911 154200 115921
rect 154440 115911 154520 115921
rect 154760 115911 154840 115921
rect 155080 115911 155160 115921
rect 155400 115911 155480 115921
rect 155720 115911 155800 115921
rect 156040 115911 156120 115921
rect 156360 115911 156440 115921
rect 156680 115911 156760 115921
rect 157000 115911 157080 115921
rect 157320 115911 157400 115921
rect 157640 115911 157720 115921
rect 157960 115911 158040 115921
rect 158280 115911 158360 115921
rect 158600 115911 158680 115921
rect 158920 115911 159000 115921
rect 159240 115911 159320 115921
rect 159560 115911 159640 115921
rect 146480 115831 146490 115911
rect 146800 115831 146810 115911
rect 147120 115831 147130 115911
rect 147440 115831 147450 115911
rect 148860 115831 148870 115911
rect 149180 115831 149190 115911
rect 149500 115831 149510 115911
rect 149820 115831 149830 115911
rect 152280 115831 152290 115911
rect 152600 115831 152610 115911
rect 152920 115831 152930 115911
rect 153240 115831 153250 115911
rect 153560 115831 153570 115911
rect 153880 115831 153890 115911
rect 154200 115831 154210 115911
rect 154520 115831 154530 115911
rect 154840 115831 154850 115911
rect 155160 115831 155170 115911
rect 155480 115831 155490 115911
rect 155800 115831 155810 115911
rect 156120 115831 156130 115911
rect 156440 115831 156450 115911
rect 156760 115831 156770 115911
rect 157080 115831 157090 115911
rect 157400 115831 157410 115911
rect 157720 115831 157730 115911
rect 158040 115831 158050 115911
rect 158360 115831 158370 115911
rect 158680 115831 158690 115911
rect 159000 115831 159010 115911
rect 159320 115831 159330 115911
rect 159640 115831 159650 115911
rect 163590 115881 163670 115891
rect 163910 115881 163990 115891
rect 164230 115881 164310 115891
rect 164550 115881 164630 115891
rect 164870 115881 164950 115891
rect 165190 115881 165270 115891
rect 165510 115881 165590 115891
rect 165830 115881 165910 115891
rect 166150 115881 166230 115891
rect 166470 115881 166550 115891
rect 166790 115881 166870 115891
rect 167110 115881 167190 115891
rect 167430 115881 167510 115891
rect 167750 115881 167830 115891
rect 168070 115881 168150 115891
rect 168390 115881 168470 115891
rect 168710 115881 168790 115891
rect 169030 115881 169110 115891
rect 169350 115881 169430 115891
rect 169670 115881 169750 115891
rect 169990 115881 170070 115891
rect 170310 115881 170390 115891
rect 170630 115881 170710 115891
rect 170950 115881 171030 115891
rect 163670 115801 163680 115881
rect 163990 115801 164000 115881
rect 164310 115801 164320 115881
rect 164630 115801 164640 115881
rect 164950 115801 164960 115881
rect 165270 115801 165280 115881
rect 165590 115801 165600 115881
rect 165910 115801 165920 115881
rect 166230 115801 166240 115881
rect 166550 115801 166560 115881
rect 166870 115801 166880 115881
rect 167190 115801 167200 115881
rect 167510 115801 167520 115881
rect 167830 115801 167840 115881
rect 168150 115801 168160 115881
rect 168470 115801 168480 115881
rect 168790 115801 168800 115881
rect 169110 115801 169120 115881
rect 169430 115801 169440 115881
rect 169750 115801 169760 115881
rect 170070 115801 170080 115881
rect 170390 115801 170400 115881
rect 170710 115801 170720 115881
rect 171030 115801 171040 115881
rect 30520 115760 30600 115770
rect 30840 115760 30920 115770
rect 31160 115760 31240 115770
rect 31480 115760 31560 115770
rect 31800 115760 31880 115770
rect 32120 115760 32200 115770
rect 32440 115760 32520 115770
rect 32760 115760 32840 115770
rect 33080 115760 33160 115770
rect 33400 115760 33480 115770
rect 33720 115760 33800 115770
rect 34040 115760 34120 115770
rect 34360 115760 34440 115770
rect 34680 115760 34760 115770
rect 35000 115760 35080 115770
rect 35320 115760 35400 115770
rect 35640 115760 35720 115770
rect 35960 115760 36040 115770
rect 36280 115760 36360 115770
rect 36600 115760 36680 115770
rect 36920 115760 37000 115770
rect 37240 115760 37320 115770
rect 37560 115760 37640 115770
rect 40340 115760 40420 115770
rect 40660 115760 40740 115770
rect 40980 115760 41060 115770
rect 42720 115760 42800 115770
rect 43040 115760 43120 115770
rect 43360 115760 43440 115770
rect 19130 115730 19210 115740
rect 19450 115730 19530 115740
rect 19770 115730 19850 115740
rect 20090 115730 20170 115740
rect 20410 115730 20490 115740
rect 20730 115730 20810 115740
rect 21050 115730 21130 115740
rect 21370 115730 21450 115740
rect 21690 115730 21770 115740
rect 22010 115730 22090 115740
rect 22330 115730 22410 115740
rect 22650 115730 22730 115740
rect 22970 115730 23050 115740
rect 23290 115730 23370 115740
rect 23610 115730 23690 115740
rect 23930 115730 24010 115740
rect 24250 115730 24330 115740
rect 24570 115730 24650 115740
rect 24890 115730 24970 115740
rect 25210 115730 25290 115740
rect 25530 115730 25610 115740
rect 25850 115730 25930 115740
rect 26170 115730 26250 115740
rect 19210 115650 19220 115730
rect 19530 115650 19540 115730
rect 19850 115650 19860 115730
rect 20170 115650 20180 115730
rect 20490 115650 20500 115730
rect 20810 115650 20820 115730
rect 21130 115650 21140 115730
rect 21450 115650 21460 115730
rect 21770 115650 21780 115730
rect 22090 115650 22100 115730
rect 22410 115650 22420 115730
rect 22730 115650 22740 115730
rect 23050 115650 23060 115730
rect 23370 115650 23380 115730
rect 23690 115650 23700 115730
rect 24010 115650 24020 115730
rect 24330 115650 24340 115730
rect 24650 115650 24660 115730
rect 24970 115650 24980 115730
rect 25290 115650 25300 115730
rect 25610 115650 25620 115730
rect 25930 115650 25940 115730
rect 26250 115650 26260 115730
rect 30600 115680 30610 115760
rect 30920 115680 30930 115760
rect 31240 115680 31250 115760
rect 31560 115680 31570 115760
rect 31880 115680 31890 115760
rect 32200 115680 32210 115760
rect 32520 115680 32530 115760
rect 32840 115680 32850 115760
rect 33160 115680 33170 115760
rect 33480 115680 33490 115760
rect 33800 115680 33810 115760
rect 34120 115680 34130 115760
rect 34440 115680 34450 115760
rect 34760 115680 34770 115760
rect 35080 115680 35090 115760
rect 35400 115680 35410 115760
rect 35720 115680 35730 115760
rect 36040 115680 36050 115760
rect 36360 115680 36370 115760
rect 36680 115680 36690 115760
rect 37000 115680 37010 115760
rect 37320 115680 37330 115760
rect 37640 115680 37650 115760
rect 40420 115680 40430 115760
rect 40740 115680 40750 115760
rect 41060 115680 41070 115760
rect 42800 115680 42810 115760
rect 43120 115680 43130 115760
rect 43440 115680 43450 115760
rect 146560 115751 146640 115761
rect 146880 115751 146960 115761
rect 147200 115751 147280 115761
rect 148940 115751 149020 115761
rect 149260 115751 149340 115761
rect 149580 115751 149660 115761
rect 152360 115751 152440 115761
rect 152680 115751 152760 115761
rect 153000 115751 153080 115761
rect 153320 115751 153400 115761
rect 153640 115751 153720 115761
rect 153960 115751 154040 115761
rect 154280 115751 154360 115761
rect 154600 115751 154680 115761
rect 154920 115751 155000 115761
rect 155240 115751 155320 115761
rect 155560 115751 155640 115761
rect 155880 115751 155960 115761
rect 156200 115751 156280 115761
rect 156520 115751 156600 115761
rect 156840 115751 156920 115761
rect 157160 115751 157240 115761
rect 157480 115751 157560 115761
rect 157800 115751 157880 115761
rect 158120 115751 158200 115761
rect 158440 115751 158520 115761
rect 158760 115751 158840 115761
rect 159080 115751 159160 115761
rect 159400 115751 159480 115761
rect 146640 115671 146650 115751
rect 146960 115671 146970 115751
rect 147280 115671 147290 115751
rect 149020 115671 149030 115751
rect 149340 115671 149350 115751
rect 149660 115671 149670 115751
rect 152440 115671 152450 115751
rect 152760 115671 152770 115751
rect 153080 115671 153090 115751
rect 153400 115671 153410 115751
rect 153720 115671 153730 115751
rect 154040 115671 154050 115751
rect 154360 115671 154370 115751
rect 154680 115671 154690 115751
rect 155000 115671 155010 115751
rect 155320 115671 155330 115751
rect 155640 115671 155650 115751
rect 155960 115671 155970 115751
rect 156280 115671 156290 115751
rect 156600 115671 156610 115751
rect 156920 115671 156930 115751
rect 157240 115671 157250 115751
rect 157560 115671 157570 115751
rect 157880 115671 157890 115751
rect 158200 115671 158210 115751
rect 158520 115671 158530 115751
rect 158840 115671 158850 115751
rect 159160 115671 159170 115751
rect 159480 115671 159490 115751
rect 163750 115721 163830 115731
rect 164070 115721 164150 115731
rect 164390 115721 164470 115731
rect 164710 115721 164790 115731
rect 165030 115721 165110 115731
rect 165350 115721 165430 115731
rect 165670 115721 165750 115731
rect 165990 115721 166070 115731
rect 166310 115721 166390 115731
rect 166630 115721 166710 115731
rect 166950 115721 167030 115731
rect 167270 115721 167350 115731
rect 167590 115721 167670 115731
rect 167910 115721 167990 115731
rect 168230 115721 168310 115731
rect 168550 115721 168630 115731
rect 168870 115721 168950 115731
rect 169190 115721 169270 115731
rect 169510 115721 169590 115731
rect 169830 115721 169910 115731
rect 170150 115721 170230 115731
rect 170470 115721 170550 115731
rect 170790 115721 170870 115731
rect 163830 115641 163840 115721
rect 164150 115641 164160 115721
rect 164470 115641 164480 115721
rect 164790 115641 164800 115721
rect 165110 115641 165120 115721
rect 165430 115641 165440 115721
rect 165750 115641 165760 115721
rect 166070 115641 166080 115721
rect 166390 115641 166400 115721
rect 166710 115641 166720 115721
rect 167030 115641 167040 115721
rect 167350 115641 167360 115721
rect 167670 115641 167680 115721
rect 167990 115641 168000 115721
rect 168310 115641 168320 115721
rect 168630 115641 168640 115721
rect 168950 115641 168960 115721
rect 169270 115641 169280 115721
rect 169590 115641 169600 115721
rect 169910 115641 169920 115721
rect 170230 115641 170240 115721
rect 170550 115641 170560 115721
rect 170870 115641 170880 115721
rect 30360 115600 30440 115610
rect 30680 115600 30760 115610
rect 31000 115600 31080 115610
rect 31320 115600 31400 115610
rect 31640 115600 31720 115610
rect 31960 115600 32040 115610
rect 32280 115600 32360 115610
rect 32600 115600 32680 115610
rect 32920 115600 33000 115610
rect 33240 115600 33320 115610
rect 33560 115600 33640 115610
rect 33880 115600 33960 115610
rect 34200 115600 34280 115610
rect 34520 115600 34600 115610
rect 34840 115600 34920 115610
rect 35160 115600 35240 115610
rect 35480 115600 35560 115610
rect 35800 115600 35880 115610
rect 36120 115600 36200 115610
rect 36440 115600 36520 115610
rect 36760 115600 36840 115610
rect 37080 115600 37160 115610
rect 37400 115600 37480 115610
rect 37720 115600 37800 115610
rect 40180 115600 40260 115610
rect 40500 115600 40580 115610
rect 40820 115600 40900 115610
rect 41140 115600 41220 115610
rect 42560 115600 42640 115610
rect 42880 115600 42960 115610
rect 43200 115600 43280 115610
rect 43520 115600 43600 115610
rect 18970 115570 19050 115580
rect 19290 115570 19370 115580
rect 19610 115570 19690 115580
rect 19930 115570 20010 115580
rect 20250 115570 20330 115580
rect 20570 115570 20650 115580
rect 20890 115570 20970 115580
rect 21210 115570 21290 115580
rect 21530 115570 21610 115580
rect 21850 115570 21930 115580
rect 22170 115570 22250 115580
rect 22490 115570 22570 115580
rect 22810 115570 22890 115580
rect 23130 115570 23210 115580
rect 23450 115570 23530 115580
rect 23770 115570 23850 115580
rect 24090 115570 24170 115580
rect 24410 115570 24490 115580
rect 24730 115570 24810 115580
rect 25050 115570 25130 115580
rect 25370 115570 25450 115580
rect 25690 115570 25770 115580
rect 26010 115570 26090 115580
rect 26330 115570 26410 115580
rect 19050 115490 19060 115570
rect 19370 115490 19380 115570
rect 19690 115490 19700 115570
rect 20010 115490 20020 115570
rect 20330 115490 20340 115570
rect 20650 115490 20660 115570
rect 20970 115490 20980 115570
rect 21290 115490 21300 115570
rect 21610 115490 21620 115570
rect 21930 115490 21940 115570
rect 22250 115490 22260 115570
rect 22570 115490 22580 115570
rect 22890 115490 22900 115570
rect 23210 115490 23220 115570
rect 23530 115490 23540 115570
rect 23850 115490 23860 115570
rect 24170 115490 24180 115570
rect 24490 115490 24500 115570
rect 24810 115490 24820 115570
rect 25130 115490 25140 115570
rect 25450 115490 25460 115570
rect 25770 115490 25780 115570
rect 26090 115490 26100 115570
rect 26410 115490 26420 115570
rect 30440 115520 30450 115600
rect 30760 115520 30770 115600
rect 31080 115520 31090 115600
rect 31400 115520 31410 115600
rect 31720 115520 31730 115600
rect 32040 115520 32050 115600
rect 32360 115520 32370 115600
rect 32680 115520 32690 115600
rect 33000 115520 33010 115600
rect 33320 115520 33330 115600
rect 33640 115520 33650 115600
rect 33960 115520 33970 115600
rect 34280 115520 34290 115600
rect 34600 115520 34610 115600
rect 34920 115520 34930 115600
rect 35240 115520 35250 115600
rect 35560 115520 35570 115600
rect 35880 115520 35890 115600
rect 36200 115520 36210 115600
rect 36520 115520 36530 115600
rect 36840 115520 36850 115600
rect 37160 115520 37170 115600
rect 37480 115520 37490 115600
rect 37800 115520 37810 115600
rect 40260 115520 40270 115600
rect 40580 115520 40590 115600
rect 40900 115520 40910 115600
rect 41220 115520 41230 115600
rect 42640 115520 42650 115600
rect 42960 115520 42970 115600
rect 43280 115520 43290 115600
rect 43600 115520 43610 115600
rect 146400 115591 146480 115601
rect 146720 115591 146800 115601
rect 147040 115591 147120 115601
rect 147360 115591 147440 115601
rect 148780 115591 148860 115601
rect 149100 115591 149180 115601
rect 149420 115591 149500 115601
rect 149740 115591 149820 115601
rect 152200 115591 152280 115601
rect 152520 115591 152600 115601
rect 152840 115591 152920 115601
rect 153160 115591 153240 115601
rect 153480 115591 153560 115601
rect 153800 115591 153880 115601
rect 154120 115591 154200 115601
rect 154440 115591 154520 115601
rect 154760 115591 154840 115601
rect 155080 115591 155160 115601
rect 155400 115591 155480 115601
rect 155720 115591 155800 115601
rect 156040 115591 156120 115601
rect 156360 115591 156440 115601
rect 156680 115591 156760 115601
rect 157000 115591 157080 115601
rect 157320 115591 157400 115601
rect 157640 115591 157720 115601
rect 157960 115591 158040 115601
rect 158280 115591 158360 115601
rect 158600 115591 158680 115601
rect 158920 115591 159000 115601
rect 159240 115591 159320 115601
rect 159560 115591 159640 115601
rect 146480 115511 146490 115591
rect 146800 115511 146810 115591
rect 147120 115511 147130 115591
rect 147440 115511 147450 115591
rect 148860 115511 148870 115591
rect 149180 115511 149190 115591
rect 149500 115511 149510 115591
rect 149820 115511 149830 115591
rect 152280 115511 152290 115591
rect 152600 115511 152610 115591
rect 152920 115511 152930 115591
rect 153240 115511 153250 115591
rect 153560 115511 153570 115591
rect 153880 115511 153890 115591
rect 154200 115511 154210 115591
rect 154520 115511 154530 115591
rect 154840 115511 154850 115591
rect 155160 115511 155170 115591
rect 155480 115511 155490 115591
rect 155800 115511 155810 115591
rect 156120 115511 156130 115591
rect 156440 115511 156450 115591
rect 156760 115511 156770 115591
rect 157080 115511 157090 115591
rect 157400 115511 157410 115591
rect 157720 115511 157730 115591
rect 158040 115511 158050 115591
rect 158360 115511 158370 115591
rect 158680 115511 158690 115591
rect 159000 115511 159010 115591
rect 159320 115511 159330 115591
rect 159640 115511 159650 115591
rect 163590 115561 163670 115571
rect 163910 115561 163990 115571
rect 164230 115561 164310 115571
rect 164550 115561 164630 115571
rect 164870 115561 164950 115571
rect 165190 115561 165270 115571
rect 165510 115561 165590 115571
rect 165830 115561 165910 115571
rect 166150 115561 166230 115571
rect 166470 115561 166550 115571
rect 166790 115561 166870 115571
rect 167110 115561 167190 115571
rect 167430 115561 167510 115571
rect 167750 115561 167830 115571
rect 168070 115561 168150 115571
rect 168390 115561 168470 115571
rect 168710 115561 168790 115571
rect 169030 115561 169110 115571
rect 169350 115561 169430 115571
rect 169670 115561 169750 115571
rect 169990 115561 170070 115571
rect 170310 115561 170390 115571
rect 170630 115561 170710 115571
rect 170950 115561 171030 115571
rect 163670 115481 163680 115561
rect 163990 115481 164000 115561
rect 164310 115481 164320 115561
rect 164630 115481 164640 115561
rect 164950 115481 164960 115561
rect 165270 115481 165280 115561
rect 165590 115481 165600 115561
rect 165910 115481 165920 115561
rect 166230 115481 166240 115561
rect 166550 115481 166560 115561
rect 166870 115481 166880 115561
rect 167190 115481 167200 115561
rect 167510 115481 167520 115561
rect 167830 115481 167840 115561
rect 168150 115481 168160 115561
rect 168470 115481 168480 115561
rect 168790 115481 168800 115561
rect 169110 115481 169120 115561
rect 169430 115481 169440 115561
rect 169750 115481 169760 115561
rect 170070 115481 170080 115561
rect 170390 115481 170400 115561
rect 170710 115481 170720 115561
rect 171030 115481 171040 115561
rect 30520 115440 30600 115450
rect 30840 115440 30920 115450
rect 31160 115440 31240 115450
rect 31480 115440 31560 115450
rect 31800 115440 31880 115450
rect 32120 115440 32200 115450
rect 32440 115440 32520 115450
rect 32760 115440 32840 115450
rect 33080 115440 33160 115450
rect 33400 115440 33480 115450
rect 33720 115440 33800 115450
rect 34040 115440 34120 115450
rect 34360 115440 34440 115450
rect 34680 115440 34760 115450
rect 35000 115440 35080 115450
rect 35320 115440 35400 115450
rect 35640 115440 35720 115450
rect 35960 115440 36040 115450
rect 36280 115440 36360 115450
rect 36600 115440 36680 115450
rect 36920 115440 37000 115450
rect 37240 115440 37320 115450
rect 37560 115440 37640 115450
rect 40340 115440 40420 115450
rect 40660 115440 40740 115450
rect 40980 115440 41060 115450
rect 42720 115440 42800 115450
rect 43040 115440 43120 115450
rect 43360 115440 43440 115450
rect 19130 115410 19210 115420
rect 19450 115410 19530 115420
rect 19770 115410 19850 115420
rect 20090 115410 20170 115420
rect 20410 115410 20490 115420
rect 20730 115410 20810 115420
rect 21050 115410 21130 115420
rect 21370 115410 21450 115420
rect 21690 115410 21770 115420
rect 22010 115410 22090 115420
rect 22330 115410 22410 115420
rect 22650 115410 22730 115420
rect 22970 115410 23050 115420
rect 23290 115410 23370 115420
rect 23610 115410 23690 115420
rect 23930 115410 24010 115420
rect 24250 115410 24330 115420
rect 24570 115410 24650 115420
rect 24890 115410 24970 115420
rect 25210 115410 25290 115420
rect 25530 115410 25610 115420
rect 25850 115410 25930 115420
rect 26170 115410 26250 115420
rect 19210 115330 19220 115410
rect 19530 115330 19540 115410
rect 19850 115330 19860 115410
rect 20170 115330 20180 115410
rect 20490 115330 20500 115410
rect 20810 115330 20820 115410
rect 21130 115330 21140 115410
rect 21450 115330 21460 115410
rect 21770 115330 21780 115410
rect 22090 115330 22100 115410
rect 22410 115330 22420 115410
rect 22730 115330 22740 115410
rect 23050 115330 23060 115410
rect 23370 115330 23380 115410
rect 23690 115330 23700 115410
rect 24010 115330 24020 115410
rect 24330 115330 24340 115410
rect 24650 115330 24660 115410
rect 24970 115330 24980 115410
rect 25290 115330 25300 115410
rect 25610 115330 25620 115410
rect 25930 115330 25940 115410
rect 26250 115330 26260 115410
rect 30600 115360 30610 115440
rect 30920 115360 30930 115440
rect 31240 115360 31250 115440
rect 31560 115360 31570 115440
rect 31880 115360 31890 115440
rect 32200 115360 32210 115440
rect 32520 115360 32530 115440
rect 32840 115360 32850 115440
rect 33160 115360 33170 115440
rect 33480 115360 33490 115440
rect 33800 115360 33810 115440
rect 34120 115360 34130 115440
rect 34440 115360 34450 115440
rect 34760 115360 34770 115440
rect 35080 115360 35090 115440
rect 35400 115360 35410 115440
rect 35720 115360 35730 115440
rect 36040 115360 36050 115440
rect 36360 115360 36370 115440
rect 36680 115360 36690 115440
rect 37000 115360 37010 115440
rect 37320 115360 37330 115440
rect 37640 115360 37650 115440
rect 40420 115360 40430 115440
rect 40740 115360 40750 115440
rect 41060 115360 41070 115440
rect 42800 115360 42810 115440
rect 43120 115360 43130 115440
rect 43440 115360 43450 115440
rect 146560 115431 146640 115441
rect 146880 115431 146960 115441
rect 147200 115431 147280 115441
rect 148940 115431 149020 115441
rect 149260 115431 149340 115441
rect 149580 115431 149660 115441
rect 152360 115431 152440 115441
rect 152680 115431 152760 115441
rect 153000 115431 153080 115441
rect 153320 115431 153400 115441
rect 153640 115431 153720 115441
rect 153960 115431 154040 115441
rect 154280 115431 154360 115441
rect 154600 115431 154680 115441
rect 154920 115431 155000 115441
rect 155240 115431 155320 115441
rect 155560 115431 155640 115441
rect 155880 115431 155960 115441
rect 156200 115431 156280 115441
rect 156520 115431 156600 115441
rect 156840 115431 156920 115441
rect 157160 115431 157240 115441
rect 157480 115431 157560 115441
rect 157800 115431 157880 115441
rect 158120 115431 158200 115441
rect 158440 115431 158520 115441
rect 158760 115431 158840 115441
rect 159080 115431 159160 115441
rect 159400 115431 159480 115441
rect 146640 115351 146650 115431
rect 146960 115351 146970 115431
rect 147280 115351 147290 115431
rect 149020 115351 149030 115431
rect 149340 115351 149350 115431
rect 149660 115351 149670 115431
rect 152440 115351 152450 115431
rect 152760 115351 152770 115431
rect 153080 115351 153090 115431
rect 153400 115351 153410 115431
rect 153720 115351 153730 115431
rect 154040 115351 154050 115431
rect 154360 115351 154370 115431
rect 154680 115351 154690 115431
rect 155000 115351 155010 115431
rect 155320 115351 155330 115431
rect 155640 115351 155650 115431
rect 155960 115351 155970 115431
rect 156280 115351 156290 115431
rect 156600 115351 156610 115431
rect 156920 115351 156930 115431
rect 157240 115351 157250 115431
rect 157560 115351 157570 115431
rect 157880 115351 157890 115431
rect 158200 115351 158210 115431
rect 158520 115351 158530 115431
rect 158840 115351 158850 115431
rect 159160 115351 159170 115431
rect 159480 115351 159490 115431
rect 163750 115401 163830 115411
rect 164070 115401 164150 115411
rect 164390 115401 164470 115411
rect 164710 115401 164790 115411
rect 165030 115401 165110 115411
rect 165350 115401 165430 115411
rect 165670 115401 165750 115411
rect 165990 115401 166070 115411
rect 166310 115401 166390 115411
rect 166630 115401 166710 115411
rect 166950 115401 167030 115411
rect 167270 115401 167350 115411
rect 167590 115401 167670 115411
rect 167910 115401 167990 115411
rect 168230 115401 168310 115411
rect 168550 115401 168630 115411
rect 168870 115401 168950 115411
rect 169190 115401 169270 115411
rect 169510 115401 169590 115411
rect 169830 115401 169910 115411
rect 170150 115401 170230 115411
rect 170470 115401 170550 115411
rect 170790 115401 170870 115411
rect 163830 115321 163840 115401
rect 164150 115321 164160 115401
rect 164470 115321 164480 115401
rect 164790 115321 164800 115401
rect 165110 115321 165120 115401
rect 165430 115321 165440 115401
rect 165750 115321 165760 115401
rect 166070 115321 166080 115401
rect 166390 115321 166400 115401
rect 166710 115321 166720 115401
rect 167030 115321 167040 115401
rect 167350 115321 167360 115401
rect 167670 115321 167680 115401
rect 167990 115321 168000 115401
rect 168310 115321 168320 115401
rect 168630 115321 168640 115401
rect 168950 115321 168960 115401
rect 169270 115321 169280 115401
rect 169590 115321 169600 115401
rect 169910 115321 169920 115401
rect 170230 115321 170240 115401
rect 170550 115321 170560 115401
rect 170870 115321 170880 115401
rect 30360 115180 30440 115190
rect 30680 115180 30760 115190
rect 31000 115180 31080 115190
rect 31320 115180 31400 115190
rect 31640 115180 31720 115190
rect 31960 115180 32040 115190
rect 32280 115180 32360 115190
rect 32600 115180 32680 115190
rect 32920 115180 33000 115190
rect 33240 115180 33320 115190
rect 33560 115180 33640 115190
rect 33880 115180 33960 115190
rect 34200 115180 34280 115190
rect 34520 115180 34600 115190
rect 34840 115180 34920 115190
rect 35160 115180 35240 115190
rect 35480 115180 35560 115190
rect 35800 115180 35880 115190
rect 36120 115180 36200 115190
rect 36440 115180 36520 115190
rect 36760 115180 36840 115190
rect 37080 115180 37160 115190
rect 37400 115180 37480 115190
rect 37720 115180 37800 115190
rect 40180 115180 40260 115190
rect 40500 115180 40580 115190
rect 40820 115180 40900 115190
rect 41140 115180 41220 115190
rect 42560 115180 42640 115190
rect 42880 115180 42960 115190
rect 43200 115180 43280 115190
rect 43520 115180 43600 115190
rect 18970 115150 19050 115160
rect 19290 115150 19370 115160
rect 19610 115150 19690 115160
rect 19930 115150 20010 115160
rect 20250 115150 20330 115160
rect 20570 115150 20650 115160
rect 20890 115150 20970 115160
rect 21210 115150 21290 115160
rect 21530 115150 21610 115160
rect 21850 115150 21930 115160
rect 22170 115150 22250 115160
rect 22490 115150 22570 115160
rect 22810 115150 22890 115160
rect 23130 115150 23210 115160
rect 23450 115150 23530 115160
rect 23770 115150 23850 115160
rect 24090 115150 24170 115160
rect 24410 115150 24490 115160
rect 24730 115150 24810 115160
rect 25050 115150 25130 115160
rect 25370 115150 25450 115160
rect 25690 115150 25770 115160
rect 26010 115150 26090 115160
rect 26330 115150 26410 115160
rect 19050 115070 19060 115150
rect 19370 115070 19380 115150
rect 19690 115070 19700 115150
rect 20010 115070 20020 115150
rect 20330 115070 20340 115150
rect 20650 115070 20660 115150
rect 20970 115070 20980 115150
rect 21290 115070 21300 115150
rect 21610 115070 21620 115150
rect 21930 115070 21940 115150
rect 22250 115070 22260 115150
rect 22570 115070 22580 115150
rect 22890 115070 22900 115150
rect 23210 115070 23220 115150
rect 23530 115070 23540 115150
rect 23850 115070 23860 115150
rect 24170 115070 24180 115150
rect 24490 115070 24500 115150
rect 24810 115070 24820 115150
rect 25130 115070 25140 115150
rect 25450 115070 25460 115150
rect 25770 115070 25780 115150
rect 26090 115070 26100 115150
rect 26410 115070 26420 115150
rect 30440 115100 30450 115180
rect 30760 115100 30770 115180
rect 31080 115100 31090 115180
rect 31400 115100 31410 115180
rect 31720 115100 31730 115180
rect 32040 115100 32050 115180
rect 32360 115100 32370 115180
rect 32680 115100 32690 115180
rect 33000 115100 33010 115180
rect 33320 115100 33330 115180
rect 33640 115100 33650 115180
rect 33960 115100 33970 115180
rect 34280 115100 34290 115180
rect 34600 115100 34610 115180
rect 34920 115100 34930 115180
rect 35240 115100 35250 115180
rect 35560 115100 35570 115180
rect 35880 115100 35890 115180
rect 36200 115100 36210 115180
rect 36520 115100 36530 115180
rect 36840 115100 36850 115180
rect 37160 115100 37170 115180
rect 37480 115100 37490 115180
rect 37800 115100 37810 115180
rect 40260 115100 40270 115180
rect 40580 115100 40590 115180
rect 40900 115100 40910 115180
rect 41220 115100 41230 115180
rect 42640 115100 42650 115180
rect 42960 115100 42970 115180
rect 43280 115100 43290 115180
rect 43600 115100 43610 115180
rect 146400 115171 146480 115181
rect 146720 115171 146800 115181
rect 147040 115171 147120 115181
rect 147360 115171 147440 115181
rect 148780 115171 148860 115181
rect 149100 115171 149180 115181
rect 149420 115171 149500 115181
rect 149740 115171 149820 115181
rect 152200 115171 152280 115181
rect 152520 115171 152600 115181
rect 152840 115171 152920 115181
rect 153160 115171 153240 115181
rect 153480 115171 153560 115181
rect 153800 115171 153880 115181
rect 154120 115171 154200 115181
rect 154440 115171 154520 115181
rect 154760 115171 154840 115181
rect 155080 115171 155160 115181
rect 155400 115171 155480 115181
rect 155720 115171 155800 115181
rect 156040 115171 156120 115181
rect 156360 115171 156440 115181
rect 156680 115171 156760 115181
rect 157000 115171 157080 115181
rect 157320 115171 157400 115181
rect 157640 115171 157720 115181
rect 157960 115171 158040 115181
rect 158280 115171 158360 115181
rect 158600 115171 158680 115181
rect 158920 115171 159000 115181
rect 159240 115171 159320 115181
rect 159560 115171 159640 115181
rect 146480 115091 146490 115171
rect 146800 115091 146810 115171
rect 147120 115091 147130 115171
rect 147440 115091 147450 115171
rect 148860 115091 148870 115171
rect 149180 115091 149190 115171
rect 149500 115091 149510 115171
rect 149820 115091 149830 115171
rect 152280 115091 152290 115171
rect 152600 115091 152610 115171
rect 152920 115091 152930 115171
rect 153240 115091 153250 115171
rect 153560 115091 153570 115171
rect 153880 115091 153890 115171
rect 154200 115091 154210 115171
rect 154520 115091 154530 115171
rect 154840 115091 154850 115171
rect 155160 115091 155170 115171
rect 155480 115091 155490 115171
rect 155800 115091 155810 115171
rect 156120 115091 156130 115171
rect 156440 115091 156450 115171
rect 156760 115091 156770 115171
rect 157080 115091 157090 115171
rect 157400 115091 157410 115171
rect 157720 115091 157730 115171
rect 158040 115091 158050 115171
rect 158360 115091 158370 115171
rect 158680 115091 158690 115171
rect 159000 115091 159010 115171
rect 159320 115091 159330 115171
rect 159640 115091 159650 115171
rect 163590 115141 163670 115151
rect 163910 115141 163990 115151
rect 164230 115141 164310 115151
rect 164550 115141 164630 115151
rect 164870 115141 164950 115151
rect 165190 115141 165270 115151
rect 165510 115141 165590 115151
rect 165830 115141 165910 115151
rect 166150 115141 166230 115151
rect 166470 115141 166550 115151
rect 166790 115141 166870 115151
rect 167110 115141 167190 115151
rect 167430 115141 167510 115151
rect 167750 115141 167830 115151
rect 168070 115141 168150 115151
rect 168390 115141 168470 115151
rect 168710 115141 168790 115151
rect 169030 115141 169110 115151
rect 169350 115141 169430 115151
rect 169670 115141 169750 115151
rect 169990 115141 170070 115151
rect 170310 115141 170390 115151
rect 170630 115141 170710 115151
rect 170950 115141 171030 115151
rect 163670 115061 163680 115141
rect 163990 115061 164000 115141
rect 164310 115061 164320 115141
rect 164630 115061 164640 115141
rect 164950 115061 164960 115141
rect 165270 115061 165280 115141
rect 165590 115061 165600 115141
rect 165910 115061 165920 115141
rect 166230 115061 166240 115141
rect 166550 115061 166560 115141
rect 166870 115061 166880 115141
rect 167190 115061 167200 115141
rect 167510 115061 167520 115141
rect 167830 115061 167840 115141
rect 168150 115061 168160 115141
rect 168470 115061 168480 115141
rect 168790 115061 168800 115141
rect 169110 115061 169120 115141
rect 169430 115061 169440 115141
rect 169750 115061 169760 115141
rect 170070 115061 170080 115141
rect 170390 115061 170400 115141
rect 170710 115061 170720 115141
rect 171030 115061 171040 115141
rect 30520 115020 30600 115030
rect 30840 115020 30920 115030
rect 31160 115020 31240 115030
rect 31480 115020 31560 115030
rect 31800 115020 31880 115030
rect 32120 115020 32200 115030
rect 32440 115020 32520 115030
rect 32760 115020 32840 115030
rect 33080 115020 33160 115030
rect 33400 115020 33480 115030
rect 33720 115020 33800 115030
rect 34040 115020 34120 115030
rect 34360 115020 34440 115030
rect 34680 115020 34760 115030
rect 35000 115020 35080 115030
rect 35320 115020 35400 115030
rect 35640 115020 35720 115030
rect 35960 115020 36040 115030
rect 36280 115020 36360 115030
rect 36600 115020 36680 115030
rect 36920 115020 37000 115030
rect 37240 115020 37320 115030
rect 37560 115020 37640 115030
rect 40340 115020 40420 115030
rect 40660 115020 40740 115030
rect 40980 115020 41060 115030
rect 42720 115020 42800 115030
rect 43040 115020 43120 115030
rect 43360 115020 43440 115030
rect 19130 114990 19210 115000
rect 19450 114990 19530 115000
rect 19770 114990 19850 115000
rect 20090 114990 20170 115000
rect 20410 114990 20490 115000
rect 20730 114990 20810 115000
rect 21050 114990 21130 115000
rect 21370 114990 21450 115000
rect 21690 114990 21770 115000
rect 22010 114990 22090 115000
rect 22330 114990 22410 115000
rect 22650 114990 22730 115000
rect 22970 114990 23050 115000
rect 23290 114990 23370 115000
rect 23610 114990 23690 115000
rect 23930 114990 24010 115000
rect 24250 114990 24330 115000
rect 24570 114990 24650 115000
rect 24890 114990 24970 115000
rect 25210 114990 25290 115000
rect 25530 114990 25610 115000
rect 25850 114990 25930 115000
rect 26170 114990 26250 115000
rect 19210 114910 19220 114990
rect 19530 114910 19540 114990
rect 19850 114910 19860 114990
rect 20170 114910 20180 114990
rect 20490 114910 20500 114990
rect 20810 114910 20820 114990
rect 21130 114910 21140 114990
rect 21450 114910 21460 114990
rect 21770 114910 21780 114990
rect 22090 114910 22100 114990
rect 22410 114910 22420 114990
rect 22730 114910 22740 114990
rect 23050 114910 23060 114990
rect 23370 114910 23380 114990
rect 23690 114910 23700 114990
rect 24010 114910 24020 114990
rect 24330 114910 24340 114990
rect 24650 114910 24660 114990
rect 24970 114910 24980 114990
rect 25290 114910 25300 114990
rect 25610 114910 25620 114990
rect 25930 114910 25940 114990
rect 26250 114910 26260 114990
rect 30600 114940 30610 115020
rect 30920 114940 30930 115020
rect 31240 114940 31250 115020
rect 31560 114940 31570 115020
rect 31880 114940 31890 115020
rect 32200 114940 32210 115020
rect 32520 114940 32530 115020
rect 32840 114940 32850 115020
rect 33160 114940 33170 115020
rect 33480 114940 33490 115020
rect 33800 114940 33810 115020
rect 34120 114940 34130 115020
rect 34440 114940 34450 115020
rect 34760 114940 34770 115020
rect 35080 114940 35090 115020
rect 35400 114940 35410 115020
rect 35720 114940 35730 115020
rect 36040 114940 36050 115020
rect 36360 114940 36370 115020
rect 36680 114940 36690 115020
rect 37000 114940 37010 115020
rect 37320 114940 37330 115020
rect 37640 114940 37650 115020
rect 40420 114940 40430 115020
rect 40740 114940 40750 115020
rect 41060 114940 41070 115020
rect 42800 114940 42810 115020
rect 43120 114940 43130 115020
rect 43440 114940 43450 115020
rect 146560 115011 146640 115021
rect 146880 115011 146960 115021
rect 147200 115011 147280 115021
rect 148940 115011 149020 115021
rect 149260 115011 149340 115021
rect 149580 115011 149660 115021
rect 152360 115011 152440 115021
rect 152680 115011 152760 115021
rect 153000 115011 153080 115021
rect 153320 115011 153400 115021
rect 153640 115011 153720 115021
rect 153960 115011 154040 115021
rect 154280 115011 154360 115021
rect 154600 115011 154680 115021
rect 154920 115011 155000 115021
rect 155240 115011 155320 115021
rect 155560 115011 155640 115021
rect 155880 115011 155960 115021
rect 156200 115011 156280 115021
rect 156520 115011 156600 115021
rect 156840 115011 156920 115021
rect 157160 115011 157240 115021
rect 157480 115011 157560 115021
rect 157800 115011 157880 115021
rect 158120 115011 158200 115021
rect 158440 115011 158520 115021
rect 158760 115011 158840 115021
rect 159080 115011 159160 115021
rect 159400 115011 159480 115021
rect 146640 114931 146650 115011
rect 146960 114931 146970 115011
rect 147280 114931 147290 115011
rect 149020 114931 149030 115011
rect 149340 114931 149350 115011
rect 149660 114931 149670 115011
rect 152440 114931 152450 115011
rect 152760 114931 152770 115011
rect 153080 114931 153090 115011
rect 153400 114931 153410 115011
rect 153720 114931 153730 115011
rect 154040 114931 154050 115011
rect 154360 114931 154370 115011
rect 154680 114931 154690 115011
rect 155000 114931 155010 115011
rect 155320 114931 155330 115011
rect 155640 114931 155650 115011
rect 155960 114931 155970 115011
rect 156280 114931 156290 115011
rect 156600 114931 156610 115011
rect 156920 114931 156930 115011
rect 157240 114931 157250 115011
rect 157560 114931 157570 115011
rect 157880 114931 157890 115011
rect 158200 114931 158210 115011
rect 158520 114931 158530 115011
rect 158840 114931 158850 115011
rect 159160 114931 159170 115011
rect 159480 114931 159490 115011
rect 163750 114981 163830 114991
rect 164070 114981 164150 114991
rect 164390 114981 164470 114991
rect 164710 114981 164790 114991
rect 165030 114981 165110 114991
rect 165350 114981 165430 114991
rect 165670 114981 165750 114991
rect 165990 114981 166070 114991
rect 166310 114981 166390 114991
rect 166630 114981 166710 114991
rect 166950 114981 167030 114991
rect 167270 114981 167350 114991
rect 167590 114981 167670 114991
rect 167910 114981 167990 114991
rect 168230 114981 168310 114991
rect 168550 114981 168630 114991
rect 168870 114981 168950 114991
rect 169190 114981 169270 114991
rect 169510 114981 169590 114991
rect 169830 114981 169910 114991
rect 170150 114981 170230 114991
rect 170470 114981 170550 114991
rect 170790 114981 170870 114991
rect 163830 114901 163840 114981
rect 164150 114901 164160 114981
rect 164470 114901 164480 114981
rect 164790 114901 164800 114981
rect 165110 114901 165120 114981
rect 165430 114901 165440 114981
rect 165750 114901 165760 114981
rect 166070 114901 166080 114981
rect 166390 114901 166400 114981
rect 166710 114901 166720 114981
rect 167030 114901 167040 114981
rect 167350 114901 167360 114981
rect 167670 114901 167680 114981
rect 167990 114901 168000 114981
rect 168310 114901 168320 114981
rect 168630 114901 168640 114981
rect 168950 114901 168960 114981
rect 169270 114901 169280 114981
rect 169590 114901 169600 114981
rect 169910 114901 169920 114981
rect 170230 114901 170240 114981
rect 170550 114901 170560 114981
rect 170870 114901 170880 114981
rect 30360 114860 30440 114870
rect 30680 114860 30760 114870
rect 31000 114860 31080 114870
rect 31320 114860 31400 114870
rect 31640 114860 31720 114870
rect 31960 114860 32040 114870
rect 32280 114860 32360 114870
rect 32600 114860 32680 114870
rect 32920 114860 33000 114870
rect 33240 114860 33320 114870
rect 33560 114860 33640 114870
rect 33880 114860 33960 114870
rect 34200 114860 34280 114870
rect 34520 114860 34600 114870
rect 34840 114860 34920 114870
rect 35160 114860 35240 114870
rect 35480 114860 35560 114870
rect 35800 114860 35880 114870
rect 36120 114860 36200 114870
rect 36440 114860 36520 114870
rect 36760 114860 36840 114870
rect 37080 114860 37160 114870
rect 37400 114860 37480 114870
rect 37720 114860 37800 114870
rect 40180 114860 40260 114870
rect 40500 114860 40580 114870
rect 40820 114860 40900 114870
rect 41140 114860 41220 114870
rect 42560 114860 42640 114870
rect 42880 114860 42960 114870
rect 43200 114860 43280 114870
rect 43520 114860 43600 114870
rect 18970 114830 19050 114840
rect 19290 114830 19370 114840
rect 19610 114830 19690 114840
rect 19930 114830 20010 114840
rect 20250 114830 20330 114840
rect 20570 114830 20650 114840
rect 20890 114830 20970 114840
rect 21210 114830 21290 114840
rect 21530 114830 21610 114840
rect 21850 114830 21930 114840
rect 22170 114830 22250 114840
rect 22490 114830 22570 114840
rect 22810 114830 22890 114840
rect 23130 114830 23210 114840
rect 23450 114830 23530 114840
rect 23770 114830 23850 114840
rect 24090 114830 24170 114840
rect 24410 114830 24490 114840
rect 24730 114830 24810 114840
rect 25050 114830 25130 114840
rect 25370 114830 25450 114840
rect 25690 114830 25770 114840
rect 26010 114830 26090 114840
rect 26330 114830 26410 114840
rect 19050 114750 19060 114830
rect 19370 114750 19380 114830
rect 19690 114750 19700 114830
rect 20010 114750 20020 114830
rect 20330 114750 20340 114830
rect 20650 114750 20660 114830
rect 20970 114750 20980 114830
rect 21290 114750 21300 114830
rect 21610 114750 21620 114830
rect 21930 114750 21940 114830
rect 22250 114750 22260 114830
rect 22570 114750 22580 114830
rect 22890 114750 22900 114830
rect 23210 114750 23220 114830
rect 23530 114750 23540 114830
rect 23850 114750 23860 114830
rect 24170 114750 24180 114830
rect 24490 114750 24500 114830
rect 24810 114750 24820 114830
rect 25130 114750 25140 114830
rect 25450 114750 25460 114830
rect 25770 114750 25780 114830
rect 26090 114750 26100 114830
rect 26410 114750 26420 114830
rect 30440 114780 30450 114860
rect 30760 114780 30770 114860
rect 31080 114780 31090 114860
rect 31400 114780 31410 114860
rect 31720 114780 31730 114860
rect 32040 114780 32050 114860
rect 32360 114780 32370 114860
rect 32680 114780 32690 114860
rect 33000 114780 33010 114860
rect 33320 114780 33330 114860
rect 33640 114780 33650 114860
rect 33960 114780 33970 114860
rect 34280 114780 34290 114860
rect 34600 114780 34610 114860
rect 34920 114780 34930 114860
rect 35240 114780 35250 114860
rect 35560 114780 35570 114860
rect 35880 114780 35890 114860
rect 36200 114780 36210 114860
rect 36520 114780 36530 114860
rect 36840 114780 36850 114860
rect 37160 114780 37170 114860
rect 37480 114780 37490 114860
rect 37800 114780 37810 114860
rect 40260 114780 40270 114860
rect 40580 114780 40590 114860
rect 40900 114780 40910 114860
rect 41220 114780 41230 114860
rect 42640 114780 42650 114860
rect 42960 114780 42970 114860
rect 43280 114780 43290 114860
rect 43600 114780 43610 114860
rect 146400 114851 146480 114861
rect 146720 114851 146800 114861
rect 147040 114851 147120 114861
rect 147360 114851 147440 114861
rect 148780 114851 148860 114861
rect 149100 114851 149180 114861
rect 149420 114851 149500 114861
rect 149740 114851 149820 114861
rect 152200 114851 152280 114861
rect 152520 114851 152600 114861
rect 152840 114851 152920 114861
rect 153160 114851 153240 114861
rect 153480 114851 153560 114861
rect 153800 114851 153880 114861
rect 154120 114851 154200 114861
rect 154440 114851 154520 114861
rect 154760 114851 154840 114861
rect 155080 114851 155160 114861
rect 155400 114851 155480 114861
rect 155720 114851 155800 114861
rect 156040 114851 156120 114861
rect 156360 114851 156440 114861
rect 156680 114851 156760 114861
rect 157000 114851 157080 114861
rect 157320 114851 157400 114861
rect 157640 114851 157720 114861
rect 157960 114851 158040 114861
rect 158280 114851 158360 114861
rect 158600 114851 158680 114861
rect 158920 114851 159000 114861
rect 159240 114851 159320 114861
rect 159560 114851 159640 114861
rect 146480 114771 146490 114851
rect 146800 114771 146810 114851
rect 147120 114771 147130 114851
rect 147440 114771 147450 114851
rect 148860 114771 148870 114851
rect 149180 114771 149190 114851
rect 149500 114771 149510 114851
rect 149820 114771 149830 114851
rect 152280 114771 152290 114851
rect 152600 114771 152610 114851
rect 152920 114771 152930 114851
rect 153240 114771 153250 114851
rect 153560 114771 153570 114851
rect 153880 114771 153890 114851
rect 154200 114771 154210 114851
rect 154520 114771 154530 114851
rect 154840 114771 154850 114851
rect 155160 114771 155170 114851
rect 155480 114771 155490 114851
rect 155800 114771 155810 114851
rect 156120 114771 156130 114851
rect 156440 114771 156450 114851
rect 156760 114771 156770 114851
rect 157080 114771 157090 114851
rect 157400 114771 157410 114851
rect 157720 114771 157730 114851
rect 158040 114771 158050 114851
rect 158360 114771 158370 114851
rect 158680 114771 158690 114851
rect 159000 114771 159010 114851
rect 159320 114771 159330 114851
rect 159640 114771 159650 114851
rect 163590 114821 163670 114831
rect 163910 114821 163990 114831
rect 164230 114821 164310 114831
rect 164550 114821 164630 114831
rect 164870 114821 164950 114831
rect 165190 114821 165270 114831
rect 165510 114821 165590 114831
rect 165830 114821 165910 114831
rect 166150 114821 166230 114831
rect 166470 114821 166550 114831
rect 166790 114821 166870 114831
rect 167110 114821 167190 114831
rect 167430 114821 167510 114831
rect 167750 114821 167830 114831
rect 168070 114821 168150 114831
rect 168390 114821 168470 114831
rect 168710 114821 168790 114831
rect 169030 114821 169110 114831
rect 169350 114821 169430 114831
rect 169670 114821 169750 114831
rect 169990 114821 170070 114831
rect 170310 114821 170390 114831
rect 170630 114821 170710 114831
rect 170950 114821 171030 114831
rect 163670 114741 163680 114821
rect 163990 114741 164000 114821
rect 164310 114741 164320 114821
rect 164630 114741 164640 114821
rect 164950 114741 164960 114821
rect 165270 114741 165280 114821
rect 165590 114741 165600 114821
rect 165910 114741 165920 114821
rect 166230 114741 166240 114821
rect 166550 114741 166560 114821
rect 166870 114741 166880 114821
rect 167190 114741 167200 114821
rect 167510 114741 167520 114821
rect 167830 114741 167840 114821
rect 168150 114741 168160 114821
rect 168470 114741 168480 114821
rect 168790 114741 168800 114821
rect 169110 114741 169120 114821
rect 169430 114741 169440 114821
rect 169750 114741 169760 114821
rect 170070 114741 170080 114821
rect 170390 114741 170400 114821
rect 170710 114741 170720 114821
rect 171030 114741 171040 114821
rect 30520 114700 30600 114710
rect 30840 114700 30920 114710
rect 31160 114700 31240 114710
rect 31480 114700 31560 114710
rect 31800 114700 31880 114710
rect 32120 114700 32200 114710
rect 32440 114700 32520 114710
rect 32760 114700 32840 114710
rect 33080 114700 33160 114710
rect 33400 114700 33480 114710
rect 33720 114700 33800 114710
rect 34040 114700 34120 114710
rect 34360 114700 34440 114710
rect 34680 114700 34760 114710
rect 35000 114700 35080 114710
rect 35320 114700 35400 114710
rect 35640 114700 35720 114710
rect 35960 114700 36040 114710
rect 36280 114700 36360 114710
rect 36600 114700 36680 114710
rect 36920 114700 37000 114710
rect 37240 114700 37320 114710
rect 37560 114700 37640 114710
rect 40340 114700 40420 114710
rect 40660 114700 40740 114710
rect 40980 114700 41060 114710
rect 42720 114700 42800 114710
rect 43040 114700 43120 114710
rect 43360 114700 43440 114710
rect 19130 114670 19210 114680
rect 19450 114670 19530 114680
rect 19770 114670 19850 114680
rect 20090 114670 20170 114680
rect 20410 114670 20490 114680
rect 20730 114670 20810 114680
rect 21050 114670 21130 114680
rect 21370 114670 21450 114680
rect 21690 114670 21770 114680
rect 22010 114670 22090 114680
rect 22330 114670 22410 114680
rect 22650 114670 22730 114680
rect 22970 114670 23050 114680
rect 23290 114670 23370 114680
rect 23610 114670 23690 114680
rect 23930 114670 24010 114680
rect 24250 114670 24330 114680
rect 24570 114670 24650 114680
rect 24890 114670 24970 114680
rect 25210 114670 25290 114680
rect 25530 114670 25610 114680
rect 25850 114670 25930 114680
rect 26170 114670 26250 114680
rect 19210 114590 19220 114670
rect 19530 114590 19540 114670
rect 19850 114590 19860 114670
rect 20170 114590 20180 114670
rect 20490 114590 20500 114670
rect 20810 114590 20820 114670
rect 21130 114590 21140 114670
rect 21450 114590 21460 114670
rect 21770 114590 21780 114670
rect 22090 114590 22100 114670
rect 22410 114590 22420 114670
rect 22730 114590 22740 114670
rect 23050 114590 23060 114670
rect 23370 114590 23380 114670
rect 23690 114590 23700 114670
rect 24010 114590 24020 114670
rect 24330 114590 24340 114670
rect 24650 114590 24660 114670
rect 24970 114590 24980 114670
rect 25290 114590 25300 114670
rect 25610 114590 25620 114670
rect 25930 114590 25940 114670
rect 26250 114590 26260 114670
rect 30600 114620 30610 114700
rect 30920 114620 30930 114700
rect 31240 114620 31250 114700
rect 31560 114620 31570 114700
rect 31880 114620 31890 114700
rect 32200 114620 32210 114700
rect 32520 114620 32530 114700
rect 32840 114620 32850 114700
rect 33160 114620 33170 114700
rect 33480 114620 33490 114700
rect 33800 114620 33810 114700
rect 34120 114620 34130 114700
rect 34440 114620 34450 114700
rect 34760 114620 34770 114700
rect 35080 114620 35090 114700
rect 35400 114620 35410 114700
rect 35720 114620 35730 114700
rect 36040 114620 36050 114700
rect 36360 114620 36370 114700
rect 36680 114620 36690 114700
rect 37000 114620 37010 114700
rect 37320 114620 37330 114700
rect 37640 114620 37650 114700
rect 40420 114620 40430 114700
rect 40740 114620 40750 114700
rect 41060 114620 41070 114700
rect 42800 114620 42810 114700
rect 43120 114620 43130 114700
rect 43440 114620 43450 114700
rect 146560 114691 146640 114701
rect 146880 114691 146960 114701
rect 147200 114691 147280 114701
rect 148940 114691 149020 114701
rect 149260 114691 149340 114701
rect 149580 114691 149660 114701
rect 152360 114691 152440 114701
rect 152680 114691 152760 114701
rect 153000 114691 153080 114701
rect 153320 114691 153400 114701
rect 153640 114691 153720 114701
rect 153960 114691 154040 114701
rect 154280 114691 154360 114701
rect 154600 114691 154680 114701
rect 154920 114691 155000 114701
rect 155240 114691 155320 114701
rect 155560 114691 155640 114701
rect 155880 114691 155960 114701
rect 156200 114691 156280 114701
rect 156520 114691 156600 114701
rect 156840 114691 156920 114701
rect 157160 114691 157240 114701
rect 157480 114691 157560 114701
rect 157800 114691 157880 114701
rect 158120 114691 158200 114701
rect 158440 114691 158520 114701
rect 158760 114691 158840 114701
rect 159080 114691 159160 114701
rect 159400 114691 159480 114701
rect 146640 114611 146650 114691
rect 146960 114611 146970 114691
rect 147280 114611 147290 114691
rect 149020 114611 149030 114691
rect 149340 114611 149350 114691
rect 149660 114611 149670 114691
rect 152440 114611 152450 114691
rect 152760 114611 152770 114691
rect 153080 114611 153090 114691
rect 153400 114611 153410 114691
rect 153720 114611 153730 114691
rect 154040 114611 154050 114691
rect 154360 114611 154370 114691
rect 154680 114611 154690 114691
rect 155000 114611 155010 114691
rect 155320 114611 155330 114691
rect 155640 114611 155650 114691
rect 155960 114611 155970 114691
rect 156280 114611 156290 114691
rect 156600 114611 156610 114691
rect 156920 114611 156930 114691
rect 157240 114611 157250 114691
rect 157560 114611 157570 114691
rect 157880 114611 157890 114691
rect 158200 114611 158210 114691
rect 158520 114611 158530 114691
rect 158840 114611 158850 114691
rect 159160 114611 159170 114691
rect 159480 114611 159490 114691
rect 163750 114661 163830 114671
rect 164070 114661 164150 114671
rect 164390 114661 164470 114671
rect 164710 114661 164790 114671
rect 165030 114661 165110 114671
rect 165350 114661 165430 114671
rect 165670 114661 165750 114671
rect 165990 114661 166070 114671
rect 166310 114661 166390 114671
rect 166630 114661 166710 114671
rect 166950 114661 167030 114671
rect 167270 114661 167350 114671
rect 167590 114661 167670 114671
rect 167910 114661 167990 114671
rect 168230 114661 168310 114671
rect 168550 114661 168630 114671
rect 168870 114661 168950 114671
rect 169190 114661 169270 114671
rect 169510 114661 169590 114671
rect 169830 114661 169910 114671
rect 170150 114661 170230 114671
rect 170470 114661 170550 114671
rect 170790 114661 170870 114671
rect 163830 114581 163840 114661
rect 164150 114581 164160 114661
rect 164470 114581 164480 114661
rect 164790 114581 164800 114661
rect 165110 114581 165120 114661
rect 165430 114581 165440 114661
rect 165750 114581 165760 114661
rect 166070 114581 166080 114661
rect 166390 114581 166400 114661
rect 166710 114581 166720 114661
rect 167030 114581 167040 114661
rect 167350 114581 167360 114661
rect 167670 114581 167680 114661
rect 167990 114581 168000 114661
rect 168310 114581 168320 114661
rect 168630 114581 168640 114661
rect 168950 114581 168960 114661
rect 169270 114581 169280 114661
rect 169590 114581 169600 114661
rect 169910 114581 169920 114661
rect 170230 114581 170240 114661
rect 170550 114581 170560 114661
rect 170870 114581 170880 114661
rect 18980 114440 19060 114450
rect 19160 114440 19240 114450
rect 19340 114440 19420 114450
rect 19520 114440 19600 114450
rect 19700 114440 19780 114450
rect 19880 114440 19960 114450
rect 20060 114440 20140 114450
rect 20240 114440 20320 114450
rect 20420 114440 20500 114450
rect 20600 114440 20680 114450
rect 20780 114440 20860 114450
rect 20960 114440 21040 114450
rect 21140 114440 21220 114450
rect 21320 114440 21400 114450
rect 21500 114440 21580 114450
rect 21680 114440 21760 114450
rect 21860 114440 21940 114450
rect 22040 114440 22120 114450
rect 22220 114440 22300 114450
rect 22400 114440 22480 114450
rect 22580 114440 22660 114450
rect 22760 114440 22840 114450
rect 22940 114440 23020 114450
rect 23120 114440 23200 114450
rect 23300 114440 23380 114450
rect 23480 114440 23560 114450
rect 23660 114440 23740 114450
rect 23840 114440 23920 114450
rect 24020 114440 24100 114450
rect 24200 114440 24280 114450
rect 24380 114440 24460 114450
rect 24560 114440 24640 114450
rect 24740 114440 24820 114450
rect 24920 114440 25000 114450
rect 25100 114440 25180 114450
rect 25280 114440 25360 114450
rect 25460 114440 25540 114450
rect 25640 114440 25720 114450
rect 25820 114440 25900 114450
rect 26000 114440 26080 114450
rect 26180 114440 26260 114450
rect 26360 114440 26440 114450
rect 26540 114440 26620 114450
rect 30280 114440 30360 114450
rect 30460 114440 30540 114450
rect 30640 114440 30720 114450
rect 30820 114440 30900 114450
rect 31000 114440 31080 114450
rect 31180 114440 31260 114450
rect 31360 114440 31440 114450
rect 31540 114440 31620 114450
rect 31720 114440 31800 114450
rect 31900 114440 31980 114450
rect 32080 114440 32160 114450
rect 32260 114440 32340 114450
rect 32440 114440 32520 114450
rect 32620 114440 32700 114450
rect 32800 114440 32880 114450
rect 32980 114440 33060 114450
rect 33160 114440 33240 114450
rect 33340 114440 33420 114450
rect 33520 114440 33600 114450
rect 33700 114440 33780 114450
rect 33880 114440 33960 114450
rect 34060 114440 34140 114450
rect 34240 114440 34320 114450
rect 34420 114440 34500 114450
rect 34600 114440 34680 114450
rect 34780 114440 34860 114450
rect 34960 114440 35040 114450
rect 35140 114440 35220 114450
rect 35320 114440 35400 114450
rect 35500 114440 35580 114450
rect 35680 114440 35760 114450
rect 35860 114440 35940 114450
rect 36040 114440 36120 114450
rect 36220 114440 36300 114450
rect 36400 114440 36480 114450
rect 36580 114440 36660 114450
rect 36760 114440 36840 114450
rect 36940 114440 37020 114450
rect 37120 114440 37200 114450
rect 37300 114440 37380 114450
rect 37480 114440 37560 114450
rect 37660 114440 37740 114450
rect 37840 114440 37920 114450
rect 40060 114440 40140 114450
rect 40200 114440 40280 114450
rect 40340 114440 40420 114450
rect 40480 114440 40560 114450
rect 40620 114440 40700 114450
rect 40760 114440 40840 114450
rect 40900 114440 40980 114450
rect 41040 114440 41120 114450
rect 41180 114440 41260 114450
rect 41320 114440 41400 114450
rect 42360 114440 42440 114450
rect 42500 114440 42580 114450
rect 42640 114440 42720 114450
rect 42780 114440 42860 114450
rect 42920 114440 43000 114450
rect 43060 114440 43140 114450
rect 43200 114440 43280 114450
rect 43340 114440 43420 114450
rect 43480 114440 43560 114450
rect 43620 114440 43700 114450
rect 146300 114440 146380 114450
rect 146440 114440 146520 114450
rect 146580 114440 146660 114450
rect 146720 114440 146800 114450
rect 146860 114440 146940 114450
rect 147000 114440 147080 114450
rect 147140 114440 147220 114450
rect 147280 114440 147360 114450
rect 147420 114440 147500 114450
rect 147560 114440 147640 114450
rect 19060 114360 19070 114440
rect 19240 114360 19250 114440
rect 19420 114360 19430 114440
rect 19600 114360 19610 114440
rect 19780 114360 19790 114440
rect 19960 114360 19970 114440
rect 20140 114360 20150 114440
rect 20320 114360 20330 114440
rect 20500 114360 20510 114440
rect 20680 114360 20690 114440
rect 20860 114360 20870 114440
rect 21040 114360 21050 114440
rect 21220 114360 21230 114440
rect 21400 114360 21410 114440
rect 21580 114360 21590 114440
rect 21760 114360 21770 114440
rect 21940 114360 21950 114440
rect 22120 114360 22130 114440
rect 22300 114360 22310 114440
rect 22480 114360 22490 114440
rect 22660 114360 22670 114440
rect 22840 114360 22850 114440
rect 23020 114360 23030 114440
rect 23200 114360 23210 114440
rect 23380 114360 23390 114440
rect 23560 114360 23570 114440
rect 23740 114360 23750 114440
rect 23920 114360 23930 114440
rect 24100 114360 24110 114440
rect 24280 114360 24290 114440
rect 24460 114360 24470 114440
rect 24640 114360 24650 114440
rect 24820 114360 24830 114440
rect 25000 114360 25010 114440
rect 25180 114360 25190 114440
rect 25360 114360 25370 114440
rect 25540 114360 25550 114440
rect 25720 114360 25730 114440
rect 25900 114360 25910 114440
rect 26080 114360 26090 114440
rect 26260 114360 26270 114440
rect 26440 114360 26450 114440
rect 26620 114360 26630 114440
rect 30360 114360 30370 114440
rect 30540 114360 30550 114440
rect 30720 114360 30730 114440
rect 30900 114360 30910 114440
rect 31080 114360 31090 114440
rect 31260 114360 31270 114440
rect 31440 114360 31450 114440
rect 31620 114360 31630 114440
rect 31800 114360 31810 114440
rect 31980 114360 31990 114440
rect 32160 114360 32170 114440
rect 32340 114360 32350 114440
rect 32520 114360 32530 114440
rect 32700 114360 32710 114440
rect 32880 114360 32890 114440
rect 33060 114360 33070 114440
rect 33240 114360 33250 114440
rect 33420 114360 33430 114440
rect 33600 114360 33610 114440
rect 33780 114360 33790 114440
rect 33960 114360 33970 114440
rect 34140 114360 34150 114440
rect 34320 114360 34330 114440
rect 34500 114360 34510 114440
rect 34680 114360 34690 114440
rect 34860 114360 34870 114440
rect 35040 114360 35050 114440
rect 35220 114360 35230 114440
rect 35400 114360 35410 114440
rect 35580 114360 35590 114440
rect 35760 114360 35770 114440
rect 35940 114360 35950 114440
rect 36120 114360 36130 114440
rect 36300 114360 36310 114440
rect 36480 114360 36490 114440
rect 36660 114360 36670 114440
rect 36840 114360 36850 114440
rect 37020 114360 37030 114440
rect 37200 114360 37210 114440
rect 37380 114360 37390 114440
rect 37560 114360 37570 114440
rect 37740 114360 37750 114440
rect 37920 114360 37930 114440
rect 40140 114360 40150 114440
rect 40280 114360 40290 114440
rect 40420 114360 40430 114440
rect 40560 114360 40570 114440
rect 40700 114360 40710 114440
rect 40840 114360 40850 114440
rect 40980 114360 40990 114440
rect 41120 114360 41130 114440
rect 41260 114360 41270 114440
rect 41400 114360 41410 114440
rect 42440 114360 42450 114440
rect 42580 114360 42590 114440
rect 42720 114360 42730 114440
rect 42860 114360 42870 114440
rect 43000 114360 43010 114440
rect 43140 114360 43150 114440
rect 43280 114360 43290 114440
rect 43420 114360 43430 114440
rect 43560 114360 43570 114440
rect 43700 114360 43710 114440
rect 146380 114360 146390 114440
rect 146520 114360 146530 114440
rect 146660 114360 146670 114440
rect 146800 114360 146810 114440
rect 146940 114360 146950 114440
rect 147080 114360 147090 114440
rect 147220 114360 147230 114440
rect 147360 114360 147370 114440
rect 147500 114360 147510 114440
rect 147640 114360 147650 114440
rect 28850 114315 28930 114325
rect 29010 114315 29090 114325
rect 29170 114315 29250 114325
rect 29330 114315 29410 114325
rect 29490 114315 29570 114325
rect 18980 114290 19060 114300
rect 19160 114290 19240 114300
rect 19340 114290 19420 114300
rect 19520 114290 19600 114300
rect 19700 114290 19780 114300
rect 19880 114290 19960 114300
rect 20060 114290 20140 114300
rect 20240 114290 20320 114300
rect 20420 114290 20500 114300
rect 20600 114290 20680 114300
rect 20780 114290 20860 114300
rect 20960 114290 21040 114300
rect 21140 114290 21220 114300
rect 21320 114290 21400 114300
rect 21500 114290 21580 114300
rect 21680 114290 21760 114300
rect 21860 114290 21940 114300
rect 22040 114290 22120 114300
rect 22220 114290 22300 114300
rect 22400 114290 22480 114300
rect 22580 114290 22660 114300
rect 22760 114290 22840 114300
rect 22940 114290 23020 114300
rect 23120 114290 23200 114300
rect 23300 114290 23380 114300
rect 23480 114290 23560 114300
rect 23660 114290 23740 114300
rect 23840 114290 23920 114300
rect 24020 114290 24100 114300
rect 24200 114290 24280 114300
rect 24380 114290 24460 114300
rect 24560 114290 24640 114300
rect 24740 114290 24820 114300
rect 24920 114290 25000 114300
rect 25100 114290 25180 114300
rect 25280 114290 25360 114300
rect 25460 114290 25540 114300
rect 25640 114290 25720 114300
rect 25820 114290 25900 114300
rect 26000 114290 26080 114300
rect 26180 114290 26260 114300
rect 26360 114290 26440 114300
rect 26540 114290 26620 114300
rect 19060 114210 19070 114290
rect 19240 114210 19250 114290
rect 19420 114210 19430 114290
rect 19600 114210 19610 114290
rect 19780 114210 19790 114290
rect 19960 114210 19970 114290
rect 20140 114210 20150 114290
rect 20320 114210 20330 114290
rect 20500 114210 20510 114290
rect 20680 114210 20690 114290
rect 20860 114210 20870 114290
rect 21040 114210 21050 114290
rect 21220 114210 21230 114290
rect 21400 114210 21410 114290
rect 21580 114210 21590 114290
rect 21760 114210 21770 114290
rect 21940 114210 21950 114290
rect 22120 114210 22130 114290
rect 22300 114210 22310 114290
rect 22480 114210 22490 114290
rect 22660 114210 22670 114290
rect 22840 114210 22850 114290
rect 23020 114210 23030 114290
rect 23200 114210 23210 114290
rect 23380 114210 23390 114290
rect 23560 114210 23570 114290
rect 23740 114210 23750 114290
rect 23920 114210 23930 114290
rect 24100 114210 24110 114290
rect 24280 114210 24290 114290
rect 24460 114210 24470 114290
rect 24640 114210 24650 114290
rect 24820 114210 24830 114290
rect 25000 114210 25010 114290
rect 25180 114210 25190 114290
rect 25360 114210 25370 114290
rect 25540 114210 25550 114290
rect 25720 114210 25730 114290
rect 25900 114210 25910 114290
rect 26080 114210 26090 114290
rect 26260 114210 26270 114290
rect 26440 114210 26450 114290
rect 26620 114210 26630 114290
rect 28930 114235 28940 114315
rect 29010 114235 29020 114315
rect 29090 114235 29100 114315
rect 29170 114235 29180 114315
rect 29250 114235 29260 114315
rect 29330 114235 29340 114315
rect 29410 114235 29420 114315
rect 29490 114235 29500 114315
rect 29570 114235 29580 114315
rect 148340 114300 150000 114570
rect 152080 114440 152160 114450
rect 152260 114440 152340 114450
rect 152440 114440 152520 114450
rect 152620 114440 152700 114450
rect 152800 114440 152880 114450
rect 152980 114440 153060 114450
rect 153160 114440 153240 114450
rect 153340 114440 153420 114450
rect 153520 114440 153600 114450
rect 153700 114440 153780 114450
rect 153880 114440 153960 114450
rect 154060 114440 154140 114450
rect 154240 114440 154320 114450
rect 154420 114440 154500 114450
rect 154600 114440 154680 114450
rect 154780 114440 154860 114450
rect 154960 114440 155040 114450
rect 155140 114440 155220 114450
rect 155320 114440 155400 114450
rect 155500 114440 155580 114450
rect 155680 114440 155760 114450
rect 155860 114440 155940 114450
rect 156040 114440 156120 114450
rect 156220 114440 156300 114450
rect 156400 114440 156480 114450
rect 156580 114440 156660 114450
rect 156760 114440 156840 114450
rect 156940 114440 157020 114450
rect 157120 114440 157200 114450
rect 157300 114440 157380 114450
rect 157480 114440 157560 114450
rect 157660 114440 157740 114450
rect 157840 114440 157920 114450
rect 158020 114440 158100 114450
rect 158200 114440 158280 114450
rect 158380 114440 158460 114450
rect 158560 114440 158640 114450
rect 158740 114440 158820 114450
rect 158920 114440 159000 114450
rect 159100 114440 159180 114450
rect 159280 114440 159360 114450
rect 159460 114440 159540 114450
rect 159640 114440 159720 114450
rect 163380 114440 163460 114450
rect 163560 114440 163640 114450
rect 163740 114440 163820 114450
rect 163920 114440 164000 114450
rect 164100 114440 164180 114450
rect 164280 114440 164360 114450
rect 164460 114440 164540 114450
rect 164640 114440 164720 114450
rect 164820 114440 164900 114450
rect 165000 114440 165080 114450
rect 165180 114440 165260 114450
rect 165360 114440 165440 114450
rect 165540 114440 165620 114450
rect 165720 114440 165800 114450
rect 165900 114440 165980 114450
rect 166080 114440 166160 114450
rect 166260 114440 166340 114450
rect 166440 114440 166520 114450
rect 166620 114440 166700 114450
rect 166800 114440 166880 114450
rect 166980 114440 167060 114450
rect 167160 114440 167240 114450
rect 167340 114440 167420 114450
rect 167520 114440 167600 114450
rect 167700 114440 167780 114450
rect 167880 114440 167960 114450
rect 168060 114440 168140 114450
rect 168240 114440 168320 114450
rect 168420 114440 168500 114450
rect 168600 114440 168680 114450
rect 168780 114440 168860 114450
rect 168960 114440 169040 114450
rect 169140 114440 169220 114450
rect 169320 114440 169400 114450
rect 169500 114440 169580 114450
rect 169680 114440 169760 114450
rect 169860 114440 169940 114450
rect 170040 114440 170120 114450
rect 170220 114440 170300 114450
rect 170400 114440 170480 114450
rect 170580 114440 170660 114450
rect 170760 114440 170840 114450
rect 170940 114440 171020 114450
rect 152160 114360 152170 114440
rect 152340 114360 152350 114440
rect 152520 114360 152530 114440
rect 152700 114360 152710 114440
rect 152880 114360 152890 114440
rect 153060 114360 153070 114440
rect 153240 114360 153250 114440
rect 153420 114360 153430 114440
rect 153600 114360 153610 114440
rect 153780 114360 153790 114440
rect 153960 114360 153970 114440
rect 154140 114360 154150 114440
rect 154320 114360 154330 114440
rect 154500 114360 154510 114440
rect 154680 114360 154690 114440
rect 154860 114360 154870 114440
rect 155040 114360 155050 114440
rect 155220 114360 155230 114440
rect 155400 114360 155410 114440
rect 155580 114360 155590 114440
rect 155760 114360 155770 114440
rect 155940 114360 155950 114440
rect 156120 114360 156130 114440
rect 156300 114360 156310 114440
rect 156480 114360 156490 114440
rect 156660 114360 156670 114440
rect 156840 114360 156850 114440
rect 157020 114360 157030 114440
rect 157200 114360 157210 114440
rect 157380 114360 157390 114440
rect 157560 114360 157570 114440
rect 157740 114360 157750 114440
rect 157920 114360 157930 114440
rect 158100 114360 158110 114440
rect 158280 114360 158290 114440
rect 158460 114360 158470 114440
rect 158640 114360 158650 114440
rect 158820 114360 158830 114440
rect 159000 114360 159010 114440
rect 159180 114360 159190 114440
rect 159360 114360 159370 114440
rect 159540 114360 159550 114440
rect 159720 114360 159730 114440
rect 163460 114360 163470 114440
rect 163640 114360 163650 114440
rect 163820 114360 163830 114440
rect 164000 114360 164010 114440
rect 164180 114360 164190 114440
rect 164360 114360 164370 114440
rect 164540 114360 164550 114440
rect 164720 114360 164730 114440
rect 164900 114360 164910 114440
rect 165080 114360 165090 114440
rect 165260 114360 165270 114440
rect 165440 114360 165450 114440
rect 165620 114360 165630 114440
rect 165800 114360 165810 114440
rect 165980 114360 165990 114440
rect 166160 114360 166170 114440
rect 166340 114360 166350 114440
rect 166520 114360 166530 114440
rect 166700 114360 166710 114440
rect 166880 114360 166890 114440
rect 167060 114360 167070 114440
rect 167240 114360 167250 114440
rect 167420 114360 167430 114440
rect 167600 114360 167610 114440
rect 167780 114360 167790 114440
rect 167960 114360 167970 114440
rect 168140 114360 168150 114440
rect 168320 114360 168330 114440
rect 168500 114360 168510 114440
rect 168680 114360 168690 114440
rect 168860 114360 168870 114440
rect 169040 114360 169050 114440
rect 169220 114360 169230 114440
rect 169400 114360 169410 114440
rect 169580 114360 169590 114440
rect 169760 114360 169770 114440
rect 169940 114360 169950 114440
rect 170120 114360 170130 114440
rect 170300 114360 170310 114440
rect 170480 114360 170490 114440
rect 170660 114360 170670 114440
rect 170840 114360 170850 114440
rect 171020 114360 171030 114440
rect 161885 114345 161965 114355
rect 162065 114345 162145 114355
rect 162245 114345 162325 114355
rect 162425 114345 162505 114355
rect 162605 114345 162685 114355
rect 30280 114290 30360 114300
rect 30460 114290 30540 114300
rect 30640 114290 30720 114300
rect 30820 114290 30900 114300
rect 31000 114290 31080 114300
rect 31180 114290 31260 114300
rect 31360 114290 31440 114300
rect 31540 114290 31620 114300
rect 31720 114290 31800 114300
rect 31900 114290 31980 114300
rect 32080 114290 32160 114300
rect 32260 114290 32340 114300
rect 32440 114290 32520 114300
rect 32620 114290 32700 114300
rect 32800 114290 32880 114300
rect 32980 114290 33060 114300
rect 33160 114290 33240 114300
rect 33340 114290 33420 114300
rect 33520 114290 33600 114300
rect 33700 114290 33780 114300
rect 33880 114290 33960 114300
rect 34060 114290 34140 114300
rect 34240 114290 34320 114300
rect 34420 114290 34500 114300
rect 34600 114290 34680 114300
rect 34780 114290 34860 114300
rect 34960 114290 35040 114300
rect 35140 114290 35220 114300
rect 35320 114290 35400 114300
rect 35500 114290 35580 114300
rect 35680 114290 35760 114300
rect 35860 114290 35940 114300
rect 36040 114290 36120 114300
rect 36220 114290 36300 114300
rect 36400 114290 36480 114300
rect 36580 114290 36660 114300
rect 36760 114290 36840 114300
rect 36940 114290 37020 114300
rect 37120 114290 37200 114300
rect 37300 114290 37380 114300
rect 37480 114290 37560 114300
rect 37660 114290 37740 114300
rect 37840 114290 37920 114300
rect 30360 114210 30370 114290
rect 30540 114210 30550 114290
rect 30720 114210 30730 114290
rect 30900 114210 30910 114290
rect 31080 114210 31090 114290
rect 31260 114210 31270 114290
rect 31440 114210 31450 114290
rect 31620 114210 31630 114290
rect 31800 114210 31810 114290
rect 31980 114210 31990 114290
rect 32160 114210 32170 114290
rect 32340 114210 32350 114290
rect 32520 114210 32530 114290
rect 32700 114210 32710 114290
rect 32880 114210 32890 114290
rect 33060 114210 33070 114290
rect 33240 114210 33250 114290
rect 33420 114210 33430 114290
rect 33600 114210 33610 114290
rect 33780 114210 33790 114290
rect 33960 114210 33970 114290
rect 34140 114210 34150 114290
rect 34320 114210 34330 114290
rect 34500 114210 34510 114290
rect 34680 114210 34690 114290
rect 34860 114210 34870 114290
rect 35040 114210 35050 114290
rect 35220 114210 35230 114290
rect 35400 114210 35410 114290
rect 35580 114210 35590 114290
rect 35760 114210 35770 114290
rect 35940 114210 35950 114290
rect 36120 114210 36130 114290
rect 36300 114210 36310 114290
rect 36480 114210 36490 114290
rect 36660 114210 36670 114290
rect 36840 114210 36850 114290
rect 37020 114210 37030 114290
rect 37200 114210 37210 114290
rect 37380 114210 37390 114290
rect 37560 114210 37570 114290
rect 37740 114210 37750 114290
rect 37920 114210 37930 114290
rect 40060 114190 40120 114220
rect 41540 114190 41600 114220
rect 42360 114190 42420 114220
rect 43840 114190 43900 114220
rect 146100 114150 146160 114180
rect 147580 114150 147640 114180
rect 148400 114150 148460 114180
rect 40060 114070 40120 114100
rect 41540 114070 41600 114100
rect 42360 114070 42420 114100
rect 43840 114070 43900 114100
rect 146100 114030 146160 114060
rect 147580 114030 147640 114060
rect 148400 114030 148460 114060
rect 40060 113950 40120 113980
rect 41540 113950 41600 113980
rect 42360 113950 42420 113980
rect 43840 113950 43900 113980
rect 19130 113910 19160 113940
rect 19250 113910 19280 113940
rect 26420 113910 26450 113940
rect 26540 113910 26570 113940
rect 30420 113910 30450 113940
rect 30540 113910 30570 113940
rect 37720 113910 37750 113940
rect 37840 113910 37870 113940
rect 146100 113910 146160 113940
rect 147580 113910 147640 113940
rect 148400 113910 148460 113940
rect 19010 113880 19070 113910
rect 19130 113880 19190 113910
rect 19250 113880 19310 113910
rect 26300 113880 26360 113910
rect 26420 113880 26480 113910
rect 26540 113880 26600 113910
rect 30300 113880 30360 113910
rect 30420 113880 30480 113910
rect 30540 113880 30600 113910
rect 37600 113880 37660 113910
rect 37720 113880 37780 113910
rect 37840 113880 37900 113910
rect 40060 113830 40120 113860
rect 41540 113830 41600 113860
rect 42360 113830 42420 113860
rect 43840 113830 43900 113860
rect 19130 113790 19160 113820
rect 19250 113790 19280 113820
rect 26420 113790 26450 113820
rect 26540 113790 26570 113820
rect 30420 113790 30450 113820
rect 30540 113790 30570 113820
rect 37720 113790 37750 113820
rect 37840 113790 37870 113820
rect 146100 113790 146160 113820
rect 147580 113790 147640 113820
rect 148400 113790 148460 113820
rect 19010 113760 19070 113790
rect 19130 113760 19190 113790
rect 19250 113760 19310 113790
rect 26300 113760 26360 113790
rect 26420 113760 26480 113790
rect 26540 113760 26600 113790
rect 30300 113760 30360 113790
rect 30420 113760 30480 113790
rect 30540 113760 30600 113790
rect 37600 113760 37660 113790
rect 37720 113760 37780 113790
rect 37840 113760 37900 113790
rect 31010 113745 37190 113760
rect 36000 113670 37190 113745
rect 40060 113710 40120 113740
rect 41540 113710 41600 113740
rect 42360 113710 42420 113740
rect 43840 113710 43900 113740
rect 148520 113736 148790 114300
rect 149820 113736 150000 114300
rect 152080 114290 152160 114300
rect 152260 114290 152340 114300
rect 152440 114290 152520 114300
rect 152620 114290 152700 114300
rect 152800 114290 152880 114300
rect 152980 114290 153060 114300
rect 153160 114290 153240 114300
rect 153340 114290 153420 114300
rect 153520 114290 153600 114300
rect 153700 114290 153780 114300
rect 153880 114290 153960 114300
rect 154060 114290 154140 114300
rect 154240 114290 154320 114300
rect 154420 114290 154500 114300
rect 154600 114290 154680 114300
rect 154780 114290 154860 114300
rect 154960 114290 155040 114300
rect 155140 114290 155220 114300
rect 155320 114290 155400 114300
rect 155500 114290 155580 114300
rect 155680 114290 155760 114300
rect 155860 114290 155940 114300
rect 156040 114290 156120 114300
rect 156220 114290 156300 114300
rect 156400 114290 156480 114300
rect 156580 114290 156660 114300
rect 156760 114290 156840 114300
rect 156940 114290 157020 114300
rect 157120 114290 157200 114300
rect 157300 114290 157380 114300
rect 157480 114290 157560 114300
rect 157660 114290 157740 114300
rect 157840 114290 157920 114300
rect 158020 114290 158100 114300
rect 158200 114290 158280 114300
rect 158380 114290 158460 114300
rect 158560 114290 158640 114300
rect 158740 114290 158820 114300
rect 158920 114290 159000 114300
rect 159100 114290 159180 114300
rect 159280 114290 159360 114300
rect 159460 114290 159540 114300
rect 159640 114290 159720 114300
rect 152160 114210 152170 114290
rect 152340 114210 152350 114290
rect 152520 114210 152530 114290
rect 152700 114210 152710 114290
rect 152880 114210 152890 114290
rect 153060 114210 153070 114290
rect 153240 114210 153250 114290
rect 153420 114210 153430 114290
rect 153600 114210 153610 114290
rect 153780 114210 153790 114290
rect 153960 114210 153970 114290
rect 154140 114210 154150 114290
rect 154320 114210 154330 114290
rect 154500 114210 154510 114290
rect 154680 114210 154690 114290
rect 154860 114210 154870 114290
rect 155040 114210 155050 114290
rect 155220 114210 155230 114290
rect 155400 114210 155410 114290
rect 155580 114210 155590 114290
rect 155760 114210 155770 114290
rect 155940 114210 155950 114290
rect 156120 114210 156130 114290
rect 156300 114210 156310 114290
rect 156480 114210 156490 114290
rect 156660 114210 156670 114290
rect 156840 114210 156850 114290
rect 157020 114210 157030 114290
rect 157200 114210 157210 114290
rect 157380 114210 157390 114290
rect 157560 114210 157570 114290
rect 157740 114210 157750 114290
rect 157920 114210 157930 114290
rect 158100 114210 158110 114290
rect 158280 114210 158290 114290
rect 158460 114210 158470 114290
rect 158640 114210 158650 114290
rect 158820 114210 158830 114290
rect 159000 114210 159010 114290
rect 159180 114210 159190 114290
rect 159360 114210 159370 114290
rect 159540 114210 159550 114290
rect 159720 114210 159730 114290
rect 161965 114265 161975 114345
rect 162145 114265 162155 114345
rect 162325 114265 162335 114345
rect 162505 114265 162515 114345
rect 162685 114265 162695 114345
rect 163380 114290 163460 114300
rect 163560 114290 163640 114300
rect 163740 114290 163820 114300
rect 163920 114290 164000 114300
rect 164100 114290 164180 114300
rect 164280 114290 164360 114300
rect 164460 114290 164540 114300
rect 164640 114290 164720 114300
rect 164820 114290 164900 114300
rect 165000 114290 165080 114300
rect 165180 114290 165260 114300
rect 165360 114290 165440 114300
rect 165540 114290 165620 114300
rect 165720 114290 165800 114300
rect 165900 114290 165980 114300
rect 166080 114290 166160 114300
rect 166260 114290 166340 114300
rect 166440 114290 166520 114300
rect 166620 114290 166700 114300
rect 166800 114290 166880 114300
rect 166980 114290 167060 114300
rect 167160 114290 167240 114300
rect 167340 114290 167420 114300
rect 167520 114290 167600 114300
rect 167700 114290 167780 114300
rect 167880 114290 167960 114300
rect 168060 114290 168140 114300
rect 168240 114290 168320 114300
rect 168420 114290 168500 114300
rect 168600 114290 168680 114300
rect 168780 114290 168860 114300
rect 168960 114290 169040 114300
rect 169140 114290 169220 114300
rect 169320 114290 169400 114300
rect 169500 114290 169580 114300
rect 169680 114290 169760 114300
rect 169860 114290 169940 114300
rect 170040 114290 170120 114300
rect 170220 114290 170300 114300
rect 170400 114290 170480 114300
rect 170580 114290 170660 114300
rect 170760 114290 170840 114300
rect 170940 114290 171020 114300
rect 163460 114210 163470 114290
rect 163640 114210 163650 114290
rect 163820 114210 163830 114290
rect 164000 114210 164010 114290
rect 164180 114210 164190 114290
rect 164360 114210 164370 114290
rect 164540 114210 164550 114290
rect 164720 114210 164730 114290
rect 164900 114210 164910 114290
rect 165080 114210 165090 114290
rect 165260 114210 165270 114290
rect 165440 114210 165450 114290
rect 165620 114210 165630 114290
rect 165800 114210 165810 114290
rect 165980 114210 165990 114290
rect 166160 114210 166170 114290
rect 166340 114210 166350 114290
rect 166520 114210 166530 114290
rect 166700 114210 166710 114290
rect 166880 114210 166890 114290
rect 167060 114210 167070 114290
rect 167240 114210 167250 114290
rect 167420 114210 167430 114290
rect 167600 114210 167610 114290
rect 167780 114210 167790 114290
rect 167960 114210 167970 114290
rect 168140 114210 168150 114290
rect 168320 114210 168330 114290
rect 168500 114210 168510 114290
rect 168680 114210 168690 114290
rect 168860 114210 168870 114290
rect 169040 114210 169050 114290
rect 169220 114210 169230 114290
rect 169400 114210 169410 114290
rect 169580 114210 169590 114290
rect 169760 114210 169770 114290
rect 169940 114210 169950 114290
rect 170120 114210 170130 114290
rect 170300 114210 170310 114290
rect 170480 114210 170490 114290
rect 170660 114210 170670 114290
rect 170840 114210 170850 114290
rect 171020 114210 171030 114290
rect 161885 114165 161965 114175
rect 162065 114165 162145 114175
rect 162245 114165 162325 114175
rect 162425 114165 162505 114175
rect 162605 114165 162685 114175
rect 152080 114140 152160 114150
rect 152260 114140 152340 114150
rect 152440 114140 152520 114150
rect 152620 114140 152700 114150
rect 152800 114140 152880 114150
rect 152980 114140 153060 114150
rect 153160 114140 153240 114150
rect 153340 114140 153420 114150
rect 153520 114140 153600 114150
rect 153700 114140 153780 114150
rect 153880 114140 153960 114150
rect 154060 114140 154140 114150
rect 154240 114140 154320 114150
rect 154420 114140 154500 114150
rect 154600 114140 154680 114150
rect 154780 114140 154860 114150
rect 154960 114140 155040 114150
rect 155140 114140 155220 114150
rect 155320 114140 155400 114150
rect 155500 114140 155580 114150
rect 155680 114140 155760 114150
rect 155860 114140 155940 114150
rect 156040 114140 156120 114150
rect 156220 114140 156300 114150
rect 156400 114140 156480 114150
rect 156580 114140 156660 114150
rect 156760 114140 156840 114150
rect 156940 114140 157020 114150
rect 157120 114140 157200 114150
rect 157300 114140 157380 114150
rect 157480 114140 157560 114150
rect 157660 114140 157740 114150
rect 157840 114140 157920 114150
rect 158020 114140 158100 114150
rect 158200 114140 158280 114150
rect 158380 114140 158460 114150
rect 158560 114140 158640 114150
rect 158740 114140 158820 114150
rect 158920 114140 159000 114150
rect 159100 114140 159180 114150
rect 159280 114140 159360 114150
rect 159460 114140 159540 114150
rect 159640 114140 159720 114150
rect 152160 114060 152170 114140
rect 152340 114060 152350 114140
rect 152520 114060 152530 114140
rect 152700 114060 152710 114140
rect 152880 114060 152890 114140
rect 153060 114060 153070 114140
rect 153240 114060 153250 114140
rect 153420 114060 153430 114140
rect 153600 114060 153610 114140
rect 153780 114060 153790 114140
rect 153960 114060 153970 114140
rect 154140 114060 154150 114140
rect 154320 114060 154330 114140
rect 154500 114060 154510 114140
rect 154680 114060 154690 114140
rect 154860 114060 154870 114140
rect 155040 114060 155050 114140
rect 155220 114060 155230 114140
rect 155400 114060 155410 114140
rect 155580 114060 155590 114140
rect 155760 114060 155770 114140
rect 155940 114060 155950 114140
rect 156120 114060 156130 114140
rect 156300 114060 156310 114140
rect 156480 114060 156490 114140
rect 156660 114060 156670 114140
rect 156840 114060 156850 114140
rect 157020 114060 157030 114140
rect 157200 114060 157210 114140
rect 157380 114060 157390 114140
rect 157560 114060 157570 114140
rect 157740 114060 157750 114140
rect 157920 114060 157930 114140
rect 158100 114060 158110 114140
rect 158280 114060 158290 114140
rect 158460 114060 158470 114140
rect 158640 114060 158650 114140
rect 158820 114060 158830 114140
rect 159000 114060 159010 114140
rect 159180 114060 159190 114140
rect 159360 114060 159370 114140
rect 159540 114060 159550 114140
rect 159720 114060 159730 114140
rect 161965 114085 161975 114165
rect 162145 114085 162155 114165
rect 162325 114085 162335 114165
rect 162505 114085 162515 114165
rect 162685 114085 162695 114165
rect 163380 114140 163460 114150
rect 163560 114140 163640 114150
rect 163740 114140 163820 114150
rect 163920 114140 164000 114150
rect 164100 114140 164180 114150
rect 164280 114140 164360 114150
rect 164460 114140 164540 114150
rect 164640 114140 164720 114150
rect 164820 114140 164900 114150
rect 165000 114140 165080 114150
rect 165180 114140 165260 114150
rect 165360 114140 165440 114150
rect 165540 114140 165620 114150
rect 165720 114140 165800 114150
rect 165900 114140 165980 114150
rect 166080 114140 166160 114150
rect 166260 114140 166340 114150
rect 166440 114140 166520 114150
rect 166620 114140 166700 114150
rect 166800 114140 166880 114150
rect 166980 114140 167060 114150
rect 167160 114140 167240 114150
rect 167340 114140 167420 114150
rect 167520 114140 167600 114150
rect 167700 114140 167780 114150
rect 167880 114140 167960 114150
rect 168060 114140 168140 114150
rect 168240 114140 168320 114150
rect 168420 114140 168500 114150
rect 168600 114140 168680 114150
rect 168780 114140 168860 114150
rect 168960 114140 169040 114150
rect 169140 114140 169220 114150
rect 169320 114140 169400 114150
rect 169500 114140 169580 114150
rect 169680 114140 169760 114150
rect 169860 114140 169940 114150
rect 170040 114140 170120 114150
rect 170220 114140 170300 114150
rect 170400 114140 170480 114150
rect 170580 114140 170660 114150
rect 170760 114140 170840 114150
rect 170940 114140 171020 114150
rect 163460 114060 163470 114140
rect 163640 114060 163650 114140
rect 163820 114060 163830 114140
rect 164000 114060 164010 114140
rect 164180 114060 164190 114140
rect 164360 114060 164370 114140
rect 164540 114060 164550 114140
rect 164720 114060 164730 114140
rect 164900 114060 164910 114140
rect 165080 114060 165090 114140
rect 165260 114060 165270 114140
rect 165440 114060 165450 114140
rect 165620 114060 165630 114140
rect 165800 114060 165810 114140
rect 165980 114060 165990 114140
rect 166160 114060 166170 114140
rect 166340 114060 166350 114140
rect 166520 114060 166530 114140
rect 166700 114060 166710 114140
rect 166880 114060 166890 114140
rect 167060 114060 167070 114140
rect 167240 114060 167250 114140
rect 167420 114060 167430 114140
rect 167600 114060 167610 114140
rect 167780 114060 167790 114140
rect 167960 114060 167970 114140
rect 168140 114060 168150 114140
rect 168320 114060 168330 114140
rect 168500 114060 168510 114140
rect 168680 114060 168690 114140
rect 168860 114060 168870 114140
rect 169040 114060 169050 114140
rect 169220 114060 169230 114140
rect 169400 114060 169410 114140
rect 169580 114060 169590 114140
rect 169760 114060 169770 114140
rect 169940 114060 169950 114140
rect 170120 114060 170130 114140
rect 170300 114060 170310 114140
rect 170480 114060 170490 114140
rect 170660 114060 170670 114140
rect 170840 114060 170850 114140
rect 171020 114060 171030 114140
rect 152220 113890 152250 113920
rect 152340 113890 152370 113920
rect 159520 113890 159550 113920
rect 159640 113890 159670 113920
rect 152100 113860 152160 113890
rect 152220 113860 152280 113890
rect 152340 113860 152400 113890
rect 159400 113860 159460 113890
rect 159520 113860 159580 113890
rect 159640 113860 159700 113890
rect 152220 113770 152250 113800
rect 152340 113770 152370 113800
rect 159520 113770 159550 113800
rect 159640 113770 159670 113800
rect 163520 113770 163550 113800
rect 163640 113770 163670 113800
rect 170810 113770 170840 113800
rect 170930 113770 170960 113800
rect 152100 113740 152160 113770
rect 152220 113740 152280 113770
rect 152340 113740 152400 113770
rect 152810 113736 158990 113760
rect 159400 113740 159460 113770
rect 159520 113740 159580 113770
rect 159640 113740 159700 113770
rect 163400 113740 163460 113770
rect 163520 113740 163580 113770
rect 163640 113740 163700 113770
rect 170690 113740 170750 113770
rect 170810 113740 170870 113770
rect 170930 113740 170990 113770
rect 164280 113736 164360 113740
rect 164460 113736 164540 113740
rect 164640 113736 164720 113740
rect 164820 113736 164900 113740
rect 165000 113736 165080 113740
rect 165180 113736 165260 113740
rect 165360 113736 165440 113740
rect 165540 113736 165620 113740
rect 165720 113736 165800 113740
rect 165900 113736 165980 113740
rect 166080 113736 166160 113740
rect 166260 113736 166340 113740
rect 166440 113736 166520 113740
rect 166620 113736 166700 113740
rect 166800 113736 166880 113740
rect 166980 113736 167060 113740
rect 167160 113736 167240 113740
rect 167340 113736 167420 113740
rect 167520 113736 167600 113740
rect 167700 113736 167780 113740
rect 167880 113736 167960 113740
rect 168060 113736 168140 113740
rect 168240 113736 168320 113740
rect 168420 113736 168500 113740
rect 168600 113736 168680 113740
rect 168780 113736 168860 113740
rect 168960 113736 169040 113740
rect 169140 113736 169220 113740
rect 169320 113736 169400 113740
rect 169500 113736 169580 113740
rect 169680 113736 169760 113740
rect 169860 113736 169940 113740
rect 170040 113736 170120 113740
rect 37720 113670 37750 113700
rect 37840 113670 37870 113700
rect 146100 113670 146160 113700
rect 36120 113650 36130 113670
rect 36300 113650 36310 113670
rect 36480 113650 36490 113670
rect 36660 113650 36670 113670
rect 36840 113650 36850 113670
rect 37020 113650 37030 113670
rect 36040 113580 36120 113590
rect 36220 113580 36300 113590
rect 36400 113580 36480 113590
rect 36580 113580 36660 113590
rect 36760 113580 36840 113590
rect 36940 113580 37020 113590
rect 36120 113500 36130 113580
rect 36300 113500 36310 113580
rect 36480 113500 36490 113580
rect 36660 113500 36670 113580
rect 36840 113500 36850 113580
rect 37020 113500 37030 113580
rect 37100 113440 37190 113670
rect 37600 113640 37660 113670
rect 37720 113640 37780 113670
rect 37840 113640 37900 113670
rect 40060 113590 40120 113620
rect 41540 113590 41600 113620
rect 42360 113590 42420 113620
rect 43840 113590 43900 113620
rect 37720 113550 37750 113580
rect 37840 113550 37870 113580
rect 146100 113550 146160 113580
rect 37600 113520 37660 113550
rect 37720 113520 37780 113550
rect 37840 113520 37900 113550
rect 40060 113470 40120 113500
rect 41540 113470 41600 113500
rect 42360 113470 42420 113500
rect 43840 113470 43900 113500
rect 36000 113410 37190 113440
rect 37720 113430 37750 113460
rect 37840 113430 37870 113460
rect 146100 113430 146160 113460
rect 36120 113350 36130 113410
rect 36300 113350 36310 113410
rect 36480 113350 36490 113410
rect 36660 113350 36670 113410
rect 36840 113350 36850 113410
rect 37020 113350 37030 113410
rect 37100 113340 37190 113410
rect 37600 113400 37660 113430
rect 37720 113400 37780 113430
rect 37840 113400 37900 113430
rect 40060 113350 40120 113380
rect 41540 113350 41600 113380
rect 42360 113350 42420 113380
rect 43840 113350 43900 113380
rect 36000 113310 37190 113340
rect 37720 113310 37750 113340
rect 37840 113310 37870 113340
rect 146100 113310 146160 113340
rect 37100 113300 37190 113310
rect 36000 113290 37190 113300
rect 36040 113110 36120 113120
rect 36220 113110 36300 113120
rect 36400 113110 36480 113120
rect 36580 113110 36660 113120
rect 36760 113110 36840 113120
rect 36940 113110 37020 113120
rect 36120 113030 36130 113110
rect 36300 113030 36310 113110
rect 36480 113030 36490 113110
rect 36660 113030 36670 113110
rect 36840 113030 36850 113110
rect 37020 113030 37030 113110
rect 36040 112790 36120 112800
rect 36220 112790 36300 112800
rect 36400 112790 36480 112800
rect 36580 112790 36660 112800
rect 36760 112790 36840 112800
rect 36940 112790 37020 112800
rect 36120 112710 36130 112790
rect 36300 112710 36310 112790
rect 36480 112710 36490 112790
rect 36660 112710 36670 112790
rect 36840 112710 36850 112790
rect 37020 112710 37030 112790
rect 37100 112620 37190 113290
rect 37600 113280 37660 113310
rect 37720 113280 37780 113310
rect 37840 113280 37900 113310
rect 40060 113230 40120 113260
rect 41540 113230 41600 113260
rect 42360 113230 42420 113260
rect 43840 113230 43900 113260
rect 37720 113190 37750 113220
rect 37840 113190 37870 113220
rect 146100 113190 146160 113220
rect 37600 113160 37660 113190
rect 37720 113160 37780 113190
rect 37840 113160 37900 113190
rect 40060 113110 40120 113140
rect 41540 113110 41600 113140
rect 42360 113110 42420 113140
rect 43840 113110 43900 113140
rect 37720 113070 37750 113100
rect 37840 113070 37870 113100
rect 37600 113040 37660 113070
rect 37720 113040 37780 113070
rect 37840 113040 37900 113070
rect 40060 112990 40120 113020
rect 41540 112990 41600 113020
rect 42360 112990 42420 113020
rect 43840 112990 43900 113020
rect 37720 112950 37750 112980
rect 37840 112950 37870 112980
rect 146100 113070 146160 113100
rect 146100 112950 146160 112980
rect 37600 112920 37660 112950
rect 37720 112920 37780 112950
rect 37840 112920 37900 112950
rect 40060 112870 40120 112900
rect 41540 112870 41600 112900
rect 42360 112870 42420 112900
rect 43840 112870 43900 112900
rect 37720 112830 37750 112860
rect 37840 112830 37870 112860
rect 146100 112830 146160 112860
rect 37600 112800 37660 112830
rect 37720 112800 37780 112830
rect 37840 112800 37900 112830
rect 40060 112750 40120 112780
rect 41540 112750 41600 112780
rect 42360 112750 42420 112780
rect 43840 112750 43900 112780
rect 37720 112710 37750 112740
rect 37840 112710 37870 112740
rect 146100 112710 146160 112740
rect 37600 112680 37660 112710
rect 37720 112680 37780 112710
rect 37840 112680 37900 112710
rect 40060 112630 40120 112660
rect 41540 112630 41600 112660
rect 42360 112630 42420 112660
rect 43840 112630 43900 112660
rect 36000 112610 37190 112620
rect 37100 112510 37190 112610
rect 37720 112590 37750 112620
rect 37840 112590 37870 112620
rect 146100 112590 146160 112620
rect 37600 112560 37660 112590
rect 37720 112560 37780 112590
rect 37840 112560 37900 112590
rect 40060 112510 40120 112540
rect 41540 112510 41600 112540
rect 42360 112510 42420 112540
rect 43840 112510 43900 112540
rect 36000 112480 37190 112510
rect 36040 112470 36120 112480
rect 36220 112470 36300 112480
rect 36400 112470 36480 112480
rect 36580 112470 36660 112480
rect 36760 112470 36840 112480
rect 36940 112470 37020 112480
rect 36120 112410 36130 112470
rect 36300 112410 36310 112470
rect 36480 112410 36490 112470
rect 36660 112410 36670 112470
rect 36840 112410 36850 112470
rect 37020 112410 37030 112470
rect 37100 112410 37190 112480
rect 37720 112470 37750 112500
rect 37840 112470 37870 112500
rect 146100 112470 146160 112500
rect 37600 112440 37660 112470
rect 37720 112440 37780 112470
rect 37840 112440 37900 112470
rect 36000 112380 37190 112410
rect 40060 112390 40120 112420
rect 41540 112390 41600 112420
rect 42360 112390 42420 112420
rect 43840 112390 43900 112420
rect 36040 112320 36120 112330
rect 36220 112320 36300 112330
rect 36400 112320 36480 112330
rect 36580 112320 36660 112330
rect 36760 112320 36840 112330
rect 36940 112320 37020 112330
rect 36120 112240 36130 112320
rect 36300 112240 36310 112320
rect 36480 112240 36490 112320
rect 36660 112240 36670 112320
rect 36840 112240 36850 112320
rect 37020 112240 37030 112320
rect 37100 112180 37190 112380
rect 37720 112350 37750 112380
rect 37840 112350 37870 112380
rect 146100 112350 146160 112380
rect 37600 112320 37660 112350
rect 37720 112320 37780 112350
rect 37840 112320 37900 112350
rect 40060 112270 40120 112300
rect 41540 112270 41600 112300
rect 42360 112270 42420 112300
rect 43840 112270 43900 112300
rect 37720 112230 37750 112260
rect 37840 112230 37870 112260
rect 146100 112230 146160 112260
rect 37600 112200 37660 112230
rect 37720 112200 37780 112230
rect 37840 112200 37900 112230
rect 36000 112150 37190 112180
rect 40060 112150 40120 112180
rect 41540 112150 41600 112180
rect 42360 112150 42420 112180
rect 43840 112150 43900 112180
rect 36120 112090 36130 112150
rect 36300 112090 36310 112150
rect 36480 112090 36490 112150
rect 36660 112090 36670 112150
rect 36840 112090 36850 112150
rect 37020 112090 37030 112150
rect 37100 112080 37190 112150
rect 37720 112110 37750 112140
rect 37840 112110 37870 112140
rect 146100 112110 146160 112140
rect 37600 112080 37660 112110
rect 37720 112080 37780 112110
rect 37840 112080 37900 112110
rect 36000 112050 37190 112080
rect 37100 112040 37190 112050
rect 36000 112030 37190 112040
rect 40060 112030 40120 112060
rect 41540 112030 41600 112060
rect 42360 112030 42420 112060
rect 43840 112030 43900 112060
rect 36040 111850 36120 111860
rect 36220 111850 36300 111860
rect 36400 111850 36480 111860
rect 36580 111850 36660 111860
rect 36760 111850 36840 111860
rect 36940 111850 37020 111860
rect 36120 111770 36130 111850
rect 36300 111770 36310 111850
rect 36480 111770 36490 111850
rect 36660 111770 36670 111850
rect 36840 111770 36850 111850
rect 37020 111770 37030 111850
rect 36040 111530 36120 111540
rect 36220 111530 36300 111540
rect 36400 111530 36480 111540
rect 36580 111530 36660 111540
rect 36760 111530 36840 111540
rect 36940 111530 37020 111540
rect 36120 111450 36130 111530
rect 36300 111450 36310 111530
rect 36480 111450 36490 111530
rect 36660 111450 36670 111530
rect 36840 111450 36850 111530
rect 37020 111450 37030 111530
rect 37100 111360 37190 112030
rect 37720 111990 37750 112020
rect 37840 111990 37870 112020
rect 146100 111990 146160 112020
rect 37600 111960 37660 111990
rect 37720 111960 37780 111990
rect 37840 111960 37900 111990
rect 40060 111910 40120 111940
rect 41540 111910 41600 111940
rect 42360 111910 42420 111940
rect 43840 111910 43900 111940
rect 37720 111870 37750 111900
rect 37840 111870 37870 111900
rect 146100 111870 146160 111900
rect 37600 111840 37660 111870
rect 37720 111840 37780 111870
rect 37840 111840 37900 111870
rect 40060 111790 40120 111820
rect 41540 111790 41600 111820
rect 42360 111790 42420 111820
rect 43840 111790 43900 111820
rect 37720 111750 37750 111780
rect 37840 111750 37870 111780
rect 146100 111750 146160 111780
rect 37600 111720 37660 111750
rect 37720 111720 37780 111750
rect 37840 111720 37900 111750
rect 40060 111670 40120 111700
rect 41540 111670 41600 111700
rect 42360 111670 42420 111700
rect 43840 111670 43900 111700
rect 37720 111630 37750 111660
rect 37840 111630 37870 111660
rect 146100 111630 146160 111660
rect 37600 111600 37660 111630
rect 37720 111600 37780 111630
rect 37840 111600 37900 111630
rect 40060 111550 40120 111580
rect 41540 111550 41600 111580
rect 42360 111550 42420 111580
rect 43840 111550 43900 111580
rect 37720 111510 37750 111540
rect 37840 111510 37870 111540
rect 146100 111510 146160 111540
rect 37600 111480 37660 111510
rect 37720 111480 37780 111510
rect 37840 111480 37900 111510
rect 40060 111430 40120 111460
rect 41540 111430 41600 111460
rect 42360 111430 42420 111460
rect 43840 111430 43900 111460
rect 37720 111390 37750 111420
rect 37840 111390 37870 111420
rect 146100 111390 146160 111420
rect 37600 111360 37660 111390
rect 37720 111360 37780 111390
rect 37840 111360 37900 111390
rect 36000 111350 37190 111360
rect 37100 111250 37190 111350
rect 40060 111310 40120 111340
rect 41540 111310 41600 111340
rect 42360 111310 42420 111340
rect 43840 111310 43900 111340
rect 37720 111270 37750 111300
rect 37840 111270 37870 111300
rect 146100 111270 146160 111300
rect 36000 111220 37190 111250
rect 37600 111240 37660 111270
rect 37720 111240 37780 111270
rect 37840 111240 37900 111270
rect 36040 111210 36120 111220
rect 36220 111210 36300 111220
rect 36400 111210 36480 111220
rect 36580 111210 36660 111220
rect 36760 111210 36840 111220
rect 36940 111210 37020 111220
rect 36120 111150 36130 111210
rect 36300 111150 36310 111210
rect 36480 111150 36490 111210
rect 36660 111150 36670 111210
rect 36840 111150 36850 111210
rect 37020 111150 37030 111210
rect 37100 111150 37190 111220
rect 40060 111190 40120 111220
rect 41540 111190 41600 111220
rect 42360 111190 42420 111220
rect 43840 111190 43900 111220
rect 37720 111150 37750 111180
rect 37840 111150 37870 111180
rect 146100 111150 146160 111180
rect 36000 111120 37190 111150
rect 37600 111120 37660 111150
rect 37720 111120 37780 111150
rect 37840 111120 37900 111150
rect 36040 111060 36120 111070
rect 36220 111060 36300 111070
rect 36400 111060 36480 111070
rect 36580 111060 36660 111070
rect 36760 111060 36840 111070
rect 36940 111060 37020 111070
rect 36120 110980 36130 111060
rect 36300 110980 36310 111060
rect 36480 110980 36490 111060
rect 36660 110980 36670 111060
rect 36840 110980 36850 111060
rect 37020 110980 37030 111060
rect 37100 110920 37190 111120
rect 40060 111070 40120 111100
rect 41540 111070 41600 111100
rect 42360 111070 42420 111100
rect 43840 111070 43900 111100
rect 37720 111030 37750 111060
rect 37840 111030 37870 111060
rect 146100 111030 146160 111060
rect 37600 111000 37660 111030
rect 37720 111000 37780 111030
rect 37840 111000 37900 111030
rect 40060 110950 40120 110980
rect 41540 110950 41600 110980
rect 42360 110950 42420 110980
rect 43840 110950 43900 110980
rect 36000 110890 37190 110920
rect 37720 110910 37750 110940
rect 37840 110910 37870 110940
rect 146100 110910 146160 110940
rect 36120 110830 36130 110890
rect 36300 110830 36310 110890
rect 36480 110830 36490 110890
rect 36660 110830 36670 110890
rect 36840 110830 36850 110890
rect 37020 110830 37030 110890
rect 37100 110820 37190 110890
rect 37600 110880 37660 110910
rect 37720 110880 37780 110910
rect 37840 110880 37900 110910
rect 40060 110830 40120 110860
rect 41540 110830 41600 110860
rect 42360 110830 42420 110860
rect 43840 110830 43900 110860
rect 36000 110790 37190 110820
rect 37720 110790 37750 110820
rect 37840 110790 37870 110820
rect 146100 110790 146160 110820
rect 37100 110780 37190 110790
rect 36000 110770 37190 110780
rect 36040 110590 36120 110600
rect 36220 110590 36300 110600
rect 36400 110590 36480 110600
rect 36580 110590 36660 110600
rect 36760 110590 36840 110600
rect 36940 110590 37020 110600
rect 36120 110510 36130 110590
rect 36300 110510 36310 110590
rect 36480 110510 36490 110590
rect 36660 110510 36670 110590
rect 36840 110510 36850 110590
rect 37020 110510 37030 110590
rect 36040 110270 36120 110280
rect 36220 110270 36300 110280
rect 36400 110270 36480 110280
rect 36580 110270 36660 110280
rect 36760 110270 36840 110280
rect 36940 110270 37020 110280
rect 36120 110190 36130 110270
rect 36300 110190 36310 110270
rect 36480 110190 36490 110270
rect 36660 110190 36670 110270
rect 36840 110190 36850 110270
rect 37020 110190 37030 110270
rect 37100 110100 37190 110770
rect 37600 110760 37660 110790
rect 37720 110760 37780 110790
rect 37840 110760 37900 110790
rect 40060 110710 40120 110740
rect 41540 110710 41600 110740
rect 42360 110710 42420 110740
rect 43840 110710 43900 110740
rect 37720 110670 37750 110700
rect 37840 110670 37870 110700
rect 146100 110670 146160 110700
rect 37600 110640 37660 110670
rect 37720 110640 37780 110670
rect 37840 110640 37900 110670
rect 40060 110590 40120 110620
rect 41540 110590 41600 110620
rect 42360 110590 42420 110620
rect 43840 110590 43900 110620
rect 37720 110550 37750 110580
rect 37840 110550 37870 110580
rect 146100 110550 146160 110580
rect 37600 110520 37660 110550
rect 37720 110520 37780 110550
rect 37840 110520 37900 110550
rect 40060 110470 40120 110500
rect 41540 110470 41600 110500
rect 42360 110470 42420 110500
rect 43840 110470 43900 110500
rect 37720 110430 37750 110460
rect 37840 110430 37870 110460
rect 146100 110430 146160 110460
rect 37600 110400 37660 110430
rect 37720 110400 37780 110430
rect 37840 110400 37900 110430
rect 40060 110350 40120 110380
rect 41540 110350 41600 110380
rect 42360 110350 42420 110380
rect 43840 110350 43900 110380
rect 37720 110310 37750 110340
rect 37840 110310 37870 110340
rect 146100 110310 146160 110340
rect 37600 110280 37660 110310
rect 37720 110280 37780 110310
rect 37840 110280 37900 110310
rect 40060 110230 40120 110260
rect 41540 110230 41600 110260
rect 42360 110230 42420 110260
rect 43840 110230 43900 110260
rect 37720 110190 37750 110220
rect 37840 110190 37870 110220
rect 146100 110190 146160 110220
rect 37600 110160 37660 110190
rect 37720 110160 37780 110190
rect 37840 110160 37900 110190
rect 40060 110110 40120 110140
rect 41540 110110 41600 110140
rect 42360 110110 42420 110140
rect 43840 110110 43900 110140
rect 36000 110090 37190 110100
rect 37100 109990 37190 110090
rect 37720 110070 37750 110100
rect 37840 110070 37870 110100
rect 146100 110070 146160 110100
rect 37600 110040 37660 110070
rect 37720 110040 37780 110070
rect 37840 110040 37900 110070
rect 40060 109990 40120 110020
rect 41540 109990 41600 110020
rect 42360 109990 42420 110020
rect 43840 109990 43900 110020
rect 36000 109960 37190 109990
rect 36040 109950 36120 109960
rect 36220 109950 36300 109960
rect 36400 109950 36480 109960
rect 36580 109950 36660 109960
rect 36760 109950 36840 109960
rect 36940 109950 37020 109960
rect 36120 109890 36130 109950
rect 36300 109890 36310 109950
rect 36480 109890 36490 109950
rect 36660 109890 36670 109950
rect 36840 109890 36850 109950
rect 37020 109890 37030 109950
rect 37100 109890 37190 109960
rect 37720 109950 37750 109980
rect 37840 109950 37870 109980
rect 146100 109950 146160 109980
rect 37600 109920 37660 109950
rect 37720 109920 37780 109950
rect 37840 109920 37900 109950
rect 36000 109860 37190 109890
rect 40060 109870 40120 109900
rect 41540 109870 41600 109900
rect 42360 109870 42420 109900
rect 43840 109870 43900 109900
rect 36040 109800 36120 109810
rect 36220 109800 36300 109810
rect 36400 109800 36480 109810
rect 36580 109800 36660 109810
rect 36760 109800 36840 109810
rect 36940 109800 37020 109810
rect 36120 109720 36130 109800
rect 36300 109720 36310 109800
rect 36480 109720 36490 109800
rect 36660 109720 36670 109800
rect 36840 109720 36850 109800
rect 37020 109720 37030 109800
rect 37100 109660 37190 109860
rect 37720 109830 37750 109860
rect 37840 109830 37870 109860
rect 146100 109830 146160 109860
rect 37600 109800 37660 109830
rect 37720 109800 37780 109830
rect 37840 109800 37900 109830
rect 40060 109750 40120 109780
rect 41540 109750 41600 109780
rect 42360 109750 42420 109780
rect 43840 109750 43900 109780
rect 37720 109710 37750 109740
rect 37840 109710 37870 109740
rect 146100 109710 146160 109740
rect 37600 109680 37660 109710
rect 37720 109680 37780 109710
rect 37840 109680 37900 109710
rect 36000 109630 37190 109660
rect 40060 109630 40120 109660
rect 41540 109630 41600 109660
rect 42360 109630 42420 109660
rect 43840 109630 43900 109660
rect 36120 109570 36130 109630
rect 36300 109570 36310 109630
rect 36480 109570 36490 109630
rect 36660 109570 36670 109630
rect 36840 109570 36850 109630
rect 37020 109570 37030 109630
rect 37100 109560 37190 109630
rect 37720 109590 37750 109620
rect 37840 109590 37870 109620
rect 146100 109590 146160 109620
rect 37600 109560 37660 109590
rect 37720 109560 37780 109590
rect 37840 109560 37900 109590
rect 36000 109530 37190 109560
rect 37100 109520 37190 109530
rect 36000 109510 37190 109520
rect 40060 109510 40120 109540
rect 41540 109510 41600 109540
rect 42360 109510 42420 109540
rect 43840 109510 43900 109540
rect 36040 109330 36120 109340
rect 36220 109330 36300 109340
rect 36400 109330 36480 109340
rect 36580 109330 36660 109340
rect 36760 109330 36840 109340
rect 36940 109330 37020 109340
rect 36120 109250 36130 109330
rect 36300 109250 36310 109330
rect 36480 109250 36490 109330
rect 36660 109250 36670 109330
rect 36840 109250 36850 109330
rect 37020 109250 37030 109330
rect 36040 109010 36120 109020
rect 36220 109010 36300 109020
rect 36400 109010 36480 109020
rect 36580 109010 36660 109020
rect 36760 109010 36840 109020
rect 36940 109010 37020 109020
rect 36120 108930 36130 109010
rect 36300 108930 36310 109010
rect 36480 108930 36490 109010
rect 36660 108930 36670 109010
rect 36840 108930 36850 109010
rect 37020 108930 37030 109010
rect 37100 108840 37190 109510
rect 37720 109470 37750 109500
rect 37840 109470 37870 109500
rect 146100 109470 146160 109500
rect 37600 109440 37660 109470
rect 37720 109440 37780 109470
rect 37840 109440 37900 109470
rect 40060 109390 40120 109420
rect 41540 109390 41600 109420
rect 42360 109390 42420 109420
rect 43840 109390 43900 109420
rect 37720 109350 37750 109380
rect 37840 109350 37870 109380
rect 146100 109350 146160 109380
rect 37600 109320 37660 109350
rect 37720 109320 37780 109350
rect 37840 109320 37900 109350
rect 40060 109270 40120 109300
rect 41540 109270 41600 109300
rect 42360 109270 42420 109300
rect 43840 109270 43900 109300
rect 37720 109230 37750 109260
rect 37840 109230 37870 109260
rect 37600 109200 37660 109230
rect 37720 109200 37780 109230
rect 37840 109200 37900 109230
rect 40060 109150 40120 109180
rect 41540 109150 41600 109180
rect 42360 109150 42420 109180
rect 43840 109150 43900 109180
rect 37720 109110 37750 109140
rect 37840 109110 37870 109140
rect 37600 109080 37660 109110
rect 37720 109080 37780 109110
rect 37840 109080 37900 109110
rect 146100 109230 146160 109260
rect 146100 109110 146160 109140
rect 40060 109030 40120 109060
rect 41540 109030 41600 109060
rect 42360 109030 42420 109060
rect 43840 109030 43900 109060
rect 37720 108990 37750 109020
rect 37840 108990 37870 109020
rect 146100 108990 146160 109020
rect 37600 108960 37660 108990
rect 37720 108960 37780 108990
rect 37840 108960 37900 108990
rect 40060 108910 40120 108940
rect 41540 108910 41600 108940
rect 42360 108910 42420 108940
rect 43840 108910 43900 108940
rect 37720 108870 37750 108900
rect 37840 108870 37870 108900
rect 146100 108870 146160 108900
rect 37600 108840 37660 108870
rect 37720 108840 37780 108870
rect 37840 108840 37900 108870
rect 36000 108830 37190 108840
rect 37100 108730 37190 108830
rect 40060 108790 40120 108820
rect 41540 108790 41600 108820
rect 42360 108790 42420 108820
rect 43840 108790 43900 108820
rect 37720 108750 37750 108780
rect 37840 108750 37870 108780
rect 146100 108750 146160 108780
rect 36000 108700 37190 108730
rect 37600 108720 37660 108750
rect 37720 108720 37780 108750
rect 37840 108720 37900 108750
rect 40685 108710 40925 108740
rect 36040 108690 36120 108700
rect 36220 108690 36300 108700
rect 36400 108690 36480 108700
rect 36580 108690 36660 108700
rect 36760 108690 36840 108700
rect 36940 108690 37020 108700
rect 36120 108630 36130 108690
rect 36300 108630 36310 108690
rect 36480 108630 36490 108690
rect 36660 108630 36670 108690
rect 36840 108630 36850 108690
rect 37020 108630 37030 108690
rect 37100 108630 37190 108700
rect 40060 108670 40120 108700
rect 37720 108630 37750 108660
rect 37840 108630 37870 108660
rect 40685 108650 40715 108710
rect 40775 108650 40865 108710
rect 40895 108650 40925 108710
rect 41540 108670 41600 108700
rect 42360 108670 42420 108700
rect 43840 108670 43900 108700
rect 36000 108600 37190 108630
rect 37600 108600 37660 108630
rect 37720 108600 37780 108630
rect 37840 108600 37900 108630
rect 40685 108620 40925 108650
rect 146100 108630 146160 108660
rect 36040 108540 36120 108550
rect 36220 108540 36300 108550
rect 36400 108540 36480 108550
rect 36580 108540 36660 108550
rect 36760 108540 36840 108550
rect 36940 108540 37020 108550
rect 36120 108460 36130 108540
rect 36300 108460 36310 108540
rect 36480 108460 36490 108540
rect 36660 108460 36670 108540
rect 36840 108460 36850 108540
rect 37020 108460 37030 108540
rect 37100 108400 37190 108600
rect 40060 108550 40120 108580
rect 41540 108550 41600 108580
rect 42360 108550 42420 108580
rect 43840 108550 43900 108580
rect 37720 108510 37750 108540
rect 37840 108510 37870 108540
rect 146100 108510 146160 108540
rect 37600 108480 37660 108510
rect 37720 108480 37780 108510
rect 37840 108480 37900 108510
rect 40060 108430 40120 108460
rect 41540 108430 41600 108460
rect 42360 108430 42420 108460
rect 43840 108430 43900 108460
rect 36000 108370 37190 108400
rect 37720 108390 37750 108420
rect 37840 108390 37870 108420
rect 146100 108390 146160 108420
rect 36120 108310 36130 108370
rect 36300 108310 36310 108370
rect 36480 108310 36490 108370
rect 36660 108310 36670 108370
rect 36840 108310 36850 108370
rect 37020 108310 37030 108370
rect 37100 108300 37190 108370
rect 37600 108360 37660 108390
rect 37720 108360 37780 108390
rect 37840 108360 37900 108390
rect 40060 108310 40120 108340
rect 41540 108310 41600 108340
rect 42360 108310 42420 108340
rect 43840 108310 43900 108340
rect 36000 108270 37190 108300
rect 37720 108270 37750 108300
rect 37840 108270 37870 108300
rect 146100 108270 146160 108300
rect 37100 108260 37190 108270
rect 36000 108250 37190 108260
rect 36040 108070 36120 108080
rect 36220 108070 36300 108080
rect 36400 108070 36480 108080
rect 36580 108070 36660 108080
rect 36760 108070 36840 108080
rect 36940 108070 37020 108080
rect 36120 107990 36130 108070
rect 36300 107990 36310 108070
rect 36480 107990 36490 108070
rect 36660 107990 36670 108070
rect 36840 107990 36850 108070
rect 37020 107990 37030 108070
rect 36040 107750 36120 107760
rect 36220 107750 36300 107760
rect 36400 107750 36480 107760
rect 36580 107750 36660 107760
rect 36760 107750 36840 107760
rect 36940 107750 37020 107760
rect 36120 107670 36130 107750
rect 36300 107670 36310 107750
rect 36480 107670 36490 107750
rect 36660 107670 36670 107750
rect 36840 107670 36850 107750
rect 37020 107670 37030 107750
rect 37100 107580 37190 108250
rect 37600 108240 37660 108270
rect 37720 108240 37780 108270
rect 37840 108240 37900 108270
rect 40060 108190 40120 108220
rect 41540 108190 41600 108220
rect 42360 108190 42420 108220
rect 43840 108190 43900 108220
rect 37720 108150 37750 108180
rect 37840 108150 37870 108180
rect 146100 108150 146160 108180
rect 37600 108120 37660 108150
rect 37720 108120 37780 108150
rect 37840 108120 37900 108150
rect 40060 108070 40120 108100
rect 41540 108070 41600 108100
rect 42360 108070 42420 108100
rect 43840 108070 43900 108100
rect 37720 108030 37750 108060
rect 37840 108030 37870 108060
rect 146100 108030 146160 108060
rect 37600 108000 37660 108030
rect 37720 108000 37780 108030
rect 37840 108000 37900 108030
rect 40678 108004 40758 108014
rect 40838 108004 40918 108014
rect 40060 107950 40120 107980
rect 37720 107910 37750 107940
rect 37840 107910 37870 107940
rect 40758 107934 40768 108004
rect 40678 107924 40768 107934
rect 40838 107934 40848 108004
rect 40918 107934 40928 108004
rect 41540 107950 41600 107980
rect 42360 107950 42420 107980
rect 43840 107950 43900 107980
rect 40838 107924 40928 107934
rect 146100 107910 146160 107940
rect 37600 107880 37660 107910
rect 37720 107880 37780 107910
rect 37840 107880 37900 107910
rect 40060 107830 40120 107860
rect 40678 107844 40758 107854
rect 40838 107844 40918 107854
rect 37720 107790 37750 107820
rect 37840 107790 37870 107820
rect 37600 107760 37660 107790
rect 37720 107760 37780 107790
rect 37840 107760 37900 107790
rect 40758 107764 40768 107844
rect 40838 107764 40848 107844
rect 40918 107764 40928 107844
rect 41540 107830 41600 107860
rect 42360 107830 42420 107860
rect 43840 107830 43900 107860
rect 146100 107790 146160 107820
rect 40060 107710 40120 107740
rect 41540 107710 41600 107740
rect 42360 107710 42420 107740
rect 43840 107710 43900 107740
rect 37720 107670 37750 107700
rect 37840 107670 37870 107700
rect 146100 107670 146160 107700
rect 37600 107640 37660 107670
rect 37720 107640 37780 107670
rect 37840 107640 37900 107670
rect 40060 107590 40120 107620
rect 41540 107590 41600 107620
rect 42360 107590 42420 107620
rect 43840 107590 43900 107620
rect 36000 107570 37190 107580
rect 37100 107470 37190 107570
rect 37720 107550 37750 107580
rect 37840 107550 37870 107580
rect 146100 107550 146160 107580
rect 37600 107520 37660 107550
rect 37720 107520 37780 107550
rect 37840 107520 37900 107550
rect 40060 107470 40120 107500
rect 41540 107470 41600 107500
rect 42360 107470 42420 107500
rect 43840 107470 43900 107500
rect 36000 107440 37190 107470
rect 36040 107430 36120 107440
rect 36220 107430 36300 107440
rect 36400 107430 36480 107440
rect 36580 107430 36660 107440
rect 36760 107430 36840 107440
rect 36940 107430 37020 107440
rect 36120 107370 36130 107430
rect 36300 107370 36310 107430
rect 36480 107370 36490 107430
rect 36660 107370 36670 107430
rect 36840 107370 36850 107430
rect 37020 107370 37030 107430
rect 37100 107370 37190 107440
rect 37720 107430 37750 107460
rect 37840 107430 37870 107460
rect 146100 107430 146160 107460
rect 37600 107400 37660 107430
rect 37720 107400 37780 107430
rect 37840 107400 37900 107430
rect 36000 107340 37190 107370
rect 40060 107350 40120 107380
rect 41540 107350 41600 107380
rect 42360 107350 42420 107380
rect 43840 107350 43900 107380
rect 36040 107280 36120 107290
rect 36220 107280 36300 107290
rect 36400 107280 36480 107290
rect 36580 107280 36660 107290
rect 36760 107280 36840 107290
rect 36940 107280 37020 107290
rect 36120 107200 36130 107280
rect 36300 107200 36310 107280
rect 36480 107200 36490 107280
rect 36660 107200 36670 107280
rect 36840 107200 36850 107280
rect 37020 107200 37030 107280
rect 37100 107140 37190 107340
rect 37720 107310 37750 107340
rect 37840 107310 37870 107340
rect 146100 107310 146160 107340
rect 37600 107280 37660 107310
rect 37720 107280 37780 107310
rect 37840 107280 37900 107310
rect 40060 107230 40120 107260
rect 41540 107230 41600 107260
rect 42360 107230 42420 107260
rect 43840 107230 43900 107260
rect 37720 107190 37750 107220
rect 37840 107190 37870 107220
rect 146100 107190 146160 107220
rect 37600 107160 37660 107190
rect 37720 107160 37780 107190
rect 37840 107160 37900 107190
rect 36000 107110 37190 107140
rect 40060 107110 40120 107140
rect 41540 107110 41600 107140
rect 42360 107110 42420 107140
rect 43840 107110 43900 107140
rect 36120 107050 36130 107110
rect 36300 107050 36310 107110
rect 36480 107050 36490 107110
rect 36660 107050 36670 107110
rect 36840 107050 36850 107110
rect 37020 107050 37030 107110
rect 37100 107040 37190 107110
rect 37720 107070 37750 107100
rect 37840 107070 37870 107100
rect 146100 107070 146160 107100
rect 37600 107040 37660 107070
rect 37720 107040 37780 107070
rect 37840 107040 37900 107070
rect 36000 107010 37190 107040
rect 37100 107000 37190 107010
rect 36000 106990 37190 107000
rect 40060 106990 40120 107020
rect 41540 106990 41600 107020
rect 42360 106990 42420 107020
rect 43840 106990 43900 107020
rect 36040 106810 36120 106820
rect 36220 106810 36300 106820
rect 36400 106810 36480 106820
rect 36580 106810 36660 106820
rect 36760 106810 36840 106820
rect 36940 106810 37020 106820
rect 36120 106730 36130 106810
rect 36300 106730 36310 106810
rect 36480 106730 36490 106810
rect 36660 106730 36670 106810
rect 36840 106730 36850 106810
rect 37020 106730 37030 106810
rect 36040 106490 36120 106500
rect 36220 106490 36300 106500
rect 36400 106490 36480 106500
rect 36580 106490 36660 106500
rect 36760 106490 36840 106500
rect 36940 106490 37020 106500
rect 36120 106410 36130 106490
rect 36300 106410 36310 106490
rect 36480 106410 36490 106490
rect 36660 106410 36670 106490
rect 36840 106410 36850 106490
rect 37020 106410 37030 106490
rect 37100 106320 37190 106990
rect 37720 106950 37750 106980
rect 37840 106950 37870 106980
rect 42595 106975 42675 106985
rect 37600 106920 37660 106950
rect 37720 106920 37780 106950
rect 37840 106920 37900 106950
rect 42675 106905 42685 106975
rect 146100 106950 146160 106980
rect 40060 106870 40120 106900
rect 41540 106870 41600 106900
rect 42360 106870 42420 106900
rect 42595 106895 42685 106905
rect 43840 106870 43900 106900
rect 37720 106830 37750 106860
rect 37840 106830 37870 106860
rect 37600 106800 37660 106830
rect 37720 106800 37780 106830
rect 37840 106800 37900 106830
rect 42595 106815 42675 106825
rect 40060 106750 40120 106780
rect 41540 106750 41600 106780
rect 42360 106750 42420 106780
rect 37720 106710 37750 106740
rect 37840 106710 37870 106740
rect 42675 106735 42685 106815
rect 43030 106800 43390 106860
rect 146100 106830 146160 106860
rect 43840 106750 43900 106780
rect 38595 106715 38675 106725
rect 38775 106715 38855 106725
rect 38955 106715 39035 106725
rect 39135 106715 39215 106725
rect 39315 106715 39395 106725
rect 37600 106680 37660 106710
rect 37720 106680 37780 106710
rect 37840 106680 37900 106710
rect 38675 106635 38685 106715
rect 38855 106635 38865 106715
rect 39035 106635 39045 106715
rect 39215 106635 39225 106715
rect 39395 106635 39405 106715
rect 43580 106670 43700 106730
rect 146100 106710 146160 106740
rect 40060 106630 40120 106660
rect 41540 106630 41600 106660
rect 42360 106630 42420 106660
rect 42950 106650 43560 106660
rect 43550 106645 43560 106650
rect 42910 106635 43560 106645
rect 37720 106590 37750 106620
rect 37840 106590 37870 106620
rect 37600 106560 37660 106590
rect 37720 106560 37780 106590
rect 37840 106560 37900 106590
rect 42900 106585 42910 106635
rect 38595 106535 38675 106545
rect 38775 106535 38855 106545
rect 38955 106535 39035 106545
rect 39135 106535 39215 106545
rect 39315 106535 39395 106545
rect 43030 106540 43390 106600
rect 37720 106470 37750 106500
rect 37840 106470 37870 106500
rect 37600 106440 37660 106470
rect 37720 106440 37780 106470
rect 37840 106440 37900 106470
rect 38675 106455 38685 106535
rect 38855 106455 38865 106535
rect 39035 106455 39045 106535
rect 39215 106455 39225 106535
rect 39395 106455 39405 106535
rect 40060 106510 40120 106540
rect 41540 106510 41600 106540
rect 42360 106510 42420 106540
rect 42682 106460 42822 106530
rect 40060 106390 40120 106420
rect 40678 106399 40758 106409
rect 40838 106399 40918 106409
rect 37720 106350 37750 106380
rect 37840 106350 37870 106380
rect 38595 106355 38675 106365
rect 38775 106355 38855 106365
rect 38955 106355 39035 106365
rect 39135 106355 39215 106365
rect 39315 106355 39395 106365
rect 37600 106320 37660 106350
rect 37720 106320 37780 106350
rect 37840 106320 37900 106350
rect 36000 106310 37190 106320
rect 37100 106210 37190 106310
rect 38675 106275 38685 106355
rect 38855 106275 38865 106355
rect 39035 106275 39045 106355
rect 39215 106275 39225 106355
rect 39395 106275 39405 106355
rect 40758 106319 40768 106399
rect 40838 106319 40848 106399
rect 40918 106319 40928 106399
rect 41540 106390 41600 106420
rect 42360 106390 42420 106420
rect 42822 106400 42892 106460
rect 42822 106390 43470 106400
rect 43550 106390 43560 106635
rect 43700 106550 43760 106670
rect 43840 106630 43900 106660
rect 146100 106590 146160 106620
rect 43840 106510 43900 106540
rect 146100 106470 146160 106500
rect 43580 106410 43700 106470
rect 42822 106320 42892 106390
rect 42910 106375 43560 106385
rect 42900 106325 42910 106375
rect 40060 106270 40120 106300
rect 37720 106230 37750 106260
rect 37840 106230 37870 106260
rect 40685 106250 40925 106280
rect 41540 106270 41600 106300
rect 42360 106270 42420 106300
rect 42682 106260 42822 106320
rect 43030 106280 43390 106340
rect 43700 106290 43760 106410
rect 43840 106390 43900 106420
rect 146100 106350 146160 106380
rect 43840 106270 43900 106300
rect 36000 106180 37190 106210
rect 37600 106200 37660 106230
rect 37720 106200 37780 106230
rect 37840 106200 37900 106230
rect 40685 106190 40715 106250
rect 40775 106190 40865 106250
rect 40895 106190 40925 106250
rect 36040 106170 36120 106180
rect 36220 106170 36300 106180
rect 36400 106170 36480 106180
rect 36580 106170 36660 106180
rect 36760 106170 36840 106180
rect 36940 106170 37020 106180
rect 36120 106110 36130 106170
rect 36300 106110 36310 106170
rect 36480 106110 36490 106170
rect 36660 106110 36670 106170
rect 36840 106110 36850 106170
rect 37020 106110 37030 106170
rect 37100 106110 37190 106180
rect 38595 106175 38675 106185
rect 38775 106175 38855 106185
rect 38955 106175 39035 106185
rect 39135 106175 39215 106185
rect 39315 106175 39395 106185
rect 37720 106110 37750 106140
rect 37840 106110 37870 106140
rect 36000 106080 37190 106110
rect 37600 106080 37660 106110
rect 37720 106080 37780 106110
rect 37840 106080 37900 106110
rect 38675 106095 38685 106175
rect 38855 106095 38865 106175
rect 39035 106095 39045 106175
rect 39215 106095 39225 106175
rect 39395 106095 39405 106175
rect 40060 106150 40120 106180
rect 40685 106160 40925 106190
rect 41540 106150 41600 106180
rect 42360 106150 42420 106180
rect 40678 106129 40758 106139
rect 40838 106129 40918 106139
rect 36040 106020 36120 106030
rect 36220 106020 36300 106030
rect 36400 106020 36480 106030
rect 36580 106020 36660 106030
rect 36760 106020 36840 106030
rect 36940 106020 37020 106030
rect 36120 105940 36130 106020
rect 36300 105940 36310 106020
rect 36480 105940 36490 106020
rect 36660 105940 36670 106020
rect 36840 105940 36850 106020
rect 37020 105940 37030 106020
rect 37100 105880 37190 106080
rect 40060 106030 40120 106060
rect 40758 106049 40768 106129
rect 40838 106049 40848 106129
rect 40918 106049 40928 106129
rect 42822 106120 42892 106260
rect 146100 106230 146160 106260
rect 43580 106150 43700 106210
rect 43840 106150 43900 106180
rect 42950 106130 43560 106140
rect 43550 106125 43560 106130
rect 42682 106060 42822 106120
rect 42910 106115 43560 106125
rect 42900 106065 42910 106115
rect 41540 106030 41600 106060
rect 42360 106030 42420 106060
rect 37720 105990 37750 106020
rect 37840 105990 37870 106020
rect 38595 105995 38675 106005
rect 38775 105995 38855 106005
rect 38955 105995 39035 106005
rect 39135 105995 39215 106005
rect 39315 105995 39395 106005
rect 37600 105960 37660 105990
rect 37720 105960 37780 105990
rect 37840 105960 37900 105990
rect 38675 105915 38685 105995
rect 38855 105915 38865 105995
rect 39035 105915 39045 105995
rect 39215 105915 39225 105995
rect 39395 105915 39405 105995
rect 40060 105910 40120 105940
rect 41540 105910 41600 105940
rect 42360 105910 42420 105940
rect 42822 105920 42892 106060
rect 43030 106020 43390 106080
rect 36000 105850 37190 105880
rect 37720 105870 37750 105900
rect 37840 105870 37870 105900
rect 36120 105790 36130 105850
rect 36300 105790 36310 105850
rect 36480 105790 36490 105850
rect 36660 105790 36670 105850
rect 36840 105790 36850 105850
rect 37020 105790 37030 105850
rect 37100 105780 37190 105850
rect 37600 105840 37660 105870
rect 37720 105840 37780 105870
rect 37840 105840 37900 105870
rect 40170 105820 40180 105910
rect 40060 105790 40120 105820
rect 36000 105750 37190 105780
rect 37720 105750 37750 105780
rect 37840 105750 37870 105780
rect 37100 105740 37190 105750
rect 36000 105730 37190 105740
rect 36040 105550 36120 105560
rect 36220 105550 36300 105560
rect 36400 105550 36480 105560
rect 36580 105550 36660 105560
rect 36760 105550 36840 105560
rect 36940 105550 37020 105560
rect 36120 105470 36130 105550
rect 36300 105470 36310 105550
rect 36480 105470 36490 105550
rect 36660 105470 36670 105550
rect 36840 105470 36850 105550
rect 37020 105470 37030 105550
rect 36040 105230 36120 105240
rect 36220 105230 36300 105240
rect 36400 105230 36480 105240
rect 36580 105230 36660 105240
rect 36760 105230 36840 105240
rect 36940 105230 37020 105240
rect 36120 105150 36130 105230
rect 36300 105150 36310 105230
rect 36480 105150 36490 105230
rect 36660 105150 36670 105230
rect 36840 105150 36850 105230
rect 37020 105150 37030 105230
rect 37100 105060 37190 105730
rect 37600 105720 37660 105750
rect 37720 105720 37780 105750
rect 37840 105720 37900 105750
rect 40060 105670 40120 105700
rect 37720 105630 37750 105660
rect 37840 105630 37870 105660
rect 37600 105600 37660 105630
rect 37720 105600 37780 105630
rect 37840 105600 37900 105630
rect 40060 105550 40120 105580
rect 37720 105510 37750 105540
rect 37840 105510 37870 105540
rect 37600 105480 37660 105510
rect 37720 105480 37780 105510
rect 37840 105480 37900 105510
rect 40060 105430 40120 105460
rect 37720 105390 37750 105420
rect 37840 105390 37870 105420
rect 37600 105360 37660 105390
rect 37720 105360 37780 105390
rect 37840 105360 37900 105390
rect 40060 105310 40120 105340
rect 37720 105270 37750 105300
rect 37840 105270 37870 105300
rect 37600 105240 37660 105270
rect 37720 105240 37780 105270
rect 37840 105240 37900 105270
rect 40060 105190 40120 105220
rect 37720 105150 37750 105180
rect 37840 105150 37870 105180
rect 37600 105120 37660 105150
rect 37720 105120 37780 105150
rect 37840 105120 37900 105150
rect 40060 105070 40120 105100
rect 36000 105050 37190 105060
rect 37100 104950 37190 105050
rect 37720 105030 37750 105060
rect 37840 105030 37870 105060
rect 40260 105030 40270 105820
rect 40380 105810 41180 105900
rect 40650 105780 40770 105810
rect 40930 105780 41050 105810
rect 41090 105780 41180 105810
rect 40650 105690 40660 105780
rect 40760 105750 40830 105780
rect 40770 105660 40830 105750
rect 40930 105690 40940 105780
rect 41050 105660 41180 105780
rect 41260 105740 41340 105750
rect 41340 105690 41350 105740
rect 41090 105625 41180 105660
rect 41230 105630 41350 105690
rect 40470 105620 41180 105625
rect 40370 105610 41180 105620
rect 40370 105530 40380 105610
rect 40470 105605 41180 105610
rect 40420 105595 41210 105605
rect 41090 105545 41180 105595
rect 40470 105530 41180 105545
rect 40460 105515 41180 105530
rect 40460 105325 40470 105515
rect 40650 105480 40770 105515
rect 40930 105480 41050 105515
rect 41090 105480 41180 105515
rect 41350 105510 41410 105630
rect 40770 105470 40830 105480
rect 40530 105460 40610 105470
rect 40670 105460 40750 105470
rect 40770 105460 40890 105470
rect 40950 105460 41030 105470
rect 40610 105380 40620 105460
rect 40750 105380 40760 105460
rect 40770 105360 40830 105460
rect 40890 105380 40900 105460
rect 41030 105380 41040 105460
rect 41050 105360 41180 105480
rect 41260 105460 41340 105470
rect 41340 105390 41350 105460
rect 41090 105325 41180 105360
rect 41230 105330 41350 105390
rect 40460 105310 41180 105325
rect 40470 105305 41180 105310
rect 40420 105295 41210 105305
rect 41090 105245 41180 105295
rect 40470 105215 41180 105245
rect 40650 105180 40770 105215
rect 40930 105180 41050 105215
rect 41090 105180 41180 105215
rect 41350 105210 41410 105330
rect 41480 105180 41490 105890
rect 42860 105870 43470 105880
rect 43550 105870 43560 106115
rect 43700 106030 43760 106150
rect 146100 106110 146160 106140
rect 43840 106030 43900 106060
rect 146100 105990 146160 106020
rect 43580 105890 43700 105950
rect 43840 105910 43900 105940
rect 42910 105855 43560 105865
rect 41540 105790 41600 105820
rect 42360 105790 42420 105820
rect 42900 105805 42910 105855
rect 43030 105760 43390 105820
rect 43700 105770 43760 105890
rect 146100 105870 146160 105900
rect 43840 105790 43900 105820
rect 146100 105750 146160 105780
rect 41540 105670 41600 105700
rect 42360 105670 42420 105700
rect 42470 105660 42480 105750
rect 43840 105670 43900 105700
rect 41540 105550 41600 105580
rect 42360 105550 42420 105580
rect 41540 105430 41600 105460
rect 42360 105430 42420 105460
rect 41540 105310 41600 105340
rect 42360 105310 42420 105340
rect 41540 105190 41600 105220
rect 42360 105190 42420 105220
rect 42560 105180 42570 105660
rect 146100 105630 146160 105660
rect 42960 105620 43460 105630
rect 42620 105600 42700 105610
rect 42700 105530 42710 105600
rect 42620 105520 42710 105530
rect 42770 105520 42780 105610
rect 43840 105550 43900 105580
rect 42620 105440 42700 105450
rect 42700 105390 42710 105440
rect 42610 105330 42730 105390
rect 42730 105305 42790 105330
rect 42860 105320 42870 105520
rect 42910 105480 43030 105540
rect 43190 105480 43310 105540
rect 146100 105510 146160 105540
rect 43030 105470 43090 105480
rect 43310 105470 43370 105480
rect 42930 105460 43010 105470
rect 43030 105460 43150 105470
rect 43210 105460 43290 105470
rect 43310 105460 43430 105470
rect 43010 105380 43020 105460
rect 43030 105360 43090 105460
rect 43150 105380 43160 105460
rect 43290 105380 43300 105460
rect 43310 105360 43370 105460
rect 43430 105380 43440 105460
rect 43840 105430 43900 105460
rect 146100 105390 146160 105420
rect 42860 105310 43500 105320
rect 43840 105310 43900 105340
rect 42730 105295 43540 105305
rect 42730 105210 42790 105295
rect 43540 105245 43550 105295
rect 42860 105180 42870 105230
rect 42910 105180 43030 105240
rect 43190 105180 43310 105240
rect 43840 105190 43900 105220
rect 46700 105195 48000 105340
rect 40770 105170 40830 105180
rect 40530 105160 40610 105170
rect 40770 105160 40890 105170
rect 40610 105080 40620 105160
rect 40770 105060 40830 105160
rect 40890 105080 40900 105160
rect 41050 105060 41180 105180
rect 43030 105170 43090 105180
rect 43310 105170 43370 105180
rect 43030 105160 43150 105170
rect 43310 105160 43430 105170
rect 46755 105160 48000 105195
rect 146100 105270 146160 105300
rect 41540 105070 41600 105100
rect 42360 105070 42420 105100
rect 43030 105060 43090 105160
rect 43150 105080 43160 105160
rect 43310 105060 43370 105160
rect 43430 105080 43440 105160
rect 146100 105150 146160 105180
rect 43840 105070 43900 105100
rect 41090 105050 41180 105060
rect 40470 105030 41180 105050
rect 146100 105030 146160 105060
rect 146210 105040 146220 105130
rect 37600 105000 37660 105030
rect 37720 105000 37780 105030
rect 37840 105000 37900 105030
rect 40060 104950 40120 104980
rect 36000 104920 37190 104950
rect 40170 104940 40180 105030
rect 40260 105020 41100 105030
rect 36040 104910 36120 104920
rect 36220 104910 36300 104920
rect 36400 104910 36480 104920
rect 36580 104910 36660 104920
rect 36760 104910 36840 104920
rect 36940 104910 37020 104920
rect 36120 104850 36130 104910
rect 36300 104850 36310 104910
rect 36480 104850 36490 104910
rect 36660 104850 36670 104910
rect 36840 104850 36850 104910
rect 37020 104850 37030 104910
rect 37100 104850 37190 104920
rect 37720 104910 37750 104940
rect 37840 104910 37870 104940
rect 37600 104880 37660 104910
rect 37720 104880 37780 104910
rect 37840 104880 37900 104910
rect 36000 104820 37190 104850
rect 40060 104830 40120 104860
rect 36040 104760 36120 104770
rect 36220 104760 36300 104770
rect 36400 104760 36480 104770
rect 36580 104760 36660 104770
rect 36760 104760 36840 104770
rect 36940 104760 37020 104770
rect 36120 104680 36130 104760
rect 36300 104680 36310 104760
rect 36480 104680 36490 104760
rect 36660 104680 36670 104760
rect 36840 104680 36850 104760
rect 37020 104680 37030 104760
rect 37100 104620 37190 104820
rect 37720 104790 37750 104820
rect 37840 104790 37870 104820
rect 37600 104760 37660 104790
rect 37720 104760 37780 104790
rect 37840 104760 37900 104790
rect 40060 104710 40120 104740
rect 37720 104670 37750 104700
rect 37840 104670 37870 104700
rect 37600 104640 37660 104670
rect 37720 104640 37780 104670
rect 37840 104640 37900 104670
rect 36000 104590 37190 104620
rect 40060 104590 40120 104620
rect 36120 104530 36130 104590
rect 36300 104530 36310 104590
rect 36480 104530 36490 104590
rect 36660 104530 36670 104590
rect 36840 104530 36850 104590
rect 37020 104530 37030 104590
rect 37100 104520 37190 104590
rect 37720 104550 37750 104580
rect 37840 104550 37870 104580
rect 37600 104520 37660 104550
rect 37720 104520 37780 104550
rect 37840 104520 37900 104550
rect 36000 104490 37190 104520
rect 37100 104480 37190 104490
rect 36000 104470 37190 104480
rect 40060 104470 40120 104500
rect 36040 104290 36120 104300
rect 36220 104290 36300 104300
rect 36400 104290 36480 104300
rect 36580 104290 36660 104300
rect 36760 104290 36840 104300
rect 36940 104290 37020 104300
rect 36120 104210 36130 104290
rect 36300 104210 36310 104290
rect 36480 104210 36490 104290
rect 36660 104210 36670 104290
rect 36840 104210 36850 104290
rect 37020 104210 37030 104290
rect 36040 103970 36120 103980
rect 36220 103970 36300 103980
rect 36400 103970 36480 103980
rect 36580 103970 36660 103980
rect 36760 103970 36840 103980
rect 36940 103970 37020 103980
rect 36120 103890 36130 103970
rect 36300 103890 36310 103970
rect 36480 103890 36490 103970
rect 36660 103890 36670 103970
rect 36840 103890 36850 103970
rect 37020 103890 37030 103970
rect 37100 103800 37190 104470
rect 37720 104430 37750 104460
rect 37840 104430 37870 104460
rect 37600 104400 37660 104430
rect 37720 104400 37780 104430
rect 37840 104400 37900 104430
rect 40060 104350 40120 104380
rect 37720 104310 37750 104340
rect 37840 104310 37870 104340
rect 37600 104280 37660 104310
rect 37720 104280 37780 104310
rect 37840 104280 37900 104310
rect 40060 104230 40120 104260
rect 37720 104190 37750 104220
rect 37840 104190 37870 104220
rect 37600 104160 37660 104190
rect 37720 104160 37780 104190
rect 37840 104160 37900 104190
rect 40060 104110 40120 104140
rect 37720 104070 37750 104100
rect 37840 104070 37870 104100
rect 37600 104040 37660 104070
rect 37720 104040 37780 104070
rect 37840 104040 37900 104070
rect 40060 103990 40120 104020
rect 37720 103950 37750 103980
rect 37840 103950 37870 103980
rect 37600 103920 37660 103950
rect 37720 103920 37780 103950
rect 37840 103920 37900 103950
rect 40060 103870 40120 103900
rect 37720 103830 37750 103860
rect 37840 103830 37870 103860
rect 37600 103800 37660 103830
rect 37720 103800 37780 103830
rect 37840 103800 37900 103830
rect 36000 103790 37190 103800
rect 37100 103690 37190 103790
rect 40060 103750 40120 103780
rect 37720 103710 37750 103740
rect 37840 103710 37870 103740
rect 36000 103660 37190 103690
rect 37600 103680 37660 103710
rect 37720 103680 37780 103710
rect 37840 103680 37900 103710
rect 36040 103650 36120 103660
rect 36220 103650 36300 103660
rect 36400 103650 36480 103660
rect 36580 103650 36660 103660
rect 36760 103650 36840 103660
rect 36940 103650 37020 103660
rect 36120 103590 36130 103650
rect 36300 103590 36310 103650
rect 36480 103590 36490 103650
rect 36660 103590 36670 103650
rect 36840 103590 36850 103650
rect 37020 103590 37030 103650
rect 37100 103590 37190 103660
rect 40060 103630 40120 103660
rect 37720 103590 37750 103620
rect 37840 103590 37870 103620
rect 36000 103560 37190 103590
rect 37600 103560 37660 103590
rect 37720 103560 37780 103590
rect 37840 103560 37900 103590
rect 36040 103500 36120 103510
rect 36220 103500 36300 103510
rect 36400 103500 36480 103510
rect 36580 103500 36660 103510
rect 36760 103500 36840 103510
rect 36940 103500 37020 103510
rect 36120 103420 36130 103500
rect 36300 103420 36310 103500
rect 36480 103420 36490 103500
rect 36660 103420 36670 103500
rect 36840 103420 36850 103500
rect 37020 103420 37030 103500
rect 36040 103350 36120 103360
rect 36220 103350 36300 103360
rect 36400 103350 36480 103360
rect 36580 103350 36660 103360
rect 36760 103350 36840 103360
rect 36940 103350 37020 103360
rect 36120 103270 36130 103350
rect 36300 103270 36310 103350
rect 36480 103270 36490 103350
rect 36660 103270 36670 103350
rect 36840 103270 36850 103350
rect 37020 103270 37030 103350
rect 37100 103330 37190 103560
rect 40060 103510 40120 103540
rect 37720 103470 37750 103500
rect 37840 103470 37870 103500
rect 37600 103440 37660 103470
rect 37720 103440 37780 103470
rect 37840 103440 37900 103470
rect 40060 103390 40120 103420
rect 37720 103350 37750 103380
rect 37840 103350 37870 103380
rect 37600 103320 37660 103350
rect 37720 103320 37780 103350
rect 37840 103320 37900 103350
rect 40060 103270 40120 103300
rect 19130 103200 19160 103255
rect 19250 103200 19280 103255
rect 26420 103200 26450 103255
rect 26540 103200 26570 103255
rect 30420 103230 30450 103255
rect 30540 103230 30570 103255
rect 37720 103230 37750 103260
rect 37840 103230 37870 103260
rect 30300 103200 30360 103230
rect 30420 103200 30480 103230
rect 30540 103200 30600 103230
rect 37600 103200 37660 103230
rect 37720 103200 37780 103230
rect 37840 103200 37900 103230
rect 40060 103150 40120 103180
rect 30420 103080 30450 103140
rect 30540 103080 30570 103140
rect 37720 103080 37750 103140
rect 37840 103080 37870 103140
rect 40060 103030 40120 103060
rect 18980 102940 19060 102950
rect 19160 102940 19240 102950
rect 19340 102940 19420 102950
rect 19520 102940 19600 102950
rect 19700 102940 19780 102950
rect 19880 102940 19960 102950
rect 20060 102940 20140 102950
rect 20240 102940 20320 102950
rect 20420 102940 20500 102950
rect 20600 102940 20680 102950
rect 20780 102940 20860 102950
rect 20960 102940 21040 102950
rect 21140 102940 21220 102950
rect 21320 102940 21400 102950
rect 21500 102940 21580 102950
rect 21680 102940 21760 102950
rect 21860 102940 21940 102950
rect 22040 102940 22120 102950
rect 22220 102940 22300 102950
rect 22400 102940 22480 102950
rect 22580 102940 22660 102950
rect 22760 102940 22840 102950
rect 22940 102940 23020 102950
rect 23120 102940 23200 102950
rect 23300 102940 23380 102950
rect 23480 102940 23560 102950
rect 23660 102940 23740 102950
rect 23840 102940 23920 102950
rect 24020 102940 24100 102950
rect 24200 102940 24280 102950
rect 24380 102940 24460 102950
rect 24560 102940 24640 102950
rect 24740 102940 24820 102950
rect 24920 102940 25000 102950
rect 25100 102940 25180 102950
rect 25280 102940 25360 102950
rect 25460 102940 25540 102950
rect 25640 102940 25720 102950
rect 25820 102940 25900 102950
rect 26000 102940 26080 102950
rect 26180 102940 26260 102950
rect 26360 102940 26440 102950
rect 26540 102940 26620 102950
rect 30280 102940 30360 102950
rect 30460 102940 30540 102950
rect 30640 102940 30720 102950
rect 30820 102940 30900 102950
rect 31000 102940 31080 102950
rect 31180 102940 31260 102950
rect 31360 102940 31440 102950
rect 31540 102940 31620 102950
rect 31720 102940 31800 102950
rect 31900 102940 31980 102950
rect 32080 102940 32160 102950
rect 32260 102940 32340 102950
rect 32440 102940 32520 102950
rect 32620 102940 32700 102950
rect 32800 102940 32880 102950
rect 32980 102940 33060 102950
rect 33160 102940 33240 102950
rect 33340 102940 33420 102950
rect 33520 102940 33600 102950
rect 33700 102940 33780 102950
rect 33880 102940 33960 102950
rect 34060 102940 34140 102950
rect 34240 102940 34320 102950
rect 34420 102940 34500 102950
rect 34600 102940 34680 102950
rect 34780 102940 34860 102950
rect 34960 102940 35040 102950
rect 35140 102940 35220 102950
rect 35320 102940 35400 102950
rect 35500 102940 35580 102950
rect 35680 102940 35760 102950
rect 35860 102940 35940 102950
rect 36040 102940 36120 102950
rect 36220 102940 36300 102950
rect 36400 102940 36480 102950
rect 36580 102940 36660 102950
rect 36760 102940 36840 102950
rect 36940 102940 37020 102950
rect 37120 102940 37200 102950
rect 37300 102940 37380 102950
rect 37480 102940 37560 102950
rect 37660 102940 37740 102950
rect 37840 102940 37920 102950
rect 40260 102940 40270 104940
rect 40380 104930 41180 105020
rect 41540 104950 41600 104980
rect 42360 104950 42420 104980
rect 43840 104950 43900 104980
rect 40650 104900 40770 104930
rect 40930 104900 41050 104930
rect 41090 104900 41180 104930
rect 146100 104910 146160 104940
rect 40650 104810 40660 104900
rect 40760 104870 40830 104900
rect 40770 104780 40830 104870
rect 40930 104810 40940 104900
rect 41050 104780 41180 104900
rect 41090 104745 41180 104780
rect 41230 104750 41350 104810
rect 40470 104740 41180 104745
rect 40370 104730 41180 104740
rect 40370 104650 40380 104730
rect 40470 104725 41180 104730
rect 40420 104715 41210 104725
rect 41090 104665 41180 104715
rect 40470 104650 41180 104665
rect 40460 104635 41180 104650
rect 40460 104445 40470 104635
rect 40650 104600 40770 104635
rect 40930 104600 41050 104635
rect 41090 104600 41180 104635
rect 41350 104630 41410 104750
rect 40770 104590 40830 104600
rect 40530 104580 40610 104590
rect 40670 104580 40750 104590
rect 40770 104580 40890 104590
rect 40950 104580 41030 104590
rect 40610 104500 40620 104580
rect 40750 104500 40760 104580
rect 40770 104480 40830 104580
rect 40890 104500 40900 104580
rect 41030 104500 41040 104580
rect 41050 104480 41180 104600
rect 41260 104580 41340 104590
rect 41340 104510 41350 104580
rect 41090 104445 41180 104480
rect 41230 104450 41350 104510
rect 40460 104430 41180 104445
rect 40470 104425 41180 104430
rect 40420 104415 41210 104425
rect 41090 104365 41180 104415
rect 40470 104335 41180 104365
rect 40650 104300 40770 104335
rect 40930 104300 41050 104335
rect 41090 104300 41180 104335
rect 41350 104330 41410 104450
rect 40650 104210 40660 104300
rect 40760 104270 40830 104300
rect 40770 104180 40830 104270
rect 40930 104210 40940 104300
rect 41050 104180 41180 104300
rect 41260 104280 41340 104290
rect 41340 104210 41350 104280
rect 41090 104145 41180 104180
rect 41230 104150 41350 104210
rect 40370 104130 40460 104140
rect 40370 104050 40380 104130
rect 40470 104125 41180 104145
rect 40420 104115 41210 104125
rect 41090 104065 41180 104115
rect 40470 104050 41180 104065
rect 40460 104035 41180 104050
rect 40460 103845 40470 104035
rect 40650 104000 40770 104035
rect 40930 104000 41050 104035
rect 41090 104000 41180 104035
rect 41350 104030 41410 104150
rect 40770 103990 40830 104000
rect 40530 103980 40610 103990
rect 40670 103980 40750 103990
rect 40770 103980 40890 103990
rect 40950 103980 41030 103990
rect 40610 103900 40620 103980
rect 40750 103900 40760 103980
rect 40770 103880 40830 103980
rect 40890 103900 40900 103980
rect 41030 103900 41040 103980
rect 41050 103880 41180 104000
rect 41260 103980 41340 103990
rect 41340 103910 41350 103980
rect 41090 103845 41180 103880
rect 41230 103850 41350 103910
rect 40460 103830 41180 103845
rect 40470 103825 41180 103830
rect 40420 103815 41210 103825
rect 41090 103765 41180 103815
rect 40470 103735 41180 103765
rect 40650 103700 40770 103735
rect 40930 103700 41050 103735
rect 41090 103700 41180 103735
rect 41350 103730 41410 103850
rect 40650 103610 40660 103700
rect 40760 103670 40830 103700
rect 40770 103580 40830 103670
rect 40930 103610 40940 103700
rect 41050 103580 41180 103700
rect 41260 103680 41340 103690
rect 41340 103610 41350 103680
rect 41090 103545 41180 103580
rect 41230 103550 41350 103610
rect 40370 103530 40460 103540
rect 40370 103450 40380 103530
rect 40470 103525 41180 103545
rect 40420 103515 41210 103525
rect 41090 103465 41180 103515
rect 40470 103450 41180 103465
rect 40460 103435 41180 103450
rect 40460 103245 40470 103435
rect 40650 103400 40770 103435
rect 40930 103400 41050 103435
rect 41090 103400 41180 103435
rect 41350 103430 41410 103550
rect 40770 103390 40830 103400
rect 40530 103380 40610 103390
rect 40670 103380 40750 103390
rect 40770 103380 40890 103390
rect 40950 103380 41030 103390
rect 40610 103300 40620 103380
rect 40750 103300 40760 103380
rect 40770 103280 40830 103380
rect 40890 103300 40900 103380
rect 41030 103300 41040 103380
rect 41050 103280 41180 103400
rect 41260 103370 41340 103380
rect 41340 103310 41350 103370
rect 41090 103245 41180 103280
rect 41230 103250 41350 103310
rect 40460 103230 41180 103245
rect 40470 103225 41180 103230
rect 40420 103215 41210 103225
rect 41090 103165 41180 103215
rect 40470 103135 41180 103165
rect 40650 103100 40770 103135
rect 40930 103100 41050 103135
rect 41090 103100 41180 103135
rect 41350 103130 41410 103250
rect 41480 103100 41490 104870
rect 41540 104830 41600 104860
rect 42360 104830 42420 104860
rect 43840 104830 43900 104860
rect 146100 104790 146160 104820
rect 41540 104710 41600 104740
rect 42360 104710 42420 104740
rect 43840 104710 43900 104740
rect 146100 104670 146160 104700
rect 41540 104590 41600 104620
rect 42360 104590 42420 104620
rect 42910 104600 43030 104660
rect 43190 104600 43310 104660
rect 43030 104590 43090 104600
rect 43310 104590 43370 104600
rect 43840 104590 43900 104620
rect 42930 104580 43010 104590
rect 43030 104580 43150 104590
rect 43210 104580 43290 104590
rect 43310 104580 43430 104590
rect 41540 104470 41600 104500
rect 42360 104470 42420 104500
rect 42470 104480 42480 104570
rect 41540 104350 41600 104380
rect 42360 104350 42420 104380
rect 41540 104230 41600 104260
rect 42360 104230 42420 104260
rect 41540 104110 41600 104140
rect 42360 104110 42420 104140
rect 41540 103990 41600 104020
rect 42360 103990 42420 104020
rect 41540 103870 41600 103900
rect 42360 103870 42420 103900
rect 41540 103750 41600 103780
rect 42360 103750 42420 103780
rect 41540 103630 41600 103660
rect 42360 103630 42420 103660
rect 41540 103510 41600 103540
rect 42360 103510 42420 103540
rect 41540 103390 41600 103420
rect 42360 103390 42420 103420
rect 41540 103270 41600 103300
rect 42360 103270 42420 103300
rect 41540 103150 41600 103180
rect 42360 103150 42420 103180
rect 42560 103120 42570 104480
rect 42610 104450 42730 104510
rect 42730 104425 42790 104450
rect 42860 104440 42870 104570
rect 43010 104500 43020 104580
rect 43030 104480 43090 104580
rect 43150 104500 43160 104580
rect 43290 104500 43300 104580
rect 43310 104480 43370 104580
rect 43430 104500 43440 104580
rect 146100 104550 146160 104580
rect 43840 104470 43900 104500
rect 42860 104430 43500 104440
rect 42730 104415 43540 104425
rect 42730 104330 42790 104415
rect 43540 104365 43550 104415
rect 42620 104240 42700 104250
rect 42700 104160 42710 104240
rect 42860 104160 42870 104350
rect 42910 104300 43030 104360
rect 43190 104300 43310 104360
rect 43020 104270 43090 104300
rect 43030 104180 43090 104270
rect 43190 104210 43200 104300
rect 43300 104270 43370 104300
rect 43310 104180 43370 104270
rect 42860 104150 43490 104160
rect 42860 104140 42870 104150
rect 42620 104060 42700 104070
rect 42700 103980 42710 104060
rect 42770 104050 42780 104140
rect 42610 103860 42730 103920
rect 42730 103835 42790 103860
rect 42860 103850 42870 104050
rect 42910 104010 43030 104070
rect 43190 104010 43310 104070
rect 43030 104000 43090 104010
rect 43310 104000 43370 104010
rect 42930 103990 43010 104000
rect 43030 103990 43150 104000
rect 43210 103990 43290 104000
rect 43310 103990 43430 104000
rect 43010 103910 43020 103990
rect 43030 103890 43090 103990
rect 43150 103910 43160 103990
rect 43290 103910 43300 103990
rect 43310 103890 43370 103990
rect 43430 103910 43440 103990
rect 42860 103840 43500 103850
rect 43580 103840 43590 104140
rect 42730 103825 43540 103835
rect 42730 103740 42790 103825
rect 43540 103775 43550 103825
rect 42620 103640 42700 103650
rect 42700 103560 42710 103640
rect 42860 103570 42870 103760
rect 42910 103710 43030 103770
rect 43190 103710 43310 103770
rect 43020 103680 43090 103710
rect 43030 103590 43090 103680
rect 43190 103620 43200 103710
rect 43300 103680 43370 103710
rect 43310 103590 43370 103680
rect 42860 103560 43490 103570
rect 42860 103550 42870 103560
rect 42620 103460 42700 103470
rect 42770 103460 42780 103550
rect 42700 103380 42710 103460
rect 42610 103270 42730 103330
rect 42730 103245 42790 103270
rect 42860 103260 42870 103460
rect 42910 103420 43030 103480
rect 43190 103420 43310 103480
rect 43030 103410 43090 103420
rect 43310 103410 43370 103420
rect 42930 103400 43010 103410
rect 43030 103400 43150 103410
rect 43210 103400 43290 103410
rect 43310 103400 43430 103410
rect 43010 103320 43020 103400
rect 43030 103300 43090 103400
rect 43150 103320 43160 103400
rect 43290 103320 43300 103400
rect 43310 103300 43370 103400
rect 43430 103320 43440 103400
rect 42860 103250 43500 103260
rect 43580 103250 43590 103550
rect 42730 103235 43540 103245
rect 42730 103150 42790 103235
rect 43540 103185 43550 103235
rect 42860 103120 42870 103170
rect 42910 103120 43030 103180
rect 43190 103120 43310 103180
rect 43030 103110 43090 103120
rect 43310 103110 43370 103120
rect 43030 103100 43150 103110
rect 43310 103100 43430 103110
rect 40770 103090 40830 103100
rect 40530 103080 40610 103090
rect 40770 103080 40890 103090
rect 40610 103000 40620 103080
rect 40770 102980 40830 103080
rect 40890 103000 40900 103080
rect 41050 102980 41180 103100
rect 41540 103030 41600 103060
rect 42360 103030 42420 103060
rect 43030 103000 43090 103100
rect 43150 103020 43160 103100
rect 43310 103000 43370 103100
rect 43430 103020 43440 103100
rect 41090 102950 41180 102980
rect 43780 102960 43790 104440
rect 146100 104430 146160 104460
rect 43840 104350 43900 104380
rect 146100 104310 146160 104340
rect 43840 104230 43900 104260
rect 146100 104190 146160 104220
rect 43840 104110 43900 104140
rect 146100 104070 146160 104100
rect 43840 103990 43900 104020
rect 146100 103950 146160 103980
rect 43840 103870 43900 103900
rect 146100 103830 146160 103860
rect 43840 103750 43900 103780
rect 146100 103710 146160 103740
rect 43840 103630 43900 103660
rect 146300 103650 146310 105040
rect 146690 105000 146810 105060
rect 146970 105000 147090 105060
rect 146810 104990 146870 105000
rect 146570 104980 146650 104990
rect 146810 104980 146930 104990
rect 146650 104900 146660 104980
rect 146810 104880 146870 104980
rect 146930 104900 146940 104980
rect 147090 104880 147150 105000
rect 146410 104830 147140 104840
rect 146410 104750 146420 104830
rect 146460 104815 147150 104825
rect 146450 104765 146460 104815
rect 146500 104560 146510 104750
rect 146690 104700 146810 104760
rect 146970 104700 147090 104760
rect 146810 104690 146870 104700
rect 146570 104680 146650 104690
rect 146710 104680 146790 104690
rect 146810 104680 146930 104690
rect 146990 104680 147070 104690
rect 146650 104600 146660 104680
rect 146790 104600 146800 104680
rect 146810 104580 146870 104680
rect 146930 104600 146940 104680
rect 147070 104600 147080 104680
rect 147090 104580 147150 104700
rect 146500 104550 147130 104560
rect 146500 104540 146510 104550
rect 146690 104410 146810 104470
rect 146970 104410 147090 104470
rect 146690 104320 146700 104410
rect 146800 104380 146870 104410
rect 146810 104290 146870 104380
rect 146970 104320 146980 104410
rect 147090 104290 147150 104410
rect 146410 104240 147140 104250
rect 146410 104160 146420 104240
rect 146460 104225 147150 104235
rect 146450 104175 146460 104225
rect 146500 103970 146510 104160
rect 146690 104110 146810 104170
rect 146970 104110 147090 104170
rect 146810 104100 146870 104110
rect 146570 104090 146650 104100
rect 146710 104090 146790 104100
rect 146810 104090 146930 104100
rect 146990 104090 147070 104100
rect 146650 104010 146660 104090
rect 146790 104010 146800 104090
rect 146810 103990 146870 104090
rect 146930 104010 146940 104090
rect 147070 104010 147080 104090
rect 147090 103990 147150 104110
rect 146500 103960 147130 103970
rect 146500 103950 146510 103960
rect 146690 103820 146810 103880
rect 146970 103820 147090 103880
rect 146690 103730 146700 103820
rect 146800 103790 146870 103820
rect 146810 103700 146870 103790
rect 146970 103730 146980 103820
rect 147090 103700 147150 103820
rect 146410 103650 147140 103660
rect 146460 103635 147150 103645
rect 146100 103590 146160 103620
rect 146450 103585 146460 103635
rect 43840 103510 43900 103540
rect 146690 103520 146810 103580
rect 146970 103520 147090 103580
rect 146810 103510 146870 103520
rect 146570 103500 146650 103510
rect 146710 103500 146790 103510
rect 146810 103500 146930 103510
rect 146990 103500 147070 103510
rect 146100 103470 146160 103500
rect 146650 103420 146660 103500
rect 146790 103420 146800 103500
rect 43840 103390 43900 103420
rect 146810 103400 146870 103500
rect 146930 103420 146940 103500
rect 147070 103420 147080 103500
rect 147090 103400 147150 103520
rect 146100 103350 146160 103380
rect 43840 103270 43900 103300
rect 146100 103230 146160 103260
rect 147580 103230 147640 103246
rect 148400 103230 148460 103246
rect 148600 103220 148610 103246
rect 148950 103220 149070 103246
rect 149230 103220 149350 103246
rect 149060 103190 149130 103220
rect 43840 103150 43900 103180
rect 146100 103110 146160 103140
rect 147580 103110 147640 103140
rect 148400 103110 148460 103140
rect 149070 103100 149130 103190
rect 149230 103130 149240 103220
rect 149340 103190 149410 103220
rect 149350 103100 149410 103190
rect 149530 103070 149620 103246
rect 149820 103060 149830 103246
rect 149880 103230 149940 103246
rect 152220 103210 152250 103240
rect 152340 103210 152370 103240
rect 159520 103210 159550 103240
rect 159640 103210 159670 103240
rect 163520 103210 163550 103240
rect 163640 103210 163670 103240
rect 163960 103235 164040 103245
rect 152100 103180 152160 103210
rect 152220 103180 152280 103210
rect 152340 103180 152400 103210
rect 159400 103180 159460 103210
rect 159520 103180 159580 103210
rect 159640 103180 159700 103210
rect 163400 103180 163460 103210
rect 163520 103180 163580 103210
rect 163640 103180 163700 103210
rect 164040 103155 164050 103235
rect 170810 103210 170840 103240
rect 170930 103210 170960 103240
rect 170690 103180 170750 103210
rect 170810 103180 170870 103210
rect 170930 103180 170990 103210
rect 149880 103110 149940 103140
rect 152220 103060 152250 103120
rect 152340 103060 152370 103120
rect 159520 103060 159550 103120
rect 159640 103060 159670 103120
rect 163520 103060 163550 103120
rect 163640 103060 163670 103120
rect 170810 103060 170840 103120
rect 170930 103060 170960 103120
rect 43840 103030 43900 103060
rect 146100 102990 146160 103020
rect 147580 102990 147640 103020
rect 148400 102990 148460 103020
rect 149880 102990 149940 103020
rect 19060 102860 19070 102940
rect 19240 102860 19250 102940
rect 19420 102860 19430 102940
rect 19600 102860 19610 102940
rect 19780 102860 19790 102940
rect 19960 102860 19970 102940
rect 20140 102860 20150 102940
rect 20320 102860 20330 102940
rect 20500 102860 20510 102940
rect 20680 102860 20690 102940
rect 20860 102860 20870 102940
rect 21040 102860 21050 102940
rect 21220 102860 21230 102940
rect 21400 102860 21410 102940
rect 21580 102860 21590 102940
rect 21760 102860 21770 102940
rect 21940 102860 21950 102940
rect 22120 102860 22130 102940
rect 22300 102860 22310 102940
rect 22480 102860 22490 102940
rect 22660 102860 22670 102940
rect 22840 102860 22850 102940
rect 23020 102860 23030 102940
rect 23200 102860 23210 102940
rect 23380 102860 23390 102940
rect 23560 102860 23570 102940
rect 23740 102860 23750 102940
rect 23920 102860 23930 102940
rect 24100 102860 24110 102940
rect 24280 102860 24290 102940
rect 24460 102860 24470 102940
rect 24640 102860 24650 102940
rect 24820 102860 24830 102940
rect 25000 102860 25010 102940
rect 25180 102860 25190 102940
rect 25360 102860 25370 102940
rect 25540 102860 25550 102940
rect 25720 102860 25730 102940
rect 25900 102860 25910 102940
rect 26080 102860 26090 102940
rect 26260 102860 26270 102940
rect 26440 102860 26450 102940
rect 26620 102860 26630 102940
rect 27315 102915 27395 102925
rect 27495 102915 27575 102925
rect 27675 102915 27755 102925
rect 27855 102915 27935 102925
rect 28035 102915 28115 102925
rect 27395 102835 27405 102915
rect 27575 102835 27585 102915
rect 27755 102835 27765 102915
rect 27935 102835 27945 102915
rect 28115 102835 28125 102915
rect 30360 102860 30370 102940
rect 30540 102860 30550 102940
rect 30720 102860 30730 102940
rect 30900 102860 30910 102940
rect 31080 102860 31090 102940
rect 31260 102860 31270 102940
rect 31440 102860 31450 102940
rect 31620 102860 31630 102940
rect 31800 102860 31810 102940
rect 31980 102860 31990 102940
rect 32160 102860 32170 102940
rect 32340 102860 32350 102940
rect 32520 102860 32530 102940
rect 32700 102860 32710 102940
rect 32880 102860 32890 102940
rect 33060 102860 33070 102940
rect 33240 102860 33250 102940
rect 33420 102860 33430 102940
rect 33600 102860 33610 102940
rect 33780 102860 33790 102940
rect 33960 102860 33970 102940
rect 34140 102860 34150 102940
rect 34320 102860 34330 102940
rect 34500 102860 34510 102940
rect 34680 102860 34690 102940
rect 34860 102860 34870 102940
rect 35040 102860 35050 102940
rect 35220 102860 35230 102940
rect 35400 102860 35410 102940
rect 35580 102860 35590 102940
rect 35760 102860 35770 102940
rect 35940 102860 35950 102940
rect 36120 102860 36130 102940
rect 36300 102860 36310 102940
rect 36480 102860 36490 102940
rect 36660 102860 36670 102940
rect 36840 102860 36850 102940
rect 37020 102860 37030 102940
rect 37200 102860 37210 102940
rect 37380 102860 37390 102940
rect 37560 102860 37570 102940
rect 37740 102860 37750 102940
rect 37920 102860 37930 102940
rect 40060 102910 40120 102940
rect 41540 102910 41600 102940
rect 42360 102910 42420 102940
rect 43840 102910 43900 102940
rect 146100 102870 146160 102900
rect 147580 102870 147640 102900
rect 148400 102870 148460 102900
rect 149880 102870 149940 102900
rect 18980 102790 19060 102800
rect 19160 102790 19240 102800
rect 19340 102790 19420 102800
rect 19520 102790 19600 102800
rect 19700 102790 19780 102800
rect 19880 102790 19960 102800
rect 20060 102790 20140 102800
rect 20240 102790 20320 102800
rect 20420 102790 20500 102800
rect 20600 102790 20680 102800
rect 20780 102790 20860 102800
rect 20960 102790 21040 102800
rect 21140 102790 21220 102800
rect 21320 102790 21400 102800
rect 21500 102790 21580 102800
rect 21680 102790 21760 102800
rect 21860 102790 21940 102800
rect 22040 102790 22120 102800
rect 22220 102790 22300 102800
rect 22400 102790 22480 102800
rect 22580 102790 22660 102800
rect 22760 102790 22840 102800
rect 22940 102790 23020 102800
rect 23120 102790 23200 102800
rect 23300 102790 23380 102800
rect 23480 102790 23560 102800
rect 23660 102790 23740 102800
rect 23840 102790 23920 102800
rect 24020 102790 24100 102800
rect 24200 102790 24280 102800
rect 24380 102790 24460 102800
rect 24560 102790 24640 102800
rect 24740 102790 24820 102800
rect 24920 102790 25000 102800
rect 25100 102790 25180 102800
rect 25280 102790 25360 102800
rect 25460 102790 25540 102800
rect 25640 102790 25720 102800
rect 25820 102790 25900 102800
rect 26000 102790 26080 102800
rect 26180 102790 26260 102800
rect 26360 102790 26440 102800
rect 26540 102790 26620 102800
rect 30280 102790 30360 102800
rect 30460 102790 30540 102800
rect 30640 102790 30720 102800
rect 30820 102790 30900 102800
rect 31000 102790 31080 102800
rect 31180 102790 31260 102800
rect 31360 102790 31440 102800
rect 31540 102790 31620 102800
rect 31720 102790 31800 102800
rect 31900 102790 31980 102800
rect 32080 102790 32160 102800
rect 32260 102790 32340 102800
rect 32440 102790 32520 102800
rect 32620 102790 32700 102800
rect 32800 102790 32880 102800
rect 32980 102790 33060 102800
rect 33160 102790 33240 102800
rect 33340 102790 33420 102800
rect 33520 102790 33600 102800
rect 33700 102790 33780 102800
rect 33880 102790 33960 102800
rect 34060 102790 34140 102800
rect 34240 102790 34320 102800
rect 34420 102790 34500 102800
rect 34600 102790 34680 102800
rect 34780 102790 34860 102800
rect 34960 102790 35040 102800
rect 35140 102790 35220 102800
rect 35320 102790 35400 102800
rect 35500 102790 35580 102800
rect 35680 102790 35760 102800
rect 35860 102790 35940 102800
rect 36040 102790 36120 102800
rect 36220 102790 36300 102800
rect 36400 102790 36480 102800
rect 36580 102790 36660 102800
rect 36760 102790 36840 102800
rect 36940 102790 37020 102800
rect 37120 102790 37200 102800
rect 37300 102790 37380 102800
rect 37480 102790 37560 102800
rect 37660 102790 37740 102800
rect 37840 102790 37920 102800
rect 152080 102790 152160 102800
rect 152260 102790 152340 102800
rect 152440 102790 152520 102800
rect 152620 102790 152700 102800
rect 152800 102790 152880 102800
rect 152980 102790 153060 102800
rect 153160 102790 153240 102800
rect 153340 102790 153420 102800
rect 153520 102790 153600 102800
rect 153700 102790 153780 102800
rect 153880 102790 153960 102800
rect 154060 102790 154140 102800
rect 154240 102790 154320 102800
rect 154420 102790 154500 102800
rect 154600 102790 154680 102800
rect 154780 102790 154860 102800
rect 154960 102790 155040 102800
rect 155140 102790 155220 102800
rect 155320 102790 155400 102800
rect 155500 102790 155580 102800
rect 155680 102790 155760 102800
rect 155860 102790 155940 102800
rect 156040 102790 156120 102800
rect 156220 102790 156300 102800
rect 156400 102790 156480 102800
rect 156580 102790 156660 102800
rect 156760 102790 156840 102800
rect 156940 102790 157020 102800
rect 157120 102790 157200 102800
rect 157300 102790 157380 102800
rect 157480 102790 157560 102800
rect 157660 102790 157740 102800
rect 157840 102790 157920 102800
rect 158020 102790 158100 102800
rect 158200 102790 158280 102800
rect 158380 102790 158460 102800
rect 158560 102790 158640 102800
rect 158740 102790 158820 102800
rect 158920 102790 159000 102800
rect 159100 102790 159180 102800
rect 159280 102790 159360 102800
rect 159460 102790 159540 102800
rect 159640 102790 159720 102800
rect 163380 102790 163460 102800
rect 163560 102790 163640 102800
rect 163740 102790 163820 102800
rect 163920 102790 164000 102800
rect 164100 102790 164180 102800
rect 164280 102790 164360 102800
rect 164460 102790 164540 102800
rect 164640 102790 164720 102800
rect 164820 102790 164900 102800
rect 165000 102790 165080 102800
rect 165180 102790 165260 102800
rect 165360 102790 165440 102800
rect 165540 102790 165620 102800
rect 165720 102790 165800 102800
rect 165900 102790 165980 102800
rect 166080 102790 166160 102800
rect 166260 102790 166340 102800
rect 166440 102790 166520 102800
rect 166620 102790 166700 102800
rect 166800 102790 166880 102800
rect 166980 102790 167060 102800
rect 167160 102790 167240 102800
rect 167340 102790 167420 102800
rect 167520 102790 167600 102800
rect 167700 102790 167780 102800
rect 167880 102790 167960 102800
rect 168060 102790 168140 102800
rect 168240 102790 168320 102800
rect 168420 102790 168500 102800
rect 168600 102790 168680 102800
rect 168780 102790 168860 102800
rect 168960 102790 169040 102800
rect 169140 102790 169220 102800
rect 169320 102790 169400 102800
rect 169500 102790 169580 102800
rect 169680 102790 169760 102800
rect 169860 102790 169940 102800
rect 170040 102790 170120 102800
rect 170220 102790 170300 102800
rect 170400 102790 170480 102800
rect 170580 102790 170660 102800
rect 170760 102790 170840 102800
rect 170940 102790 171020 102800
rect 19060 102710 19070 102790
rect 19240 102710 19250 102790
rect 19420 102710 19430 102790
rect 19600 102710 19610 102790
rect 19780 102710 19790 102790
rect 19960 102710 19970 102790
rect 20140 102710 20150 102790
rect 20320 102710 20330 102790
rect 20500 102710 20510 102790
rect 20680 102710 20690 102790
rect 20860 102710 20870 102790
rect 21040 102710 21050 102790
rect 21220 102710 21230 102790
rect 21400 102710 21410 102790
rect 21580 102710 21590 102790
rect 21760 102710 21770 102790
rect 21940 102710 21950 102790
rect 22120 102710 22130 102790
rect 22300 102710 22310 102790
rect 22480 102710 22490 102790
rect 22660 102710 22670 102790
rect 22840 102710 22850 102790
rect 23020 102710 23030 102790
rect 23200 102710 23210 102790
rect 23380 102710 23390 102790
rect 23560 102710 23570 102790
rect 23740 102710 23750 102790
rect 23920 102710 23930 102790
rect 24100 102710 24110 102790
rect 24280 102710 24290 102790
rect 24460 102710 24470 102790
rect 24640 102710 24650 102790
rect 24820 102710 24830 102790
rect 25000 102710 25010 102790
rect 25180 102710 25190 102790
rect 25360 102710 25370 102790
rect 25540 102710 25550 102790
rect 25720 102710 25730 102790
rect 25900 102710 25910 102790
rect 26080 102710 26090 102790
rect 26260 102710 26270 102790
rect 26440 102710 26450 102790
rect 26620 102710 26630 102790
rect 27315 102735 27395 102745
rect 27495 102735 27575 102745
rect 27675 102735 27755 102745
rect 27855 102735 27935 102745
rect 28035 102735 28115 102745
rect 27395 102655 27405 102735
rect 27575 102655 27585 102735
rect 27755 102655 27765 102735
rect 27935 102655 27945 102735
rect 28115 102655 28125 102735
rect 30360 102710 30370 102790
rect 30540 102710 30550 102790
rect 30720 102710 30730 102790
rect 30900 102710 30910 102790
rect 31080 102710 31090 102790
rect 31260 102710 31270 102790
rect 31440 102710 31450 102790
rect 31620 102710 31630 102790
rect 31800 102710 31810 102790
rect 31980 102710 31990 102790
rect 32160 102710 32170 102790
rect 32340 102710 32350 102790
rect 32520 102710 32530 102790
rect 32700 102710 32710 102790
rect 32880 102710 32890 102790
rect 33060 102710 33070 102790
rect 33240 102710 33250 102790
rect 33420 102710 33430 102790
rect 33600 102710 33610 102790
rect 33780 102710 33790 102790
rect 33960 102710 33970 102790
rect 34140 102710 34150 102790
rect 34320 102710 34330 102790
rect 34500 102710 34510 102790
rect 34680 102710 34690 102790
rect 34860 102710 34870 102790
rect 35040 102710 35050 102790
rect 35220 102710 35230 102790
rect 35400 102710 35410 102790
rect 35580 102710 35590 102790
rect 35760 102710 35770 102790
rect 35940 102710 35950 102790
rect 36120 102710 36130 102790
rect 36300 102710 36310 102790
rect 36480 102710 36490 102790
rect 36660 102710 36670 102790
rect 36840 102710 36850 102790
rect 37020 102710 37030 102790
rect 37200 102710 37210 102790
rect 37380 102710 37390 102790
rect 37560 102710 37570 102790
rect 37740 102710 37750 102790
rect 37920 102710 37930 102790
rect 152160 102710 152170 102790
rect 152340 102710 152350 102790
rect 152520 102710 152530 102790
rect 152700 102710 152710 102790
rect 152880 102710 152890 102790
rect 153060 102710 153070 102790
rect 153240 102710 153250 102790
rect 153420 102710 153430 102790
rect 153600 102710 153610 102790
rect 153780 102710 153790 102790
rect 153960 102710 153970 102790
rect 154140 102710 154150 102790
rect 154320 102710 154330 102790
rect 154500 102710 154510 102790
rect 154680 102710 154690 102790
rect 154860 102710 154870 102790
rect 155040 102710 155050 102790
rect 155220 102710 155230 102790
rect 155400 102710 155410 102790
rect 155580 102710 155590 102790
rect 155760 102710 155770 102790
rect 155940 102710 155950 102790
rect 156120 102710 156130 102790
rect 156300 102710 156310 102790
rect 156480 102710 156490 102790
rect 156660 102710 156670 102790
rect 156840 102710 156850 102790
rect 157020 102710 157030 102790
rect 157200 102710 157210 102790
rect 157380 102710 157390 102790
rect 157560 102710 157570 102790
rect 157740 102710 157750 102790
rect 157920 102710 157930 102790
rect 158100 102710 158110 102790
rect 158280 102710 158290 102790
rect 158460 102710 158470 102790
rect 158640 102710 158650 102790
rect 158820 102710 158830 102790
rect 159000 102710 159010 102790
rect 159180 102710 159190 102790
rect 159360 102710 159370 102790
rect 159540 102710 159550 102790
rect 159720 102710 159730 102790
rect 160430 102765 160510 102775
rect 160590 102765 160670 102775
rect 160750 102765 160830 102775
rect 160910 102765 160990 102775
rect 161070 102765 161150 102775
rect 160510 102685 160520 102765
rect 160590 102685 160600 102765
rect 160670 102685 160680 102765
rect 160750 102685 160760 102765
rect 160830 102685 160840 102765
rect 160910 102685 160920 102765
rect 160990 102685 161000 102765
rect 161070 102685 161080 102765
rect 161150 102685 161160 102765
rect 163460 102710 163470 102790
rect 163640 102710 163650 102790
rect 163820 102710 163830 102790
rect 164000 102710 164010 102790
rect 164180 102710 164190 102790
rect 164360 102710 164370 102790
rect 164540 102710 164550 102790
rect 164720 102710 164730 102790
rect 164900 102710 164910 102790
rect 165080 102710 165090 102790
rect 165260 102710 165270 102790
rect 165440 102710 165450 102790
rect 165620 102710 165630 102790
rect 165800 102710 165810 102790
rect 165980 102710 165990 102790
rect 166160 102710 166170 102790
rect 166340 102710 166350 102790
rect 166520 102710 166530 102790
rect 166700 102710 166710 102790
rect 166880 102710 166890 102790
rect 167060 102710 167070 102790
rect 167240 102710 167250 102790
rect 167420 102710 167430 102790
rect 167600 102710 167610 102790
rect 167780 102710 167790 102790
rect 167960 102710 167970 102790
rect 168140 102710 168150 102790
rect 168320 102710 168330 102790
rect 168500 102710 168510 102790
rect 168680 102710 168690 102790
rect 168860 102710 168870 102790
rect 169040 102710 169050 102790
rect 169220 102710 169230 102790
rect 169400 102710 169410 102790
rect 169580 102710 169590 102790
rect 169760 102710 169770 102790
rect 169940 102710 169950 102790
rect 170120 102710 170130 102790
rect 170300 102710 170310 102790
rect 170480 102710 170490 102790
rect 170660 102710 170670 102790
rect 170840 102710 170850 102790
rect 171020 102710 171030 102790
rect 18980 102640 19060 102650
rect 19160 102640 19240 102650
rect 19340 102640 19420 102650
rect 19520 102640 19600 102650
rect 19700 102640 19780 102650
rect 19880 102640 19960 102650
rect 20060 102640 20140 102650
rect 20240 102640 20320 102650
rect 20420 102640 20500 102650
rect 20600 102640 20680 102650
rect 20780 102640 20860 102650
rect 20960 102640 21040 102650
rect 21140 102640 21220 102650
rect 21320 102640 21400 102650
rect 21500 102640 21580 102650
rect 21680 102640 21760 102650
rect 21860 102640 21940 102650
rect 22040 102640 22120 102650
rect 22220 102640 22300 102650
rect 22400 102640 22480 102650
rect 22580 102640 22660 102650
rect 22760 102640 22840 102650
rect 22940 102640 23020 102650
rect 23120 102640 23200 102650
rect 23300 102640 23380 102650
rect 23480 102640 23560 102650
rect 23660 102640 23740 102650
rect 23840 102640 23920 102650
rect 24020 102640 24100 102650
rect 24200 102640 24280 102650
rect 24380 102640 24460 102650
rect 24560 102640 24640 102650
rect 24740 102640 24820 102650
rect 24920 102640 25000 102650
rect 25100 102640 25180 102650
rect 25280 102640 25360 102650
rect 25460 102640 25540 102650
rect 25640 102640 25720 102650
rect 25820 102640 25900 102650
rect 26000 102640 26080 102650
rect 26180 102640 26260 102650
rect 26360 102640 26440 102650
rect 26540 102640 26620 102650
rect 30280 102640 30360 102650
rect 30460 102640 30540 102650
rect 30640 102640 30720 102650
rect 30820 102640 30900 102650
rect 31000 102640 31080 102650
rect 31180 102640 31260 102650
rect 31360 102640 31440 102650
rect 31540 102640 31620 102650
rect 31720 102640 31800 102650
rect 31900 102640 31980 102650
rect 32080 102640 32160 102650
rect 32260 102640 32340 102650
rect 32440 102640 32520 102650
rect 32620 102640 32700 102650
rect 32800 102640 32880 102650
rect 32980 102640 33060 102650
rect 33160 102640 33240 102650
rect 33340 102640 33420 102650
rect 33520 102640 33600 102650
rect 33700 102640 33780 102650
rect 33880 102640 33960 102650
rect 34060 102640 34140 102650
rect 34240 102640 34320 102650
rect 34420 102640 34500 102650
rect 34600 102640 34680 102650
rect 34780 102640 34860 102650
rect 34960 102640 35040 102650
rect 35140 102640 35220 102650
rect 35320 102640 35400 102650
rect 35500 102640 35580 102650
rect 35680 102640 35760 102650
rect 35860 102640 35940 102650
rect 36040 102640 36120 102650
rect 36220 102640 36300 102650
rect 36400 102640 36480 102650
rect 36580 102640 36660 102650
rect 36760 102640 36840 102650
rect 36940 102640 37020 102650
rect 37120 102640 37200 102650
rect 37300 102640 37380 102650
rect 37480 102640 37560 102650
rect 37660 102640 37740 102650
rect 37840 102640 37920 102650
rect 40060 102640 40140 102650
rect 40200 102640 40280 102650
rect 40340 102640 40420 102650
rect 40480 102640 40560 102650
rect 40620 102640 40700 102650
rect 40760 102640 40840 102650
rect 40900 102640 40980 102650
rect 41040 102640 41120 102650
rect 41180 102640 41260 102650
rect 41320 102640 41400 102650
rect 42360 102640 42440 102650
rect 42500 102640 42580 102650
rect 42640 102640 42720 102650
rect 42780 102640 42860 102650
rect 42920 102640 43000 102650
rect 43060 102640 43140 102650
rect 43200 102640 43280 102650
rect 43340 102640 43420 102650
rect 43480 102640 43560 102650
rect 43620 102640 43700 102650
rect 146300 102640 146380 102650
rect 146440 102640 146520 102650
rect 146580 102640 146660 102650
rect 146720 102640 146800 102650
rect 146860 102640 146940 102650
rect 147000 102640 147080 102650
rect 147140 102640 147220 102650
rect 147280 102640 147360 102650
rect 147420 102640 147500 102650
rect 147560 102640 147640 102650
rect 148600 102640 148680 102650
rect 148740 102640 148820 102650
rect 148880 102640 148960 102650
rect 149020 102640 149100 102650
rect 149160 102640 149240 102650
rect 149300 102640 149380 102650
rect 149440 102640 149520 102650
rect 149580 102640 149660 102650
rect 149720 102640 149800 102650
rect 149860 102640 149940 102650
rect 152080 102640 152160 102650
rect 152260 102640 152340 102650
rect 152440 102640 152520 102650
rect 152620 102640 152700 102650
rect 152800 102640 152880 102650
rect 152980 102640 153060 102650
rect 153160 102640 153240 102650
rect 153340 102640 153420 102650
rect 153520 102640 153600 102650
rect 153700 102640 153780 102650
rect 153880 102640 153960 102650
rect 154060 102640 154140 102650
rect 154240 102640 154320 102650
rect 154420 102640 154500 102650
rect 154600 102640 154680 102650
rect 154780 102640 154860 102650
rect 154960 102640 155040 102650
rect 155140 102640 155220 102650
rect 155320 102640 155400 102650
rect 155500 102640 155580 102650
rect 155680 102640 155760 102650
rect 155860 102640 155940 102650
rect 156040 102640 156120 102650
rect 156220 102640 156300 102650
rect 156400 102640 156480 102650
rect 156580 102640 156660 102650
rect 156760 102640 156840 102650
rect 156940 102640 157020 102650
rect 157120 102640 157200 102650
rect 157300 102640 157380 102650
rect 157480 102640 157560 102650
rect 157660 102640 157740 102650
rect 157840 102640 157920 102650
rect 158020 102640 158100 102650
rect 158200 102640 158280 102650
rect 158380 102640 158460 102650
rect 158560 102640 158640 102650
rect 158740 102640 158820 102650
rect 158920 102640 159000 102650
rect 159100 102640 159180 102650
rect 159280 102640 159360 102650
rect 159460 102640 159540 102650
rect 159640 102640 159720 102650
rect 163380 102640 163460 102650
rect 163560 102640 163640 102650
rect 163740 102640 163820 102650
rect 163920 102640 164000 102650
rect 164100 102640 164180 102650
rect 164280 102640 164360 102650
rect 164460 102640 164540 102650
rect 164640 102640 164720 102650
rect 164820 102640 164900 102650
rect 165000 102640 165080 102650
rect 165180 102640 165260 102650
rect 165360 102640 165440 102650
rect 165540 102640 165620 102650
rect 165720 102640 165800 102650
rect 165900 102640 165980 102650
rect 166080 102640 166160 102650
rect 166260 102640 166340 102650
rect 166440 102640 166520 102650
rect 166620 102640 166700 102650
rect 166800 102640 166880 102650
rect 166980 102640 167060 102650
rect 167160 102640 167240 102650
rect 167340 102640 167420 102650
rect 167520 102640 167600 102650
rect 167700 102640 167780 102650
rect 167880 102640 167960 102650
rect 168060 102640 168140 102650
rect 168240 102640 168320 102650
rect 168420 102640 168500 102650
rect 168600 102640 168680 102650
rect 168780 102640 168860 102650
rect 168960 102640 169040 102650
rect 169140 102640 169220 102650
rect 169320 102640 169400 102650
rect 169500 102640 169580 102650
rect 169680 102640 169760 102650
rect 169860 102640 169940 102650
rect 170040 102640 170120 102650
rect 170220 102640 170300 102650
rect 170400 102640 170480 102650
rect 170580 102640 170660 102650
rect 170760 102640 170840 102650
rect 170940 102640 171020 102650
rect 19060 102560 19070 102640
rect 19240 102560 19250 102640
rect 19420 102560 19430 102640
rect 19600 102560 19610 102640
rect 19780 102560 19790 102640
rect 19960 102560 19970 102640
rect 20140 102560 20150 102640
rect 20320 102560 20330 102640
rect 20500 102560 20510 102640
rect 20680 102560 20690 102640
rect 20860 102560 20870 102640
rect 21040 102560 21050 102640
rect 21220 102560 21230 102640
rect 21400 102560 21410 102640
rect 21580 102560 21590 102640
rect 21760 102560 21770 102640
rect 21940 102560 21950 102640
rect 22120 102560 22130 102640
rect 22300 102560 22310 102640
rect 22480 102560 22490 102640
rect 22660 102560 22670 102640
rect 22840 102560 22850 102640
rect 23020 102560 23030 102640
rect 23200 102560 23210 102640
rect 23380 102560 23390 102640
rect 23560 102560 23570 102640
rect 23740 102560 23750 102640
rect 23920 102560 23930 102640
rect 24100 102560 24110 102640
rect 24280 102560 24290 102640
rect 24460 102560 24470 102640
rect 24640 102560 24650 102640
rect 24820 102560 24830 102640
rect 25000 102560 25010 102640
rect 25180 102560 25190 102640
rect 25360 102560 25370 102640
rect 25540 102560 25550 102640
rect 25720 102560 25730 102640
rect 25900 102560 25910 102640
rect 26080 102560 26090 102640
rect 26260 102560 26270 102640
rect 26440 102560 26450 102640
rect 26620 102560 26630 102640
rect 30360 102560 30370 102640
rect 30540 102560 30550 102640
rect 30720 102560 30730 102640
rect 30900 102560 30910 102640
rect 31080 102560 31090 102640
rect 31260 102560 31270 102640
rect 31440 102560 31450 102640
rect 31620 102560 31630 102640
rect 31800 102560 31810 102640
rect 31980 102560 31990 102640
rect 32160 102560 32170 102640
rect 32340 102560 32350 102640
rect 32520 102560 32530 102640
rect 32700 102560 32710 102640
rect 32880 102560 32890 102640
rect 33060 102560 33070 102640
rect 33240 102560 33250 102640
rect 33420 102560 33430 102640
rect 33600 102560 33610 102640
rect 33780 102560 33790 102640
rect 33960 102560 33970 102640
rect 34140 102560 34150 102640
rect 34320 102560 34330 102640
rect 34500 102560 34510 102640
rect 34680 102560 34690 102640
rect 34860 102560 34870 102640
rect 35040 102560 35050 102640
rect 35220 102560 35230 102640
rect 35400 102560 35410 102640
rect 35580 102560 35590 102640
rect 35760 102560 35770 102640
rect 35940 102560 35950 102640
rect 36120 102560 36130 102640
rect 36300 102560 36310 102640
rect 36480 102560 36490 102640
rect 36660 102560 36670 102640
rect 36840 102560 36850 102640
rect 37020 102560 37030 102640
rect 37200 102560 37210 102640
rect 37380 102560 37390 102640
rect 37560 102560 37570 102640
rect 37740 102560 37750 102640
rect 37920 102560 37930 102640
rect 40140 102560 40150 102640
rect 40280 102560 40290 102640
rect 40420 102560 40430 102640
rect 40560 102560 40570 102640
rect 40700 102560 40710 102640
rect 40840 102560 40850 102640
rect 40980 102560 40990 102640
rect 41120 102560 41130 102640
rect 41260 102560 41270 102640
rect 41400 102560 41410 102640
rect 42440 102560 42450 102640
rect 42580 102560 42590 102640
rect 42720 102560 42730 102640
rect 42860 102560 42870 102640
rect 43000 102560 43010 102640
rect 43140 102560 43150 102640
rect 43280 102560 43290 102640
rect 43420 102560 43430 102640
rect 43560 102560 43570 102640
rect 43700 102560 43710 102640
rect 146380 102581 146390 102640
rect 146520 102581 146530 102640
rect 146660 102581 146670 102640
rect 146800 102581 146810 102640
rect 146940 102581 146950 102640
rect 147080 102581 147090 102640
rect 147220 102581 147230 102640
rect 147360 102581 147370 102640
rect 147500 102581 147510 102640
rect 147640 102581 147650 102640
rect 148680 102581 148690 102640
rect 148820 102581 148830 102640
rect 148960 102581 148970 102640
rect 149100 102581 149110 102640
rect 149240 102581 149250 102640
rect 149380 102581 149390 102640
rect 149520 102581 149530 102640
rect 149660 102581 149670 102640
rect 149800 102581 149810 102640
rect 149940 102581 149950 102640
rect 152160 102581 152170 102640
rect 152340 102581 152350 102640
rect 152520 102581 152530 102640
rect 152700 102581 152710 102640
rect 152880 102581 152890 102640
rect 153060 102581 153070 102640
rect 153240 102581 153250 102640
rect 153420 102581 153430 102640
rect 153600 102581 153610 102640
rect 153780 102581 153790 102640
rect 153960 102581 153970 102640
rect 154140 102581 154150 102640
rect 154320 102581 154330 102640
rect 154500 102581 154510 102640
rect 154680 102581 154690 102640
rect 154860 102581 154870 102640
rect 155040 102581 155050 102640
rect 155220 102581 155230 102640
rect 155400 102581 155410 102640
rect 155580 102581 155590 102640
rect 155760 102581 155770 102640
rect 155940 102581 155950 102640
rect 156120 102581 156130 102640
rect 156300 102581 156310 102640
rect 156480 102581 156490 102640
rect 156660 102581 156670 102640
rect 156840 102581 156850 102640
rect 157020 102581 157030 102640
rect 157200 102581 157210 102640
rect 157380 102581 157390 102640
rect 157560 102581 157570 102640
rect 157740 102581 157750 102640
rect 157920 102581 157930 102640
rect 158100 102581 158110 102640
rect 158280 102581 158290 102640
rect 158460 102581 158470 102640
rect 158640 102581 158650 102640
rect 158820 102581 158830 102640
rect 159000 102581 159010 102640
rect 159180 102581 159190 102640
rect 159360 102581 159370 102640
rect 159540 102581 159550 102640
rect 159720 102581 159730 102640
rect 163460 102581 163470 102640
rect 163640 102581 163650 102640
rect 163820 102581 163830 102640
rect 164000 102581 164010 102640
rect 164180 102581 164190 102640
rect 164360 102581 164370 102640
rect 164540 102581 164550 102640
rect 164720 102581 164730 102640
rect 164900 102581 164910 102640
rect 165080 102581 165090 102640
rect 165260 102581 165270 102640
rect 165440 102581 165450 102640
rect 165620 102581 165630 102640
rect 165800 102581 165810 102640
rect 165980 102581 165990 102640
rect 166160 102581 166170 102640
rect 166340 102581 166350 102640
rect 166520 102581 166530 102640
rect 166700 102581 166710 102640
rect 166880 102581 166890 102640
rect 167060 102581 167070 102640
rect 167240 102581 167250 102640
rect 167420 102581 167430 102640
rect 167600 102581 167610 102640
rect 167780 102581 167790 102640
rect 167960 102581 167970 102640
rect 168140 102581 168150 102640
rect 168320 102581 168330 102640
rect 168500 102581 168510 102640
rect 168680 102581 168690 102640
rect 168860 102581 168870 102640
rect 169040 102581 169050 102640
rect 169220 102581 169230 102640
rect 169400 102581 169410 102640
rect 169580 102581 169590 102640
rect 169760 102581 169770 102640
rect 169940 102581 169950 102640
rect 170120 102581 170130 102640
rect 170300 102581 170310 102640
rect 170480 102581 170490 102640
rect 170660 102581 170670 102640
rect 170840 102581 170850 102640
rect 171020 102581 171030 102640
rect 146040 102500 147700 102581
rect 148340 102500 150000 102581
rect 152000 102500 159800 102581
rect 163210 102560 171100 102581
rect 163300 102500 171100 102560
rect 30360 102420 30440 102430
rect 30680 102420 30760 102430
rect 31000 102420 31080 102430
rect 31320 102420 31400 102430
rect 31640 102420 31720 102430
rect 31960 102420 32040 102430
rect 32280 102420 32360 102430
rect 32600 102420 32680 102430
rect 32920 102420 33000 102430
rect 33240 102420 33320 102430
rect 33560 102420 33640 102430
rect 33880 102420 33960 102430
rect 34200 102420 34280 102430
rect 34520 102420 34600 102430
rect 34840 102420 34920 102430
rect 35160 102420 35240 102430
rect 35480 102420 35560 102430
rect 35800 102420 35880 102430
rect 36120 102420 36200 102430
rect 36440 102420 36520 102430
rect 36760 102420 36840 102430
rect 37080 102420 37160 102430
rect 37400 102420 37480 102430
rect 37720 102420 37800 102430
rect 40180 102420 40260 102430
rect 40500 102420 40580 102430
rect 40820 102420 40900 102430
rect 41140 102420 41220 102430
rect 42560 102420 42640 102430
rect 42880 102420 42960 102430
rect 43200 102420 43280 102430
rect 43520 102420 43600 102430
rect 18970 102390 19050 102400
rect 19290 102390 19370 102400
rect 19610 102390 19690 102400
rect 19930 102390 20010 102400
rect 20250 102390 20330 102400
rect 20570 102390 20650 102400
rect 20890 102390 20970 102400
rect 21210 102390 21290 102400
rect 21530 102390 21610 102400
rect 21850 102390 21930 102400
rect 22170 102390 22250 102400
rect 22490 102390 22570 102400
rect 22810 102390 22890 102400
rect 23130 102390 23210 102400
rect 23450 102390 23530 102400
rect 23770 102390 23850 102400
rect 24090 102390 24170 102400
rect 24410 102390 24490 102400
rect 24730 102390 24810 102400
rect 25050 102390 25130 102400
rect 25370 102390 25450 102400
rect 25690 102390 25770 102400
rect 26010 102390 26090 102400
rect 26330 102390 26410 102400
rect 19050 102310 19060 102390
rect 19370 102310 19380 102390
rect 19690 102310 19700 102390
rect 20010 102310 20020 102390
rect 20330 102310 20340 102390
rect 20650 102310 20660 102390
rect 20970 102310 20980 102390
rect 21290 102310 21300 102390
rect 21610 102310 21620 102390
rect 21930 102310 21940 102390
rect 22250 102310 22260 102390
rect 22570 102310 22580 102390
rect 22890 102310 22900 102390
rect 23210 102310 23220 102390
rect 23530 102310 23540 102390
rect 23850 102310 23860 102390
rect 24170 102310 24180 102390
rect 24490 102310 24500 102390
rect 24810 102310 24820 102390
rect 25130 102310 25140 102390
rect 25450 102310 25460 102390
rect 25770 102310 25780 102390
rect 26090 102310 26100 102390
rect 26410 102310 26420 102390
rect 30440 102340 30450 102420
rect 30760 102340 30770 102420
rect 31080 102340 31090 102420
rect 31400 102340 31410 102420
rect 31720 102340 31730 102420
rect 32040 102340 32050 102420
rect 32360 102340 32370 102420
rect 32680 102340 32690 102420
rect 33000 102340 33010 102420
rect 33320 102340 33330 102420
rect 33640 102340 33650 102420
rect 33960 102340 33970 102420
rect 34280 102340 34290 102420
rect 34600 102340 34610 102420
rect 34920 102340 34930 102420
rect 35240 102340 35250 102420
rect 35560 102340 35570 102420
rect 35880 102340 35890 102420
rect 36200 102340 36210 102420
rect 36520 102340 36530 102420
rect 36840 102340 36850 102420
rect 37160 102340 37170 102420
rect 37480 102340 37490 102420
rect 37800 102340 37810 102420
rect 40260 102340 40270 102420
rect 40580 102340 40590 102420
rect 40900 102340 40910 102420
rect 41220 102340 41230 102420
rect 42640 102340 42650 102420
rect 42960 102340 42970 102420
rect 43280 102340 43290 102420
rect 43600 102340 43610 102420
rect 146400 102411 146480 102421
rect 146720 102411 146800 102421
rect 147040 102411 147120 102421
rect 147360 102411 147440 102421
rect 148780 102411 148860 102421
rect 149100 102411 149180 102421
rect 149420 102411 149500 102421
rect 149740 102411 149820 102421
rect 152200 102411 152280 102421
rect 152520 102411 152600 102421
rect 152840 102411 152920 102421
rect 153160 102411 153240 102421
rect 153480 102411 153560 102421
rect 153800 102411 153880 102421
rect 154120 102411 154200 102421
rect 154440 102411 154520 102421
rect 154760 102411 154840 102421
rect 155080 102411 155160 102421
rect 155400 102411 155480 102421
rect 155720 102411 155800 102421
rect 156040 102411 156120 102421
rect 156360 102411 156440 102421
rect 156680 102411 156760 102421
rect 157000 102411 157080 102421
rect 157320 102411 157400 102421
rect 157640 102411 157720 102421
rect 157960 102411 158040 102421
rect 158280 102411 158360 102421
rect 158600 102411 158680 102421
rect 158920 102411 159000 102421
rect 159240 102411 159320 102421
rect 159560 102411 159640 102421
rect 146480 102331 146490 102411
rect 146800 102331 146810 102411
rect 147120 102331 147130 102411
rect 147440 102331 147450 102411
rect 148860 102331 148870 102411
rect 149180 102331 149190 102411
rect 149500 102331 149510 102411
rect 149820 102331 149830 102411
rect 152280 102331 152290 102411
rect 152600 102331 152610 102411
rect 152920 102331 152930 102411
rect 153240 102331 153250 102411
rect 153560 102331 153570 102411
rect 153880 102331 153890 102411
rect 154200 102331 154210 102411
rect 154520 102331 154530 102411
rect 154840 102331 154850 102411
rect 155160 102331 155170 102411
rect 155480 102331 155490 102411
rect 155800 102331 155810 102411
rect 156120 102331 156130 102411
rect 156440 102331 156450 102411
rect 156760 102331 156770 102411
rect 157080 102331 157090 102411
rect 157400 102331 157410 102411
rect 157720 102331 157730 102411
rect 158040 102331 158050 102411
rect 158360 102331 158370 102411
rect 158680 102331 158690 102411
rect 159000 102331 159010 102411
rect 159320 102331 159330 102411
rect 159640 102331 159650 102411
rect 163590 102381 163670 102391
rect 163910 102381 163990 102391
rect 164230 102381 164310 102391
rect 164550 102381 164630 102391
rect 164870 102381 164950 102391
rect 165190 102381 165270 102391
rect 165510 102381 165590 102391
rect 165830 102381 165910 102391
rect 166150 102381 166230 102391
rect 166470 102381 166550 102391
rect 166790 102381 166870 102391
rect 167110 102381 167190 102391
rect 167430 102381 167510 102391
rect 167750 102381 167830 102391
rect 168070 102381 168150 102391
rect 168390 102381 168470 102391
rect 168710 102381 168790 102391
rect 169030 102381 169110 102391
rect 169350 102381 169430 102391
rect 169670 102381 169750 102391
rect 169990 102381 170070 102391
rect 170310 102381 170390 102391
rect 170630 102381 170710 102391
rect 170950 102381 171030 102391
rect 163670 102301 163680 102381
rect 163990 102301 164000 102381
rect 164310 102301 164320 102381
rect 164630 102301 164640 102381
rect 164950 102301 164960 102381
rect 165270 102301 165280 102381
rect 165590 102301 165600 102381
rect 165910 102301 165920 102381
rect 166230 102301 166240 102381
rect 166550 102301 166560 102381
rect 166870 102301 166880 102381
rect 167190 102301 167200 102381
rect 167510 102301 167520 102381
rect 167830 102301 167840 102381
rect 168150 102301 168160 102381
rect 168470 102301 168480 102381
rect 168790 102301 168800 102381
rect 169110 102301 169120 102381
rect 169430 102301 169440 102381
rect 169750 102301 169760 102381
rect 170070 102301 170080 102381
rect 170390 102301 170400 102381
rect 170710 102301 170720 102381
rect 171030 102301 171040 102381
rect 30520 102260 30600 102270
rect 30840 102260 30920 102270
rect 31160 102260 31240 102270
rect 31480 102260 31560 102270
rect 31800 102260 31880 102270
rect 32120 102260 32200 102270
rect 32440 102260 32520 102270
rect 32760 102260 32840 102270
rect 33080 102260 33160 102270
rect 33400 102260 33480 102270
rect 33720 102260 33800 102270
rect 34040 102260 34120 102270
rect 34360 102260 34440 102270
rect 34680 102260 34760 102270
rect 35000 102260 35080 102270
rect 35320 102260 35400 102270
rect 35640 102260 35720 102270
rect 35960 102260 36040 102270
rect 36280 102260 36360 102270
rect 36600 102260 36680 102270
rect 36920 102260 37000 102270
rect 37240 102260 37320 102270
rect 37560 102260 37640 102270
rect 40340 102260 40420 102270
rect 40660 102260 40740 102270
rect 40980 102260 41060 102270
rect 42720 102260 42800 102270
rect 43040 102260 43120 102270
rect 43360 102260 43440 102270
rect 19130 102230 19210 102240
rect 19450 102230 19530 102240
rect 19770 102230 19850 102240
rect 20090 102230 20170 102240
rect 20410 102230 20490 102240
rect 20730 102230 20810 102240
rect 21050 102230 21130 102240
rect 21370 102230 21450 102240
rect 21690 102230 21770 102240
rect 22010 102230 22090 102240
rect 22330 102230 22410 102240
rect 22650 102230 22730 102240
rect 22970 102230 23050 102240
rect 23290 102230 23370 102240
rect 23610 102230 23690 102240
rect 23930 102230 24010 102240
rect 24250 102230 24330 102240
rect 24570 102230 24650 102240
rect 24890 102230 24970 102240
rect 25210 102230 25290 102240
rect 25530 102230 25610 102240
rect 25850 102230 25930 102240
rect 26170 102230 26250 102240
rect 19210 102150 19220 102230
rect 19530 102150 19540 102230
rect 19850 102150 19860 102230
rect 20170 102150 20180 102230
rect 20490 102150 20500 102230
rect 20810 102150 20820 102230
rect 21130 102150 21140 102230
rect 21450 102150 21460 102230
rect 21770 102150 21780 102230
rect 22090 102150 22100 102230
rect 22410 102150 22420 102230
rect 22730 102150 22740 102230
rect 23050 102150 23060 102230
rect 23370 102150 23380 102230
rect 23690 102150 23700 102230
rect 24010 102150 24020 102230
rect 24330 102150 24340 102230
rect 24650 102150 24660 102230
rect 24970 102150 24980 102230
rect 25290 102150 25300 102230
rect 25610 102150 25620 102230
rect 25930 102150 25940 102230
rect 26250 102150 26260 102230
rect 30600 102180 30610 102260
rect 30920 102180 30930 102260
rect 31240 102180 31250 102260
rect 31560 102180 31570 102260
rect 31880 102180 31890 102260
rect 32200 102180 32210 102260
rect 32520 102180 32530 102260
rect 32840 102180 32850 102260
rect 33160 102180 33170 102260
rect 33480 102180 33490 102260
rect 33800 102180 33810 102260
rect 34120 102180 34130 102260
rect 34440 102180 34450 102260
rect 34760 102180 34770 102260
rect 35080 102180 35090 102260
rect 35400 102180 35410 102260
rect 35720 102180 35730 102260
rect 36040 102180 36050 102260
rect 36360 102180 36370 102260
rect 36680 102180 36690 102260
rect 37000 102180 37010 102260
rect 37320 102180 37330 102260
rect 37640 102180 37650 102260
rect 40420 102180 40430 102260
rect 40740 102180 40750 102260
rect 41060 102180 41070 102260
rect 42800 102180 42810 102260
rect 43120 102180 43130 102260
rect 43440 102180 43450 102260
rect 146560 102251 146640 102261
rect 146880 102251 146960 102261
rect 147200 102251 147280 102261
rect 148940 102251 149020 102261
rect 149260 102251 149340 102261
rect 149580 102251 149660 102261
rect 152360 102251 152440 102261
rect 152680 102251 152760 102261
rect 153000 102251 153080 102261
rect 153320 102251 153400 102261
rect 153640 102251 153720 102261
rect 153960 102251 154040 102261
rect 154280 102251 154360 102261
rect 154600 102251 154680 102261
rect 154920 102251 155000 102261
rect 155240 102251 155320 102261
rect 155560 102251 155640 102261
rect 155880 102251 155960 102261
rect 156200 102251 156280 102261
rect 156520 102251 156600 102261
rect 156840 102251 156920 102261
rect 157160 102251 157240 102261
rect 157480 102251 157560 102261
rect 157800 102251 157880 102261
rect 158120 102251 158200 102261
rect 158440 102251 158520 102261
rect 158760 102251 158840 102261
rect 159080 102251 159160 102261
rect 159400 102251 159480 102261
rect 146640 102171 146650 102251
rect 146960 102171 146970 102251
rect 147280 102171 147290 102251
rect 149020 102171 149030 102251
rect 149340 102171 149350 102251
rect 149660 102171 149670 102251
rect 152440 102171 152450 102251
rect 152760 102171 152770 102251
rect 153080 102171 153090 102251
rect 153400 102171 153410 102251
rect 153720 102171 153730 102251
rect 154040 102171 154050 102251
rect 154360 102171 154370 102251
rect 154680 102171 154690 102251
rect 155000 102171 155010 102251
rect 155320 102171 155330 102251
rect 155640 102171 155650 102251
rect 155960 102171 155970 102251
rect 156280 102171 156290 102251
rect 156600 102171 156610 102251
rect 156920 102171 156930 102251
rect 157240 102171 157250 102251
rect 157560 102171 157570 102251
rect 157880 102171 157890 102251
rect 158200 102171 158210 102251
rect 158520 102171 158530 102251
rect 158840 102171 158850 102251
rect 159160 102171 159170 102251
rect 159480 102171 159490 102251
rect 163750 102221 163830 102231
rect 164070 102221 164150 102231
rect 164390 102221 164470 102231
rect 164710 102221 164790 102231
rect 165030 102221 165110 102231
rect 165350 102221 165430 102231
rect 165670 102221 165750 102231
rect 165990 102221 166070 102231
rect 166310 102221 166390 102231
rect 166630 102221 166710 102231
rect 166950 102221 167030 102231
rect 167270 102221 167350 102231
rect 167590 102221 167670 102231
rect 167910 102221 167990 102231
rect 168230 102221 168310 102231
rect 168550 102221 168630 102231
rect 168870 102221 168950 102231
rect 169190 102221 169270 102231
rect 169510 102221 169590 102231
rect 169830 102221 169910 102231
rect 170150 102221 170230 102231
rect 170470 102221 170550 102231
rect 170790 102221 170870 102231
rect 163830 102141 163840 102221
rect 164150 102141 164160 102221
rect 164470 102141 164480 102221
rect 164790 102141 164800 102221
rect 165110 102141 165120 102221
rect 165430 102141 165440 102221
rect 165750 102141 165760 102221
rect 166070 102141 166080 102221
rect 166390 102141 166400 102221
rect 166710 102141 166720 102221
rect 167030 102141 167040 102221
rect 167350 102141 167360 102221
rect 167670 102141 167680 102221
rect 167990 102141 168000 102221
rect 168310 102141 168320 102221
rect 168630 102141 168640 102221
rect 168950 102141 168960 102221
rect 169270 102141 169280 102221
rect 169590 102141 169600 102221
rect 169910 102141 169920 102221
rect 170230 102141 170240 102221
rect 170550 102141 170560 102221
rect 170870 102141 170880 102221
rect 30360 102100 30440 102110
rect 30680 102100 30760 102110
rect 31000 102100 31080 102110
rect 31320 102100 31400 102110
rect 31640 102100 31720 102110
rect 31960 102100 32040 102110
rect 32280 102100 32360 102110
rect 32600 102100 32680 102110
rect 32920 102100 33000 102110
rect 33240 102100 33320 102110
rect 33560 102100 33640 102110
rect 33880 102100 33960 102110
rect 34200 102100 34280 102110
rect 34520 102100 34600 102110
rect 34840 102100 34920 102110
rect 35160 102100 35240 102110
rect 35480 102100 35560 102110
rect 35800 102100 35880 102110
rect 36120 102100 36200 102110
rect 36440 102100 36520 102110
rect 36760 102100 36840 102110
rect 37080 102100 37160 102110
rect 37400 102100 37480 102110
rect 37720 102100 37800 102110
rect 40180 102100 40260 102110
rect 40500 102100 40580 102110
rect 40820 102100 40900 102110
rect 41140 102100 41220 102110
rect 42560 102100 42640 102110
rect 42880 102100 42960 102110
rect 43200 102100 43280 102110
rect 43520 102100 43600 102110
rect 18970 102070 19050 102080
rect 19290 102070 19370 102080
rect 19610 102070 19690 102080
rect 19930 102070 20010 102080
rect 20250 102070 20330 102080
rect 20570 102070 20650 102080
rect 20890 102070 20970 102080
rect 21210 102070 21290 102080
rect 21530 102070 21610 102080
rect 21850 102070 21930 102080
rect 22170 102070 22250 102080
rect 22490 102070 22570 102080
rect 22810 102070 22890 102080
rect 23130 102070 23210 102080
rect 23450 102070 23530 102080
rect 23770 102070 23850 102080
rect 24090 102070 24170 102080
rect 24410 102070 24490 102080
rect 24730 102070 24810 102080
rect 25050 102070 25130 102080
rect 25370 102070 25450 102080
rect 25690 102070 25770 102080
rect 26010 102070 26090 102080
rect 26330 102070 26410 102080
rect 19050 101990 19060 102070
rect 19370 101990 19380 102070
rect 19690 101990 19700 102070
rect 20010 101990 20020 102070
rect 20330 101990 20340 102070
rect 20650 101990 20660 102070
rect 20970 101990 20980 102070
rect 21290 101990 21300 102070
rect 21610 101990 21620 102070
rect 21930 101990 21940 102070
rect 22250 101990 22260 102070
rect 22570 101990 22580 102070
rect 22890 101990 22900 102070
rect 23210 101990 23220 102070
rect 23530 101990 23540 102070
rect 23850 101990 23860 102070
rect 24170 101990 24180 102070
rect 24490 101990 24500 102070
rect 24810 101990 24820 102070
rect 25130 101990 25140 102070
rect 25450 101990 25460 102070
rect 25770 101990 25780 102070
rect 26090 101990 26100 102070
rect 26410 101990 26420 102070
rect 30440 102020 30450 102100
rect 30760 102020 30770 102100
rect 31080 102020 31090 102100
rect 31400 102020 31410 102100
rect 31720 102020 31730 102100
rect 32040 102020 32050 102100
rect 32360 102020 32370 102100
rect 32680 102020 32690 102100
rect 33000 102020 33010 102100
rect 33320 102020 33330 102100
rect 33640 102020 33650 102100
rect 33960 102020 33970 102100
rect 34280 102020 34290 102100
rect 34600 102020 34610 102100
rect 34920 102020 34930 102100
rect 35240 102020 35250 102100
rect 35560 102020 35570 102100
rect 35880 102020 35890 102100
rect 36200 102020 36210 102100
rect 36520 102020 36530 102100
rect 36840 102020 36850 102100
rect 37160 102020 37170 102100
rect 37480 102020 37490 102100
rect 37800 102020 37810 102100
rect 40260 102020 40270 102100
rect 40580 102020 40590 102100
rect 40900 102020 40910 102100
rect 41220 102020 41230 102100
rect 42640 102020 42650 102100
rect 42960 102020 42970 102100
rect 43280 102020 43290 102100
rect 43600 102020 43610 102100
rect 146400 102091 146480 102101
rect 146720 102091 146800 102101
rect 147040 102091 147120 102101
rect 147360 102091 147440 102101
rect 148780 102091 148860 102101
rect 149100 102091 149180 102101
rect 149420 102091 149500 102101
rect 149740 102091 149820 102101
rect 152200 102091 152280 102101
rect 152520 102091 152600 102101
rect 152840 102091 152920 102101
rect 153160 102091 153240 102101
rect 153480 102091 153560 102101
rect 153800 102091 153880 102101
rect 154120 102091 154200 102101
rect 154440 102091 154520 102101
rect 154760 102091 154840 102101
rect 155080 102091 155160 102101
rect 155400 102091 155480 102101
rect 155720 102091 155800 102101
rect 156040 102091 156120 102101
rect 156360 102091 156440 102101
rect 156680 102091 156760 102101
rect 157000 102091 157080 102101
rect 157320 102091 157400 102101
rect 157640 102091 157720 102101
rect 157960 102091 158040 102101
rect 158280 102091 158360 102101
rect 158600 102091 158680 102101
rect 158920 102091 159000 102101
rect 159240 102091 159320 102101
rect 159560 102091 159640 102101
rect 146480 102011 146490 102091
rect 146800 102011 146810 102091
rect 147120 102011 147130 102091
rect 147440 102011 147450 102091
rect 148860 102011 148870 102091
rect 149180 102011 149190 102091
rect 149500 102011 149510 102091
rect 149820 102011 149830 102091
rect 152280 102011 152290 102091
rect 152600 102011 152610 102091
rect 152920 102011 152930 102091
rect 153240 102011 153250 102091
rect 153560 102011 153570 102091
rect 153880 102011 153890 102091
rect 154200 102011 154210 102091
rect 154520 102011 154530 102091
rect 154840 102011 154850 102091
rect 155160 102011 155170 102091
rect 155480 102011 155490 102091
rect 155800 102011 155810 102091
rect 156120 102011 156130 102091
rect 156440 102011 156450 102091
rect 156760 102011 156770 102091
rect 157080 102011 157090 102091
rect 157400 102011 157410 102091
rect 157720 102011 157730 102091
rect 158040 102011 158050 102091
rect 158360 102011 158370 102091
rect 158680 102011 158690 102091
rect 159000 102011 159010 102091
rect 159320 102011 159330 102091
rect 159640 102011 159650 102091
rect 163590 102061 163670 102071
rect 163910 102061 163990 102071
rect 164230 102061 164310 102071
rect 164550 102061 164630 102071
rect 164870 102061 164950 102071
rect 165190 102061 165270 102071
rect 165510 102061 165590 102071
rect 165830 102061 165910 102071
rect 166150 102061 166230 102071
rect 166470 102061 166550 102071
rect 166790 102061 166870 102071
rect 167110 102061 167190 102071
rect 167430 102061 167510 102071
rect 167750 102061 167830 102071
rect 168070 102061 168150 102071
rect 168390 102061 168470 102071
rect 168710 102061 168790 102071
rect 169030 102061 169110 102071
rect 169350 102061 169430 102071
rect 169670 102061 169750 102071
rect 169990 102061 170070 102071
rect 170310 102061 170390 102071
rect 170630 102061 170710 102071
rect 170950 102061 171030 102071
rect 163670 101981 163680 102061
rect 163990 101981 164000 102061
rect 164310 101981 164320 102061
rect 164630 101981 164640 102061
rect 164950 101981 164960 102061
rect 165270 101981 165280 102061
rect 165590 101981 165600 102061
rect 165910 101981 165920 102061
rect 166230 101981 166240 102061
rect 166550 101981 166560 102061
rect 166870 101981 166880 102061
rect 167190 101981 167200 102061
rect 167510 101981 167520 102061
rect 167830 101981 167840 102061
rect 168150 101981 168160 102061
rect 168470 101981 168480 102061
rect 168790 101981 168800 102061
rect 169110 101981 169120 102061
rect 169430 101981 169440 102061
rect 169750 101981 169760 102061
rect 170070 101981 170080 102061
rect 170390 101981 170400 102061
rect 170710 101981 170720 102061
rect 171030 101981 171040 102061
rect 30520 101940 30600 101950
rect 30840 101940 30920 101950
rect 31160 101940 31240 101950
rect 31480 101940 31560 101950
rect 31800 101940 31880 101950
rect 32120 101940 32200 101950
rect 32440 101940 32520 101950
rect 32760 101940 32840 101950
rect 33080 101940 33160 101950
rect 33400 101940 33480 101950
rect 33720 101940 33800 101950
rect 34040 101940 34120 101950
rect 34360 101940 34440 101950
rect 34680 101940 34760 101950
rect 35000 101940 35080 101950
rect 35320 101940 35400 101950
rect 35640 101940 35720 101950
rect 35960 101940 36040 101950
rect 36280 101940 36360 101950
rect 36600 101940 36680 101950
rect 36920 101940 37000 101950
rect 37240 101940 37320 101950
rect 37560 101940 37640 101950
rect 40340 101940 40420 101950
rect 40660 101940 40740 101950
rect 40980 101940 41060 101950
rect 42720 101940 42800 101950
rect 43040 101940 43120 101950
rect 43360 101940 43440 101950
rect 19130 101910 19210 101920
rect 19450 101910 19530 101920
rect 19770 101910 19850 101920
rect 20090 101910 20170 101920
rect 20410 101910 20490 101920
rect 20730 101910 20810 101920
rect 21050 101910 21130 101920
rect 21370 101910 21450 101920
rect 21690 101910 21770 101920
rect 22010 101910 22090 101920
rect 22330 101910 22410 101920
rect 22650 101910 22730 101920
rect 22970 101910 23050 101920
rect 23290 101910 23370 101920
rect 23610 101910 23690 101920
rect 23930 101910 24010 101920
rect 24250 101910 24330 101920
rect 24570 101910 24650 101920
rect 24890 101910 24970 101920
rect 25210 101910 25290 101920
rect 25530 101910 25610 101920
rect 25850 101910 25930 101920
rect 26170 101910 26250 101920
rect 19210 101830 19220 101910
rect 19530 101830 19540 101910
rect 19850 101830 19860 101910
rect 20170 101830 20180 101910
rect 20490 101830 20500 101910
rect 20810 101830 20820 101910
rect 21130 101830 21140 101910
rect 21450 101830 21460 101910
rect 21770 101830 21780 101910
rect 22090 101830 22100 101910
rect 22410 101830 22420 101910
rect 22730 101830 22740 101910
rect 23050 101830 23060 101910
rect 23370 101830 23380 101910
rect 23690 101830 23700 101910
rect 24010 101830 24020 101910
rect 24330 101830 24340 101910
rect 24650 101830 24660 101910
rect 24970 101830 24980 101910
rect 25290 101830 25300 101910
rect 25610 101830 25620 101910
rect 25930 101830 25940 101910
rect 26250 101830 26260 101910
rect 30600 101860 30610 101940
rect 30920 101860 30930 101940
rect 31240 101860 31250 101940
rect 31560 101860 31570 101940
rect 31880 101860 31890 101940
rect 32200 101860 32210 101940
rect 32520 101860 32530 101940
rect 32840 101860 32850 101940
rect 33160 101860 33170 101940
rect 33480 101860 33490 101940
rect 33800 101860 33810 101940
rect 34120 101860 34130 101940
rect 34440 101860 34450 101940
rect 34760 101860 34770 101940
rect 35080 101860 35090 101940
rect 35400 101860 35410 101940
rect 35720 101860 35730 101940
rect 36040 101860 36050 101940
rect 36360 101860 36370 101940
rect 36680 101860 36690 101940
rect 37000 101860 37010 101940
rect 37320 101860 37330 101940
rect 37640 101860 37650 101940
rect 40420 101860 40430 101940
rect 40740 101860 40750 101940
rect 41060 101860 41070 101940
rect 42800 101860 42810 101940
rect 43120 101860 43130 101940
rect 43440 101860 43450 101940
rect 146560 101931 146640 101941
rect 146880 101931 146960 101941
rect 147200 101931 147280 101941
rect 148940 101931 149020 101941
rect 149260 101931 149340 101941
rect 149580 101931 149660 101941
rect 152360 101931 152440 101941
rect 152680 101931 152760 101941
rect 153000 101931 153080 101941
rect 153320 101931 153400 101941
rect 153640 101931 153720 101941
rect 153960 101931 154040 101941
rect 154280 101931 154360 101941
rect 154600 101931 154680 101941
rect 154920 101931 155000 101941
rect 155240 101931 155320 101941
rect 155560 101931 155640 101941
rect 155880 101931 155960 101941
rect 156200 101931 156280 101941
rect 156520 101931 156600 101941
rect 156840 101931 156920 101941
rect 157160 101931 157240 101941
rect 157480 101931 157560 101941
rect 157800 101931 157880 101941
rect 158120 101931 158200 101941
rect 158440 101931 158520 101941
rect 158760 101931 158840 101941
rect 159080 101931 159160 101941
rect 159400 101931 159480 101941
rect 146640 101851 146650 101931
rect 146960 101851 146970 101931
rect 147280 101851 147290 101931
rect 149020 101851 149030 101931
rect 149340 101851 149350 101931
rect 149660 101851 149670 101931
rect 152440 101851 152450 101931
rect 152760 101851 152770 101931
rect 153080 101851 153090 101931
rect 153400 101851 153410 101931
rect 153720 101851 153730 101931
rect 154040 101851 154050 101931
rect 154360 101851 154370 101931
rect 154680 101851 154690 101931
rect 155000 101851 155010 101931
rect 155320 101851 155330 101931
rect 155640 101851 155650 101931
rect 155960 101851 155970 101931
rect 156280 101851 156290 101931
rect 156600 101851 156610 101931
rect 156920 101851 156930 101931
rect 157240 101851 157250 101931
rect 157560 101851 157570 101931
rect 157880 101851 157890 101931
rect 158200 101851 158210 101931
rect 158520 101851 158530 101931
rect 158840 101851 158850 101931
rect 159160 101851 159170 101931
rect 159480 101851 159490 101931
rect 163750 101901 163830 101911
rect 164070 101901 164150 101911
rect 164390 101901 164470 101911
rect 164710 101901 164790 101911
rect 165030 101901 165110 101911
rect 165350 101901 165430 101911
rect 165670 101901 165750 101911
rect 165990 101901 166070 101911
rect 166310 101901 166390 101911
rect 166630 101901 166710 101911
rect 166950 101901 167030 101911
rect 167270 101901 167350 101911
rect 167590 101901 167670 101911
rect 167910 101901 167990 101911
rect 168230 101901 168310 101911
rect 168550 101901 168630 101911
rect 168870 101901 168950 101911
rect 169190 101901 169270 101911
rect 169510 101901 169590 101911
rect 169830 101901 169910 101911
rect 170150 101901 170230 101911
rect 170470 101901 170550 101911
rect 170790 101901 170870 101911
rect 163830 101821 163840 101901
rect 164150 101821 164160 101901
rect 164470 101821 164480 101901
rect 164790 101821 164800 101901
rect 165110 101821 165120 101901
rect 165430 101821 165440 101901
rect 165750 101821 165760 101901
rect 166070 101821 166080 101901
rect 166390 101821 166400 101901
rect 166710 101821 166720 101901
rect 167030 101821 167040 101901
rect 167350 101821 167360 101901
rect 167670 101821 167680 101901
rect 167990 101821 168000 101901
rect 168310 101821 168320 101901
rect 168630 101821 168640 101901
rect 168950 101821 168960 101901
rect 169270 101821 169280 101901
rect 169590 101821 169600 101901
rect 169910 101821 169920 101901
rect 170230 101821 170240 101901
rect 170550 101821 170560 101901
rect 170870 101821 170880 101901
rect 30360 101680 30440 101690
rect 30680 101680 30760 101690
rect 31000 101680 31080 101690
rect 31320 101680 31400 101690
rect 31640 101680 31720 101690
rect 31960 101680 32040 101690
rect 32280 101680 32360 101690
rect 32600 101680 32680 101690
rect 32920 101680 33000 101690
rect 33240 101680 33320 101690
rect 33560 101680 33640 101690
rect 33880 101680 33960 101690
rect 34200 101680 34280 101690
rect 34520 101680 34600 101690
rect 34840 101680 34920 101690
rect 35160 101680 35240 101690
rect 35480 101680 35560 101690
rect 35800 101680 35880 101690
rect 36120 101680 36200 101690
rect 36440 101680 36520 101690
rect 36760 101680 36840 101690
rect 37080 101680 37160 101690
rect 37400 101680 37480 101690
rect 37720 101680 37800 101690
rect 40180 101680 40260 101690
rect 40500 101680 40580 101690
rect 40820 101680 40900 101690
rect 41140 101680 41220 101690
rect 42560 101680 42640 101690
rect 42880 101680 42960 101690
rect 43200 101680 43280 101690
rect 43520 101680 43600 101690
rect 18970 101650 19050 101660
rect 19290 101650 19370 101660
rect 19610 101650 19690 101660
rect 19930 101650 20010 101660
rect 20250 101650 20330 101660
rect 20570 101650 20650 101660
rect 20890 101650 20970 101660
rect 21210 101650 21290 101660
rect 21530 101650 21610 101660
rect 21850 101650 21930 101660
rect 22170 101650 22250 101660
rect 22490 101650 22570 101660
rect 22810 101650 22890 101660
rect 23130 101650 23210 101660
rect 23450 101650 23530 101660
rect 23770 101650 23850 101660
rect 24090 101650 24170 101660
rect 24410 101650 24490 101660
rect 24730 101650 24810 101660
rect 25050 101650 25130 101660
rect 25370 101650 25450 101660
rect 25690 101650 25770 101660
rect 26010 101650 26090 101660
rect 26330 101650 26410 101660
rect 19050 101570 19060 101650
rect 19370 101570 19380 101650
rect 19690 101570 19700 101650
rect 20010 101570 20020 101650
rect 20330 101570 20340 101650
rect 20650 101570 20660 101650
rect 20970 101570 20980 101650
rect 21290 101570 21300 101650
rect 21610 101570 21620 101650
rect 21930 101570 21940 101650
rect 22250 101570 22260 101650
rect 22570 101570 22580 101650
rect 22890 101570 22900 101650
rect 23210 101570 23220 101650
rect 23530 101570 23540 101650
rect 23850 101570 23860 101650
rect 24170 101570 24180 101650
rect 24490 101570 24500 101650
rect 24810 101570 24820 101650
rect 25130 101570 25140 101650
rect 25450 101570 25460 101650
rect 25770 101570 25780 101650
rect 26090 101570 26100 101650
rect 26410 101570 26420 101650
rect 30440 101600 30450 101680
rect 30760 101600 30770 101680
rect 31080 101600 31090 101680
rect 31400 101600 31410 101680
rect 31720 101600 31730 101680
rect 32040 101600 32050 101680
rect 32360 101600 32370 101680
rect 32680 101600 32690 101680
rect 33000 101600 33010 101680
rect 33320 101600 33330 101680
rect 33640 101600 33650 101680
rect 33960 101600 33970 101680
rect 34280 101600 34290 101680
rect 34600 101600 34610 101680
rect 34920 101600 34930 101680
rect 35240 101600 35250 101680
rect 35560 101600 35570 101680
rect 35880 101600 35890 101680
rect 36200 101600 36210 101680
rect 36520 101600 36530 101680
rect 36840 101600 36850 101680
rect 37160 101600 37170 101680
rect 37480 101600 37490 101680
rect 37800 101600 37810 101680
rect 40260 101600 40270 101680
rect 40580 101600 40590 101680
rect 40900 101600 40910 101680
rect 41220 101600 41230 101680
rect 42640 101600 42650 101680
rect 42960 101600 42970 101680
rect 43280 101600 43290 101680
rect 43600 101600 43610 101680
rect 146400 101671 146480 101681
rect 146720 101671 146800 101681
rect 147040 101671 147120 101681
rect 147360 101671 147440 101681
rect 148780 101671 148860 101681
rect 149100 101671 149180 101681
rect 149420 101671 149500 101681
rect 149740 101671 149820 101681
rect 152200 101671 152280 101681
rect 152520 101671 152600 101681
rect 152840 101671 152920 101681
rect 153160 101671 153240 101681
rect 153480 101671 153560 101681
rect 153800 101671 153880 101681
rect 154120 101671 154200 101681
rect 154440 101671 154520 101681
rect 154760 101671 154840 101681
rect 155080 101671 155160 101681
rect 155400 101671 155480 101681
rect 155720 101671 155800 101681
rect 156040 101671 156120 101681
rect 156360 101671 156440 101681
rect 156680 101671 156760 101681
rect 157000 101671 157080 101681
rect 157320 101671 157400 101681
rect 157640 101671 157720 101681
rect 157960 101671 158040 101681
rect 158280 101671 158360 101681
rect 158600 101671 158680 101681
rect 158920 101671 159000 101681
rect 159240 101671 159320 101681
rect 159560 101671 159640 101681
rect 146480 101591 146490 101671
rect 146800 101591 146810 101671
rect 147120 101591 147130 101671
rect 147440 101591 147450 101671
rect 148860 101591 148870 101671
rect 149180 101591 149190 101671
rect 149500 101591 149510 101671
rect 149820 101591 149830 101671
rect 152280 101591 152290 101671
rect 152600 101591 152610 101671
rect 152920 101591 152930 101671
rect 153240 101591 153250 101671
rect 153560 101591 153570 101671
rect 153880 101591 153890 101671
rect 154200 101591 154210 101671
rect 154520 101591 154530 101671
rect 154840 101591 154850 101671
rect 155160 101591 155170 101671
rect 155480 101591 155490 101671
rect 155800 101591 155810 101671
rect 156120 101591 156130 101671
rect 156440 101591 156450 101671
rect 156760 101591 156770 101671
rect 157080 101591 157090 101671
rect 157400 101591 157410 101671
rect 157720 101591 157730 101671
rect 158040 101591 158050 101671
rect 158360 101591 158370 101671
rect 158680 101591 158690 101671
rect 159000 101591 159010 101671
rect 159320 101591 159330 101671
rect 159640 101591 159650 101671
rect 163590 101641 163670 101651
rect 163910 101641 163990 101651
rect 164230 101641 164310 101651
rect 164550 101641 164630 101651
rect 164870 101641 164950 101651
rect 165190 101641 165270 101651
rect 165510 101641 165590 101651
rect 165830 101641 165910 101651
rect 166150 101641 166230 101651
rect 166470 101641 166550 101651
rect 166790 101641 166870 101651
rect 167110 101641 167190 101651
rect 167430 101641 167510 101651
rect 167750 101641 167830 101651
rect 168070 101641 168150 101651
rect 168390 101641 168470 101651
rect 168710 101641 168790 101651
rect 169030 101641 169110 101651
rect 169350 101641 169430 101651
rect 169670 101641 169750 101651
rect 169990 101641 170070 101651
rect 170310 101641 170390 101651
rect 170630 101641 170710 101651
rect 170950 101641 171030 101651
rect 163670 101561 163680 101641
rect 163990 101561 164000 101641
rect 164310 101561 164320 101641
rect 164630 101561 164640 101641
rect 164950 101561 164960 101641
rect 165270 101561 165280 101641
rect 165590 101561 165600 101641
rect 165910 101561 165920 101641
rect 166230 101561 166240 101641
rect 166550 101561 166560 101641
rect 166870 101561 166880 101641
rect 167190 101561 167200 101641
rect 167510 101561 167520 101641
rect 167830 101561 167840 101641
rect 168150 101561 168160 101641
rect 168470 101561 168480 101641
rect 168790 101561 168800 101641
rect 169110 101561 169120 101641
rect 169430 101561 169440 101641
rect 169750 101561 169760 101641
rect 170070 101561 170080 101641
rect 170390 101561 170400 101641
rect 170710 101561 170720 101641
rect 171030 101561 171040 101641
rect 30520 101520 30600 101530
rect 30840 101520 30920 101530
rect 31160 101520 31240 101530
rect 31480 101520 31560 101530
rect 31800 101520 31880 101530
rect 32120 101520 32200 101530
rect 32440 101520 32520 101530
rect 32760 101520 32840 101530
rect 33080 101520 33160 101530
rect 33400 101520 33480 101530
rect 33720 101520 33800 101530
rect 34040 101520 34120 101530
rect 34360 101520 34440 101530
rect 34680 101520 34760 101530
rect 35000 101520 35080 101530
rect 35320 101520 35400 101530
rect 35640 101520 35720 101530
rect 35960 101520 36040 101530
rect 36280 101520 36360 101530
rect 36600 101520 36680 101530
rect 36920 101520 37000 101530
rect 37240 101520 37320 101530
rect 37560 101520 37640 101530
rect 40340 101520 40420 101530
rect 40660 101520 40740 101530
rect 40980 101520 41060 101530
rect 42720 101520 42800 101530
rect 43040 101520 43120 101530
rect 43360 101520 43440 101530
rect 19130 101490 19210 101500
rect 19450 101490 19530 101500
rect 19770 101490 19850 101500
rect 20090 101490 20170 101500
rect 20410 101490 20490 101500
rect 20730 101490 20810 101500
rect 21050 101490 21130 101500
rect 21370 101490 21450 101500
rect 21690 101490 21770 101500
rect 22010 101490 22090 101500
rect 22330 101490 22410 101500
rect 22650 101490 22730 101500
rect 22970 101490 23050 101500
rect 23290 101490 23370 101500
rect 23610 101490 23690 101500
rect 23930 101490 24010 101500
rect 24250 101490 24330 101500
rect 24570 101490 24650 101500
rect 24890 101490 24970 101500
rect 25210 101490 25290 101500
rect 25530 101490 25610 101500
rect 25850 101490 25930 101500
rect 26170 101490 26250 101500
rect 19210 101410 19220 101490
rect 19530 101410 19540 101490
rect 19850 101410 19860 101490
rect 20170 101410 20180 101490
rect 20490 101410 20500 101490
rect 20810 101410 20820 101490
rect 21130 101410 21140 101490
rect 21450 101410 21460 101490
rect 21770 101410 21780 101490
rect 22090 101410 22100 101490
rect 22410 101410 22420 101490
rect 22730 101410 22740 101490
rect 23050 101410 23060 101490
rect 23370 101410 23380 101490
rect 23690 101410 23700 101490
rect 24010 101410 24020 101490
rect 24330 101410 24340 101490
rect 24650 101410 24660 101490
rect 24970 101410 24980 101490
rect 25290 101410 25300 101490
rect 25610 101410 25620 101490
rect 25930 101410 25940 101490
rect 26250 101410 26260 101490
rect 30600 101440 30610 101520
rect 30920 101440 30930 101520
rect 31240 101440 31250 101520
rect 31560 101440 31570 101520
rect 31880 101440 31890 101520
rect 32200 101440 32210 101520
rect 32520 101440 32530 101520
rect 32840 101440 32850 101520
rect 33160 101440 33170 101520
rect 33480 101440 33490 101520
rect 33800 101440 33810 101520
rect 34120 101440 34130 101520
rect 34440 101440 34450 101520
rect 34760 101440 34770 101520
rect 35080 101440 35090 101520
rect 35400 101440 35410 101520
rect 35720 101440 35730 101520
rect 36040 101440 36050 101520
rect 36360 101440 36370 101520
rect 36680 101440 36690 101520
rect 37000 101440 37010 101520
rect 37320 101440 37330 101520
rect 37640 101440 37650 101520
rect 40420 101440 40430 101520
rect 40740 101440 40750 101520
rect 41060 101440 41070 101520
rect 42800 101440 42810 101520
rect 43120 101440 43130 101520
rect 43440 101440 43450 101520
rect 146560 101511 146640 101521
rect 146880 101511 146960 101521
rect 147200 101511 147280 101521
rect 148940 101511 149020 101521
rect 149260 101511 149340 101521
rect 149580 101511 149660 101521
rect 152360 101511 152440 101521
rect 152680 101511 152760 101521
rect 153000 101511 153080 101521
rect 153320 101511 153400 101521
rect 153640 101511 153720 101521
rect 153960 101511 154040 101521
rect 154280 101511 154360 101521
rect 154600 101511 154680 101521
rect 154920 101511 155000 101521
rect 155240 101511 155320 101521
rect 155560 101511 155640 101521
rect 155880 101511 155960 101521
rect 156200 101511 156280 101521
rect 156520 101511 156600 101521
rect 156840 101511 156920 101521
rect 157160 101511 157240 101521
rect 157480 101511 157560 101521
rect 157800 101511 157880 101521
rect 158120 101511 158200 101521
rect 158440 101511 158520 101521
rect 158760 101511 158840 101521
rect 159080 101511 159160 101521
rect 159400 101511 159480 101521
rect 30360 101360 30440 101370
rect 30680 101360 30760 101370
rect 31000 101360 31080 101370
rect 31320 101360 31400 101370
rect 31640 101360 31720 101370
rect 31960 101360 32040 101370
rect 32280 101360 32360 101370
rect 32600 101360 32680 101370
rect 32920 101360 33000 101370
rect 33240 101360 33320 101370
rect 33560 101360 33640 101370
rect 33880 101360 33960 101370
rect 34200 101360 34280 101370
rect 34520 101360 34600 101370
rect 34840 101360 34920 101370
rect 35160 101360 35240 101370
rect 35480 101360 35560 101370
rect 35800 101360 35880 101370
rect 36120 101360 36200 101370
rect 36440 101360 36520 101370
rect 36760 101360 36840 101370
rect 37080 101360 37160 101370
rect 37400 101360 37480 101370
rect 37720 101360 37800 101370
rect 40180 101360 40260 101370
rect 40500 101360 40580 101370
rect 40820 101360 40900 101370
rect 41140 101360 41220 101370
rect 42560 101360 42640 101370
rect 42880 101360 42960 101370
rect 43200 101360 43280 101370
rect 43520 101360 43600 101370
rect 18970 101330 19050 101340
rect 19290 101330 19370 101340
rect 19610 101330 19690 101340
rect 19930 101330 20010 101340
rect 20250 101330 20330 101340
rect 20570 101330 20650 101340
rect 20890 101330 20970 101340
rect 21210 101330 21290 101340
rect 21530 101330 21610 101340
rect 21850 101330 21930 101340
rect 22170 101330 22250 101340
rect 22490 101330 22570 101340
rect 22810 101330 22890 101340
rect 23130 101330 23210 101340
rect 23450 101330 23530 101340
rect 23770 101330 23850 101340
rect 24090 101330 24170 101340
rect 24410 101330 24490 101340
rect 24730 101330 24810 101340
rect 25050 101330 25130 101340
rect 25370 101330 25450 101340
rect 25690 101330 25770 101340
rect 26010 101330 26090 101340
rect 26330 101330 26410 101340
rect 19050 101250 19060 101330
rect 19370 101250 19380 101330
rect 19690 101250 19700 101330
rect 20010 101250 20020 101330
rect 20330 101250 20340 101330
rect 20650 101250 20660 101330
rect 20970 101250 20980 101330
rect 21290 101250 21300 101330
rect 21610 101250 21620 101330
rect 21930 101250 21940 101330
rect 22250 101250 22260 101330
rect 22570 101250 22580 101330
rect 22890 101250 22900 101330
rect 23210 101250 23220 101330
rect 23530 101250 23540 101330
rect 23850 101250 23860 101330
rect 24170 101250 24180 101330
rect 24490 101250 24500 101330
rect 24810 101250 24820 101330
rect 25130 101250 25140 101330
rect 25450 101250 25460 101330
rect 25770 101250 25780 101330
rect 26090 101250 26100 101330
rect 26410 101250 26420 101330
rect 30440 101280 30450 101360
rect 30760 101280 30770 101360
rect 31080 101280 31090 101360
rect 31400 101280 31410 101360
rect 31720 101280 31730 101360
rect 32040 101280 32050 101360
rect 32360 101280 32370 101360
rect 32680 101280 32690 101360
rect 33000 101280 33010 101360
rect 33320 101280 33330 101360
rect 33640 101280 33650 101360
rect 33960 101280 33970 101360
rect 34280 101280 34290 101360
rect 34600 101280 34610 101360
rect 34920 101280 34930 101360
rect 35240 101280 35250 101360
rect 35560 101280 35570 101360
rect 35880 101280 35890 101360
rect 36200 101280 36210 101360
rect 36520 101280 36530 101360
rect 36840 101280 36850 101360
rect 37160 101280 37170 101360
rect 37480 101280 37490 101360
rect 37800 101280 37810 101360
rect 40260 101280 40270 101360
rect 40580 101280 40590 101360
rect 40900 101280 40910 101360
rect 41220 101280 41230 101360
rect 42640 101280 42650 101360
rect 42960 101280 42970 101360
rect 43280 101280 43290 101360
rect 43600 101280 43610 101360
rect 46660 101260 48570 101440
rect 146640 101431 146650 101511
rect 146960 101431 146970 101511
rect 147280 101431 147290 101511
rect 149020 101431 149030 101511
rect 149340 101431 149350 101511
rect 149660 101431 149670 101511
rect 152440 101431 152450 101511
rect 152760 101431 152770 101511
rect 153080 101431 153090 101511
rect 153400 101431 153410 101511
rect 153720 101431 153730 101511
rect 154040 101431 154050 101511
rect 154360 101431 154370 101511
rect 154680 101431 154690 101511
rect 155000 101431 155010 101511
rect 155320 101431 155330 101511
rect 155640 101431 155650 101511
rect 155960 101431 155970 101511
rect 156280 101431 156290 101511
rect 156600 101431 156610 101511
rect 156920 101431 156930 101511
rect 157240 101431 157250 101511
rect 157560 101431 157570 101511
rect 157880 101431 157890 101511
rect 158200 101431 158210 101511
rect 158520 101431 158530 101511
rect 158840 101431 158850 101511
rect 159160 101431 159170 101511
rect 159480 101431 159490 101511
rect 163750 101481 163830 101491
rect 164070 101481 164150 101491
rect 164390 101481 164470 101491
rect 164710 101481 164790 101491
rect 165030 101481 165110 101491
rect 165350 101481 165430 101491
rect 165670 101481 165750 101491
rect 165990 101481 166070 101491
rect 166310 101481 166390 101491
rect 166630 101481 166710 101491
rect 166950 101481 167030 101491
rect 167270 101481 167350 101491
rect 167590 101481 167670 101491
rect 167910 101481 167990 101491
rect 168230 101481 168310 101491
rect 168550 101481 168630 101491
rect 168870 101481 168950 101491
rect 169190 101481 169270 101491
rect 169510 101481 169590 101491
rect 169830 101481 169910 101491
rect 170150 101481 170230 101491
rect 170470 101481 170550 101491
rect 170790 101481 170870 101491
rect 163830 101401 163840 101481
rect 164150 101401 164160 101481
rect 164470 101401 164480 101481
rect 164790 101401 164800 101481
rect 165110 101401 165120 101481
rect 165430 101401 165440 101481
rect 165750 101401 165760 101481
rect 166070 101401 166080 101481
rect 166390 101401 166400 101481
rect 166710 101401 166720 101481
rect 167030 101401 167040 101481
rect 167350 101401 167360 101481
rect 167670 101401 167680 101481
rect 167990 101401 168000 101481
rect 168310 101401 168320 101481
rect 168630 101401 168640 101481
rect 168950 101401 168960 101481
rect 169270 101401 169280 101481
rect 169590 101401 169600 101481
rect 169910 101401 169920 101481
rect 170230 101401 170240 101481
rect 170550 101401 170560 101481
rect 170870 101401 170880 101481
rect 146400 101351 146480 101361
rect 146720 101351 146800 101361
rect 147040 101351 147120 101361
rect 147360 101351 147440 101361
rect 148780 101351 148860 101361
rect 149100 101351 149180 101361
rect 149420 101351 149500 101361
rect 149740 101351 149820 101361
rect 152200 101351 152280 101361
rect 152520 101351 152600 101361
rect 152840 101351 152920 101361
rect 153160 101351 153240 101361
rect 153480 101351 153560 101361
rect 153800 101351 153880 101361
rect 154120 101351 154200 101361
rect 154440 101351 154520 101361
rect 154760 101351 154840 101361
rect 155080 101351 155160 101361
rect 155400 101351 155480 101361
rect 155720 101351 155800 101361
rect 156040 101351 156120 101361
rect 156360 101351 156440 101361
rect 156680 101351 156760 101361
rect 157000 101351 157080 101361
rect 157320 101351 157400 101361
rect 157640 101351 157720 101361
rect 157960 101351 158040 101361
rect 158280 101351 158360 101361
rect 158600 101351 158680 101361
rect 158920 101351 159000 101361
rect 159240 101351 159320 101361
rect 159560 101351 159640 101361
rect 146480 101271 146490 101351
rect 146800 101271 146810 101351
rect 147120 101271 147130 101351
rect 147440 101271 147450 101351
rect 148860 101271 148870 101351
rect 149180 101271 149190 101351
rect 149500 101271 149510 101351
rect 149820 101271 149830 101351
rect 152280 101271 152290 101351
rect 152600 101271 152610 101351
rect 152920 101271 152930 101351
rect 153240 101271 153250 101351
rect 153560 101271 153570 101351
rect 153880 101271 153890 101351
rect 154200 101271 154210 101351
rect 154520 101271 154530 101351
rect 154840 101271 154850 101351
rect 155160 101271 155170 101351
rect 155480 101271 155490 101351
rect 155800 101271 155810 101351
rect 156120 101271 156130 101351
rect 156440 101271 156450 101351
rect 156760 101271 156770 101351
rect 157080 101271 157090 101351
rect 157400 101271 157410 101351
rect 157720 101271 157730 101351
rect 158040 101271 158050 101351
rect 158360 101271 158370 101351
rect 158680 101271 158690 101351
rect 159000 101271 159010 101351
rect 159320 101271 159330 101351
rect 159640 101271 159650 101351
rect 163590 101321 163670 101331
rect 163910 101321 163990 101331
rect 164230 101321 164310 101331
rect 164550 101321 164630 101331
rect 164870 101321 164950 101331
rect 165190 101321 165270 101331
rect 165510 101321 165590 101331
rect 165830 101321 165910 101331
rect 166150 101321 166230 101331
rect 166470 101321 166550 101331
rect 166790 101321 166870 101331
rect 167110 101321 167190 101331
rect 167430 101321 167510 101331
rect 167750 101321 167830 101331
rect 168070 101321 168150 101331
rect 168390 101321 168470 101331
rect 168710 101321 168790 101331
rect 169030 101321 169110 101331
rect 169350 101321 169430 101331
rect 169670 101321 169750 101331
rect 169990 101321 170070 101331
rect 170310 101321 170390 101331
rect 170630 101321 170710 101331
rect 170950 101321 171030 101331
rect 163670 101241 163680 101321
rect 163990 101241 164000 101321
rect 164310 101241 164320 101321
rect 164630 101241 164640 101321
rect 164950 101241 164960 101321
rect 165270 101241 165280 101321
rect 165590 101241 165600 101321
rect 165910 101241 165920 101321
rect 166230 101241 166240 101321
rect 166550 101241 166560 101321
rect 166870 101241 166880 101321
rect 167190 101241 167200 101321
rect 167510 101241 167520 101321
rect 167830 101241 167840 101321
rect 168150 101241 168160 101321
rect 168470 101241 168480 101321
rect 168790 101241 168800 101321
rect 169110 101241 169120 101321
rect 169430 101241 169440 101321
rect 169750 101241 169760 101321
rect 170070 101241 170080 101321
rect 170390 101241 170400 101321
rect 170710 101241 170720 101321
rect 171030 101241 171040 101321
rect 30520 101200 30600 101210
rect 30840 101200 30920 101210
rect 31160 101200 31240 101210
rect 31480 101200 31560 101210
rect 31800 101200 31880 101210
rect 32120 101200 32200 101210
rect 32440 101200 32520 101210
rect 32760 101200 32840 101210
rect 33080 101200 33160 101210
rect 33400 101200 33480 101210
rect 33720 101200 33800 101210
rect 34040 101200 34120 101210
rect 34360 101200 34440 101210
rect 34680 101200 34760 101210
rect 35000 101200 35080 101210
rect 35320 101200 35400 101210
rect 35640 101200 35720 101210
rect 35960 101200 36040 101210
rect 36280 101200 36360 101210
rect 36600 101200 36680 101210
rect 36920 101200 37000 101210
rect 37240 101200 37320 101210
rect 37560 101200 37640 101210
rect 40340 101200 40420 101210
rect 40660 101200 40740 101210
rect 40980 101200 41060 101210
rect 42720 101200 42800 101210
rect 43040 101200 43120 101210
rect 43360 101200 43440 101210
rect 19130 101170 19210 101180
rect 19450 101170 19530 101180
rect 19770 101170 19850 101180
rect 20090 101170 20170 101180
rect 20410 101170 20490 101180
rect 20730 101170 20810 101180
rect 21050 101170 21130 101180
rect 21370 101170 21450 101180
rect 21690 101170 21770 101180
rect 22010 101170 22090 101180
rect 22330 101170 22410 101180
rect 22650 101170 22730 101180
rect 22970 101170 23050 101180
rect 23290 101170 23370 101180
rect 23610 101170 23690 101180
rect 23930 101170 24010 101180
rect 24250 101170 24330 101180
rect 24570 101170 24650 101180
rect 24890 101170 24970 101180
rect 25210 101170 25290 101180
rect 25530 101170 25610 101180
rect 25850 101170 25930 101180
rect 26170 101170 26250 101180
rect 19210 101090 19220 101170
rect 19530 101090 19540 101170
rect 19850 101090 19860 101170
rect 20170 101090 20180 101170
rect 20490 101090 20500 101170
rect 20810 101090 20820 101170
rect 21130 101090 21140 101170
rect 21450 101090 21460 101170
rect 21770 101090 21780 101170
rect 22090 101090 22100 101170
rect 22410 101090 22420 101170
rect 22730 101090 22740 101170
rect 23050 101090 23060 101170
rect 23370 101090 23380 101170
rect 23690 101090 23700 101170
rect 24010 101090 24020 101170
rect 24330 101090 24340 101170
rect 24650 101090 24660 101170
rect 24970 101090 24980 101170
rect 25290 101090 25300 101170
rect 25610 101090 25620 101170
rect 25930 101090 25940 101170
rect 26250 101090 26260 101170
rect 30600 101120 30610 101200
rect 30920 101120 30930 101200
rect 31240 101120 31250 101200
rect 31560 101120 31570 101200
rect 31880 101120 31890 101200
rect 32200 101120 32210 101200
rect 32520 101120 32530 101200
rect 32840 101120 32850 101200
rect 33160 101120 33170 101200
rect 33480 101120 33490 101200
rect 33800 101120 33810 101200
rect 34120 101120 34130 101200
rect 34440 101120 34450 101200
rect 34760 101120 34770 101200
rect 35080 101120 35090 101200
rect 35400 101120 35410 101200
rect 35720 101120 35730 101200
rect 36040 101120 36050 101200
rect 36360 101120 36370 101200
rect 36680 101120 36690 101200
rect 37000 101120 37010 101200
rect 37320 101120 37330 101200
rect 37640 101120 37650 101200
rect 40420 101120 40430 101200
rect 40740 101120 40750 101200
rect 41060 101120 41070 101200
rect 42800 101120 42810 101200
rect 43120 101120 43130 101200
rect 43440 101120 43450 101200
rect 146560 101191 146640 101201
rect 146880 101191 146960 101201
rect 147200 101191 147280 101201
rect 148940 101191 149020 101201
rect 149260 101191 149340 101201
rect 149580 101191 149660 101201
rect 152360 101191 152440 101201
rect 152680 101191 152760 101201
rect 153000 101191 153080 101201
rect 153320 101191 153400 101201
rect 153640 101191 153720 101201
rect 153960 101191 154040 101201
rect 154280 101191 154360 101201
rect 154600 101191 154680 101201
rect 154920 101191 155000 101201
rect 155240 101191 155320 101201
rect 155560 101191 155640 101201
rect 155880 101191 155960 101201
rect 156200 101191 156280 101201
rect 156520 101191 156600 101201
rect 156840 101191 156920 101201
rect 157160 101191 157240 101201
rect 157480 101191 157560 101201
rect 157800 101191 157880 101201
rect 158120 101191 158200 101201
rect 158440 101191 158520 101201
rect 158760 101191 158840 101201
rect 159080 101191 159160 101201
rect 159400 101191 159480 101201
rect 146640 101111 146650 101191
rect 146960 101111 146970 101191
rect 147280 101111 147290 101191
rect 149020 101111 149030 101191
rect 149340 101111 149350 101191
rect 149660 101111 149670 101191
rect 152440 101111 152450 101191
rect 152760 101111 152770 101191
rect 153080 101111 153090 101191
rect 153400 101111 153410 101191
rect 153720 101111 153730 101191
rect 154040 101111 154050 101191
rect 154360 101111 154370 101191
rect 154680 101111 154690 101191
rect 155000 101111 155010 101191
rect 155320 101111 155330 101191
rect 155640 101111 155650 101191
rect 155960 101111 155970 101191
rect 156280 101111 156290 101191
rect 156600 101111 156610 101191
rect 156920 101111 156930 101191
rect 157240 101111 157250 101191
rect 157560 101111 157570 101191
rect 157880 101111 157890 101191
rect 158200 101111 158210 101191
rect 158520 101111 158530 101191
rect 158840 101111 158850 101191
rect 159160 101111 159170 101191
rect 159480 101111 159490 101191
rect 163750 101161 163830 101171
rect 164070 101161 164150 101171
rect 164390 101161 164470 101171
rect 164710 101161 164790 101171
rect 165030 101161 165110 101171
rect 165350 101161 165430 101171
rect 165670 101161 165750 101171
rect 165990 101161 166070 101171
rect 166310 101161 166390 101171
rect 166630 101161 166710 101171
rect 166950 101161 167030 101171
rect 167270 101161 167350 101171
rect 167590 101161 167670 101171
rect 167910 101161 167990 101171
rect 168230 101161 168310 101171
rect 168550 101161 168630 101171
rect 168870 101161 168950 101171
rect 169190 101161 169270 101171
rect 169510 101161 169590 101171
rect 169830 101161 169910 101171
rect 170150 101161 170230 101171
rect 170470 101161 170550 101171
rect 170790 101161 170870 101171
rect 163830 101081 163840 101161
rect 164150 101081 164160 101161
rect 164470 101081 164480 101161
rect 164790 101081 164800 101161
rect 165110 101081 165120 101161
rect 165430 101081 165440 101161
rect 165750 101081 165760 101161
rect 166070 101081 166080 101161
rect 166390 101081 166400 101161
rect 166710 101081 166720 101161
rect 167030 101081 167040 101161
rect 167350 101081 167360 101161
rect 167670 101081 167680 101161
rect 167990 101081 168000 101161
rect 168310 101081 168320 101161
rect 168630 101081 168640 101161
rect 168950 101081 168960 101161
rect 169270 101081 169280 101161
rect 169590 101081 169600 101161
rect 169910 101081 169920 101161
rect 170230 101081 170240 101161
rect 170550 101081 170560 101161
rect 170870 101081 170880 101161
rect 18980 100940 19060 100950
rect 19160 100940 19240 100950
rect 19340 100940 19420 100950
rect 19520 100940 19600 100950
rect 19700 100940 19780 100950
rect 19880 100940 19960 100950
rect 20060 100940 20140 100950
rect 20240 100940 20320 100950
rect 20420 100940 20500 100950
rect 20600 100940 20680 100950
rect 20780 100940 20860 100950
rect 20960 100940 21040 100950
rect 21140 100940 21220 100950
rect 21320 100940 21400 100950
rect 21500 100940 21580 100950
rect 21680 100940 21760 100950
rect 21860 100940 21940 100950
rect 22040 100940 22120 100950
rect 22220 100940 22300 100950
rect 22400 100940 22480 100950
rect 22580 100940 22660 100950
rect 22760 100940 22840 100950
rect 22940 100940 23020 100950
rect 23120 100940 23200 100950
rect 23300 100940 23380 100950
rect 23480 100940 23560 100950
rect 23660 100940 23740 100950
rect 23840 100940 23920 100950
rect 24020 100940 24100 100950
rect 24200 100940 24280 100950
rect 24380 100940 24460 100950
rect 24560 100940 24640 100950
rect 24740 100940 24820 100950
rect 24920 100940 25000 100950
rect 25100 100940 25180 100950
rect 25280 100940 25360 100950
rect 25460 100940 25540 100950
rect 25640 100940 25720 100950
rect 25820 100940 25900 100950
rect 26000 100940 26080 100950
rect 26180 100940 26260 100950
rect 26360 100940 26440 100950
rect 26540 100940 26620 100950
rect 30280 100940 30360 100950
rect 30460 100940 30540 100950
rect 30640 100940 30720 100950
rect 30820 100940 30900 100950
rect 31000 100940 31080 100950
rect 31180 100940 31260 100950
rect 31360 100940 31440 100950
rect 31540 100940 31620 100950
rect 31720 100940 31800 100950
rect 31900 100940 31980 100950
rect 32080 100940 32160 100950
rect 32260 100940 32340 100950
rect 32440 100940 32520 100950
rect 32620 100940 32700 100950
rect 32800 100940 32880 100950
rect 32980 100940 33060 100950
rect 33160 100940 33240 100950
rect 33340 100940 33420 100950
rect 33520 100940 33600 100950
rect 33700 100940 33780 100950
rect 33880 100940 33960 100950
rect 34060 100940 34140 100950
rect 34240 100940 34320 100950
rect 34420 100940 34500 100950
rect 34600 100940 34680 100950
rect 34780 100940 34860 100950
rect 34960 100940 35040 100950
rect 35140 100940 35220 100950
rect 35320 100940 35400 100950
rect 35500 100940 35580 100950
rect 35680 100940 35760 100950
rect 35860 100940 35940 100950
rect 36040 100940 36120 100950
rect 36220 100940 36300 100950
rect 36400 100940 36480 100950
rect 36580 100940 36660 100950
rect 36760 100940 36840 100950
rect 36940 100940 37020 100950
rect 37120 100940 37200 100950
rect 37300 100940 37380 100950
rect 37480 100940 37560 100950
rect 37660 100940 37740 100950
rect 37840 100940 37920 100950
rect 40060 100940 40140 100950
rect 40200 100940 40280 100950
rect 40340 100940 40420 100950
rect 40480 100940 40560 100950
rect 40620 100940 40700 100950
rect 40760 100940 40840 100950
rect 40900 100940 40980 100950
rect 41040 100940 41120 100950
rect 41180 100940 41260 100950
rect 41320 100940 41400 100950
rect 42360 100940 42440 100950
rect 42500 100940 42580 100950
rect 42640 100940 42720 100950
rect 42780 100940 42860 100950
rect 42920 100940 43000 100950
rect 43060 100940 43140 100950
rect 43200 100940 43280 100950
rect 43340 100940 43420 100950
rect 43480 100940 43560 100950
rect 43620 100940 43700 100950
rect 146300 100940 146380 100950
rect 146440 100940 146520 100950
rect 146580 100940 146660 100950
rect 146720 100940 146800 100950
rect 146860 100940 146940 100950
rect 147000 100940 147080 100950
rect 147140 100940 147220 100950
rect 147280 100940 147360 100950
rect 147420 100940 147500 100950
rect 147560 100940 147640 100950
rect 148600 100940 148680 100950
rect 148740 100940 148820 100950
rect 148880 100940 148960 100950
rect 149020 100940 149100 100950
rect 149160 100940 149240 100950
rect 149300 100940 149380 100950
rect 149440 100940 149520 100950
rect 149580 100940 149660 100950
rect 149720 100940 149800 100950
rect 149860 100940 149940 100950
rect 152080 100940 152160 100950
rect 152260 100940 152340 100950
rect 152440 100940 152520 100950
rect 152620 100940 152700 100950
rect 152800 100940 152880 100950
rect 152980 100940 153060 100950
rect 153160 100940 153240 100950
rect 153340 100940 153420 100950
rect 153520 100940 153600 100950
rect 153700 100940 153780 100950
rect 153880 100940 153960 100950
rect 154060 100940 154140 100950
rect 154240 100940 154320 100950
rect 154420 100940 154500 100950
rect 154600 100940 154680 100950
rect 154780 100940 154860 100950
rect 154960 100940 155040 100950
rect 155140 100940 155220 100950
rect 155320 100940 155400 100950
rect 155500 100940 155580 100950
rect 155680 100940 155760 100950
rect 155860 100940 155940 100950
rect 156040 100940 156120 100950
rect 156220 100940 156300 100950
rect 156400 100940 156480 100950
rect 156580 100940 156660 100950
rect 156760 100940 156840 100950
rect 156940 100940 157020 100950
rect 157120 100940 157200 100950
rect 157300 100940 157380 100950
rect 157480 100940 157560 100950
rect 157660 100940 157740 100950
rect 157840 100940 157920 100950
rect 158020 100940 158100 100950
rect 158200 100940 158280 100950
rect 158380 100940 158460 100950
rect 158560 100940 158640 100950
rect 158740 100940 158820 100950
rect 158920 100940 159000 100950
rect 159100 100940 159180 100950
rect 159280 100940 159360 100950
rect 159460 100940 159540 100950
rect 159640 100940 159720 100950
rect 163380 100940 163460 100950
rect 163560 100940 163640 100950
rect 163740 100940 163820 100950
rect 163920 100940 164000 100950
rect 164100 100940 164180 100950
rect 164280 100940 164360 100950
rect 164460 100940 164540 100950
rect 164640 100940 164720 100950
rect 164820 100940 164900 100950
rect 165000 100940 165080 100950
rect 165180 100940 165260 100950
rect 165360 100940 165440 100950
rect 165540 100940 165620 100950
rect 165720 100940 165800 100950
rect 165900 100940 165980 100950
rect 166080 100940 166160 100950
rect 166260 100940 166340 100950
rect 166440 100940 166520 100950
rect 166620 100940 166700 100950
rect 166800 100940 166880 100950
rect 166980 100940 167060 100950
rect 167160 100940 167240 100950
rect 167340 100940 167420 100950
rect 167520 100940 167600 100950
rect 167700 100940 167780 100950
rect 167880 100940 167960 100950
rect 168060 100940 168140 100950
rect 168240 100940 168320 100950
rect 168420 100940 168500 100950
rect 168600 100940 168680 100950
rect 168780 100940 168860 100950
rect 168960 100940 169040 100950
rect 169140 100940 169220 100950
rect 169320 100940 169400 100950
rect 169500 100940 169580 100950
rect 169680 100940 169760 100950
rect 169860 100940 169940 100950
rect 170040 100940 170120 100950
rect 170220 100940 170300 100950
rect 170400 100940 170480 100950
rect 170580 100940 170660 100950
rect 170760 100940 170840 100950
rect 170940 100940 171020 100950
rect 19060 100860 19070 100940
rect 19240 100860 19250 100940
rect 19420 100860 19430 100940
rect 19600 100860 19610 100940
rect 19780 100860 19790 100940
rect 19960 100860 19970 100940
rect 20140 100860 20150 100940
rect 20320 100860 20330 100940
rect 20500 100860 20510 100940
rect 20680 100860 20690 100940
rect 20860 100860 20870 100940
rect 21040 100860 21050 100940
rect 21220 100860 21230 100940
rect 21400 100860 21410 100940
rect 21580 100860 21590 100940
rect 21760 100860 21770 100940
rect 21940 100860 21950 100940
rect 22120 100860 22130 100940
rect 22300 100860 22310 100940
rect 22480 100860 22490 100940
rect 22660 100860 22670 100940
rect 22840 100860 22850 100940
rect 23020 100860 23030 100940
rect 23200 100860 23210 100940
rect 23380 100860 23390 100940
rect 23560 100860 23570 100940
rect 23740 100860 23750 100940
rect 23920 100860 23930 100940
rect 24100 100860 24110 100940
rect 24280 100860 24290 100940
rect 24460 100860 24470 100940
rect 24640 100860 24650 100940
rect 24820 100860 24830 100940
rect 25000 100860 25010 100940
rect 25180 100860 25190 100940
rect 25360 100860 25370 100940
rect 25540 100860 25550 100940
rect 25720 100860 25730 100940
rect 25900 100860 25910 100940
rect 26080 100860 26090 100940
rect 26260 100860 26270 100940
rect 26440 100860 26450 100940
rect 26620 100860 26630 100940
rect 30360 100860 30370 100940
rect 30540 100860 30550 100940
rect 30720 100860 30730 100940
rect 30900 100860 30910 100940
rect 31080 100860 31090 100940
rect 31260 100860 31270 100940
rect 31440 100860 31450 100940
rect 31620 100860 31630 100940
rect 31800 100860 31810 100940
rect 31980 100860 31990 100940
rect 32160 100860 32170 100940
rect 32340 100860 32350 100940
rect 32520 100860 32530 100940
rect 32700 100860 32710 100940
rect 32880 100860 32890 100940
rect 33060 100860 33070 100940
rect 33240 100860 33250 100940
rect 33420 100860 33430 100940
rect 33600 100860 33610 100940
rect 33780 100860 33790 100940
rect 33960 100860 33970 100940
rect 34140 100860 34150 100940
rect 34320 100860 34330 100940
rect 34500 100860 34510 100940
rect 34680 100860 34690 100940
rect 34860 100860 34870 100940
rect 35040 100860 35050 100940
rect 35220 100860 35230 100940
rect 35400 100860 35410 100940
rect 35580 100860 35590 100940
rect 35760 100860 35770 100940
rect 35940 100860 35950 100940
rect 36120 100860 36130 100940
rect 36300 100860 36310 100940
rect 36480 100860 36490 100940
rect 36660 100860 36670 100940
rect 36840 100860 36850 100940
rect 37020 100860 37030 100940
rect 37200 100860 37210 100940
rect 37380 100860 37390 100940
rect 37560 100860 37570 100940
rect 37740 100860 37750 100940
rect 37920 100860 37930 100940
rect 40140 100860 40150 100940
rect 40280 100860 40290 100940
rect 40420 100860 40430 100940
rect 40560 100860 40570 100940
rect 40700 100860 40710 100940
rect 40840 100860 40850 100940
rect 40980 100860 40990 100940
rect 41120 100860 41130 100940
rect 41260 100860 41270 100940
rect 41400 100860 41410 100940
rect 42440 100860 42450 100940
rect 42580 100860 42590 100940
rect 42720 100860 42730 100940
rect 42860 100860 42870 100940
rect 43000 100860 43010 100940
rect 43140 100860 43150 100940
rect 43280 100860 43290 100940
rect 43420 100860 43430 100940
rect 43560 100860 43570 100940
rect 43700 100860 43710 100940
rect 146380 100860 146390 100940
rect 146520 100860 146530 100940
rect 146660 100860 146670 100940
rect 146800 100860 146810 100940
rect 146940 100860 146950 100940
rect 147080 100860 147090 100940
rect 147220 100860 147230 100940
rect 147360 100860 147370 100940
rect 147500 100860 147510 100940
rect 147640 100860 147650 100940
rect 148680 100860 148690 100940
rect 148820 100860 148830 100940
rect 148960 100860 148970 100940
rect 149100 100860 149110 100940
rect 149240 100860 149250 100940
rect 149380 100860 149390 100940
rect 149520 100860 149530 100940
rect 149660 100860 149670 100940
rect 149800 100860 149810 100940
rect 149940 100860 149950 100940
rect 152160 100860 152170 100940
rect 152340 100860 152350 100940
rect 152520 100860 152530 100940
rect 152700 100860 152710 100940
rect 152880 100860 152890 100940
rect 153060 100860 153070 100940
rect 153240 100860 153250 100940
rect 153420 100860 153430 100940
rect 153600 100860 153610 100940
rect 153780 100860 153790 100940
rect 153960 100860 153970 100940
rect 154140 100860 154150 100940
rect 154320 100860 154330 100940
rect 154500 100860 154510 100940
rect 154680 100860 154690 100940
rect 154860 100860 154870 100940
rect 155040 100860 155050 100940
rect 155220 100860 155230 100940
rect 155400 100860 155410 100940
rect 155580 100860 155590 100940
rect 155760 100860 155770 100940
rect 155940 100860 155950 100940
rect 156120 100860 156130 100940
rect 156300 100860 156310 100940
rect 156480 100860 156490 100940
rect 156660 100860 156670 100940
rect 156840 100860 156850 100940
rect 157020 100860 157030 100940
rect 157200 100860 157210 100940
rect 157380 100860 157390 100940
rect 157560 100860 157570 100940
rect 157740 100860 157750 100940
rect 157920 100860 157930 100940
rect 158100 100860 158110 100940
rect 158280 100860 158290 100940
rect 158460 100860 158470 100940
rect 158640 100860 158650 100940
rect 158820 100860 158830 100940
rect 159000 100860 159010 100940
rect 159180 100860 159190 100940
rect 159360 100860 159370 100940
rect 159540 100860 159550 100940
rect 159720 100860 159730 100940
rect 163460 100860 163470 100940
rect 163640 100860 163650 100940
rect 163820 100860 163830 100940
rect 164000 100860 164010 100940
rect 164180 100860 164190 100940
rect 164360 100860 164370 100940
rect 164540 100860 164550 100940
rect 164720 100860 164730 100940
rect 164900 100860 164910 100940
rect 165080 100860 165090 100940
rect 165260 100860 165270 100940
rect 165440 100860 165450 100940
rect 165620 100860 165630 100940
rect 165800 100860 165810 100940
rect 165980 100860 165990 100940
rect 166160 100860 166170 100940
rect 166340 100860 166350 100940
rect 166520 100860 166530 100940
rect 166700 100860 166710 100940
rect 166880 100860 166890 100940
rect 167060 100860 167070 100940
rect 167240 100860 167250 100940
rect 167420 100860 167430 100940
rect 167600 100860 167610 100940
rect 167780 100860 167790 100940
rect 167960 100860 167970 100940
rect 168140 100860 168150 100940
rect 168320 100860 168330 100940
rect 168500 100860 168510 100940
rect 168680 100860 168690 100940
rect 168860 100860 168870 100940
rect 169040 100860 169050 100940
rect 169220 100860 169230 100940
rect 169400 100860 169410 100940
rect 169580 100860 169590 100940
rect 169760 100860 169770 100940
rect 169940 100860 169950 100940
rect 170120 100860 170130 100940
rect 170300 100860 170310 100940
rect 170480 100860 170490 100940
rect 170660 100860 170670 100940
rect 170840 100860 170850 100940
rect 171020 100860 171030 100940
rect 161885 100845 161965 100855
rect 162065 100845 162145 100855
rect 162245 100845 162325 100855
rect 162425 100845 162505 100855
rect 162605 100845 162685 100855
rect 28850 100815 28930 100825
rect 29010 100815 29090 100825
rect 29170 100815 29250 100825
rect 29330 100815 29410 100825
rect 29490 100815 29570 100825
rect 18980 100790 19060 100800
rect 19160 100790 19240 100800
rect 19340 100790 19420 100800
rect 19520 100790 19600 100800
rect 19700 100790 19780 100800
rect 19880 100790 19960 100800
rect 20060 100790 20140 100800
rect 20240 100790 20320 100800
rect 20420 100790 20500 100800
rect 20600 100790 20680 100800
rect 20780 100790 20860 100800
rect 20960 100790 21040 100800
rect 21140 100790 21220 100800
rect 21320 100790 21400 100800
rect 21500 100790 21580 100800
rect 21680 100790 21760 100800
rect 21860 100790 21940 100800
rect 22040 100790 22120 100800
rect 22220 100790 22300 100800
rect 22400 100790 22480 100800
rect 22580 100790 22660 100800
rect 22760 100790 22840 100800
rect 22940 100790 23020 100800
rect 23120 100790 23200 100800
rect 23300 100790 23380 100800
rect 23480 100790 23560 100800
rect 23660 100790 23740 100800
rect 23840 100790 23920 100800
rect 24020 100790 24100 100800
rect 24200 100790 24280 100800
rect 24380 100790 24460 100800
rect 24560 100790 24640 100800
rect 24740 100790 24820 100800
rect 24920 100790 25000 100800
rect 25100 100790 25180 100800
rect 25280 100790 25360 100800
rect 25460 100790 25540 100800
rect 25640 100790 25720 100800
rect 25820 100790 25900 100800
rect 26000 100790 26080 100800
rect 26180 100790 26260 100800
rect 26360 100790 26440 100800
rect 26540 100790 26620 100800
rect 19060 100710 19070 100790
rect 19240 100710 19250 100790
rect 19420 100710 19430 100790
rect 19600 100710 19610 100790
rect 19780 100710 19790 100790
rect 19960 100710 19970 100790
rect 20140 100710 20150 100790
rect 20320 100710 20330 100790
rect 20500 100710 20510 100790
rect 20680 100710 20690 100790
rect 20860 100710 20870 100790
rect 21040 100710 21050 100790
rect 21220 100710 21230 100790
rect 21400 100710 21410 100790
rect 21580 100710 21590 100790
rect 21760 100710 21770 100790
rect 21940 100710 21950 100790
rect 22120 100710 22130 100790
rect 22300 100710 22310 100790
rect 22480 100710 22490 100790
rect 22660 100710 22670 100790
rect 22840 100710 22850 100790
rect 23020 100710 23030 100790
rect 23200 100710 23210 100790
rect 23380 100710 23390 100790
rect 23560 100710 23570 100790
rect 23740 100710 23750 100790
rect 23920 100710 23930 100790
rect 24100 100710 24110 100790
rect 24280 100710 24290 100790
rect 24460 100710 24470 100790
rect 24640 100710 24650 100790
rect 24820 100710 24830 100790
rect 25000 100710 25010 100790
rect 25180 100710 25190 100790
rect 25360 100710 25370 100790
rect 25540 100710 25550 100790
rect 25720 100710 25730 100790
rect 25900 100710 25910 100790
rect 26080 100710 26090 100790
rect 26260 100710 26270 100790
rect 26440 100710 26450 100790
rect 26620 100710 26630 100790
rect 28930 100735 28940 100815
rect 29010 100735 29020 100815
rect 29090 100735 29100 100815
rect 29170 100735 29180 100815
rect 29250 100735 29260 100815
rect 29330 100735 29340 100815
rect 29410 100735 29420 100815
rect 29490 100735 29500 100815
rect 29570 100735 29580 100815
rect 30280 100790 30360 100800
rect 30460 100790 30540 100800
rect 30640 100790 30720 100800
rect 30820 100790 30900 100800
rect 31000 100790 31080 100800
rect 31180 100790 31260 100800
rect 31360 100790 31440 100800
rect 31540 100790 31620 100800
rect 31720 100790 31800 100800
rect 31900 100790 31980 100800
rect 32080 100790 32160 100800
rect 32260 100790 32340 100800
rect 32440 100790 32520 100800
rect 32620 100790 32700 100800
rect 32800 100790 32880 100800
rect 32980 100790 33060 100800
rect 33160 100790 33240 100800
rect 33340 100790 33420 100800
rect 33520 100790 33600 100800
rect 33700 100790 33780 100800
rect 33880 100790 33960 100800
rect 34060 100790 34140 100800
rect 34240 100790 34320 100800
rect 34420 100790 34500 100800
rect 34600 100790 34680 100800
rect 34780 100790 34860 100800
rect 34960 100790 35040 100800
rect 35140 100790 35220 100800
rect 35320 100790 35400 100800
rect 35500 100790 35580 100800
rect 35680 100790 35760 100800
rect 35860 100790 35940 100800
rect 36040 100790 36120 100800
rect 36220 100790 36300 100800
rect 36400 100790 36480 100800
rect 36580 100790 36660 100800
rect 36760 100790 36840 100800
rect 36940 100790 37020 100800
rect 37120 100790 37200 100800
rect 37300 100790 37380 100800
rect 37480 100790 37560 100800
rect 37660 100790 37740 100800
rect 37840 100790 37920 100800
rect 152080 100790 152160 100800
rect 152260 100790 152340 100800
rect 152440 100790 152520 100800
rect 152620 100790 152700 100800
rect 152800 100790 152880 100800
rect 152980 100790 153060 100800
rect 153160 100790 153240 100800
rect 153340 100790 153420 100800
rect 153520 100790 153600 100800
rect 153700 100790 153780 100800
rect 153880 100790 153960 100800
rect 154060 100790 154140 100800
rect 154240 100790 154320 100800
rect 154420 100790 154500 100800
rect 154600 100790 154680 100800
rect 154780 100790 154860 100800
rect 154960 100790 155040 100800
rect 155140 100790 155220 100800
rect 155320 100790 155400 100800
rect 155500 100790 155580 100800
rect 155680 100790 155760 100800
rect 155860 100790 155940 100800
rect 156040 100790 156120 100800
rect 156220 100790 156300 100800
rect 156400 100790 156480 100800
rect 156580 100790 156660 100800
rect 156760 100790 156840 100800
rect 156940 100790 157020 100800
rect 157120 100790 157200 100800
rect 157300 100790 157380 100800
rect 157480 100790 157560 100800
rect 157660 100790 157740 100800
rect 157840 100790 157920 100800
rect 158020 100790 158100 100800
rect 158200 100790 158280 100800
rect 158380 100790 158460 100800
rect 158560 100790 158640 100800
rect 158740 100790 158820 100800
rect 158920 100790 159000 100800
rect 159100 100790 159180 100800
rect 159280 100790 159360 100800
rect 159460 100790 159540 100800
rect 159640 100790 159720 100800
rect 30360 100710 30370 100790
rect 30540 100710 30550 100790
rect 30720 100710 30730 100790
rect 30900 100710 30910 100790
rect 31080 100710 31090 100790
rect 31260 100710 31270 100790
rect 31440 100710 31450 100790
rect 31620 100710 31630 100790
rect 31800 100710 31810 100790
rect 31980 100710 31990 100790
rect 32160 100710 32170 100790
rect 32340 100710 32350 100790
rect 32520 100710 32530 100790
rect 32700 100710 32710 100790
rect 32880 100710 32890 100790
rect 33060 100710 33070 100790
rect 33240 100710 33250 100790
rect 33420 100710 33430 100790
rect 33600 100710 33610 100790
rect 33780 100710 33790 100790
rect 33960 100710 33970 100790
rect 34140 100710 34150 100790
rect 34320 100710 34330 100790
rect 34500 100710 34510 100790
rect 34680 100710 34690 100790
rect 34860 100710 34870 100790
rect 35040 100710 35050 100790
rect 35220 100710 35230 100790
rect 35400 100710 35410 100790
rect 35580 100710 35590 100790
rect 35760 100710 35770 100790
rect 35940 100710 35950 100790
rect 36120 100710 36130 100790
rect 36300 100710 36310 100790
rect 36480 100710 36490 100790
rect 36660 100710 36670 100790
rect 36840 100710 36850 100790
rect 37020 100710 37030 100790
rect 37200 100710 37210 100790
rect 37380 100710 37390 100790
rect 37560 100710 37570 100790
rect 37740 100710 37750 100790
rect 37920 100710 37930 100790
rect 40060 100690 40120 100720
rect 41540 100690 41600 100720
rect 42360 100690 42420 100720
rect 43840 100690 43900 100720
rect 152160 100710 152170 100790
rect 152340 100710 152350 100790
rect 152520 100710 152530 100790
rect 152700 100710 152710 100790
rect 152880 100710 152890 100790
rect 153060 100710 153070 100790
rect 153240 100710 153250 100790
rect 153420 100710 153430 100790
rect 153600 100710 153610 100790
rect 153780 100710 153790 100790
rect 153960 100710 153970 100790
rect 154140 100710 154150 100790
rect 154320 100710 154330 100790
rect 154500 100710 154510 100790
rect 154680 100710 154690 100790
rect 154860 100710 154870 100790
rect 155040 100710 155050 100790
rect 155220 100710 155230 100790
rect 155400 100710 155410 100790
rect 155580 100710 155590 100790
rect 155760 100710 155770 100790
rect 155940 100710 155950 100790
rect 156120 100710 156130 100790
rect 156300 100710 156310 100790
rect 156480 100710 156490 100790
rect 156660 100710 156670 100790
rect 156840 100710 156850 100790
rect 157020 100710 157030 100790
rect 157200 100710 157210 100790
rect 157380 100710 157390 100790
rect 157560 100710 157570 100790
rect 157740 100710 157750 100790
rect 157920 100710 157930 100790
rect 158100 100710 158110 100790
rect 158280 100710 158290 100790
rect 158460 100710 158470 100790
rect 158640 100710 158650 100790
rect 158820 100710 158830 100790
rect 159000 100710 159010 100790
rect 159180 100710 159190 100790
rect 159360 100710 159370 100790
rect 159540 100710 159550 100790
rect 159720 100710 159730 100790
rect 161965 100765 161975 100845
rect 162145 100765 162155 100845
rect 162325 100765 162335 100845
rect 162505 100765 162515 100845
rect 162685 100765 162695 100845
rect 163380 100790 163460 100800
rect 163560 100790 163640 100800
rect 163740 100790 163820 100800
rect 163920 100790 164000 100800
rect 164100 100790 164180 100800
rect 164280 100790 164360 100800
rect 164460 100790 164540 100800
rect 164640 100790 164720 100800
rect 164820 100790 164900 100800
rect 165000 100790 165080 100800
rect 165180 100790 165260 100800
rect 165360 100790 165440 100800
rect 165540 100790 165620 100800
rect 165720 100790 165800 100800
rect 165900 100790 165980 100800
rect 166080 100790 166160 100800
rect 166260 100790 166340 100800
rect 166440 100790 166520 100800
rect 166620 100790 166700 100800
rect 166800 100790 166880 100800
rect 166980 100790 167060 100800
rect 167160 100790 167240 100800
rect 167340 100790 167420 100800
rect 167520 100790 167600 100800
rect 167700 100790 167780 100800
rect 167880 100790 167960 100800
rect 168060 100790 168140 100800
rect 168240 100790 168320 100800
rect 168420 100790 168500 100800
rect 168600 100790 168680 100800
rect 168780 100790 168860 100800
rect 168960 100790 169040 100800
rect 169140 100790 169220 100800
rect 169320 100790 169400 100800
rect 169500 100790 169580 100800
rect 169680 100790 169760 100800
rect 169860 100790 169940 100800
rect 170040 100790 170120 100800
rect 170220 100790 170300 100800
rect 170400 100790 170480 100800
rect 170580 100790 170660 100800
rect 170760 100790 170840 100800
rect 170940 100790 171020 100800
rect 163460 100710 163470 100790
rect 163640 100710 163650 100790
rect 163820 100710 163830 100790
rect 164000 100710 164010 100790
rect 164180 100710 164190 100790
rect 164360 100710 164370 100790
rect 164540 100710 164550 100790
rect 164720 100710 164730 100790
rect 164900 100710 164910 100790
rect 165080 100710 165090 100790
rect 165260 100710 165270 100790
rect 165440 100710 165450 100790
rect 165620 100710 165630 100790
rect 165800 100710 165810 100790
rect 165980 100710 165990 100790
rect 166160 100710 166170 100790
rect 166340 100710 166350 100790
rect 166520 100710 166530 100790
rect 166700 100710 166710 100790
rect 166880 100710 166890 100790
rect 167060 100710 167070 100790
rect 167240 100710 167250 100790
rect 167420 100710 167430 100790
rect 167600 100710 167610 100790
rect 167780 100710 167790 100790
rect 167960 100710 167970 100790
rect 168140 100710 168150 100790
rect 168320 100710 168330 100790
rect 168500 100710 168510 100790
rect 168680 100710 168690 100790
rect 168860 100710 168870 100790
rect 169040 100710 169050 100790
rect 169220 100710 169230 100790
rect 169400 100710 169410 100790
rect 169580 100710 169590 100790
rect 169760 100710 169770 100790
rect 169940 100710 169950 100790
rect 170120 100710 170130 100790
rect 170300 100710 170310 100790
rect 170480 100710 170490 100790
rect 170660 100710 170670 100790
rect 170840 100710 170850 100790
rect 171020 100710 171030 100790
rect 146100 100650 146160 100680
rect 147580 100650 147640 100680
rect 148400 100650 148460 100680
rect 149880 100650 149940 100680
rect 161885 100665 161965 100675
rect 162065 100665 162145 100675
rect 162245 100665 162325 100675
rect 162425 100665 162505 100675
rect 162605 100665 162685 100675
rect 40060 100570 40120 100600
rect 41540 100570 41600 100600
rect 42360 100570 42420 100600
rect 43840 100570 43900 100600
rect 146100 100530 146160 100560
rect 146210 100540 146220 100630
rect 40060 100450 40120 100480
rect 41540 100450 41600 100480
rect 42360 100450 42420 100480
rect 43840 100450 43900 100480
rect 19130 100410 19160 100440
rect 19250 100410 19280 100440
rect 26420 100410 26450 100440
rect 26540 100410 26570 100440
rect 30420 100410 30450 100440
rect 30540 100410 30570 100440
rect 37720 100410 37750 100440
rect 37840 100410 37870 100440
rect 146100 100410 146160 100440
rect 19010 100380 19070 100410
rect 19130 100380 19190 100410
rect 19250 100380 19310 100410
rect 26300 100380 26360 100410
rect 26420 100380 26480 100410
rect 26540 100380 26600 100410
rect 30300 100380 30360 100410
rect 30420 100380 30480 100410
rect 30540 100380 30600 100410
rect 37600 100380 37660 100410
rect 37720 100380 37780 100410
rect 37840 100380 37900 100410
rect 40060 100330 40120 100360
rect 41540 100330 41600 100360
rect 42360 100330 42420 100360
rect 43840 100330 43900 100360
rect 19130 100290 19160 100320
rect 19250 100290 19280 100320
rect 26420 100290 26450 100320
rect 26540 100290 26570 100320
rect 30420 100290 30450 100320
rect 30540 100290 30570 100320
rect 37720 100290 37750 100320
rect 37840 100290 37870 100320
rect 146100 100290 146160 100320
rect 19010 100260 19070 100290
rect 19130 100260 19190 100290
rect 19250 100260 19310 100290
rect 26300 100260 26360 100290
rect 26420 100260 26480 100290
rect 26540 100260 26600 100290
rect 30300 100260 30360 100290
rect 30420 100260 30480 100290
rect 30540 100260 30600 100290
rect 37600 100260 37660 100290
rect 37720 100260 37780 100290
rect 37840 100260 37900 100290
rect 31010 100245 37190 100260
rect 36000 100170 37190 100245
rect 40060 100210 40120 100240
rect 41540 100210 41600 100240
rect 42360 100210 42420 100240
rect 43840 100210 43900 100240
rect 37720 100170 37750 100200
rect 37840 100170 37870 100200
rect 146100 100170 146160 100200
rect 36120 100150 36130 100170
rect 36300 100150 36310 100170
rect 36480 100150 36490 100170
rect 36660 100150 36670 100170
rect 36840 100150 36850 100170
rect 37020 100150 37030 100170
rect 36040 100080 36120 100090
rect 36220 100080 36300 100090
rect 36400 100080 36480 100090
rect 36580 100080 36660 100090
rect 36760 100080 36840 100090
rect 36940 100080 37020 100090
rect 36120 100000 36130 100080
rect 36300 100000 36310 100080
rect 36480 100000 36490 100080
rect 36660 100000 36670 100080
rect 36840 100000 36850 100080
rect 37020 100000 37030 100080
rect 37100 99940 37190 100170
rect 37600 100140 37660 100170
rect 37720 100140 37780 100170
rect 37840 100140 37900 100170
rect 40060 100090 40120 100120
rect 41540 100090 41600 100120
rect 42360 100090 42420 100120
rect 43840 100090 43900 100120
rect 37720 100050 37750 100080
rect 37840 100050 37870 100080
rect 146100 100050 146160 100080
rect 37600 100020 37660 100050
rect 37720 100020 37780 100050
rect 37840 100020 37900 100050
rect 40060 99970 40120 100000
rect 41540 99970 41600 100000
rect 42360 99970 42420 100000
rect 43840 99970 43900 100000
rect 36000 99910 37190 99940
rect 37720 99930 37750 99960
rect 37840 99930 37870 99960
rect 146100 99930 146160 99960
rect 36120 99850 36130 99910
rect 36300 99850 36310 99910
rect 36480 99850 36490 99910
rect 36660 99850 36670 99910
rect 36840 99850 36850 99910
rect 37020 99850 37030 99910
rect 37100 99840 37190 99910
rect 37600 99900 37660 99930
rect 37720 99900 37780 99930
rect 37840 99900 37900 99930
rect 40060 99850 40120 99880
rect 41540 99850 41600 99880
rect 42360 99850 42420 99880
rect 43840 99850 43900 99880
rect 36000 99810 37190 99840
rect 37720 99810 37750 99840
rect 37840 99810 37870 99840
rect 146100 99810 146160 99840
rect 37100 99800 37190 99810
rect 36000 99790 37190 99800
rect 36040 99610 36120 99620
rect 36220 99610 36300 99620
rect 36400 99610 36480 99620
rect 36580 99610 36660 99620
rect 36760 99610 36840 99620
rect 36940 99610 37020 99620
rect 36120 99530 36130 99610
rect 36300 99530 36310 99610
rect 36480 99530 36490 99610
rect 36660 99530 36670 99610
rect 36840 99530 36850 99610
rect 37020 99530 37030 99610
rect 36040 99290 36120 99300
rect 36220 99290 36300 99300
rect 36400 99290 36480 99300
rect 36580 99290 36660 99300
rect 36760 99290 36840 99300
rect 36940 99290 37020 99300
rect 36120 99210 36130 99290
rect 36300 99210 36310 99290
rect 36480 99210 36490 99290
rect 36660 99210 36670 99290
rect 36840 99210 36850 99290
rect 37020 99210 37030 99290
rect 37100 99120 37190 99790
rect 37600 99780 37660 99810
rect 37720 99780 37780 99810
rect 37840 99780 37900 99810
rect 40060 99730 40120 99760
rect 41540 99730 41600 99760
rect 42360 99730 42420 99760
rect 43840 99730 43900 99760
rect 37720 99690 37750 99720
rect 37840 99690 37870 99720
rect 146100 99690 146160 99720
rect 37600 99660 37660 99690
rect 37720 99660 37780 99690
rect 37840 99660 37900 99690
rect 40060 99610 40120 99640
rect 41540 99610 41600 99640
rect 42360 99610 42420 99640
rect 43840 99610 43900 99640
rect 37720 99570 37750 99600
rect 37840 99570 37870 99600
rect 146100 99570 146160 99600
rect 37600 99540 37660 99570
rect 37720 99540 37780 99570
rect 37840 99540 37900 99570
rect 40060 99490 40120 99520
rect 41540 99490 41600 99520
rect 42360 99490 42420 99520
rect 43840 99490 43900 99520
rect 37720 99450 37750 99480
rect 37840 99450 37870 99480
rect 146100 99450 146160 99480
rect 37600 99420 37660 99450
rect 37720 99420 37780 99450
rect 37840 99420 37900 99450
rect 40060 99370 40120 99400
rect 41540 99370 41600 99400
rect 42360 99370 42420 99400
rect 43840 99370 43900 99400
rect 37720 99330 37750 99360
rect 37840 99330 37870 99360
rect 146100 99330 146160 99360
rect 37600 99300 37660 99330
rect 37720 99300 37780 99330
rect 37840 99300 37900 99330
rect 40060 99250 40120 99280
rect 41540 99250 41600 99280
rect 42360 99250 42420 99280
rect 43840 99250 43900 99280
rect 37720 99210 37750 99240
rect 37840 99210 37870 99240
rect 146100 99210 146160 99240
rect 37600 99180 37660 99210
rect 37720 99180 37780 99210
rect 37840 99180 37900 99210
rect 40060 99130 40120 99160
rect 41540 99130 41600 99160
rect 42360 99130 42420 99160
rect 43840 99130 43900 99160
rect 146300 99150 146310 100540
rect 146690 100500 146810 100560
rect 146970 100500 147090 100560
rect 147580 100530 147640 100560
rect 148400 100530 148460 100560
rect 148820 100550 149620 100640
rect 148950 100520 149070 100550
rect 149230 100520 149350 100550
rect 149070 100510 149130 100520
rect 149350 100510 149410 100520
rect 149070 100500 149190 100510
rect 149350 100500 149470 100510
rect 146810 100490 146870 100500
rect 146570 100480 146650 100490
rect 146810 100480 146930 100490
rect 146650 100400 146660 100480
rect 146810 100380 146870 100480
rect 146930 100400 146940 100480
rect 147090 100380 147150 100500
rect 146410 100330 147140 100340
rect 146410 100250 146420 100330
rect 147220 100325 147230 100380
rect 147270 100350 147390 100410
rect 146460 100315 147250 100325
rect 146450 100265 146460 100315
rect 146500 100060 146510 100250
rect 146690 100200 146810 100260
rect 146970 100200 147090 100260
rect 147220 100236 147230 100315
rect 147390 100236 147450 100350
rect 147520 100236 147530 100470
rect 147580 100410 147640 100440
rect 148400 100410 148460 100440
rect 148510 100400 148520 100490
rect 147580 100290 147640 100320
rect 148400 100290 148460 100320
rect 148600 100236 148610 100400
rect 148650 100370 148770 100430
rect 149070 100400 149130 100500
rect 149190 100420 149200 100500
rect 149350 100400 149410 100500
rect 149470 100420 149480 100500
rect 148770 100345 148830 100370
rect 149530 100365 149620 100550
rect 148910 100360 149620 100365
rect 148900 100350 149630 100360
rect 148910 100345 149630 100350
rect 148770 100335 149630 100345
rect 148770 100250 148830 100335
rect 149530 100285 149630 100335
rect 148910 100255 149630 100285
rect 148950 100236 149070 100255
rect 149230 100236 149350 100255
rect 149530 100236 149630 100255
rect 149820 100236 149830 100650
rect 152080 100640 152160 100650
rect 152260 100640 152340 100650
rect 152440 100640 152520 100650
rect 152620 100640 152700 100650
rect 152800 100640 152880 100650
rect 152980 100640 153060 100650
rect 153160 100640 153240 100650
rect 153340 100640 153420 100650
rect 153520 100640 153600 100650
rect 153700 100640 153780 100650
rect 153880 100640 153960 100650
rect 154060 100640 154140 100650
rect 154240 100640 154320 100650
rect 154420 100640 154500 100650
rect 154600 100640 154680 100650
rect 154780 100640 154860 100650
rect 154960 100640 155040 100650
rect 155140 100640 155220 100650
rect 155320 100640 155400 100650
rect 155500 100640 155580 100650
rect 155680 100640 155760 100650
rect 155860 100640 155940 100650
rect 156040 100640 156120 100650
rect 156220 100640 156300 100650
rect 156400 100640 156480 100650
rect 156580 100640 156660 100650
rect 156760 100640 156840 100650
rect 156940 100640 157020 100650
rect 157120 100640 157200 100650
rect 157300 100640 157380 100650
rect 157480 100640 157560 100650
rect 157660 100640 157740 100650
rect 157840 100640 157920 100650
rect 158020 100640 158100 100650
rect 158200 100640 158280 100650
rect 158380 100640 158460 100650
rect 158560 100640 158640 100650
rect 158740 100640 158820 100650
rect 158920 100640 159000 100650
rect 159100 100640 159180 100650
rect 159280 100640 159360 100650
rect 159460 100640 159540 100650
rect 159640 100640 159720 100650
rect 152160 100560 152170 100640
rect 152340 100560 152350 100640
rect 152520 100560 152530 100640
rect 152700 100560 152710 100640
rect 152880 100560 152890 100640
rect 153060 100560 153070 100640
rect 153240 100560 153250 100640
rect 153420 100560 153430 100640
rect 153600 100560 153610 100640
rect 153780 100560 153790 100640
rect 153960 100560 153970 100640
rect 154140 100560 154150 100640
rect 154320 100560 154330 100640
rect 154500 100560 154510 100640
rect 154680 100560 154690 100640
rect 154860 100560 154870 100640
rect 155040 100560 155050 100640
rect 155220 100560 155230 100640
rect 155400 100560 155410 100640
rect 155580 100560 155590 100640
rect 155760 100560 155770 100640
rect 155940 100560 155950 100640
rect 156120 100560 156130 100640
rect 156300 100560 156310 100640
rect 156480 100560 156490 100640
rect 156660 100560 156670 100640
rect 156840 100560 156850 100640
rect 157020 100560 157030 100640
rect 157200 100560 157210 100640
rect 157380 100560 157390 100640
rect 157560 100560 157570 100640
rect 157740 100560 157750 100640
rect 157920 100560 157930 100640
rect 158100 100560 158110 100640
rect 158280 100560 158290 100640
rect 158460 100560 158470 100640
rect 158640 100560 158650 100640
rect 158820 100560 158830 100640
rect 159000 100560 159010 100640
rect 159180 100560 159190 100640
rect 159360 100560 159370 100640
rect 159540 100560 159550 100640
rect 159720 100560 159730 100640
rect 161965 100585 161975 100665
rect 162145 100585 162155 100665
rect 162325 100585 162335 100665
rect 162505 100585 162515 100665
rect 162685 100585 162695 100665
rect 163380 100640 163460 100650
rect 163560 100640 163640 100650
rect 163740 100640 163820 100650
rect 163920 100640 164000 100650
rect 164100 100640 164180 100650
rect 164280 100640 164360 100650
rect 164460 100640 164540 100650
rect 164640 100640 164720 100650
rect 164820 100640 164900 100650
rect 165000 100640 165080 100650
rect 165180 100640 165260 100650
rect 165360 100640 165440 100650
rect 165540 100640 165620 100650
rect 165720 100640 165800 100650
rect 165900 100640 165980 100650
rect 166080 100640 166160 100650
rect 166260 100640 166340 100650
rect 166440 100640 166520 100650
rect 166620 100640 166700 100650
rect 166800 100640 166880 100650
rect 166980 100640 167060 100650
rect 167160 100640 167240 100650
rect 167340 100640 167420 100650
rect 167520 100640 167600 100650
rect 167700 100640 167780 100650
rect 167880 100640 167960 100650
rect 168060 100640 168140 100650
rect 168240 100640 168320 100650
rect 168420 100640 168500 100650
rect 168600 100640 168680 100650
rect 168780 100640 168860 100650
rect 168960 100640 169040 100650
rect 169140 100640 169220 100650
rect 169320 100640 169400 100650
rect 169500 100640 169580 100650
rect 169680 100640 169760 100650
rect 169860 100640 169940 100650
rect 170040 100640 170120 100650
rect 170220 100640 170300 100650
rect 170400 100640 170480 100650
rect 170580 100640 170660 100650
rect 170760 100640 170840 100650
rect 170940 100640 171020 100650
rect 163460 100560 163470 100640
rect 163640 100560 163650 100640
rect 163820 100560 163830 100640
rect 164000 100560 164010 100640
rect 164180 100560 164190 100640
rect 164360 100560 164370 100640
rect 164540 100560 164550 100640
rect 164720 100560 164730 100640
rect 164900 100560 164910 100640
rect 165080 100560 165090 100640
rect 165260 100560 165270 100640
rect 165440 100560 165450 100640
rect 165620 100560 165630 100640
rect 165800 100560 165810 100640
rect 165980 100560 165990 100640
rect 166160 100560 166170 100640
rect 166340 100560 166350 100640
rect 166520 100560 166530 100640
rect 166700 100560 166710 100640
rect 166880 100560 166890 100640
rect 167060 100560 167070 100640
rect 167240 100560 167250 100640
rect 167420 100560 167430 100640
rect 167600 100560 167610 100640
rect 167780 100560 167790 100640
rect 167960 100560 167970 100640
rect 168140 100560 168150 100640
rect 168320 100560 168330 100640
rect 168500 100560 168510 100640
rect 168680 100560 168690 100640
rect 168860 100560 168870 100640
rect 169040 100560 169050 100640
rect 169220 100560 169230 100640
rect 169400 100560 169410 100640
rect 169580 100560 169590 100640
rect 169760 100560 169770 100640
rect 169940 100560 169950 100640
rect 170120 100560 170130 100640
rect 170300 100560 170310 100640
rect 170480 100560 170490 100640
rect 170660 100560 170670 100640
rect 170840 100560 170850 100640
rect 171020 100560 171030 100640
rect 149880 100530 149940 100560
rect 149880 100410 149940 100440
rect 152220 100390 152250 100420
rect 152340 100390 152370 100420
rect 159520 100390 159550 100420
rect 159640 100390 159670 100420
rect 152100 100360 152160 100390
rect 152220 100360 152280 100390
rect 152340 100360 152400 100390
rect 159400 100360 159460 100390
rect 159520 100360 159580 100390
rect 159640 100360 159700 100390
rect 149880 100290 149940 100320
rect 152220 100270 152250 100300
rect 152340 100270 152370 100300
rect 159520 100270 159550 100300
rect 159640 100270 159670 100300
rect 163520 100270 163550 100300
rect 163640 100270 163670 100300
rect 170810 100270 170840 100300
rect 170930 100270 170960 100300
rect 152100 100240 152160 100270
rect 152220 100240 152280 100270
rect 152340 100240 152400 100270
rect 152810 100236 158990 100260
rect 159400 100240 159460 100270
rect 159520 100240 159580 100270
rect 159640 100240 159700 100270
rect 163400 100240 163460 100270
rect 163520 100240 163580 100270
rect 163640 100240 163700 100270
rect 170690 100240 170750 100270
rect 170810 100240 170870 100270
rect 170930 100240 170990 100270
rect 164280 100236 164360 100240
rect 164460 100236 164540 100240
rect 164640 100236 164720 100240
rect 164820 100236 164900 100240
rect 165000 100236 165080 100240
rect 165180 100236 165260 100240
rect 165360 100236 165440 100240
rect 165540 100236 165620 100240
rect 165720 100236 165800 100240
rect 165900 100236 165980 100240
rect 166080 100236 166160 100240
rect 166260 100236 166340 100240
rect 166440 100236 166520 100240
rect 166620 100236 166700 100240
rect 166800 100236 166880 100240
rect 166980 100236 167060 100240
rect 167160 100236 167240 100240
rect 167340 100236 167420 100240
rect 167520 100236 167600 100240
rect 167700 100236 167780 100240
rect 167880 100236 167960 100240
rect 168060 100236 168140 100240
rect 168240 100236 168320 100240
rect 168420 100236 168500 100240
rect 168600 100236 168680 100240
rect 168780 100236 168860 100240
rect 168960 100236 169040 100240
rect 169140 100236 169220 100240
rect 169320 100236 169400 100240
rect 169500 100236 169580 100240
rect 169680 100236 169760 100240
rect 169860 100236 169940 100240
rect 170040 100236 170120 100240
rect 146810 100190 146870 100200
rect 146570 100180 146650 100190
rect 146710 100180 146790 100190
rect 146810 100180 146930 100190
rect 146990 100180 147070 100190
rect 146650 100100 146660 100180
rect 146790 100100 146800 100180
rect 146810 100080 146870 100180
rect 146930 100100 146940 100180
rect 147070 100100 147080 100180
rect 147090 100080 147150 100200
rect 146500 100050 147130 100060
rect 146500 100040 146510 100050
rect 146690 99910 146810 99970
rect 146970 99910 147090 99970
rect 146690 99820 146700 99910
rect 146800 99880 146870 99910
rect 146810 99790 146870 99880
rect 146970 99820 146980 99910
rect 147090 99790 147150 99910
rect 146410 99740 147140 99750
rect 146410 99660 146420 99740
rect 146460 99725 147150 99735
rect 146450 99675 146460 99725
rect 146500 99470 146510 99660
rect 146690 99610 146810 99670
rect 146970 99610 147090 99670
rect 146810 99600 146870 99610
rect 146570 99590 146650 99600
rect 146710 99590 146790 99600
rect 146810 99590 146930 99600
rect 146990 99590 147070 99600
rect 146650 99510 146660 99590
rect 146790 99510 146800 99590
rect 146810 99490 146870 99590
rect 146930 99510 146940 99590
rect 147070 99510 147080 99590
rect 147090 99490 147150 99610
rect 146500 99460 147130 99470
rect 146500 99450 146510 99460
rect 146690 99320 146810 99380
rect 146970 99320 147090 99380
rect 146690 99230 146700 99320
rect 146800 99290 146870 99320
rect 146810 99200 146870 99290
rect 146970 99230 146980 99320
rect 147090 99200 147150 99320
rect 146410 99150 147140 99160
rect 146460 99135 147150 99145
rect 36000 99110 37190 99120
rect 37100 99010 37190 99110
rect 37720 99090 37750 99120
rect 37840 99090 37870 99120
rect 146100 99090 146160 99120
rect 37600 99060 37660 99090
rect 37720 99060 37780 99090
rect 37840 99060 37900 99090
rect 146450 99085 146460 99135
rect 40060 99010 40120 99040
rect 41540 99010 41600 99040
rect 42360 99010 42420 99040
rect 43840 99010 43900 99040
rect 146690 99020 146810 99080
rect 146970 99020 147090 99080
rect 146810 99010 146870 99020
rect 36000 98980 37190 99010
rect 146570 99000 146650 99010
rect 146710 99000 146790 99010
rect 146810 99000 146930 99010
rect 146990 99000 147070 99010
rect 36040 98970 36120 98980
rect 36220 98970 36300 98980
rect 36400 98970 36480 98980
rect 36580 98970 36660 98980
rect 36760 98970 36840 98980
rect 36940 98970 37020 98980
rect 36120 98910 36130 98970
rect 36300 98910 36310 98970
rect 36480 98910 36490 98970
rect 36660 98910 36670 98970
rect 36840 98910 36850 98970
rect 37020 98910 37030 98970
rect 37100 98910 37190 98980
rect 37720 98970 37750 99000
rect 37840 98970 37870 99000
rect 146100 98970 146160 99000
rect 37600 98940 37660 98970
rect 37720 98940 37780 98970
rect 37840 98940 37900 98970
rect 146650 98920 146660 99000
rect 146790 98920 146800 99000
rect 36000 98880 37190 98910
rect 40060 98890 40120 98920
rect 41540 98890 41600 98920
rect 42360 98890 42420 98920
rect 43840 98890 43900 98920
rect 146810 98900 146870 99000
rect 146930 98920 146940 99000
rect 147070 98920 147080 99000
rect 147090 98900 147150 99020
rect 36040 98820 36120 98830
rect 36220 98820 36300 98830
rect 36400 98820 36480 98830
rect 36580 98820 36660 98830
rect 36760 98820 36840 98830
rect 36940 98820 37020 98830
rect 36120 98740 36130 98820
rect 36300 98740 36310 98820
rect 36480 98740 36490 98820
rect 36660 98740 36670 98820
rect 36840 98740 36850 98820
rect 37020 98740 37030 98820
rect 37100 98680 37190 98880
rect 37720 98850 37750 98880
rect 37840 98850 37870 98880
rect 146100 98850 146160 98880
rect 37600 98820 37660 98850
rect 37720 98820 37780 98850
rect 37840 98820 37900 98850
rect 40060 98770 40120 98800
rect 41540 98770 41600 98800
rect 42360 98770 42420 98800
rect 43840 98770 43900 98800
rect 37720 98730 37750 98760
rect 37840 98730 37870 98760
rect 146100 98730 146160 98760
rect 37600 98700 37660 98730
rect 37720 98700 37780 98730
rect 37840 98700 37900 98730
rect 36000 98650 37190 98680
rect 40060 98650 40120 98680
rect 41540 98650 41600 98680
rect 42360 98650 42420 98680
rect 43840 98650 43900 98680
rect 36120 98590 36130 98650
rect 36300 98590 36310 98650
rect 36480 98590 36490 98650
rect 36660 98590 36670 98650
rect 36840 98590 36850 98650
rect 37020 98590 37030 98650
rect 37100 98580 37190 98650
rect 37720 98610 37750 98640
rect 37840 98610 37870 98640
rect 146100 98610 146160 98640
rect 37600 98580 37660 98610
rect 37720 98580 37780 98610
rect 37840 98580 37900 98610
rect 36000 98550 37190 98580
rect 37100 98540 37190 98550
rect 36000 98530 37190 98540
rect 40060 98530 40120 98560
rect 41540 98530 41600 98560
rect 42360 98530 42420 98560
rect 43840 98530 43900 98560
rect 36040 98350 36120 98360
rect 36220 98350 36300 98360
rect 36400 98350 36480 98360
rect 36580 98350 36660 98360
rect 36760 98350 36840 98360
rect 36940 98350 37020 98360
rect 36120 98270 36130 98350
rect 36300 98270 36310 98350
rect 36480 98270 36490 98350
rect 36660 98270 36670 98350
rect 36840 98270 36850 98350
rect 37020 98270 37030 98350
rect 36040 98030 36120 98040
rect 36220 98030 36300 98040
rect 36400 98030 36480 98040
rect 36580 98030 36660 98040
rect 36760 98030 36840 98040
rect 36940 98030 37020 98040
rect 36120 97950 36130 98030
rect 36300 97950 36310 98030
rect 36480 97950 36490 98030
rect 36660 97950 36670 98030
rect 36840 97950 36850 98030
rect 37020 97950 37030 98030
rect 37100 97860 37190 98530
rect 37720 98490 37750 98520
rect 37840 98490 37870 98520
rect 146100 98490 146160 98520
rect 37600 98460 37660 98490
rect 37720 98460 37780 98490
rect 37840 98460 37900 98490
rect 146690 98440 146810 98500
rect 146970 98440 147090 98500
rect 40060 98410 40120 98440
rect 41540 98410 41600 98440
rect 42360 98410 42420 98440
rect 43840 98410 43900 98440
rect 146810 98430 146870 98440
rect 146570 98420 146650 98430
rect 146810 98420 146930 98430
rect 37720 98370 37750 98400
rect 37840 98370 37870 98400
rect 146100 98370 146160 98400
rect 37600 98340 37660 98370
rect 37720 98340 37780 98370
rect 37840 98340 37900 98370
rect 146650 98340 146660 98420
rect 146810 98320 146870 98420
rect 146930 98340 146940 98420
rect 147090 98320 147150 98440
rect 40060 98290 40120 98320
rect 41540 98290 41600 98320
rect 42360 98290 42420 98320
rect 43840 98290 43900 98320
rect 37720 98250 37750 98280
rect 37840 98250 37870 98280
rect 146100 98250 146160 98280
rect 146500 98270 147140 98280
rect 146460 98255 147150 98265
rect 37600 98220 37660 98250
rect 37720 98220 37780 98250
rect 37840 98220 37900 98250
rect 146450 98205 146460 98255
rect 40060 98170 40120 98200
rect 41540 98170 41600 98200
rect 42360 98170 42420 98200
rect 43840 98170 43900 98200
rect 37720 98130 37750 98160
rect 37840 98130 37870 98160
rect 146100 98130 146160 98160
rect 146690 98140 146810 98200
rect 146970 98140 147090 98200
rect 146810 98130 146870 98140
rect 37600 98100 37660 98130
rect 37720 98100 37780 98130
rect 37840 98100 37900 98130
rect 146570 98120 146650 98130
rect 146710 98120 146790 98130
rect 146810 98120 146930 98130
rect 146990 98120 147070 98130
rect 40060 98050 40120 98080
rect 41540 98050 41600 98080
rect 42360 98050 42420 98080
rect 43840 98050 43900 98080
rect 146650 98040 146660 98120
rect 146790 98040 146800 98120
rect 37720 98010 37750 98040
rect 37840 98010 37870 98040
rect 146100 98010 146160 98040
rect 146810 98020 146870 98120
rect 146930 98040 146940 98120
rect 147070 98040 147080 98120
rect 147090 98020 147150 98140
rect 37600 97980 37660 98010
rect 37720 97980 37780 98010
rect 37840 97980 37900 98010
rect 146510 97990 147130 98000
rect 40060 97930 40120 97960
rect 41540 97930 41600 97960
rect 42360 97930 42420 97960
rect 43840 97930 43900 97960
rect 37720 97890 37750 97920
rect 37840 97890 37870 97920
rect 146100 97890 146160 97920
rect 37600 97860 37660 97890
rect 37720 97860 37780 97890
rect 37840 97860 37900 97890
rect 146610 97860 146970 97920
rect 36000 97850 37190 97860
rect 37100 97750 37190 97850
rect 40060 97810 40120 97840
rect 41540 97810 41600 97840
rect 42360 97810 42420 97840
rect 43840 97810 43900 97840
rect 37720 97770 37750 97800
rect 37840 97770 37870 97800
rect 146100 97770 146160 97800
rect 36000 97720 37190 97750
rect 37600 97740 37660 97770
rect 37720 97740 37780 97770
rect 37840 97740 37900 97770
rect 146300 97730 146420 97790
rect 146420 97720 146480 97730
rect 36040 97710 36120 97720
rect 36220 97710 36300 97720
rect 36400 97710 36480 97720
rect 36580 97710 36660 97720
rect 36760 97710 36840 97720
rect 36940 97710 37020 97720
rect 36120 97650 36130 97710
rect 36300 97650 36310 97710
rect 36480 97650 36490 97710
rect 36660 97650 36670 97710
rect 36840 97650 36850 97710
rect 37020 97650 37030 97710
rect 37100 97650 37190 97720
rect 40060 97690 40120 97720
rect 41540 97690 41600 97720
rect 42360 97690 42420 97720
rect 43840 97690 43900 97720
rect 146420 97710 147050 97720
rect 146420 97705 146480 97710
rect 146420 97695 147090 97705
rect 37720 97650 37750 97680
rect 37840 97650 37870 97680
rect 146100 97650 146160 97680
rect 36000 97620 37190 97650
rect 37600 97620 37660 97650
rect 37720 97620 37780 97650
rect 37840 97620 37900 97650
rect 36040 97560 36120 97570
rect 36220 97560 36300 97570
rect 36400 97560 36480 97570
rect 36580 97560 36660 97570
rect 36760 97560 36840 97570
rect 36940 97560 37020 97570
rect 36120 97480 36130 97560
rect 36300 97480 36310 97560
rect 36480 97480 36490 97560
rect 36660 97480 36670 97560
rect 36840 97480 36850 97560
rect 37020 97480 37030 97560
rect 37100 97420 37190 97620
rect 146420 97610 146480 97695
rect 40060 97570 40120 97600
rect 41540 97570 41600 97600
rect 42360 97570 42420 97600
rect 43840 97570 43900 97600
rect 37720 97530 37750 97560
rect 37840 97530 37870 97560
rect 37600 97500 37660 97530
rect 37720 97500 37780 97530
rect 37840 97500 37900 97530
rect 40060 97450 40120 97480
rect 41540 97450 41600 97480
rect 42360 97450 42420 97480
rect 43840 97450 43900 97480
rect 36000 97390 37190 97420
rect 37720 97410 37750 97440
rect 37840 97410 37870 97440
rect 36120 97330 36130 97390
rect 36300 97330 36310 97390
rect 36480 97330 36490 97390
rect 36660 97330 36670 97390
rect 36840 97330 36850 97390
rect 37020 97330 37030 97390
rect 37100 97320 37190 97390
rect 37600 97380 37660 97410
rect 37720 97380 37780 97410
rect 37840 97380 37900 97410
rect 46660 97360 48000 97540
rect 146100 97530 146160 97560
rect 146300 97470 146420 97530
rect 146420 97445 146480 97470
rect 146530 97460 146540 97630
rect 146610 97600 146970 97660
rect 147090 97645 147100 97695
rect 146530 97450 147140 97460
rect 146100 97410 146160 97440
rect 146420 97435 147090 97445
rect 40060 97330 40120 97360
rect 41540 97330 41600 97360
rect 42360 97330 42420 97360
rect 43840 97330 43900 97360
rect 146420 97350 146480 97435
rect 146610 97340 146970 97400
rect 147090 97385 147100 97435
rect 36000 97290 37190 97320
rect 37720 97290 37750 97320
rect 37840 97290 37870 97320
rect 146100 97290 146160 97320
rect 37100 97280 37190 97290
rect 36000 97270 37190 97280
rect 36040 97090 36120 97100
rect 36220 97090 36300 97100
rect 36400 97090 36480 97100
rect 36580 97090 36660 97100
rect 36760 97090 36840 97100
rect 36940 97090 37020 97100
rect 36120 97010 36130 97090
rect 36300 97010 36310 97090
rect 36480 97010 36490 97090
rect 36660 97010 36670 97090
rect 36840 97010 36850 97090
rect 37020 97010 37030 97090
rect 36040 96770 36120 96780
rect 36220 96770 36300 96780
rect 36400 96770 36480 96780
rect 36580 96770 36660 96780
rect 36760 96770 36840 96780
rect 36940 96770 37020 96780
rect 36120 96690 36130 96770
rect 36300 96690 36310 96770
rect 36480 96690 36490 96770
rect 36660 96690 36670 96770
rect 36840 96690 36850 96770
rect 37020 96690 37030 96770
rect 37100 96600 37190 97270
rect 37600 97260 37660 97290
rect 37720 97260 37780 97290
rect 37840 97260 37900 97290
rect 40060 97210 40120 97240
rect 41540 97210 41600 97240
rect 42360 97210 42420 97240
rect 43840 97210 43900 97240
rect 146300 97210 146420 97270
rect 146420 97200 146480 97210
rect 37720 97170 37750 97200
rect 37840 97170 37870 97200
rect 146100 97170 146160 97200
rect 146420 97190 147050 97200
rect 146420 97185 146480 97190
rect 146420 97175 147090 97185
rect 37600 97140 37660 97170
rect 37720 97140 37780 97170
rect 37840 97140 37900 97170
rect 40060 97090 40120 97120
rect 41540 97090 41600 97120
rect 42360 97090 42420 97120
rect 43840 97090 43900 97120
rect 146420 97090 146480 97175
rect 37720 97050 37750 97080
rect 37840 97050 37870 97080
rect 146100 97050 146160 97080
rect 37600 97020 37660 97050
rect 37720 97020 37780 97050
rect 37840 97020 37900 97050
rect 40060 96970 40120 97000
rect 41540 96970 41600 97000
rect 42360 96970 42420 97000
rect 43840 96970 43900 97000
rect 37720 96930 37750 96960
rect 37840 96930 37870 96960
rect 146100 96930 146160 96960
rect 146300 96950 146420 97010
rect 37600 96900 37660 96930
rect 37720 96900 37780 96930
rect 37840 96900 37900 96930
rect 146420 96925 146480 96950
rect 146530 96940 146540 97110
rect 146610 97080 146970 97140
rect 147090 97125 147100 97175
rect 146530 96930 147140 96940
rect 146420 96915 147090 96925
rect 40060 96850 40120 96880
rect 41540 96850 41600 96880
rect 42360 96850 42420 96880
rect 43840 96850 43900 96880
rect 37720 96810 37750 96840
rect 37840 96810 37870 96840
rect 146100 96810 146160 96840
rect 146420 96830 146480 96915
rect 146610 96820 146970 96880
rect 147090 96865 147100 96915
rect 37600 96780 37660 96810
rect 37720 96780 37780 96810
rect 37840 96780 37900 96810
rect 40060 96730 40120 96760
rect 41540 96730 41600 96760
rect 42360 96730 42420 96760
rect 43840 96730 43900 96760
rect 37720 96690 37750 96720
rect 37840 96690 37870 96720
rect 146100 96690 146160 96720
rect 37600 96660 37660 96690
rect 37720 96660 37780 96690
rect 37840 96660 37900 96690
rect 40060 96610 40120 96640
rect 41540 96610 41600 96640
rect 42360 96610 42420 96640
rect 43840 96610 43900 96640
rect 36000 96590 37190 96600
rect 37100 96490 37190 96590
rect 37720 96570 37750 96600
rect 37840 96570 37870 96600
rect 146100 96570 146160 96600
rect 37600 96540 37660 96570
rect 37720 96540 37780 96570
rect 37840 96540 37900 96570
rect 40060 96490 40120 96520
rect 41540 96490 41600 96520
rect 42360 96490 42420 96520
rect 43840 96490 43900 96520
rect 36000 96460 37190 96490
rect 36040 96450 36120 96460
rect 36220 96450 36300 96460
rect 36400 96450 36480 96460
rect 36580 96450 36660 96460
rect 36760 96450 36840 96460
rect 36940 96450 37020 96460
rect 36120 96390 36130 96450
rect 36300 96390 36310 96450
rect 36480 96390 36490 96450
rect 36660 96390 36670 96450
rect 36840 96390 36850 96450
rect 37020 96390 37030 96450
rect 37100 96390 37190 96460
rect 37720 96450 37750 96480
rect 37840 96450 37870 96480
rect 146100 96450 146160 96480
rect 37600 96420 37660 96450
rect 37720 96420 37780 96450
rect 37840 96420 37900 96450
rect 36000 96360 37190 96390
rect 40060 96370 40120 96400
rect 41540 96370 41600 96400
rect 42360 96370 42420 96400
rect 43840 96370 43900 96400
rect 36040 96300 36120 96310
rect 36220 96300 36300 96310
rect 36400 96300 36480 96310
rect 36580 96300 36660 96310
rect 36760 96300 36840 96310
rect 36940 96300 37020 96310
rect 36120 96220 36130 96300
rect 36300 96220 36310 96300
rect 36480 96220 36490 96300
rect 36660 96220 36670 96300
rect 36840 96220 36850 96300
rect 37020 96220 37030 96300
rect 37100 96160 37190 96360
rect 37720 96330 37750 96360
rect 37840 96330 37870 96360
rect 146100 96330 146160 96360
rect 37600 96300 37660 96330
rect 37720 96300 37780 96330
rect 37840 96300 37900 96330
rect 40060 96250 40120 96280
rect 41540 96250 41600 96280
rect 42360 96250 42420 96280
rect 43840 96250 43900 96280
rect 37720 96210 37750 96240
rect 37840 96210 37870 96240
rect 146100 96210 146160 96240
rect 37600 96180 37660 96210
rect 37720 96180 37780 96210
rect 37840 96180 37900 96210
rect 36000 96130 37190 96160
rect 40060 96130 40120 96160
rect 41540 96130 41600 96160
rect 42360 96130 42420 96160
rect 43840 96130 43900 96160
rect 36120 96070 36130 96130
rect 36300 96070 36310 96130
rect 36480 96070 36490 96130
rect 36660 96070 36670 96130
rect 36840 96070 36850 96130
rect 37020 96070 37030 96130
rect 37100 96060 37190 96130
rect 37720 96090 37750 96120
rect 37840 96090 37870 96120
rect 146100 96090 146160 96120
rect 37600 96060 37660 96090
rect 37720 96060 37780 96090
rect 37840 96060 37900 96090
rect 36000 96030 37190 96060
rect 37100 96020 37190 96030
rect 36000 96010 37190 96020
rect 40060 96010 40120 96040
rect 41540 96010 41600 96040
rect 42360 96010 42420 96040
rect 43840 96010 43900 96040
rect 36040 95830 36120 95840
rect 36220 95830 36300 95840
rect 36400 95830 36480 95840
rect 36580 95830 36660 95840
rect 36760 95830 36840 95840
rect 36940 95830 37020 95840
rect 36120 95750 36130 95830
rect 36300 95750 36310 95830
rect 36480 95750 36490 95830
rect 36660 95750 36670 95830
rect 36840 95750 36850 95830
rect 37020 95750 37030 95830
rect 36040 95510 36120 95520
rect 36220 95510 36300 95520
rect 36400 95510 36480 95520
rect 36580 95510 36660 95520
rect 36760 95510 36840 95520
rect 36940 95510 37020 95520
rect 36120 95430 36130 95510
rect 36300 95430 36310 95510
rect 36480 95430 36490 95510
rect 36660 95430 36670 95510
rect 36840 95430 36850 95510
rect 37020 95430 37030 95510
rect 37100 95340 37190 96010
rect 37720 95970 37750 96000
rect 37840 95970 37870 96000
rect 146100 95970 146160 96000
rect 37600 95940 37660 95970
rect 37720 95940 37780 95970
rect 37840 95940 37900 95970
rect 40060 95890 40120 95920
rect 41540 95890 41600 95920
rect 42360 95890 42420 95920
rect 43840 95890 43900 95920
rect 37720 95850 37750 95880
rect 37840 95850 37870 95880
rect 146100 95850 146160 95880
rect 37600 95820 37660 95850
rect 37720 95820 37780 95850
rect 37840 95820 37900 95850
rect 40060 95770 40120 95800
rect 41540 95770 41600 95800
rect 42360 95770 42420 95800
rect 43840 95770 43900 95800
rect 37720 95730 37750 95760
rect 37840 95730 37870 95760
rect 146100 95730 146160 95760
rect 37600 95700 37660 95730
rect 37720 95700 37780 95730
rect 37840 95700 37900 95730
rect 40060 95650 40120 95680
rect 41540 95650 41600 95680
rect 42360 95650 42420 95680
rect 43840 95650 43900 95680
rect 37720 95610 37750 95640
rect 37840 95610 37870 95640
rect 146100 95610 146160 95640
rect 37600 95580 37660 95610
rect 37720 95580 37780 95610
rect 37840 95580 37900 95610
rect 40060 95530 40120 95560
rect 41540 95530 41600 95560
rect 42360 95530 42420 95560
rect 43840 95530 43900 95560
rect 37720 95490 37750 95520
rect 37840 95490 37870 95520
rect 146100 95490 146160 95520
rect 37600 95460 37660 95490
rect 37720 95460 37780 95490
rect 37840 95460 37900 95490
rect 40060 95410 40120 95440
rect 41540 95410 41600 95440
rect 42360 95410 42420 95440
rect 43840 95410 43900 95440
rect 37720 95370 37750 95400
rect 37840 95370 37870 95400
rect 146100 95370 146160 95400
rect 37600 95340 37660 95370
rect 37720 95340 37780 95370
rect 37840 95340 37900 95370
rect 36000 95330 37190 95340
rect 37100 95230 37190 95330
rect 40060 95290 40120 95320
rect 41540 95290 41600 95320
rect 42360 95290 42420 95320
rect 43840 95290 43900 95320
rect 37720 95250 37750 95280
rect 37840 95250 37870 95280
rect 146100 95250 146160 95280
rect 36000 95200 37190 95230
rect 37600 95220 37660 95250
rect 37720 95220 37780 95250
rect 37840 95220 37900 95250
rect 40685 95210 40925 95240
rect 36040 95190 36120 95200
rect 36220 95190 36300 95200
rect 36400 95190 36480 95200
rect 36580 95190 36660 95200
rect 36760 95190 36840 95200
rect 36940 95190 37020 95200
rect 36120 95130 36130 95190
rect 36300 95130 36310 95190
rect 36480 95130 36490 95190
rect 36660 95130 36670 95190
rect 36840 95130 36850 95190
rect 37020 95130 37030 95190
rect 37100 95130 37190 95200
rect 40060 95170 40120 95200
rect 37720 95130 37750 95160
rect 37840 95130 37870 95160
rect 40685 95150 40715 95210
rect 40775 95150 40865 95210
rect 40895 95150 40925 95210
rect 41540 95170 41600 95200
rect 42360 95170 42420 95200
rect 43840 95170 43900 95200
rect 36000 95100 37190 95130
rect 37600 95100 37660 95130
rect 37720 95100 37780 95130
rect 37840 95100 37900 95130
rect 40685 95120 40925 95150
rect 146100 95130 146160 95160
rect 36040 95040 36120 95050
rect 36220 95040 36300 95050
rect 36400 95040 36480 95050
rect 36580 95040 36660 95050
rect 36760 95040 36840 95050
rect 36940 95040 37020 95050
rect 36120 94960 36130 95040
rect 36300 94960 36310 95040
rect 36480 94960 36490 95040
rect 36660 94960 36670 95040
rect 36840 94960 36850 95040
rect 37020 94960 37030 95040
rect 37100 94900 37190 95100
rect 40060 95050 40120 95080
rect 41540 95050 41600 95080
rect 42360 95050 42420 95080
rect 43840 95050 43900 95080
rect 37720 95010 37750 95040
rect 37840 95010 37870 95040
rect 146100 95010 146160 95040
rect 37600 94980 37660 95010
rect 37720 94980 37780 95010
rect 37840 94980 37900 95010
rect 40060 94930 40120 94960
rect 41540 94930 41600 94960
rect 42360 94930 42420 94960
rect 43840 94930 43900 94960
rect 36000 94870 37190 94900
rect 37720 94890 37750 94920
rect 37840 94890 37870 94920
rect 146100 94890 146160 94920
rect 36120 94810 36130 94870
rect 36300 94810 36310 94870
rect 36480 94810 36490 94870
rect 36660 94810 36670 94870
rect 36840 94810 36850 94870
rect 37020 94810 37030 94870
rect 37100 94800 37190 94870
rect 37600 94860 37660 94890
rect 37720 94860 37780 94890
rect 37840 94860 37900 94890
rect 40060 94810 40120 94840
rect 41540 94810 41600 94840
rect 42360 94810 42420 94840
rect 43840 94810 43900 94840
rect 36000 94770 37190 94800
rect 37720 94770 37750 94800
rect 37840 94770 37870 94800
rect 146100 94770 146160 94800
rect 37100 94760 37190 94770
rect 36000 94750 37190 94760
rect 36040 94570 36120 94580
rect 36220 94570 36300 94580
rect 36400 94570 36480 94580
rect 36580 94570 36660 94580
rect 36760 94570 36840 94580
rect 36940 94570 37020 94580
rect 36120 94490 36130 94570
rect 36300 94490 36310 94570
rect 36480 94490 36490 94570
rect 36660 94490 36670 94570
rect 36840 94490 36850 94570
rect 37020 94490 37030 94570
rect 36040 94250 36120 94260
rect 36220 94250 36300 94260
rect 36400 94250 36480 94260
rect 36580 94250 36660 94260
rect 36760 94250 36840 94260
rect 36940 94250 37020 94260
rect 36120 94170 36130 94250
rect 36300 94170 36310 94250
rect 36480 94170 36490 94250
rect 36660 94170 36670 94250
rect 36840 94170 36850 94250
rect 37020 94170 37030 94250
rect 37100 94080 37190 94750
rect 37600 94740 37660 94770
rect 37720 94740 37780 94770
rect 37840 94740 37900 94770
rect 40060 94690 40120 94720
rect 41540 94690 41600 94720
rect 42360 94690 42420 94720
rect 43840 94690 43900 94720
rect 37720 94650 37750 94680
rect 37840 94650 37870 94680
rect 146100 94650 146160 94680
rect 37600 94620 37660 94650
rect 37720 94620 37780 94650
rect 37840 94620 37900 94650
rect 40060 94570 40120 94600
rect 41540 94570 41600 94600
rect 42360 94570 42420 94600
rect 43840 94570 43900 94600
rect 37720 94530 37750 94560
rect 37840 94530 37870 94560
rect 146100 94530 146160 94560
rect 37600 94500 37660 94530
rect 37720 94500 37780 94530
rect 37840 94500 37900 94530
rect 40678 94504 40758 94514
rect 40838 94504 40918 94514
rect 40060 94450 40120 94480
rect 37720 94410 37750 94440
rect 37840 94410 37870 94440
rect 40758 94434 40768 94504
rect 40678 94424 40768 94434
rect 40838 94434 40848 94504
rect 40918 94434 40928 94504
rect 41540 94450 41600 94480
rect 42360 94450 42420 94480
rect 43840 94450 43900 94480
rect 40838 94424 40928 94434
rect 146100 94410 146160 94440
rect 37600 94380 37660 94410
rect 37720 94380 37780 94410
rect 37840 94380 37900 94410
rect 40060 94330 40120 94360
rect 40678 94344 40758 94354
rect 40838 94344 40918 94354
rect 37720 94290 37750 94320
rect 37840 94290 37870 94320
rect 37600 94260 37660 94290
rect 37720 94260 37780 94290
rect 37840 94260 37900 94290
rect 40758 94264 40768 94344
rect 40838 94264 40848 94344
rect 40918 94264 40928 94344
rect 41540 94330 41600 94360
rect 42360 94330 42420 94360
rect 43840 94330 43900 94360
rect 146100 94290 146160 94320
rect 40060 94210 40120 94240
rect 41540 94210 41600 94240
rect 42360 94210 42420 94240
rect 43840 94210 43900 94240
rect 37720 94170 37750 94200
rect 37840 94170 37870 94200
rect 146100 94170 146160 94200
rect 37600 94140 37660 94170
rect 37720 94140 37780 94170
rect 37840 94140 37900 94170
rect 40060 94090 40120 94120
rect 41540 94090 41600 94120
rect 42360 94090 42420 94120
rect 43840 94090 43900 94120
rect 36000 94070 37190 94080
rect 37100 93970 37190 94070
rect 37720 94050 37750 94080
rect 37840 94050 37870 94080
rect 146100 94050 146160 94080
rect 37600 94020 37660 94050
rect 37720 94020 37780 94050
rect 37840 94020 37900 94050
rect 40060 93970 40120 94000
rect 41540 93970 41600 94000
rect 42360 93970 42420 94000
rect 43840 93970 43900 94000
rect 36000 93940 37190 93970
rect 36040 93930 36120 93940
rect 36220 93930 36300 93940
rect 36400 93930 36480 93940
rect 36580 93930 36660 93940
rect 36760 93930 36840 93940
rect 36940 93930 37020 93940
rect 36120 93870 36130 93930
rect 36300 93870 36310 93930
rect 36480 93870 36490 93930
rect 36660 93870 36670 93930
rect 36840 93870 36850 93930
rect 37020 93870 37030 93930
rect 37100 93870 37190 93940
rect 37720 93930 37750 93960
rect 37840 93930 37870 93960
rect 146100 93930 146160 93960
rect 37600 93900 37660 93930
rect 37720 93900 37780 93930
rect 37840 93900 37900 93930
rect 36000 93840 37190 93870
rect 40060 93850 40120 93880
rect 41540 93850 41600 93880
rect 42360 93850 42420 93880
rect 43840 93850 43900 93880
rect 36040 93780 36120 93790
rect 36220 93780 36300 93790
rect 36400 93780 36480 93790
rect 36580 93780 36660 93790
rect 36760 93780 36840 93790
rect 36940 93780 37020 93790
rect 36120 93700 36130 93780
rect 36300 93700 36310 93780
rect 36480 93700 36490 93780
rect 36660 93700 36670 93780
rect 36840 93700 36850 93780
rect 37020 93700 37030 93780
rect 37100 93640 37190 93840
rect 37720 93810 37750 93840
rect 37840 93810 37870 93840
rect 146100 93810 146160 93840
rect 37600 93780 37660 93810
rect 37720 93780 37780 93810
rect 37840 93780 37900 93810
rect 40060 93730 40120 93760
rect 41540 93730 41600 93760
rect 42360 93730 42420 93760
rect 43840 93730 43900 93760
rect 37720 93690 37750 93720
rect 37840 93690 37870 93720
rect 146100 93690 146160 93720
rect 37600 93660 37660 93690
rect 37720 93660 37780 93690
rect 37840 93660 37900 93690
rect 36000 93610 37190 93640
rect 40060 93610 40120 93640
rect 41540 93610 41600 93640
rect 42360 93610 42420 93640
rect 43840 93610 43900 93640
rect 36120 93550 36130 93610
rect 36300 93550 36310 93610
rect 36480 93550 36490 93610
rect 36660 93550 36670 93610
rect 36840 93550 36850 93610
rect 37020 93550 37030 93610
rect 37100 93540 37190 93610
rect 37720 93570 37750 93600
rect 37840 93570 37870 93600
rect 37600 93540 37660 93570
rect 37720 93540 37780 93570
rect 37840 93540 37900 93570
rect 36000 93510 37190 93540
rect 37100 93500 37190 93510
rect 36000 93490 37190 93500
rect 40060 93490 40120 93520
rect 41540 93490 41600 93520
rect 42360 93490 42420 93520
rect 43840 93490 43900 93520
rect 36040 93310 36120 93320
rect 36220 93310 36300 93320
rect 36400 93310 36480 93320
rect 36580 93310 36660 93320
rect 36760 93310 36840 93320
rect 36940 93310 37020 93320
rect 36120 93230 36130 93310
rect 36300 93230 36310 93310
rect 36480 93230 36490 93310
rect 36660 93230 36670 93310
rect 36840 93230 36850 93310
rect 37020 93230 37030 93310
rect 36040 92990 36120 93000
rect 36220 92990 36300 93000
rect 36400 92990 36480 93000
rect 36580 92990 36660 93000
rect 36760 92990 36840 93000
rect 36940 92990 37020 93000
rect 36120 92910 36130 92990
rect 36300 92910 36310 92990
rect 36480 92910 36490 92990
rect 36660 92910 36670 92990
rect 36840 92910 36850 92990
rect 37020 92910 37030 92990
rect 37100 92820 37190 93490
rect 37720 93450 37750 93480
rect 37840 93450 37870 93480
rect 42595 93475 42675 93485
rect 37600 93420 37660 93450
rect 37720 93420 37780 93450
rect 37840 93420 37900 93450
rect 42675 93405 42685 93475
rect 46660 93460 47160 93640
rect 146100 93570 146160 93600
rect 146100 93450 146160 93480
rect 40060 93370 40120 93400
rect 41540 93370 41600 93400
rect 42360 93370 42420 93400
rect 42595 93395 42685 93405
rect 43840 93370 43900 93400
rect 37720 93330 37750 93360
rect 37840 93330 37870 93360
rect 37600 93300 37660 93330
rect 37720 93300 37780 93330
rect 37840 93300 37900 93330
rect 42595 93315 42675 93325
rect 40060 93250 40120 93280
rect 41540 93250 41600 93280
rect 42360 93250 42420 93280
rect 37720 93210 37750 93240
rect 37840 93210 37870 93240
rect 42675 93235 42685 93315
rect 43030 93300 43390 93360
rect 146100 93330 146160 93360
rect 43840 93250 43900 93280
rect 38595 93215 38675 93225
rect 38775 93215 38855 93225
rect 38955 93215 39035 93225
rect 39135 93215 39215 93225
rect 39315 93215 39395 93225
rect 37600 93180 37660 93210
rect 37720 93180 37780 93210
rect 37840 93180 37900 93210
rect 38675 93135 38685 93215
rect 38855 93135 38865 93215
rect 39035 93135 39045 93215
rect 39215 93135 39225 93215
rect 39395 93135 39405 93215
rect 43580 93170 43700 93230
rect 146100 93210 146160 93240
rect 40060 93130 40120 93160
rect 41540 93130 41600 93160
rect 42360 93130 42420 93160
rect 42950 93150 43560 93160
rect 43550 93145 43560 93150
rect 42910 93135 43560 93145
rect 37720 93090 37750 93120
rect 37840 93090 37870 93120
rect 37600 93060 37660 93090
rect 37720 93060 37780 93090
rect 37840 93060 37900 93090
rect 42900 93085 42910 93135
rect 38595 93035 38675 93045
rect 38775 93035 38855 93045
rect 38955 93035 39035 93045
rect 39135 93035 39215 93045
rect 39315 93035 39395 93045
rect 43030 93040 43390 93100
rect 37720 92970 37750 93000
rect 37840 92970 37870 93000
rect 37600 92940 37660 92970
rect 37720 92940 37780 92970
rect 37840 92940 37900 92970
rect 38675 92955 38685 93035
rect 38855 92955 38865 93035
rect 39035 92955 39045 93035
rect 39215 92955 39225 93035
rect 39395 92955 39405 93035
rect 40060 93010 40120 93040
rect 41540 93010 41600 93040
rect 42360 93010 42420 93040
rect 42682 92960 42822 93030
rect 40060 92890 40120 92920
rect 40678 92899 40758 92909
rect 40838 92899 40918 92909
rect 37720 92850 37750 92880
rect 37840 92850 37870 92880
rect 38595 92855 38675 92865
rect 38775 92855 38855 92865
rect 38955 92855 39035 92865
rect 39135 92855 39215 92865
rect 39315 92855 39395 92865
rect 37600 92820 37660 92850
rect 37720 92820 37780 92850
rect 37840 92820 37900 92850
rect 36000 92810 37190 92820
rect 37100 92710 37190 92810
rect 38675 92775 38685 92855
rect 38855 92775 38865 92855
rect 39035 92775 39045 92855
rect 39215 92775 39225 92855
rect 39395 92775 39405 92855
rect 40758 92819 40768 92899
rect 40838 92819 40848 92899
rect 40918 92819 40928 92899
rect 41540 92890 41600 92920
rect 42360 92890 42420 92920
rect 42822 92900 42892 92960
rect 42822 92890 43470 92900
rect 43550 92890 43560 93135
rect 43700 93050 43760 93170
rect 43840 93130 43900 93160
rect 146100 93090 146160 93120
rect 43840 93010 43900 93040
rect 146100 92970 146160 93000
rect 43580 92910 43700 92970
rect 42822 92820 42892 92890
rect 42910 92875 43560 92885
rect 42900 92825 42910 92875
rect 40060 92770 40120 92800
rect 37720 92730 37750 92760
rect 37840 92730 37870 92760
rect 40685 92750 40925 92780
rect 41540 92770 41600 92800
rect 42360 92770 42420 92800
rect 42682 92760 42822 92820
rect 43030 92780 43390 92840
rect 43700 92790 43760 92910
rect 43840 92890 43900 92920
rect 146100 92850 146160 92880
rect 43840 92770 43900 92800
rect 36000 92680 37190 92710
rect 37600 92700 37660 92730
rect 37720 92700 37780 92730
rect 37840 92700 37900 92730
rect 40685 92690 40715 92750
rect 40775 92690 40865 92750
rect 40895 92690 40925 92750
rect 36040 92670 36120 92680
rect 36220 92670 36300 92680
rect 36400 92670 36480 92680
rect 36580 92670 36660 92680
rect 36760 92670 36840 92680
rect 36940 92670 37020 92680
rect 36120 92610 36130 92670
rect 36300 92610 36310 92670
rect 36480 92610 36490 92670
rect 36660 92610 36670 92670
rect 36840 92610 36850 92670
rect 37020 92610 37030 92670
rect 37100 92610 37190 92680
rect 38595 92675 38675 92685
rect 38775 92675 38855 92685
rect 38955 92675 39035 92685
rect 39135 92675 39215 92685
rect 39315 92675 39395 92685
rect 37720 92610 37750 92640
rect 37840 92610 37870 92640
rect 36000 92580 37190 92610
rect 37600 92580 37660 92610
rect 37720 92580 37780 92610
rect 37840 92580 37900 92610
rect 38675 92595 38685 92675
rect 38855 92595 38865 92675
rect 39035 92595 39045 92675
rect 39215 92595 39225 92675
rect 39395 92595 39405 92675
rect 40060 92650 40120 92680
rect 40685 92660 40925 92690
rect 41540 92650 41600 92680
rect 42360 92650 42420 92680
rect 40678 92629 40758 92639
rect 40838 92629 40918 92639
rect 36040 92520 36120 92530
rect 36220 92520 36300 92530
rect 36400 92520 36480 92530
rect 36580 92520 36660 92530
rect 36760 92520 36840 92530
rect 36940 92520 37020 92530
rect 36120 92440 36130 92520
rect 36300 92440 36310 92520
rect 36480 92440 36490 92520
rect 36660 92440 36670 92520
rect 36840 92440 36850 92520
rect 37020 92440 37030 92520
rect 37100 92380 37190 92580
rect 40060 92530 40120 92560
rect 40758 92549 40768 92629
rect 40838 92549 40848 92629
rect 40918 92549 40928 92629
rect 42822 92620 42892 92760
rect 146100 92730 146160 92760
rect 43580 92650 43700 92710
rect 43840 92650 43900 92680
rect 42950 92630 43560 92640
rect 43550 92625 43560 92630
rect 42682 92560 42822 92620
rect 42910 92615 43560 92625
rect 42900 92565 42910 92615
rect 41540 92530 41600 92560
rect 42360 92530 42420 92560
rect 37720 92490 37750 92520
rect 37840 92490 37870 92520
rect 38595 92495 38675 92505
rect 38775 92495 38855 92505
rect 38955 92495 39035 92505
rect 39135 92495 39215 92505
rect 39315 92495 39395 92505
rect 37600 92460 37660 92490
rect 37720 92460 37780 92490
rect 37840 92460 37900 92490
rect 38675 92415 38685 92495
rect 38855 92415 38865 92495
rect 39035 92415 39045 92495
rect 39215 92415 39225 92495
rect 39395 92415 39405 92495
rect 40060 92410 40120 92440
rect 41540 92410 41600 92440
rect 42360 92410 42420 92440
rect 42822 92420 42892 92560
rect 43030 92520 43390 92580
rect 36000 92350 37190 92380
rect 37720 92370 37750 92400
rect 37840 92370 37870 92400
rect 36120 92290 36130 92350
rect 36300 92290 36310 92350
rect 36480 92290 36490 92350
rect 36660 92290 36670 92350
rect 36840 92290 36850 92350
rect 37020 92290 37030 92350
rect 37100 92280 37190 92350
rect 37600 92340 37660 92370
rect 37720 92340 37780 92370
rect 37840 92340 37900 92370
rect 40170 92320 40180 92410
rect 40060 92290 40120 92320
rect 36000 92250 37190 92280
rect 37720 92250 37750 92280
rect 37840 92250 37870 92280
rect 37100 92240 37190 92250
rect 36000 92230 37190 92240
rect 36040 92050 36120 92060
rect 36220 92050 36300 92060
rect 36400 92050 36480 92060
rect 36580 92050 36660 92060
rect 36760 92050 36840 92060
rect 36940 92050 37020 92060
rect 36120 91970 36130 92050
rect 36300 91970 36310 92050
rect 36480 91970 36490 92050
rect 36660 91970 36670 92050
rect 36840 91970 36850 92050
rect 37020 91970 37030 92050
rect 36040 91730 36120 91740
rect 36220 91730 36300 91740
rect 36400 91730 36480 91740
rect 36580 91730 36660 91740
rect 36760 91730 36840 91740
rect 36940 91730 37020 91740
rect 36120 91650 36130 91730
rect 36300 91650 36310 91730
rect 36480 91650 36490 91730
rect 36660 91650 36670 91730
rect 36840 91650 36850 91730
rect 37020 91650 37030 91730
rect 37100 91560 37190 92230
rect 37600 92220 37660 92250
rect 37720 92220 37780 92250
rect 37840 92220 37900 92250
rect 40060 92170 40120 92200
rect 37720 92130 37750 92160
rect 37840 92130 37870 92160
rect 37600 92100 37660 92130
rect 37720 92100 37780 92130
rect 37840 92100 37900 92130
rect 40060 92050 40120 92080
rect 37720 92010 37750 92040
rect 37840 92010 37870 92040
rect 37600 91980 37660 92010
rect 37720 91980 37780 92010
rect 37840 91980 37900 92010
rect 40060 91930 40120 91960
rect 37720 91890 37750 91920
rect 37840 91890 37870 91920
rect 37600 91860 37660 91890
rect 37720 91860 37780 91890
rect 37840 91860 37900 91890
rect 40060 91810 40120 91840
rect 37720 91770 37750 91800
rect 37840 91770 37870 91800
rect 37600 91740 37660 91770
rect 37720 91740 37780 91770
rect 37840 91740 37900 91770
rect 40060 91690 40120 91720
rect 37720 91650 37750 91680
rect 37840 91650 37870 91680
rect 37600 91620 37660 91650
rect 37720 91620 37780 91650
rect 37840 91620 37900 91650
rect 40060 91570 40120 91600
rect 36000 91550 37190 91560
rect 37100 91450 37190 91550
rect 37720 91530 37750 91560
rect 37840 91530 37870 91560
rect 40260 91530 40270 92320
rect 40380 92310 41180 92400
rect 40650 92280 40770 92310
rect 40930 92280 41050 92310
rect 41090 92280 41180 92310
rect 40650 92190 40660 92280
rect 40760 92250 40830 92280
rect 40770 92160 40830 92250
rect 40930 92190 40940 92280
rect 41050 92160 41180 92280
rect 41260 92240 41340 92250
rect 41340 92190 41350 92240
rect 41090 92125 41180 92160
rect 41230 92130 41350 92190
rect 40470 92120 41180 92125
rect 40370 92110 41180 92120
rect 40370 92030 40380 92110
rect 40470 92105 41180 92110
rect 40420 92095 41210 92105
rect 41090 92045 41180 92095
rect 40470 92030 41180 92045
rect 40460 92015 41180 92030
rect 40460 91825 40470 92015
rect 40650 91980 40770 92015
rect 40930 91980 41050 92015
rect 41090 91980 41180 92015
rect 41350 92010 41410 92130
rect 40770 91970 40830 91980
rect 40530 91960 40610 91970
rect 40670 91960 40750 91970
rect 40770 91960 40890 91970
rect 40950 91960 41030 91970
rect 40610 91880 40620 91960
rect 40750 91880 40760 91960
rect 40770 91860 40830 91960
rect 40890 91880 40900 91960
rect 41030 91880 41040 91960
rect 41050 91860 41180 91980
rect 41260 91960 41340 91970
rect 41340 91890 41350 91960
rect 41090 91825 41180 91860
rect 41230 91830 41350 91890
rect 40460 91810 41180 91825
rect 40470 91805 41180 91810
rect 40420 91795 41210 91805
rect 41090 91745 41180 91795
rect 40470 91715 41180 91745
rect 40650 91680 40770 91715
rect 40930 91680 41050 91715
rect 41090 91680 41180 91715
rect 41350 91710 41410 91830
rect 41480 91680 41490 92390
rect 42860 92370 43470 92380
rect 43550 92370 43560 92615
rect 43700 92530 43760 92650
rect 146100 92610 146160 92640
rect 43840 92530 43900 92560
rect 146100 92490 146160 92520
rect 43580 92390 43700 92450
rect 43840 92410 43900 92440
rect 42910 92355 43560 92365
rect 41540 92290 41600 92320
rect 42360 92290 42420 92320
rect 42900 92305 42910 92355
rect 43030 92260 43390 92320
rect 43700 92270 43760 92390
rect 146100 92370 146160 92400
rect 43840 92290 43900 92320
rect 146100 92250 146160 92280
rect 41540 92170 41600 92200
rect 42360 92170 42420 92200
rect 42470 92160 42480 92250
rect 43840 92170 43900 92200
rect 41540 92050 41600 92080
rect 42360 92050 42420 92080
rect 41540 91930 41600 91960
rect 42360 91930 42420 91960
rect 41540 91810 41600 91840
rect 42360 91810 42420 91840
rect 41540 91690 41600 91720
rect 42360 91690 42420 91720
rect 42560 91680 42570 92160
rect 146100 92130 146160 92160
rect 42960 92120 43460 92130
rect 42620 92100 42700 92110
rect 42700 92030 42710 92100
rect 42620 92020 42710 92030
rect 42770 92020 42780 92110
rect 43840 92050 43900 92080
rect 42620 91940 42700 91950
rect 42700 91890 42710 91940
rect 42610 91830 42730 91890
rect 42730 91805 42790 91830
rect 42860 91820 42870 92020
rect 42910 91980 43030 92040
rect 43190 91980 43310 92040
rect 146100 92010 146160 92040
rect 43030 91970 43090 91980
rect 43310 91970 43370 91980
rect 42930 91960 43010 91970
rect 43030 91960 43150 91970
rect 43210 91960 43290 91970
rect 43310 91960 43430 91970
rect 43010 91880 43020 91960
rect 43030 91860 43090 91960
rect 43150 91880 43160 91960
rect 43290 91880 43300 91960
rect 43310 91860 43370 91960
rect 43430 91880 43440 91960
rect 43840 91930 43900 91960
rect 146100 91890 146160 91920
rect 42860 91810 43500 91820
rect 43840 91810 43900 91840
rect 42730 91795 43540 91805
rect 42730 91710 42790 91795
rect 43540 91745 43550 91795
rect 146100 91770 146160 91800
rect 42860 91680 42870 91730
rect 42910 91680 43030 91740
rect 43190 91680 43310 91740
rect 43840 91690 43900 91720
rect 40770 91670 40830 91680
rect 40530 91660 40610 91670
rect 40770 91660 40890 91670
rect 40610 91580 40620 91660
rect 40770 91560 40830 91660
rect 40890 91580 40900 91660
rect 41050 91560 41180 91680
rect 43030 91670 43090 91680
rect 43310 91670 43370 91680
rect 43030 91660 43150 91670
rect 43310 91660 43430 91670
rect 41540 91570 41600 91600
rect 42360 91570 42420 91600
rect 43030 91560 43090 91660
rect 43150 91580 43160 91660
rect 43310 91560 43370 91660
rect 43430 91580 43440 91660
rect 146100 91650 146160 91680
rect 43840 91570 43900 91600
rect 41090 91550 41180 91560
rect 40470 91530 41180 91550
rect 146100 91530 146160 91560
rect 37600 91500 37660 91530
rect 37720 91500 37780 91530
rect 37840 91500 37900 91530
rect 40060 91450 40120 91480
rect 36000 91420 37190 91450
rect 40170 91440 40180 91530
rect 40260 91520 41100 91530
rect 36040 91410 36120 91420
rect 36220 91410 36300 91420
rect 36400 91410 36480 91420
rect 36580 91410 36660 91420
rect 36760 91410 36840 91420
rect 36940 91410 37020 91420
rect 36120 91350 36130 91410
rect 36300 91350 36310 91410
rect 36480 91350 36490 91410
rect 36660 91350 36670 91410
rect 36840 91350 36850 91410
rect 37020 91350 37030 91410
rect 37100 91350 37190 91420
rect 37720 91410 37750 91440
rect 37840 91410 37870 91440
rect 37600 91380 37660 91410
rect 37720 91380 37780 91410
rect 37840 91380 37900 91410
rect 36000 91320 37190 91350
rect 40060 91330 40120 91360
rect 36040 91260 36120 91270
rect 36220 91260 36300 91270
rect 36400 91260 36480 91270
rect 36580 91260 36660 91270
rect 36760 91260 36840 91270
rect 36940 91260 37020 91270
rect 36120 91180 36130 91260
rect 36300 91180 36310 91260
rect 36480 91180 36490 91260
rect 36660 91180 36670 91260
rect 36840 91180 36850 91260
rect 37020 91180 37030 91260
rect 37100 91120 37190 91320
rect 37720 91290 37750 91320
rect 37840 91290 37870 91320
rect 37600 91260 37660 91290
rect 37720 91260 37780 91290
rect 37840 91260 37900 91290
rect 40060 91210 40120 91240
rect 37720 91170 37750 91200
rect 37840 91170 37870 91200
rect 37600 91140 37660 91170
rect 37720 91140 37780 91170
rect 37840 91140 37900 91170
rect 36000 91090 37190 91120
rect 40060 91090 40120 91120
rect 36120 91030 36130 91090
rect 36300 91030 36310 91090
rect 36480 91030 36490 91090
rect 36660 91030 36670 91090
rect 36840 91030 36850 91090
rect 37020 91030 37030 91090
rect 37100 91020 37190 91090
rect 37720 91050 37750 91080
rect 37840 91050 37870 91080
rect 37600 91020 37660 91050
rect 37720 91020 37780 91050
rect 37840 91020 37900 91050
rect 36000 90990 37190 91020
rect 37100 90980 37190 90990
rect 36000 90970 37190 90980
rect 40060 90970 40120 91000
rect 36040 90790 36120 90800
rect 36220 90790 36300 90800
rect 36400 90790 36480 90800
rect 36580 90790 36660 90800
rect 36760 90790 36840 90800
rect 36940 90790 37020 90800
rect 36120 90710 36130 90790
rect 36300 90710 36310 90790
rect 36480 90710 36490 90790
rect 36660 90710 36670 90790
rect 36840 90710 36850 90790
rect 37020 90710 37030 90790
rect 36040 90470 36120 90480
rect 36220 90470 36300 90480
rect 36400 90470 36480 90480
rect 36580 90470 36660 90480
rect 36760 90470 36840 90480
rect 36940 90470 37020 90480
rect 36120 90390 36130 90470
rect 36300 90390 36310 90470
rect 36480 90390 36490 90470
rect 36660 90390 36670 90470
rect 36840 90390 36850 90470
rect 37020 90390 37030 90470
rect 37100 90300 37190 90970
rect 37720 90930 37750 90960
rect 37840 90930 37870 90960
rect 37600 90900 37660 90930
rect 37720 90900 37780 90930
rect 37840 90900 37900 90930
rect 40060 90850 40120 90880
rect 37720 90810 37750 90840
rect 37840 90810 37870 90840
rect 37600 90780 37660 90810
rect 37720 90780 37780 90810
rect 37840 90780 37900 90810
rect 40060 90730 40120 90760
rect 37720 90690 37750 90720
rect 37840 90690 37870 90720
rect 37600 90660 37660 90690
rect 37720 90660 37780 90690
rect 37840 90660 37900 90690
rect 40060 90610 40120 90640
rect 37720 90570 37750 90600
rect 37840 90570 37870 90600
rect 37600 90540 37660 90570
rect 37720 90540 37780 90570
rect 37840 90540 37900 90570
rect 40060 90490 40120 90520
rect 37720 90450 37750 90480
rect 37840 90450 37870 90480
rect 37600 90420 37660 90450
rect 37720 90420 37780 90450
rect 37840 90420 37900 90450
rect 40060 90370 40120 90400
rect 37720 90330 37750 90360
rect 37840 90330 37870 90360
rect 37600 90300 37660 90330
rect 37720 90300 37780 90330
rect 37840 90300 37900 90330
rect 36000 90290 37190 90300
rect 37100 90190 37190 90290
rect 40060 90250 40120 90280
rect 37720 90210 37750 90240
rect 37840 90210 37870 90240
rect 36000 90160 37190 90190
rect 37600 90180 37660 90210
rect 37720 90180 37780 90210
rect 37840 90180 37900 90210
rect 36040 90150 36120 90160
rect 36220 90150 36300 90160
rect 36400 90150 36480 90160
rect 36580 90150 36660 90160
rect 36760 90150 36840 90160
rect 36940 90150 37020 90160
rect 36120 90090 36130 90150
rect 36300 90090 36310 90150
rect 36480 90090 36490 90150
rect 36660 90090 36670 90150
rect 36840 90090 36850 90150
rect 37020 90090 37030 90150
rect 37100 90090 37190 90160
rect 40060 90130 40120 90160
rect 37720 90090 37750 90120
rect 37840 90090 37870 90120
rect 36000 90060 37190 90090
rect 37600 90060 37660 90090
rect 37720 90060 37780 90090
rect 37840 90060 37900 90090
rect 36040 90000 36120 90010
rect 36220 90000 36300 90010
rect 36400 90000 36480 90010
rect 36580 90000 36660 90010
rect 36760 90000 36840 90010
rect 36940 90000 37020 90010
rect 36120 89920 36130 90000
rect 36300 89920 36310 90000
rect 36480 89920 36490 90000
rect 36660 89920 36670 90000
rect 36840 89920 36850 90000
rect 37020 89920 37030 90000
rect 36040 89850 36120 89860
rect 36220 89850 36300 89860
rect 36400 89850 36480 89860
rect 36580 89850 36660 89860
rect 36760 89850 36840 89860
rect 36940 89850 37020 89860
rect 36120 89770 36130 89850
rect 36300 89770 36310 89850
rect 36480 89770 36490 89850
rect 36660 89770 36670 89850
rect 36840 89770 36850 89850
rect 37020 89770 37030 89850
rect 37100 89830 37190 90060
rect 40060 90010 40120 90040
rect 37720 89970 37750 90000
rect 37840 89970 37870 90000
rect 37600 89940 37660 89970
rect 37720 89940 37780 89970
rect 37840 89940 37900 89970
rect 40060 89890 40120 89920
rect 37720 89850 37750 89880
rect 37840 89850 37870 89880
rect 37600 89820 37660 89850
rect 37720 89820 37780 89850
rect 37840 89820 37900 89850
rect 40060 89770 40120 89800
rect 19130 89700 19160 89755
rect 19250 89700 19280 89755
rect 26420 89700 26450 89755
rect 26540 89700 26570 89755
rect 30420 89730 30450 89755
rect 30540 89730 30570 89755
rect 37720 89730 37750 89760
rect 37840 89730 37870 89760
rect 30300 89700 30360 89730
rect 30420 89700 30480 89730
rect 30540 89700 30600 89730
rect 37600 89700 37660 89730
rect 37720 89700 37780 89730
rect 37840 89700 37900 89730
rect 40060 89650 40120 89680
rect 30420 89580 30450 89640
rect 30540 89580 30570 89640
rect 37720 89580 37750 89640
rect 37840 89580 37870 89640
rect 40060 89530 40120 89560
rect 18980 89440 19060 89450
rect 19160 89440 19240 89450
rect 19340 89440 19420 89450
rect 19520 89440 19600 89450
rect 19700 89440 19780 89450
rect 19880 89440 19960 89450
rect 20060 89440 20140 89450
rect 20240 89440 20320 89450
rect 20420 89440 20500 89450
rect 20600 89440 20680 89450
rect 20780 89440 20860 89450
rect 20960 89440 21040 89450
rect 21140 89440 21220 89450
rect 21320 89440 21400 89450
rect 21500 89440 21580 89450
rect 21680 89440 21760 89450
rect 21860 89440 21940 89450
rect 22040 89440 22120 89450
rect 22220 89440 22300 89450
rect 22400 89440 22480 89450
rect 22580 89440 22660 89450
rect 22760 89440 22840 89450
rect 22940 89440 23020 89450
rect 23120 89440 23200 89450
rect 23300 89440 23380 89450
rect 23480 89440 23560 89450
rect 23660 89440 23740 89450
rect 23840 89440 23920 89450
rect 24020 89440 24100 89450
rect 24200 89440 24280 89450
rect 24380 89440 24460 89450
rect 24560 89440 24640 89450
rect 24740 89440 24820 89450
rect 24920 89440 25000 89450
rect 25100 89440 25180 89450
rect 25280 89440 25360 89450
rect 25460 89440 25540 89450
rect 25640 89440 25720 89450
rect 25820 89440 25900 89450
rect 26000 89440 26080 89450
rect 26180 89440 26260 89450
rect 26360 89440 26440 89450
rect 26540 89440 26620 89450
rect 30280 89440 30360 89450
rect 30460 89440 30540 89450
rect 30640 89440 30720 89450
rect 30820 89440 30900 89450
rect 31000 89440 31080 89450
rect 31180 89440 31260 89450
rect 31360 89440 31440 89450
rect 31540 89440 31620 89450
rect 31720 89440 31800 89450
rect 31900 89440 31980 89450
rect 32080 89440 32160 89450
rect 32260 89440 32340 89450
rect 32440 89440 32520 89450
rect 32620 89440 32700 89450
rect 32800 89440 32880 89450
rect 32980 89440 33060 89450
rect 33160 89440 33240 89450
rect 33340 89440 33420 89450
rect 33520 89440 33600 89450
rect 33700 89440 33780 89450
rect 33880 89440 33960 89450
rect 34060 89440 34140 89450
rect 34240 89440 34320 89450
rect 34420 89440 34500 89450
rect 34600 89440 34680 89450
rect 34780 89440 34860 89450
rect 34960 89440 35040 89450
rect 35140 89440 35220 89450
rect 35320 89440 35400 89450
rect 35500 89440 35580 89450
rect 35680 89440 35760 89450
rect 35860 89440 35940 89450
rect 36040 89440 36120 89450
rect 36220 89440 36300 89450
rect 36400 89440 36480 89450
rect 36580 89440 36660 89450
rect 36760 89440 36840 89450
rect 36940 89440 37020 89450
rect 37120 89440 37200 89450
rect 37300 89440 37380 89450
rect 37480 89440 37560 89450
rect 37660 89440 37740 89450
rect 37840 89440 37920 89450
rect 40260 89440 40270 91440
rect 40380 91430 41180 91520
rect 41540 91450 41600 91480
rect 42360 91450 42420 91480
rect 43840 91450 43900 91480
rect 40650 91400 40770 91430
rect 40930 91400 41050 91430
rect 41090 91400 41180 91430
rect 146100 91410 146160 91440
rect 40650 91310 40660 91400
rect 40760 91370 40830 91400
rect 40770 91280 40830 91370
rect 40930 91310 40940 91400
rect 41050 91280 41180 91400
rect 41090 91245 41180 91280
rect 41230 91250 41350 91310
rect 40470 91240 41180 91245
rect 40370 91230 41180 91240
rect 40370 91150 40380 91230
rect 40470 91225 41180 91230
rect 40420 91215 41210 91225
rect 41090 91165 41180 91215
rect 40470 91150 41180 91165
rect 40460 91135 41180 91150
rect 40460 90945 40470 91135
rect 40650 91100 40770 91135
rect 40930 91100 41050 91135
rect 41090 91100 41180 91135
rect 41350 91130 41410 91250
rect 40770 91090 40830 91100
rect 40530 91080 40610 91090
rect 40670 91080 40750 91090
rect 40770 91080 40890 91090
rect 40950 91080 41030 91090
rect 40610 91000 40620 91080
rect 40750 91000 40760 91080
rect 40770 90980 40830 91080
rect 40890 91000 40900 91080
rect 41030 91000 41040 91080
rect 41050 90980 41180 91100
rect 41260 91080 41340 91090
rect 41340 91010 41350 91080
rect 41090 90945 41180 90980
rect 41230 90950 41350 91010
rect 40460 90930 41180 90945
rect 40470 90925 41180 90930
rect 40420 90915 41210 90925
rect 41090 90865 41180 90915
rect 40470 90835 41180 90865
rect 40650 90800 40770 90835
rect 40930 90800 41050 90835
rect 41090 90800 41180 90835
rect 41350 90830 41410 90950
rect 40650 90710 40660 90800
rect 40760 90770 40830 90800
rect 40770 90680 40830 90770
rect 40930 90710 40940 90800
rect 41050 90680 41180 90800
rect 41260 90780 41340 90790
rect 41340 90710 41350 90780
rect 41090 90645 41180 90680
rect 41230 90650 41350 90710
rect 40370 90630 40460 90640
rect 40370 90550 40380 90630
rect 40470 90625 41180 90645
rect 40420 90615 41210 90625
rect 41090 90565 41180 90615
rect 40470 90550 41180 90565
rect 40460 90535 41180 90550
rect 40460 90345 40470 90535
rect 40650 90500 40770 90535
rect 40930 90500 41050 90535
rect 41090 90500 41180 90535
rect 41350 90530 41410 90650
rect 40770 90490 40830 90500
rect 40530 90480 40610 90490
rect 40670 90480 40750 90490
rect 40770 90480 40890 90490
rect 40950 90480 41030 90490
rect 40610 90400 40620 90480
rect 40750 90400 40760 90480
rect 40770 90380 40830 90480
rect 40890 90400 40900 90480
rect 41030 90400 41040 90480
rect 41050 90380 41180 90500
rect 41260 90480 41340 90490
rect 41340 90410 41350 90480
rect 41090 90345 41180 90380
rect 41230 90350 41350 90410
rect 40460 90330 41180 90345
rect 40470 90325 41180 90330
rect 40420 90315 41210 90325
rect 41090 90265 41180 90315
rect 40470 90235 41180 90265
rect 40650 90200 40770 90235
rect 40930 90200 41050 90235
rect 41090 90200 41180 90235
rect 41350 90230 41410 90350
rect 40650 90110 40660 90200
rect 40760 90170 40830 90200
rect 40770 90080 40830 90170
rect 40930 90110 40940 90200
rect 41050 90080 41180 90200
rect 41260 90180 41340 90190
rect 41340 90110 41350 90180
rect 41090 90045 41180 90080
rect 41230 90050 41350 90110
rect 40370 90030 40460 90040
rect 40370 89950 40380 90030
rect 40470 90025 41180 90045
rect 40420 90015 41210 90025
rect 41090 89965 41180 90015
rect 40470 89950 41180 89965
rect 40460 89935 41180 89950
rect 40460 89745 40470 89935
rect 40650 89900 40770 89935
rect 40930 89900 41050 89935
rect 41090 89900 41180 89935
rect 41350 89930 41410 90050
rect 40770 89890 40830 89900
rect 40530 89880 40610 89890
rect 40670 89880 40750 89890
rect 40770 89880 40890 89890
rect 40950 89880 41030 89890
rect 40610 89800 40620 89880
rect 40750 89800 40760 89880
rect 40770 89780 40830 89880
rect 40890 89800 40900 89880
rect 41030 89800 41040 89880
rect 41050 89780 41180 89900
rect 41260 89870 41340 89880
rect 41340 89810 41350 89870
rect 41090 89745 41180 89780
rect 41230 89750 41350 89810
rect 40460 89730 41180 89745
rect 40470 89725 41180 89730
rect 40420 89715 41210 89725
rect 41090 89665 41180 89715
rect 40470 89635 41180 89665
rect 40650 89600 40770 89635
rect 40930 89600 41050 89635
rect 41090 89600 41180 89635
rect 41350 89630 41410 89750
rect 41480 89600 41490 91370
rect 41540 91330 41600 91360
rect 42360 91330 42420 91360
rect 43840 91330 43900 91360
rect 146100 91290 146160 91320
rect 41540 91210 41600 91240
rect 42360 91210 42420 91240
rect 43840 91210 43900 91240
rect 146100 91170 146160 91200
rect 41540 91090 41600 91120
rect 42360 91090 42420 91120
rect 42910 91100 43030 91160
rect 43190 91100 43310 91160
rect 43030 91090 43090 91100
rect 43310 91090 43370 91100
rect 43840 91090 43900 91120
rect 42930 91080 43010 91090
rect 43030 91080 43150 91090
rect 43210 91080 43290 91090
rect 43310 91080 43430 91090
rect 41540 90970 41600 91000
rect 42360 90970 42420 91000
rect 42470 90980 42480 91070
rect 41540 90850 41600 90880
rect 42360 90850 42420 90880
rect 41540 90730 41600 90760
rect 42360 90730 42420 90760
rect 41540 90610 41600 90640
rect 42360 90610 42420 90640
rect 41540 90490 41600 90520
rect 42360 90490 42420 90520
rect 41540 90370 41600 90400
rect 42360 90370 42420 90400
rect 41540 90250 41600 90280
rect 42360 90250 42420 90280
rect 41540 90130 41600 90160
rect 42360 90130 42420 90160
rect 41540 90010 41600 90040
rect 42360 90010 42420 90040
rect 41540 89890 41600 89920
rect 42360 89890 42420 89920
rect 41540 89770 41600 89800
rect 42360 89770 42420 89800
rect 41540 89650 41600 89680
rect 42360 89650 42420 89680
rect 42560 89620 42570 90980
rect 42610 90950 42730 91010
rect 42730 90925 42790 90950
rect 42860 90940 42870 91070
rect 43010 91000 43020 91080
rect 43030 90980 43090 91080
rect 43150 91000 43160 91080
rect 43290 91000 43300 91080
rect 43310 90980 43370 91080
rect 43430 91000 43440 91080
rect 146100 91050 146160 91080
rect 43840 90970 43900 91000
rect 42860 90930 43500 90940
rect 42730 90915 43540 90925
rect 42730 90830 42790 90915
rect 43540 90865 43550 90915
rect 42620 90740 42700 90750
rect 42700 90660 42710 90740
rect 42860 90660 42870 90850
rect 42910 90800 43030 90860
rect 43190 90800 43310 90860
rect 43020 90770 43090 90800
rect 43030 90680 43090 90770
rect 43190 90710 43200 90800
rect 43300 90770 43370 90800
rect 43310 90680 43370 90770
rect 42860 90650 43490 90660
rect 42860 90640 42870 90650
rect 42620 90560 42700 90570
rect 42700 90480 42710 90560
rect 42770 90550 42780 90640
rect 42610 90360 42730 90420
rect 42730 90335 42790 90360
rect 42860 90350 42870 90550
rect 42910 90510 43030 90570
rect 43190 90510 43310 90570
rect 43030 90500 43090 90510
rect 43310 90500 43370 90510
rect 42930 90490 43010 90500
rect 43030 90490 43150 90500
rect 43210 90490 43290 90500
rect 43310 90490 43430 90500
rect 43010 90410 43020 90490
rect 43030 90390 43090 90490
rect 43150 90410 43160 90490
rect 43290 90410 43300 90490
rect 43310 90390 43370 90490
rect 43430 90410 43440 90490
rect 42860 90340 43500 90350
rect 43580 90340 43590 90640
rect 42730 90325 43540 90335
rect 42730 90240 42790 90325
rect 43540 90275 43550 90325
rect 42620 90140 42700 90150
rect 42700 90060 42710 90140
rect 42860 90070 42870 90260
rect 42910 90210 43030 90270
rect 43190 90210 43310 90270
rect 43020 90180 43090 90210
rect 43030 90090 43090 90180
rect 43190 90120 43200 90210
rect 43300 90180 43370 90210
rect 43310 90090 43370 90180
rect 42860 90060 43490 90070
rect 42860 90050 42870 90060
rect 42620 89960 42700 89970
rect 42770 89960 42780 90050
rect 42700 89880 42710 89960
rect 42610 89770 42730 89830
rect 42730 89745 42790 89770
rect 42860 89760 42870 89960
rect 42910 89920 43030 89980
rect 43190 89920 43310 89980
rect 43030 89910 43090 89920
rect 43310 89910 43370 89920
rect 42930 89900 43010 89910
rect 43030 89900 43150 89910
rect 43210 89900 43290 89910
rect 43310 89900 43430 89910
rect 43010 89820 43020 89900
rect 43030 89800 43090 89900
rect 43150 89820 43160 89900
rect 43290 89820 43300 89900
rect 43310 89800 43370 89900
rect 43430 89820 43440 89900
rect 42860 89750 43500 89760
rect 43580 89750 43590 90050
rect 42730 89735 43540 89745
rect 42730 89650 42790 89735
rect 43540 89685 43550 89735
rect 42860 89620 42870 89670
rect 42910 89620 43030 89680
rect 43190 89620 43310 89680
rect 43030 89610 43090 89620
rect 43310 89610 43370 89620
rect 43030 89600 43150 89610
rect 43310 89600 43430 89610
rect 40770 89590 40830 89600
rect 40530 89580 40610 89590
rect 40770 89580 40890 89590
rect 40610 89500 40620 89580
rect 40770 89480 40830 89580
rect 40890 89500 40900 89580
rect 41050 89480 41180 89600
rect 41540 89530 41600 89560
rect 42360 89530 42420 89560
rect 43030 89500 43090 89600
rect 43150 89520 43160 89600
rect 43310 89500 43370 89600
rect 43430 89520 43440 89600
rect 41090 89450 41180 89480
rect 43780 89460 43790 90940
rect 146100 90930 146160 90960
rect 43840 90850 43900 90880
rect 146100 90810 146160 90840
rect 43840 90730 43900 90760
rect 146100 90690 146160 90720
rect 43840 90610 43900 90640
rect 146100 90570 146160 90600
rect 43840 90490 43900 90520
rect 146100 90450 146160 90480
rect 43840 90370 43900 90400
rect 146100 90330 146160 90360
rect 43840 90250 43900 90280
rect 146100 90210 146160 90240
rect 43840 90130 43900 90160
rect 146100 90090 146160 90120
rect 43840 90010 43900 90040
rect 146100 89970 146160 90000
rect 43840 89890 43900 89920
rect 146100 89850 146160 89880
rect 43840 89770 43900 89800
rect 43840 89650 43900 89680
rect 46660 89560 47160 89740
rect 146100 89730 146160 89760
rect 147580 89730 147640 89746
rect 148400 89730 148460 89746
rect 149880 89730 149940 89746
rect 152220 89710 152250 89740
rect 152340 89710 152370 89740
rect 159520 89710 159550 89740
rect 159640 89710 159670 89740
rect 163520 89710 163550 89740
rect 163640 89710 163670 89740
rect 170810 89710 170840 89740
rect 170930 89710 170960 89740
rect 152100 89680 152160 89710
rect 152220 89680 152280 89710
rect 152340 89680 152400 89710
rect 159400 89680 159460 89710
rect 159520 89680 159580 89710
rect 159640 89680 159700 89710
rect 163400 89680 163460 89710
rect 163520 89680 163580 89710
rect 163640 89680 163700 89710
rect 170690 89680 170750 89710
rect 170810 89680 170870 89710
rect 170930 89680 170990 89710
rect 146100 89610 146160 89640
rect 147580 89610 147640 89640
rect 148400 89610 148460 89640
rect 149880 89610 149940 89640
rect 152220 89560 152250 89620
rect 152340 89560 152370 89620
rect 159520 89560 159550 89620
rect 159640 89560 159670 89620
rect 163520 89560 163550 89620
rect 163640 89560 163670 89620
rect 170810 89560 170840 89620
rect 170930 89560 170960 89620
rect 43840 89530 43900 89560
rect 146100 89490 146160 89520
rect 147580 89490 147640 89520
rect 148400 89490 148460 89520
rect 149880 89490 149940 89520
rect 19060 89360 19070 89440
rect 19240 89360 19250 89440
rect 19420 89360 19430 89440
rect 19600 89360 19610 89440
rect 19780 89360 19790 89440
rect 19960 89360 19970 89440
rect 20140 89360 20150 89440
rect 20320 89360 20330 89440
rect 20500 89360 20510 89440
rect 20680 89360 20690 89440
rect 20860 89360 20870 89440
rect 21040 89360 21050 89440
rect 21220 89360 21230 89440
rect 21400 89360 21410 89440
rect 21580 89360 21590 89440
rect 21760 89360 21770 89440
rect 21940 89360 21950 89440
rect 22120 89360 22130 89440
rect 22300 89360 22310 89440
rect 22480 89360 22490 89440
rect 22660 89360 22670 89440
rect 22840 89360 22850 89440
rect 23020 89360 23030 89440
rect 23200 89360 23210 89440
rect 23380 89360 23390 89440
rect 23560 89360 23570 89440
rect 23740 89360 23750 89440
rect 23920 89360 23930 89440
rect 24100 89360 24110 89440
rect 24280 89360 24290 89440
rect 24460 89360 24470 89440
rect 24640 89360 24650 89440
rect 24820 89360 24830 89440
rect 25000 89360 25010 89440
rect 25180 89360 25190 89440
rect 25360 89360 25370 89440
rect 25540 89360 25550 89440
rect 25720 89360 25730 89440
rect 25900 89360 25910 89440
rect 26080 89360 26090 89440
rect 26260 89360 26270 89440
rect 26440 89360 26450 89440
rect 26620 89360 26630 89440
rect 27315 89415 27395 89425
rect 27495 89415 27575 89425
rect 27675 89415 27755 89425
rect 27855 89415 27935 89425
rect 28035 89415 28115 89425
rect 27395 89335 27405 89415
rect 27575 89335 27585 89415
rect 27755 89335 27765 89415
rect 27935 89335 27945 89415
rect 28115 89335 28125 89415
rect 30360 89360 30370 89440
rect 30540 89360 30550 89440
rect 30720 89360 30730 89440
rect 30900 89360 30910 89440
rect 31080 89360 31090 89440
rect 31260 89360 31270 89440
rect 31440 89360 31450 89440
rect 31620 89360 31630 89440
rect 31800 89360 31810 89440
rect 31980 89360 31990 89440
rect 32160 89360 32170 89440
rect 32340 89360 32350 89440
rect 32520 89360 32530 89440
rect 32700 89360 32710 89440
rect 32880 89360 32890 89440
rect 33060 89360 33070 89440
rect 33240 89360 33250 89440
rect 33420 89360 33430 89440
rect 33600 89360 33610 89440
rect 33780 89360 33790 89440
rect 33960 89360 33970 89440
rect 34140 89360 34150 89440
rect 34320 89360 34330 89440
rect 34500 89360 34510 89440
rect 34680 89360 34690 89440
rect 34860 89360 34870 89440
rect 35040 89360 35050 89440
rect 35220 89360 35230 89440
rect 35400 89360 35410 89440
rect 35580 89360 35590 89440
rect 35760 89360 35770 89440
rect 35940 89360 35950 89440
rect 36120 89360 36130 89440
rect 36300 89360 36310 89440
rect 36480 89360 36490 89440
rect 36660 89360 36670 89440
rect 36840 89360 36850 89440
rect 37020 89360 37030 89440
rect 37200 89360 37210 89440
rect 37380 89360 37390 89440
rect 37560 89360 37570 89440
rect 37740 89360 37750 89440
rect 37920 89360 37930 89440
rect 40060 89410 40120 89440
rect 41540 89410 41600 89440
rect 42360 89410 42420 89440
rect 43840 89410 43900 89440
rect 146100 89370 146160 89400
rect 147580 89370 147640 89400
rect 148400 89370 148460 89400
rect 149880 89370 149940 89400
rect 18980 89290 19060 89300
rect 19160 89290 19240 89300
rect 19340 89290 19420 89300
rect 19520 89290 19600 89300
rect 19700 89290 19780 89300
rect 19880 89290 19960 89300
rect 20060 89290 20140 89300
rect 20240 89290 20320 89300
rect 20420 89290 20500 89300
rect 20600 89290 20680 89300
rect 20780 89290 20860 89300
rect 20960 89290 21040 89300
rect 21140 89290 21220 89300
rect 21320 89290 21400 89300
rect 21500 89290 21580 89300
rect 21680 89290 21760 89300
rect 21860 89290 21940 89300
rect 22040 89290 22120 89300
rect 22220 89290 22300 89300
rect 22400 89290 22480 89300
rect 22580 89290 22660 89300
rect 22760 89290 22840 89300
rect 22940 89290 23020 89300
rect 23120 89290 23200 89300
rect 23300 89290 23380 89300
rect 23480 89290 23560 89300
rect 23660 89290 23740 89300
rect 23840 89290 23920 89300
rect 24020 89290 24100 89300
rect 24200 89290 24280 89300
rect 24380 89290 24460 89300
rect 24560 89290 24640 89300
rect 24740 89290 24820 89300
rect 24920 89290 25000 89300
rect 25100 89290 25180 89300
rect 25280 89290 25360 89300
rect 25460 89290 25540 89300
rect 25640 89290 25720 89300
rect 25820 89290 25900 89300
rect 26000 89290 26080 89300
rect 26180 89290 26260 89300
rect 26360 89290 26440 89300
rect 26540 89290 26620 89300
rect 30280 89290 30360 89300
rect 30460 89290 30540 89300
rect 30640 89290 30720 89300
rect 30820 89290 30900 89300
rect 31000 89290 31080 89300
rect 31180 89290 31260 89300
rect 31360 89290 31440 89300
rect 31540 89290 31620 89300
rect 31720 89290 31800 89300
rect 31900 89290 31980 89300
rect 32080 89290 32160 89300
rect 32260 89290 32340 89300
rect 32440 89290 32520 89300
rect 32620 89290 32700 89300
rect 32800 89290 32880 89300
rect 32980 89290 33060 89300
rect 33160 89290 33240 89300
rect 33340 89290 33420 89300
rect 33520 89290 33600 89300
rect 33700 89290 33780 89300
rect 33880 89290 33960 89300
rect 34060 89290 34140 89300
rect 34240 89290 34320 89300
rect 34420 89290 34500 89300
rect 34600 89290 34680 89300
rect 34780 89290 34860 89300
rect 34960 89290 35040 89300
rect 35140 89290 35220 89300
rect 35320 89290 35400 89300
rect 35500 89290 35580 89300
rect 35680 89290 35760 89300
rect 35860 89290 35940 89300
rect 36040 89290 36120 89300
rect 36220 89290 36300 89300
rect 36400 89290 36480 89300
rect 36580 89290 36660 89300
rect 36760 89290 36840 89300
rect 36940 89290 37020 89300
rect 37120 89290 37200 89300
rect 37300 89290 37380 89300
rect 37480 89290 37560 89300
rect 37660 89290 37740 89300
rect 37840 89290 37920 89300
rect 152080 89290 152160 89300
rect 152260 89290 152340 89300
rect 152440 89290 152520 89300
rect 152620 89290 152700 89300
rect 152800 89290 152880 89300
rect 152980 89290 153060 89300
rect 153160 89290 153240 89300
rect 153340 89290 153420 89300
rect 153520 89290 153600 89300
rect 153700 89290 153780 89300
rect 153880 89290 153960 89300
rect 154060 89290 154140 89300
rect 154240 89290 154320 89300
rect 154420 89290 154500 89300
rect 154600 89290 154680 89300
rect 154780 89290 154860 89300
rect 154960 89290 155040 89300
rect 155140 89290 155220 89300
rect 155320 89290 155400 89300
rect 155500 89290 155580 89300
rect 155680 89290 155760 89300
rect 155860 89290 155940 89300
rect 156040 89290 156120 89300
rect 156220 89290 156300 89300
rect 156400 89290 156480 89300
rect 156580 89290 156660 89300
rect 156760 89290 156840 89300
rect 156940 89290 157020 89300
rect 157120 89290 157200 89300
rect 157300 89290 157380 89300
rect 157480 89290 157560 89300
rect 157660 89290 157740 89300
rect 157840 89290 157920 89300
rect 158020 89290 158100 89300
rect 158200 89290 158280 89300
rect 158380 89290 158460 89300
rect 158560 89290 158640 89300
rect 158740 89290 158820 89300
rect 158920 89290 159000 89300
rect 159100 89290 159180 89300
rect 159280 89290 159360 89300
rect 159460 89290 159540 89300
rect 159640 89290 159720 89300
rect 163380 89290 163460 89300
rect 163560 89290 163640 89300
rect 163740 89290 163820 89300
rect 163920 89290 164000 89300
rect 164100 89290 164180 89300
rect 164280 89290 164360 89300
rect 164460 89290 164540 89300
rect 164640 89290 164720 89300
rect 164820 89290 164900 89300
rect 165000 89290 165080 89300
rect 165180 89290 165260 89300
rect 165360 89290 165440 89300
rect 165540 89290 165620 89300
rect 165720 89290 165800 89300
rect 165900 89290 165980 89300
rect 166080 89290 166160 89300
rect 166260 89290 166340 89300
rect 166440 89290 166520 89300
rect 166620 89290 166700 89300
rect 166800 89290 166880 89300
rect 166980 89290 167060 89300
rect 167160 89290 167240 89300
rect 167340 89290 167420 89300
rect 167520 89290 167600 89300
rect 167700 89290 167780 89300
rect 167880 89290 167960 89300
rect 168060 89290 168140 89300
rect 168240 89290 168320 89300
rect 168420 89290 168500 89300
rect 168600 89290 168680 89300
rect 168780 89290 168860 89300
rect 168960 89290 169040 89300
rect 169140 89290 169220 89300
rect 169320 89290 169400 89300
rect 169500 89290 169580 89300
rect 169680 89290 169760 89300
rect 169860 89290 169940 89300
rect 170040 89290 170120 89300
rect 170220 89290 170300 89300
rect 170400 89290 170480 89300
rect 170580 89290 170660 89300
rect 170760 89290 170840 89300
rect 170940 89290 171020 89300
rect 19060 89210 19070 89290
rect 19240 89210 19250 89290
rect 19420 89210 19430 89290
rect 19600 89210 19610 89290
rect 19780 89210 19790 89290
rect 19960 89210 19970 89290
rect 20140 89210 20150 89290
rect 20320 89210 20330 89290
rect 20500 89210 20510 89290
rect 20680 89210 20690 89290
rect 20860 89210 20870 89290
rect 21040 89210 21050 89290
rect 21220 89210 21230 89290
rect 21400 89210 21410 89290
rect 21580 89210 21590 89290
rect 21760 89210 21770 89290
rect 21940 89210 21950 89290
rect 22120 89210 22130 89290
rect 22300 89210 22310 89290
rect 22480 89210 22490 89290
rect 22660 89210 22670 89290
rect 22840 89210 22850 89290
rect 23020 89210 23030 89290
rect 23200 89210 23210 89290
rect 23380 89210 23390 89290
rect 23560 89210 23570 89290
rect 23740 89210 23750 89290
rect 23920 89210 23930 89290
rect 24100 89210 24110 89290
rect 24280 89210 24290 89290
rect 24460 89210 24470 89290
rect 24640 89210 24650 89290
rect 24820 89210 24830 89290
rect 25000 89210 25010 89290
rect 25180 89210 25190 89290
rect 25360 89210 25370 89290
rect 25540 89210 25550 89290
rect 25720 89210 25730 89290
rect 25900 89210 25910 89290
rect 26080 89210 26090 89290
rect 26260 89210 26270 89290
rect 26440 89210 26450 89290
rect 26620 89210 26630 89290
rect 27315 89235 27395 89245
rect 27495 89235 27575 89245
rect 27675 89235 27755 89245
rect 27855 89235 27935 89245
rect 28035 89235 28115 89245
rect 27395 89155 27405 89235
rect 27575 89155 27585 89235
rect 27755 89155 27765 89235
rect 27935 89155 27945 89235
rect 28115 89155 28125 89235
rect 30360 89210 30370 89290
rect 30540 89210 30550 89290
rect 30720 89210 30730 89290
rect 30900 89210 30910 89290
rect 31080 89210 31090 89290
rect 31260 89210 31270 89290
rect 31440 89210 31450 89290
rect 31620 89210 31630 89290
rect 31800 89210 31810 89290
rect 31980 89210 31990 89290
rect 32160 89210 32170 89290
rect 32340 89210 32350 89290
rect 32520 89210 32530 89290
rect 32700 89210 32710 89290
rect 32880 89210 32890 89290
rect 33060 89210 33070 89290
rect 33240 89210 33250 89290
rect 33420 89210 33430 89290
rect 33600 89210 33610 89290
rect 33780 89210 33790 89290
rect 33960 89210 33970 89290
rect 34140 89210 34150 89290
rect 34320 89210 34330 89290
rect 34500 89210 34510 89290
rect 34680 89210 34690 89290
rect 34860 89210 34870 89290
rect 35040 89210 35050 89290
rect 35220 89210 35230 89290
rect 35400 89210 35410 89290
rect 35580 89210 35590 89290
rect 35760 89210 35770 89290
rect 35940 89210 35950 89290
rect 36120 89210 36130 89290
rect 36300 89210 36310 89290
rect 36480 89210 36490 89290
rect 36660 89210 36670 89290
rect 36840 89210 36850 89290
rect 37020 89210 37030 89290
rect 37200 89210 37210 89290
rect 37380 89210 37390 89290
rect 37560 89210 37570 89290
rect 37740 89210 37750 89290
rect 37920 89210 37930 89290
rect 152160 89210 152170 89290
rect 152340 89210 152350 89290
rect 152520 89210 152530 89290
rect 152700 89210 152710 89290
rect 152880 89210 152890 89290
rect 153060 89210 153070 89290
rect 153240 89210 153250 89290
rect 153420 89210 153430 89290
rect 153600 89210 153610 89290
rect 153780 89210 153790 89290
rect 153960 89210 153970 89290
rect 154140 89210 154150 89290
rect 154320 89210 154330 89290
rect 154500 89210 154510 89290
rect 154680 89210 154690 89290
rect 154860 89210 154870 89290
rect 155040 89210 155050 89290
rect 155220 89210 155230 89290
rect 155400 89210 155410 89290
rect 155580 89210 155590 89290
rect 155760 89210 155770 89290
rect 155940 89210 155950 89290
rect 156120 89210 156130 89290
rect 156300 89210 156310 89290
rect 156480 89210 156490 89290
rect 156660 89210 156670 89290
rect 156840 89210 156850 89290
rect 157020 89210 157030 89290
rect 157200 89210 157210 89290
rect 157380 89210 157390 89290
rect 157560 89210 157570 89290
rect 157740 89210 157750 89290
rect 157920 89210 157930 89290
rect 158100 89210 158110 89290
rect 158280 89210 158290 89290
rect 158460 89210 158470 89290
rect 158640 89210 158650 89290
rect 158820 89210 158830 89290
rect 159000 89210 159010 89290
rect 159180 89210 159190 89290
rect 159360 89210 159370 89290
rect 159540 89210 159550 89290
rect 159720 89210 159730 89290
rect 160430 89265 160510 89275
rect 160590 89265 160670 89275
rect 160750 89265 160830 89275
rect 160910 89265 160990 89275
rect 161070 89265 161150 89275
rect 160510 89185 160520 89265
rect 160590 89185 160600 89265
rect 160670 89185 160680 89265
rect 160750 89185 160760 89265
rect 160830 89185 160840 89265
rect 160910 89185 160920 89265
rect 160990 89185 161000 89265
rect 161070 89185 161080 89265
rect 161150 89185 161160 89265
rect 163460 89210 163470 89290
rect 163640 89210 163650 89290
rect 163820 89210 163830 89290
rect 164000 89210 164010 89290
rect 164180 89210 164190 89290
rect 164360 89210 164370 89290
rect 164540 89210 164550 89290
rect 164720 89210 164730 89290
rect 164900 89210 164910 89290
rect 165080 89210 165090 89290
rect 165260 89210 165270 89290
rect 165440 89210 165450 89290
rect 165620 89210 165630 89290
rect 165800 89210 165810 89290
rect 165980 89210 165990 89290
rect 166160 89210 166170 89290
rect 166340 89210 166350 89290
rect 166520 89210 166530 89290
rect 166700 89210 166710 89290
rect 166880 89210 166890 89290
rect 167060 89210 167070 89290
rect 167240 89210 167250 89290
rect 167420 89210 167430 89290
rect 167600 89210 167610 89290
rect 167780 89210 167790 89290
rect 167960 89210 167970 89290
rect 168140 89210 168150 89290
rect 168320 89210 168330 89290
rect 168500 89210 168510 89290
rect 168680 89210 168690 89290
rect 168860 89210 168870 89290
rect 169040 89210 169050 89290
rect 169220 89210 169230 89290
rect 169400 89210 169410 89290
rect 169580 89210 169590 89290
rect 169760 89210 169770 89290
rect 169940 89210 169950 89290
rect 170120 89210 170130 89290
rect 170300 89210 170310 89290
rect 170480 89210 170490 89290
rect 170660 89210 170670 89290
rect 170840 89210 170850 89290
rect 171020 89210 171030 89290
rect 18980 89140 19060 89150
rect 19160 89140 19240 89150
rect 19340 89140 19420 89150
rect 19520 89140 19600 89150
rect 19700 89140 19780 89150
rect 19880 89140 19960 89150
rect 20060 89140 20140 89150
rect 20240 89140 20320 89150
rect 20420 89140 20500 89150
rect 20600 89140 20680 89150
rect 20780 89140 20860 89150
rect 20960 89140 21040 89150
rect 21140 89140 21220 89150
rect 21320 89140 21400 89150
rect 21500 89140 21580 89150
rect 21680 89140 21760 89150
rect 21860 89140 21940 89150
rect 22040 89140 22120 89150
rect 22220 89140 22300 89150
rect 22400 89140 22480 89150
rect 22580 89140 22660 89150
rect 22760 89140 22840 89150
rect 22940 89140 23020 89150
rect 23120 89140 23200 89150
rect 23300 89140 23380 89150
rect 23480 89140 23560 89150
rect 23660 89140 23740 89150
rect 23840 89140 23920 89150
rect 24020 89140 24100 89150
rect 24200 89140 24280 89150
rect 24380 89140 24460 89150
rect 24560 89140 24640 89150
rect 24740 89140 24820 89150
rect 24920 89140 25000 89150
rect 25100 89140 25180 89150
rect 25280 89140 25360 89150
rect 25460 89140 25540 89150
rect 25640 89140 25720 89150
rect 25820 89140 25900 89150
rect 26000 89140 26080 89150
rect 26180 89140 26260 89150
rect 26360 89140 26440 89150
rect 26540 89140 26620 89150
rect 30280 89140 30360 89150
rect 30460 89140 30540 89150
rect 30640 89140 30720 89150
rect 30820 89140 30900 89150
rect 31000 89140 31080 89150
rect 31180 89140 31260 89150
rect 31360 89140 31440 89150
rect 31540 89140 31620 89150
rect 31720 89140 31800 89150
rect 31900 89140 31980 89150
rect 32080 89140 32160 89150
rect 32260 89140 32340 89150
rect 32440 89140 32520 89150
rect 32620 89140 32700 89150
rect 32800 89140 32880 89150
rect 32980 89140 33060 89150
rect 33160 89140 33240 89150
rect 33340 89140 33420 89150
rect 33520 89140 33600 89150
rect 33700 89140 33780 89150
rect 33880 89140 33960 89150
rect 34060 89140 34140 89150
rect 34240 89140 34320 89150
rect 34420 89140 34500 89150
rect 34600 89140 34680 89150
rect 34780 89140 34860 89150
rect 34960 89140 35040 89150
rect 35140 89140 35220 89150
rect 35320 89140 35400 89150
rect 35500 89140 35580 89150
rect 35680 89140 35760 89150
rect 35860 89140 35940 89150
rect 36040 89140 36120 89150
rect 36220 89140 36300 89150
rect 36400 89140 36480 89150
rect 36580 89140 36660 89150
rect 36760 89140 36840 89150
rect 36940 89140 37020 89150
rect 37120 89140 37200 89150
rect 37300 89140 37380 89150
rect 37480 89140 37560 89150
rect 37660 89140 37740 89150
rect 37840 89140 37920 89150
rect 40060 89140 40140 89150
rect 40200 89140 40280 89150
rect 40340 89140 40420 89150
rect 40480 89140 40560 89150
rect 40620 89140 40700 89150
rect 40760 89140 40840 89150
rect 40900 89140 40980 89150
rect 41040 89140 41120 89150
rect 41180 89140 41260 89150
rect 41320 89140 41400 89150
rect 42360 89140 42440 89150
rect 42500 89140 42580 89150
rect 42640 89140 42720 89150
rect 42780 89140 42860 89150
rect 42920 89140 43000 89150
rect 43060 89140 43140 89150
rect 43200 89140 43280 89150
rect 43340 89140 43420 89150
rect 43480 89140 43560 89150
rect 43620 89140 43700 89150
rect 146300 89140 146380 89150
rect 146440 89140 146520 89150
rect 146580 89140 146660 89150
rect 146720 89140 146800 89150
rect 146860 89140 146940 89150
rect 147000 89140 147080 89150
rect 147140 89140 147220 89150
rect 147280 89140 147360 89150
rect 147420 89140 147500 89150
rect 147560 89140 147640 89150
rect 148600 89140 148680 89150
rect 148740 89140 148820 89150
rect 148880 89140 148960 89150
rect 149020 89140 149100 89150
rect 149160 89140 149240 89150
rect 149300 89140 149380 89150
rect 149440 89140 149520 89150
rect 149580 89140 149660 89150
rect 149720 89140 149800 89150
rect 149860 89140 149940 89150
rect 152080 89140 152160 89150
rect 152260 89140 152340 89150
rect 152440 89140 152520 89150
rect 152620 89140 152700 89150
rect 152800 89140 152880 89150
rect 152980 89140 153060 89150
rect 153160 89140 153240 89150
rect 153340 89140 153420 89150
rect 153520 89140 153600 89150
rect 153700 89140 153780 89150
rect 153880 89140 153960 89150
rect 154060 89140 154140 89150
rect 154240 89140 154320 89150
rect 154420 89140 154500 89150
rect 154600 89140 154680 89150
rect 154780 89140 154860 89150
rect 154960 89140 155040 89150
rect 155140 89140 155220 89150
rect 155320 89140 155400 89150
rect 155500 89140 155580 89150
rect 155680 89140 155760 89150
rect 155860 89140 155940 89150
rect 156040 89140 156120 89150
rect 156220 89140 156300 89150
rect 156400 89140 156480 89150
rect 156580 89140 156660 89150
rect 156760 89140 156840 89150
rect 156940 89140 157020 89150
rect 157120 89140 157200 89150
rect 157300 89140 157380 89150
rect 157480 89140 157560 89150
rect 157660 89140 157740 89150
rect 157840 89140 157920 89150
rect 158020 89140 158100 89150
rect 158200 89140 158280 89150
rect 158380 89140 158460 89150
rect 158560 89140 158640 89150
rect 158740 89140 158820 89150
rect 158920 89140 159000 89150
rect 159100 89140 159180 89150
rect 159280 89140 159360 89150
rect 159460 89140 159540 89150
rect 159640 89140 159720 89150
rect 163380 89140 163460 89150
rect 163560 89140 163640 89150
rect 163740 89140 163820 89150
rect 163920 89140 164000 89150
rect 164100 89140 164180 89150
rect 164280 89140 164360 89150
rect 164460 89140 164540 89150
rect 164640 89140 164720 89150
rect 164820 89140 164900 89150
rect 165000 89140 165080 89150
rect 165180 89140 165260 89150
rect 165360 89140 165440 89150
rect 165540 89140 165620 89150
rect 165720 89140 165800 89150
rect 165900 89140 165980 89150
rect 166080 89140 166160 89150
rect 166260 89140 166340 89150
rect 166440 89140 166520 89150
rect 166620 89140 166700 89150
rect 166800 89140 166880 89150
rect 166980 89140 167060 89150
rect 167160 89140 167240 89150
rect 167340 89140 167420 89150
rect 167520 89140 167600 89150
rect 167700 89140 167780 89150
rect 167880 89140 167960 89150
rect 168060 89140 168140 89150
rect 168240 89140 168320 89150
rect 168420 89140 168500 89150
rect 168600 89140 168680 89150
rect 168780 89140 168860 89150
rect 168960 89140 169040 89150
rect 169140 89140 169220 89150
rect 169320 89140 169400 89150
rect 169500 89140 169580 89150
rect 169680 89140 169760 89150
rect 169860 89140 169940 89150
rect 170040 89140 170120 89150
rect 170220 89140 170300 89150
rect 170400 89140 170480 89150
rect 170580 89140 170660 89150
rect 170760 89140 170840 89150
rect 170940 89140 171020 89150
rect 19060 89060 19070 89140
rect 19240 89060 19250 89140
rect 19420 89060 19430 89140
rect 19600 89060 19610 89140
rect 19780 89060 19790 89140
rect 19960 89060 19970 89140
rect 20140 89060 20150 89140
rect 20320 89060 20330 89140
rect 20500 89060 20510 89140
rect 20680 89060 20690 89140
rect 20860 89060 20870 89140
rect 21040 89060 21050 89140
rect 21220 89060 21230 89140
rect 21400 89060 21410 89140
rect 21580 89060 21590 89140
rect 21760 89060 21770 89140
rect 21940 89060 21950 89140
rect 22120 89060 22130 89140
rect 22300 89060 22310 89140
rect 22480 89060 22490 89140
rect 22660 89060 22670 89140
rect 22840 89060 22850 89140
rect 23020 89060 23030 89140
rect 23200 89060 23210 89140
rect 23380 89060 23390 89140
rect 23560 89060 23570 89140
rect 23740 89060 23750 89140
rect 23920 89060 23930 89140
rect 24100 89060 24110 89140
rect 24280 89060 24290 89140
rect 24460 89060 24470 89140
rect 24640 89060 24650 89140
rect 24820 89060 24830 89140
rect 25000 89060 25010 89140
rect 25180 89060 25190 89140
rect 25360 89060 25370 89140
rect 25540 89060 25550 89140
rect 25720 89060 25730 89140
rect 25900 89060 25910 89140
rect 26080 89060 26090 89140
rect 26260 89060 26270 89140
rect 26440 89060 26450 89140
rect 26620 89060 26630 89140
rect 30360 89060 30370 89140
rect 30540 89060 30550 89140
rect 30720 89060 30730 89140
rect 30900 89060 30910 89140
rect 31080 89060 31090 89140
rect 31260 89060 31270 89140
rect 31440 89060 31450 89140
rect 31620 89060 31630 89140
rect 31800 89060 31810 89140
rect 31980 89060 31990 89140
rect 32160 89060 32170 89140
rect 32340 89060 32350 89140
rect 32520 89060 32530 89140
rect 32700 89060 32710 89140
rect 32880 89060 32890 89140
rect 33060 89060 33070 89140
rect 33240 89060 33250 89140
rect 33420 89060 33430 89140
rect 33600 89060 33610 89140
rect 33780 89060 33790 89140
rect 33960 89060 33970 89140
rect 34140 89060 34150 89140
rect 34320 89060 34330 89140
rect 34500 89060 34510 89140
rect 34680 89060 34690 89140
rect 34860 89060 34870 89140
rect 35040 89060 35050 89140
rect 35220 89060 35230 89140
rect 35400 89060 35410 89140
rect 35580 89060 35590 89140
rect 35760 89060 35770 89140
rect 35940 89060 35950 89140
rect 36120 89060 36130 89140
rect 36300 89060 36310 89140
rect 36480 89060 36490 89140
rect 36660 89060 36670 89140
rect 36840 89060 36850 89140
rect 37020 89060 37030 89140
rect 37200 89060 37210 89140
rect 37380 89060 37390 89140
rect 37560 89060 37570 89140
rect 37740 89060 37750 89140
rect 37920 89060 37930 89140
rect 40140 89060 40150 89140
rect 40280 89060 40290 89140
rect 40420 89060 40430 89140
rect 40560 89060 40570 89140
rect 40700 89060 40710 89140
rect 40840 89060 40850 89140
rect 40980 89060 40990 89140
rect 41120 89060 41130 89140
rect 41260 89060 41270 89140
rect 41400 89060 41410 89140
rect 42440 89060 42450 89140
rect 42580 89060 42590 89140
rect 42720 89060 42730 89140
rect 42860 89060 42870 89140
rect 43000 89060 43010 89140
rect 43140 89060 43150 89140
rect 43280 89060 43290 89140
rect 43420 89060 43430 89140
rect 43560 89060 43570 89140
rect 43700 89060 43710 89140
rect 146380 89081 146390 89140
rect 146520 89081 146530 89140
rect 146660 89081 146670 89140
rect 146800 89081 146810 89140
rect 146940 89081 146950 89140
rect 147080 89081 147090 89140
rect 147220 89081 147230 89140
rect 147360 89081 147370 89140
rect 147500 89081 147510 89140
rect 147640 89081 147650 89140
rect 148680 89081 148690 89140
rect 148820 89081 148830 89140
rect 148960 89081 148970 89140
rect 149100 89081 149110 89140
rect 149240 89081 149250 89140
rect 149380 89081 149390 89140
rect 149520 89081 149530 89140
rect 149660 89081 149670 89140
rect 149800 89081 149810 89140
rect 149940 89081 149950 89140
rect 152160 89081 152170 89140
rect 152340 89081 152350 89140
rect 152520 89081 152530 89140
rect 152700 89081 152710 89140
rect 152880 89081 152890 89140
rect 153060 89081 153070 89140
rect 153240 89081 153250 89140
rect 153420 89081 153430 89140
rect 153600 89081 153610 89140
rect 153780 89081 153790 89140
rect 153960 89081 153970 89140
rect 154140 89081 154150 89140
rect 154320 89081 154330 89140
rect 154500 89081 154510 89140
rect 154680 89081 154690 89140
rect 154860 89081 154870 89140
rect 155040 89081 155050 89140
rect 155220 89081 155230 89140
rect 155400 89081 155410 89140
rect 155580 89081 155590 89140
rect 155760 89081 155770 89140
rect 155940 89081 155950 89140
rect 156120 89081 156130 89140
rect 156300 89081 156310 89140
rect 156480 89081 156490 89140
rect 156660 89081 156670 89140
rect 156840 89081 156850 89140
rect 157020 89081 157030 89140
rect 157200 89081 157210 89140
rect 157380 89081 157390 89140
rect 157560 89081 157570 89140
rect 157740 89081 157750 89140
rect 157920 89081 157930 89140
rect 158100 89081 158110 89140
rect 158280 89081 158290 89140
rect 158460 89081 158470 89140
rect 158640 89081 158650 89140
rect 158820 89081 158830 89140
rect 159000 89081 159010 89140
rect 159180 89081 159190 89140
rect 159360 89081 159370 89140
rect 159540 89081 159550 89140
rect 159720 89081 159730 89140
rect 163460 89081 163470 89140
rect 163640 89081 163650 89140
rect 163820 89081 163830 89140
rect 164000 89081 164010 89140
rect 164180 89081 164190 89140
rect 164360 89081 164370 89140
rect 164540 89081 164550 89140
rect 164720 89081 164730 89140
rect 164900 89081 164910 89140
rect 165080 89081 165090 89140
rect 165260 89081 165270 89140
rect 165440 89081 165450 89140
rect 165620 89081 165630 89140
rect 165800 89081 165810 89140
rect 165980 89081 165990 89140
rect 166160 89081 166170 89140
rect 166340 89081 166350 89140
rect 166520 89081 166530 89140
rect 166700 89081 166710 89140
rect 166880 89081 166890 89140
rect 167060 89081 167070 89140
rect 167240 89081 167250 89140
rect 167420 89081 167430 89140
rect 167600 89081 167610 89140
rect 167780 89081 167790 89140
rect 167960 89081 167970 89140
rect 168140 89081 168150 89140
rect 168320 89081 168330 89140
rect 168500 89081 168510 89140
rect 168680 89081 168690 89140
rect 168860 89081 168870 89140
rect 169040 89081 169050 89140
rect 169220 89081 169230 89140
rect 169400 89081 169410 89140
rect 169580 89081 169590 89140
rect 169760 89081 169770 89140
rect 169940 89081 169950 89140
rect 170120 89081 170130 89140
rect 170300 89081 170310 89140
rect 170480 89081 170490 89140
rect 170660 89081 170670 89140
rect 170840 89081 170850 89140
rect 171020 89081 171030 89140
rect 146040 89000 147700 89081
rect 148340 89000 150000 89081
rect 152000 89000 159800 89081
rect 163210 89060 171100 89081
rect 163300 89000 171100 89060
rect 30360 88920 30440 88930
rect 30680 88920 30760 88930
rect 31000 88920 31080 88930
rect 31320 88920 31400 88930
rect 31640 88920 31720 88930
rect 31960 88920 32040 88930
rect 32280 88920 32360 88930
rect 32600 88920 32680 88930
rect 32920 88920 33000 88930
rect 33240 88920 33320 88930
rect 33560 88920 33640 88930
rect 33880 88920 33960 88930
rect 34200 88920 34280 88930
rect 34520 88920 34600 88930
rect 34840 88920 34920 88930
rect 35160 88920 35240 88930
rect 35480 88920 35560 88930
rect 35800 88920 35880 88930
rect 36120 88920 36200 88930
rect 36440 88920 36520 88930
rect 36760 88920 36840 88930
rect 37080 88920 37160 88930
rect 37400 88920 37480 88930
rect 37720 88920 37800 88930
rect 40180 88920 40260 88930
rect 40500 88920 40580 88930
rect 40820 88920 40900 88930
rect 41140 88920 41220 88930
rect 42560 88920 42640 88930
rect 42880 88920 42960 88930
rect 43200 88920 43280 88930
rect 43520 88920 43600 88930
rect 18970 88890 19050 88900
rect 19290 88890 19370 88900
rect 19610 88890 19690 88900
rect 19930 88890 20010 88900
rect 20250 88890 20330 88900
rect 20570 88890 20650 88900
rect 20890 88890 20970 88900
rect 21210 88890 21290 88900
rect 21530 88890 21610 88900
rect 21850 88890 21930 88900
rect 22170 88890 22250 88900
rect 22490 88890 22570 88900
rect 22810 88890 22890 88900
rect 23130 88890 23210 88900
rect 23450 88890 23530 88900
rect 23770 88890 23850 88900
rect 24090 88890 24170 88900
rect 24410 88890 24490 88900
rect 24730 88890 24810 88900
rect 25050 88890 25130 88900
rect 25370 88890 25450 88900
rect 25690 88890 25770 88900
rect 26010 88890 26090 88900
rect 26330 88890 26410 88900
rect 19050 88810 19060 88890
rect 19370 88810 19380 88890
rect 19690 88810 19700 88890
rect 20010 88810 20020 88890
rect 20330 88810 20340 88890
rect 20650 88810 20660 88890
rect 20970 88810 20980 88890
rect 21290 88810 21300 88890
rect 21610 88810 21620 88890
rect 21930 88810 21940 88890
rect 22250 88810 22260 88890
rect 22570 88810 22580 88890
rect 22890 88810 22900 88890
rect 23210 88810 23220 88890
rect 23530 88810 23540 88890
rect 23850 88810 23860 88890
rect 24170 88810 24180 88890
rect 24490 88810 24500 88890
rect 24810 88810 24820 88890
rect 25130 88810 25140 88890
rect 25450 88810 25460 88890
rect 25770 88810 25780 88890
rect 26090 88810 26100 88890
rect 26410 88810 26420 88890
rect 30440 88840 30450 88920
rect 30760 88840 30770 88920
rect 31080 88840 31090 88920
rect 31400 88840 31410 88920
rect 31720 88840 31730 88920
rect 32040 88840 32050 88920
rect 32360 88840 32370 88920
rect 32680 88840 32690 88920
rect 33000 88840 33010 88920
rect 33320 88840 33330 88920
rect 33640 88840 33650 88920
rect 33960 88840 33970 88920
rect 34280 88840 34290 88920
rect 34600 88840 34610 88920
rect 34920 88840 34930 88920
rect 35240 88840 35250 88920
rect 35560 88840 35570 88920
rect 35880 88840 35890 88920
rect 36200 88840 36210 88920
rect 36520 88840 36530 88920
rect 36840 88840 36850 88920
rect 37160 88840 37170 88920
rect 37480 88840 37490 88920
rect 37800 88840 37810 88920
rect 40260 88840 40270 88920
rect 40580 88840 40590 88920
rect 40900 88840 40910 88920
rect 41220 88840 41230 88920
rect 42640 88840 42650 88920
rect 42960 88840 42970 88920
rect 43280 88840 43290 88920
rect 43600 88840 43610 88920
rect 146400 88911 146480 88921
rect 146720 88911 146800 88921
rect 147040 88911 147120 88921
rect 147360 88911 147440 88921
rect 148780 88911 148860 88921
rect 149100 88911 149180 88921
rect 149420 88911 149500 88921
rect 149740 88911 149820 88921
rect 152200 88911 152280 88921
rect 152520 88911 152600 88921
rect 152840 88911 152920 88921
rect 153160 88911 153240 88921
rect 153480 88911 153560 88921
rect 153800 88911 153880 88921
rect 154120 88911 154200 88921
rect 154440 88911 154520 88921
rect 154760 88911 154840 88921
rect 155080 88911 155160 88921
rect 155400 88911 155480 88921
rect 155720 88911 155800 88921
rect 156040 88911 156120 88921
rect 156360 88911 156440 88921
rect 156680 88911 156760 88921
rect 157000 88911 157080 88921
rect 157320 88911 157400 88921
rect 157640 88911 157720 88921
rect 157960 88911 158040 88921
rect 158280 88911 158360 88921
rect 158600 88911 158680 88921
rect 158920 88911 159000 88921
rect 159240 88911 159320 88921
rect 159560 88911 159640 88921
rect 146480 88831 146490 88911
rect 146800 88831 146810 88911
rect 147120 88831 147130 88911
rect 147440 88831 147450 88911
rect 148860 88831 148870 88911
rect 149180 88831 149190 88911
rect 149500 88831 149510 88911
rect 149820 88831 149830 88911
rect 152280 88831 152290 88911
rect 152600 88831 152610 88911
rect 152920 88831 152930 88911
rect 153240 88831 153250 88911
rect 153560 88831 153570 88911
rect 153880 88831 153890 88911
rect 154200 88831 154210 88911
rect 154520 88831 154530 88911
rect 154840 88831 154850 88911
rect 155160 88831 155170 88911
rect 155480 88831 155490 88911
rect 155800 88831 155810 88911
rect 156120 88831 156130 88911
rect 156440 88831 156450 88911
rect 156760 88831 156770 88911
rect 157080 88831 157090 88911
rect 157400 88831 157410 88911
rect 157720 88831 157730 88911
rect 158040 88831 158050 88911
rect 158360 88831 158370 88911
rect 158680 88831 158690 88911
rect 159000 88831 159010 88911
rect 159320 88831 159330 88911
rect 159640 88831 159650 88911
rect 163590 88881 163670 88891
rect 163910 88881 163990 88891
rect 164230 88881 164310 88891
rect 164550 88881 164630 88891
rect 164870 88881 164950 88891
rect 165190 88881 165270 88891
rect 165510 88881 165590 88891
rect 165830 88881 165910 88891
rect 166150 88881 166230 88891
rect 166470 88881 166550 88891
rect 166790 88881 166870 88891
rect 167110 88881 167190 88891
rect 167430 88881 167510 88891
rect 167750 88881 167830 88891
rect 168070 88881 168150 88891
rect 168390 88881 168470 88891
rect 168710 88881 168790 88891
rect 169030 88881 169110 88891
rect 169350 88881 169430 88891
rect 169670 88881 169750 88891
rect 169990 88881 170070 88891
rect 170310 88881 170390 88891
rect 170630 88881 170710 88891
rect 170950 88881 171030 88891
rect 163670 88801 163680 88881
rect 163990 88801 164000 88881
rect 164310 88801 164320 88881
rect 164630 88801 164640 88881
rect 164950 88801 164960 88881
rect 165270 88801 165280 88881
rect 165590 88801 165600 88881
rect 165910 88801 165920 88881
rect 166230 88801 166240 88881
rect 166550 88801 166560 88881
rect 166870 88801 166880 88881
rect 167190 88801 167200 88881
rect 167510 88801 167520 88881
rect 167830 88801 167840 88881
rect 168150 88801 168160 88881
rect 168470 88801 168480 88881
rect 168790 88801 168800 88881
rect 169110 88801 169120 88881
rect 169430 88801 169440 88881
rect 169750 88801 169760 88881
rect 170070 88801 170080 88881
rect 170390 88801 170400 88881
rect 170710 88801 170720 88881
rect 171030 88801 171040 88881
rect 30520 88760 30600 88770
rect 30840 88760 30920 88770
rect 31160 88760 31240 88770
rect 31480 88760 31560 88770
rect 31800 88760 31880 88770
rect 32120 88760 32200 88770
rect 32440 88760 32520 88770
rect 32760 88760 32840 88770
rect 33080 88760 33160 88770
rect 33400 88760 33480 88770
rect 33720 88760 33800 88770
rect 34040 88760 34120 88770
rect 34360 88760 34440 88770
rect 34680 88760 34760 88770
rect 35000 88760 35080 88770
rect 35320 88760 35400 88770
rect 35640 88760 35720 88770
rect 35960 88760 36040 88770
rect 36280 88760 36360 88770
rect 36600 88760 36680 88770
rect 36920 88760 37000 88770
rect 37240 88760 37320 88770
rect 37560 88760 37640 88770
rect 40340 88760 40420 88770
rect 40660 88760 40740 88770
rect 40980 88760 41060 88770
rect 42720 88760 42800 88770
rect 43040 88760 43120 88770
rect 43360 88760 43440 88770
rect 19130 88730 19210 88740
rect 19450 88730 19530 88740
rect 19770 88730 19850 88740
rect 20090 88730 20170 88740
rect 20410 88730 20490 88740
rect 20730 88730 20810 88740
rect 21050 88730 21130 88740
rect 21370 88730 21450 88740
rect 21690 88730 21770 88740
rect 22010 88730 22090 88740
rect 22330 88730 22410 88740
rect 22650 88730 22730 88740
rect 22970 88730 23050 88740
rect 23290 88730 23370 88740
rect 23610 88730 23690 88740
rect 23930 88730 24010 88740
rect 24250 88730 24330 88740
rect 24570 88730 24650 88740
rect 24890 88730 24970 88740
rect 25210 88730 25290 88740
rect 25530 88730 25610 88740
rect 25850 88730 25930 88740
rect 26170 88730 26250 88740
rect 19210 88650 19220 88730
rect 19530 88650 19540 88730
rect 19850 88650 19860 88730
rect 20170 88650 20180 88730
rect 20490 88650 20500 88730
rect 20810 88650 20820 88730
rect 21130 88650 21140 88730
rect 21450 88650 21460 88730
rect 21770 88650 21780 88730
rect 22090 88650 22100 88730
rect 22410 88650 22420 88730
rect 22730 88650 22740 88730
rect 23050 88650 23060 88730
rect 23370 88650 23380 88730
rect 23690 88650 23700 88730
rect 24010 88650 24020 88730
rect 24330 88650 24340 88730
rect 24650 88650 24660 88730
rect 24970 88650 24980 88730
rect 25290 88650 25300 88730
rect 25610 88650 25620 88730
rect 25930 88650 25940 88730
rect 26250 88650 26260 88730
rect 30600 88680 30610 88760
rect 30920 88680 30930 88760
rect 31240 88680 31250 88760
rect 31560 88680 31570 88760
rect 31880 88680 31890 88760
rect 32200 88680 32210 88760
rect 32520 88680 32530 88760
rect 32840 88680 32850 88760
rect 33160 88680 33170 88760
rect 33480 88680 33490 88760
rect 33800 88680 33810 88760
rect 34120 88680 34130 88760
rect 34440 88680 34450 88760
rect 34760 88680 34770 88760
rect 35080 88680 35090 88760
rect 35400 88680 35410 88760
rect 35720 88680 35730 88760
rect 36040 88680 36050 88760
rect 36360 88680 36370 88760
rect 36680 88680 36690 88760
rect 37000 88680 37010 88760
rect 37320 88680 37330 88760
rect 37640 88680 37650 88760
rect 40420 88680 40430 88760
rect 40740 88680 40750 88760
rect 41060 88680 41070 88760
rect 42800 88680 42810 88760
rect 43120 88680 43130 88760
rect 43440 88680 43450 88760
rect 146560 88751 146640 88761
rect 146880 88751 146960 88761
rect 147200 88751 147280 88761
rect 148940 88751 149020 88761
rect 149260 88751 149340 88761
rect 149580 88751 149660 88761
rect 152360 88751 152440 88761
rect 152680 88751 152760 88761
rect 153000 88751 153080 88761
rect 153320 88751 153400 88761
rect 153640 88751 153720 88761
rect 153960 88751 154040 88761
rect 154280 88751 154360 88761
rect 154600 88751 154680 88761
rect 154920 88751 155000 88761
rect 155240 88751 155320 88761
rect 155560 88751 155640 88761
rect 155880 88751 155960 88761
rect 156200 88751 156280 88761
rect 156520 88751 156600 88761
rect 156840 88751 156920 88761
rect 157160 88751 157240 88761
rect 157480 88751 157560 88761
rect 157800 88751 157880 88761
rect 158120 88751 158200 88761
rect 158440 88751 158520 88761
rect 158760 88751 158840 88761
rect 159080 88751 159160 88761
rect 159400 88751 159480 88761
rect 146640 88671 146650 88751
rect 146960 88671 146970 88751
rect 147280 88671 147290 88751
rect 149020 88671 149030 88751
rect 149340 88671 149350 88751
rect 149660 88671 149670 88751
rect 152440 88671 152450 88751
rect 152760 88671 152770 88751
rect 153080 88671 153090 88751
rect 153400 88671 153410 88751
rect 153720 88671 153730 88751
rect 154040 88671 154050 88751
rect 154360 88671 154370 88751
rect 154680 88671 154690 88751
rect 155000 88671 155010 88751
rect 155320 88671 155330 88751
rect 155640 88671 155650 88751
rect 155960 88671 155970 88751
rect 156280 88671 156290 88751
rect 156600 88671 156610 88751
rect 156920 88671 156930 88751
rect 157240 88671 157250 88751
rect 157560 88671 157570 88751
rect 157880 88671 157890 88751
rect 158200 88671 158210 88751
rect 158520 88671 158530 88751
rect 158840 88671 158850 88751
rect 159160 88671 159170 88751
rect 159480 88671 159490 88751
rect 163750 88721 163830 88731
rect 164070 88721 164150 88731
rect 164390 88721 164470 88731
rect 164710 88721 164790 88731
rect 165030 88721 165110 88731
rect 165350 88721 165430 88731
rect 165670 88721 165750 88731
rect 165990 88721 166070 88731
rect 166310 88721 166390 88731
rect 166630 88721 166710 88731
rect 166950 88721 167030 88731
rect 167270 88721 167350 88731
rect 167590 88721 167670 88731
rect 167910 88721 167990 88731
rect 168230 88721 168310 88731
rect 168550 88721 168630 88731
rect 168870 88721 168950 88731
rect 169190 88721 169270 88731
rect 169510 88721 169590 88731
rect 169830 88721 169910 88731
rect 170150 88721 170230 88731
rect 170470 88721 170550 88731
rect 170790 88721 170870 88731
rect 163830 88641 163840 88721
rect 164150 88641 164160 88721
rect 164470 88641 164480 88721
rect 164790 88641 164800 88721
rect 165110 88641 165120 88721
rect 165430 88641 165440 88721
rect 165750 88641 165760 88721
rect 166070 88641 166080 88721
rect 166390 88641 166400 88721
rect 166710 88641 166720 88721
rect 167030 88641 167040 88721
rect 167350 88641 167360 88721
rect 167670 88641 167680 88721
rect 167990 88641 168000 88721
rect 168310 88641 168320 88721
rect 168630 88641 168640 88721
rect 168950 88641 168960 88721
rect 169270 88641 169280 88721
rect 169590 88641 169600 88721
rect 169910 88641 169920 88721
rect 170230 88641 170240 88721
rect 170550 88641 170560 88721
rect 170870 88641 170880 88721
rect 30360 88600 30440 88610
rect 30680 88600 30760 88610
rect 31000 88600 31080 88610
rect 31320 88600 31400 88610
rect 31640 88600 31720 88610
rect 31960 88600 32040 88610
rect 32280 88600 32360 88610
rect 32600 88600 32680 88610
rect 32920 88600 33000 88610
rect 33240 88600 33320 88610
rect 33560 88600 33640 88610
rect 33880 88600 33960 88610
rect 34200 88600 34280 88610
rect 34520 88600 34600 88610
rect 34840 88600 34920 88610
rect 35160 88600 35240 88610
rect 35480 88600 35560 88610
rect 35800 88600 35880 88610
rect 36120 88600 36200 88610
rect 36440 88600 36520 88610
rect 36760 88600 36840 88610
rect 37080 88600 37160 88610
rect 37400 88600 37480 88610
rect 37720 88600 37800 88610
rect 40180 88600 40260 88610
rect 40500 88600 40580 88610
rect 40820 88600 40900 88610
rect 41140 88600 41220 88610
rect 42560 88600 42640 88610
rect 42880 88600 42960 88610
rect 43200 88600 43280 88610
rect 43520 88600 43600 88610
rect 18970 88570 19050 88580
rect 19290 88570 19370 88580
rect 19610 88570 19690 88580
rect 19930 88570 20010 88580
rect 20250 88570 20330 88580
rect 20570 88570 20650 88580
rect 20890 88570 20970 88580
rect 21210 88570 21290 88580
rect 21530 88570 21610 88580
rect 21850 88570 21930 88580
rect 22170 88570 22250 88580
rect 22490 88570 22570 88580
rect 22810 88570 22890 88580
rect 23130 88570 23210 88580
rect 23450 88570 23530 88580
rect 23770 88570 23850 88580
rect 24090 88570 24170 88580
rect 24410 88570 24490 88580
rect 24730 88570 24810 88580
rect 25050 88570 25130 88580
rect 25370 88570 25450 88580
rect 25690 88570 25770 88580
rect 26010 88570 26090 88580
rect 26330 88570 26410 88580
rect 19050 88490 19060 88570
rect 19370 88490 19380 88570
rect 19690 88490 19700 88570
rect 20010 88490 20020 88570
rect 20330 88490 20340 88570
rect 20650 88490 20660 88570
rect 20970 88490 20980 88570
rect 21290 88490 21300 88570
rect 21610 88490 21620 88570
rect 21930 88490 21940 88570
rect 22250 88490 22260 88570
rect 22570 88490 22580 88570
rect 22890 88490 22900 88570
rect 23210 88490 23220 88570
rect 23530 88490 23540 88570
rect 23850 88490 23860 88570
rect 24170 88490 24180 88570
rect 24490 88490 24500 88570
rect 24810 88490 24820 88570
rect 25130 88490 25140 88570
rect 25450 88490 25460 88570
rect 25770 88490 25780 88570
rect 26090 88490 26100 88570
rect 26410 88490 26420 88570
rect 30440 88520 30450 88600
rect 30760 88520 30770 88600
rect 31080 88520 31090 88600
rect 31400 88520 31410 88600
rect 31720 88520 31730 88600
rect 32040 88520 32050 88600
rect 32360 88520 32370 88600
rect 32680 88520 32690 88600
rect 33000 88520 33010 88600
rect 33320 88520 33330 88600
rect 33640 88520 33650 88600
rect 33960 88520 33970 88600
rect 34280 88520 34290 88600
rect 34600 88520 34610 88600
rect 34920 88520 34930 88600
rect 35240 88520 35250 88600
rect 35560 88520 35570 88600
rect 35880 88520 35890 88600
rect 36200 88520 36210 88600
rect 36520 88520 36530 88600
rect 36840 88520 36850 88600
rect 37160 88520 37170 88600
rect 37480 88520 37490 88600
rect 37800 88520 37810 88600
rect 40260 88520 40270 88600
rect 40580 88520 40590 88600
rect 40900 88520 40910 88600
rect 41220 88520 41230 88600
rect 42640 88520 42650 88600
rect 42960 88520 42970 88600
rect 43280 88520 43290 88600
rect 43600 88520 43610 88600
rect 146400 88591 146480 88601
rect 146720 88591 146800 88601
rect 147040 88591 147120 88601
rect 147360 88591 147440 88601
rect 148780 88591 148860 88601
rect 149100 88591 149180 88601
rect 149420 88591 149500 88601
rect 149740 88591 149820 88601
rect 152200 88591 152280 88601
rect 152520 88591 152600 88601
rect 152840 88591 152920 88601
rect 153160 88591 153240 88601
rect 153480 88591 153560 88601
rect 153800 88591 153880 88601
rect 154120 88591 154200 88601
rect 154440 88591 154520 88601
rect 154760 88591 154840 88601
rect 155080 88591 155160 88601
rect 155400 88591 155480 88601
rect 155720 88591 155800 88601
rect 156040 88591 156120 88601
rect 156360 88591 156440 88601
rect 156680 88591 156760 88601
rect 157000 88591 157080 88601
rect 157320 88591 157400 88601
rect 157640 88591 157720 88601
rect 157960 88591 158040 88601
rect 158280 88591 158360 88601
rect 158600 88591 158680 88601
rect 158920 88591 159000 88601
rect 159240 88591 159320 88601
rect 159560 88591 159640 88601
rect 146480 88511 146490 88591
rect 146800 88511 146810 88591
rect 147120 88511 147130 88591
rect 147440 88511 147450 88591
rect 148860 88511 148870 88591
rect 149180 88511 149190 88591
rect 149500 88511 149510 88591
rect 149820 88511 149830 88591
rect 152280 88511 152290 88591
rect 152600 88511 152610 88591
rect 152920 88511 152930 88591
rect 153240 88511 153250 88591
rect 153560 88511 153570 88591
rect 153880 88511 153890 88591
rect 154200 88511 154210 88591
rect 154520 88511 154530 88591
rect 154840 88511 154850 88591
rect 155160 88511 155170 88591
rect 155480 88511 155490 88591
rect 155800 88511 155810 88591
rect 156120 88511 156130 88591
rect 156440 88511 156450 88591
rect 156760 88511 156770 88591
rect 157080 88511 157090 88591
rect 157400 88511 157410 88591
rect 157720 88511 157730 88591
rect 158040 88511 158050 88591
rect 158360 88511 158370 88591
rect 158680 88511 158690 88591
rect 159000 88511 159010 88591
rect 159320 88511 159330 88591
rect 159640 88511 159650 88591
rect 163590 88561 163670 88571
rect 163910 88561 163990 88571
rect 164230 88561 164310 88571
rect 164550 88561 164630 88571
rect 164870 88561 164950 88571
rect 165190 88561 165270 88571
rect 165510 88561 165590 88571
rect 165830 88561 165910 88571
rect 166150 88561 166230 88571
rect 166470 88561 166550 88571
rect 166790 88561 166870 88571
rect 167110 88561 167190 88571
rect 167430 88561 167510 88571
rect 167750 88561 167830 88571
rect 168070 88561 168150 88571
rect 168390 88561 168470 88571
rect 168710 88561 168790 88571
rect 169030 88561 169110 88571
rect 169350 88561 169430 88571
rect 169670 88561 169750 88571
rect 169990 88561 170070 88571
rect 170310 88561 170390 88571
rect 170630 88561 170710 88571
rect 170950 88561 171030 88571
rect 163670 88481 163680 88561
rect 163990 88481 164000 88561
rect 164310 88481 164320 88561
rect 164630 88481 164640 88561
rect 164950 88481 164960 88561
rect 165270 88481 165280 88561
rect 165590 88481 165600 88561
rect 165910 88481 165920 88561
rect 166230 88481 166240 88561
rect 166550 88481 166560 88561
rect 166870 88481 166880 88561
rect 167190 88481 167200 88561
rect 167510 88481 167520 88561
rect 167830 88481 167840 88561
rect 168150 88481 168160 88561
rect 168470 88481 168480 88561
rect 168790 88481 168800 88561
rect 169110 88481 169120 88561
rect 169430 88481 169440 88561
rect 169750 88481 169760 88561
rect 170070 88481 170080 88561
rect 170390 88481 170400 88561
rect 170710 88481 170720 88561
rect 171030 88481 171040 88561
rect 30520 88440 30600 88450
rect 30840 88440 30920 88450
rect 31160 88440 31240 88450
rect 31480 88440 31560 88450
rect 31800 88440 31880 88450
rect 32120 88440 32200 88450
rect 32440 88440 32520 88450
rect 32760 88440 32840 88450
rect 33080 88440 33160 88450
rect 33400 88440 33480 88450
rect 33720 88440 33800 88450
rect 34040 88440 34120 88450
rect 34360 88440 34440 88450
rect 34680 88440 34760 88450
rect 35000 88440 35080 88450
rect 35320 88440 35400 88450
rect 35640 88440 35720 88450
rect 35960 88440 36040 88450
rect 36280 88440 36360 88450
rect 36600 88440 36680 88450
rect 36920 88440 37000 88450
rect 37240 88440 37320 88450
rect 37560 88440 37640 88450
rect 40340 88440 40420 88450
rect 40660 88440 40740 88450
rect 40980 88440 41060 88450
rect 42720 88440 42800 88450
rect 43040 88440 43120 88450
rect 43360 88440 43440 88450
rect 19130 88410 19210 88420
rect 19450 88410 19530 88420
rect 19770 88410 19850 88420
rect 20090 88410 20170 88420
rect 20410 88410 20490 88420
rect 20730 88410 20810 88420
rect 21050 88410 21130 88420
rect 21370 88410 21450 88420
rect 21690 88410 21770 88420
rect 22010 88410 22090 88420
rect 22330 88410 22410 88420
rect 22650 88410 22730 88420
rect 22970 88410 23050 88420
rect 23290 88410 23370 88420
rect 23610 88410 23690 88420
rect 23930 88410 24010 88420
rect 24250 88410 24330 88420
rect 24570 88410 24650 88420
rect 24890 88410 24970 88420
rect 25210 88410 25290 88420
rect 25530 88410 25610 88420
rect 25850 88410 25930 88420
rect 26170 88410 26250 88420
rect 19210 88330 19220 88410
rect 19530 88330 19540 88410
rect 19850 88330 19860 88410
rect 20170 88330 20180 88410
rect 20490 88330 20500 88410
rect 20810 88330 20820 88410
rect 21130 88330 21140 88410
rect 21450 88330 21460 88410
rect 21770 88330 21780 88410
rect 22090 88330 22100 88410
rect 22410 88330 22420 88410
rect 22730 88330 22740 88410
rect 23050 88330 23060 88410
rect 23370 88330 23380 88410
rect 23690 88330 23700 88410
rect 24010 88330 24020 88410
rect 24330 88330 24340 88410
rect 24650 88330 24660 88410
rect 24970 88330 24980 88410
rect 25290 88330 25300 88410
rect 25610 88330 25620 88410
rect 25930 88330 25940 88410
rect 26250 88330 26260 88410
rect 30600 88360 30610 88440
rect 30920 88360 30930 88440
rect 31240 88360 31250 88440
rect 31560 88360 31570 88440
rect 31880 88360 31890 88440
rect 32200 88360 32210 88440
rect 32520 88360 32530 88440
rect 32840 88360 32850 88440
rect 33160 88360 33170 88440
rect 33480 88360 33490 88440
rect 33800 88360 33810 88440
rect 34120 88360 34130 88440
rect 34440 88360 34450 88440
rect 34760 88360 34770 88440
rect 35080 88360 35090 88440
rect 35400 88360 35410 88440
rect 35720 88360 35730 88440
rect 36040 88360 36050 88440
rect 36360 88360 36370 88440
rect 36680 88360 36690 88440
rect 37000 88360 37010 88440
rect 37320 88360 37330 88440
rect 37640 88360 37650 88440
rect 40420 88360 40430 88440
rect 40740 88360 40750 88440
rect 41060 88360 41070 88440
rect 42800 88360 42810 88440
rect 43120 88360 43130 88440
rect 43440 88360 43450 88440
rect 146560 88431 146640 88441
rect 146880 88431 146960 88441
rect 147200 88431 147280 88441
rect 148940 88431 149020 88441
rect 149260 88431 149340 88441
rect 149580 88431 149660 88441
rect 152360 88431 152440 88441
rect 152680 88431 152760 88441
rect 153000 88431 153080 88441
rect 153320 88431 153400 88441
rect 153640 88431 153720 88441
rect 153960 88431 154040 88441
rect 154280 88431 154360 88441
rect 154600 88431 154680 88441
rect 154920 88431 155000 88441
rect 155240 88431 155320 88441
rect 155560 88431 155640 88441
rect 155880 88431 155960 88441
rect 156200 88431 156280 88441
rect 156520 88431 156600 88441
rect 156840 88431 156920 88441
rect 157160 88431 157240 88441
rect 157480 88431 157560 88441
rect 157800 88431 157880 88441
rect 158120 88431 158200 88441
rect 158440 88431 158520 88441
rect 158760 88431 158840 88441
rect 159080 88431 159160 88441
rect 159400 88431 159480 88441
rect 146640 88351 146650 88431
rect 146960 88351 146970 88431
rect 147280 88351 147290 88431
rect 149020 88351 149030 88431
rect 149340 88351 149350 88431
rect 149660 88351 149670 88431
rect 152440 88351 152450 88431
rect 152760 88351 152770 88431
rect 153080 88351 153090 88431
rect 153400 88351 153410 88431
rect 153720 88351 153730 88431
rect 154040 88351 154050 88431
rect 154360 88351 154370 88431
rect 154680 88351 154690 88431
rect 155000 88351 155010 88431
rect 155320 88351 155330 88431
rect 155640 88351 155650 88431
rect 155960 88351 155970 88431
rect 156280 88351 156290 88431
rect 156600 88351 156610 88431
rect 156920 88351 156930 88431
rect 157240 88351 157250 88431
rect 157560 88351 157570 88431
rect 157880 88351 157890 88431
rect 158200 88351 158210 88431
rect 158520 88351 158530 88431
rect 158840 88351 158850 88431
rect 159160 88351 159170 88431
rect 159480 88351 159490 88431
rect 163750 88401 163830 88411
rect 164070 88401 164150 88411
rect 164390 88401 164470 88411
rect 164710 88401 164790 88411
rect 165030 88401 165110 88411
rect 165350 88401 165430 88411
rect 165670 88401 165750 88411
rect 165990 88401 166070 88411
rect 166310 88401 166390 88411
rect 166630 88401 166710 88411
rect 166950 88401 167030 88411
rect 167270 88401 167350 88411
rect 167590 88401 167670 88411
rect 167910 88401 167990 88411
rect 168230 88401 168310 88411
rect 168550 88401 168630 88411
rect 168870 88401 168950 88411
rect 169190 88401 169270 88411
rect 169510 88401 169590 88411
rect 169830 88401 169910 88411
rect 170150 88401 170230 88411
rect 170470 88401 170550 88411
rect 170790 88401 170870 88411
rect 163830 88321 163840 88401
rect 164150 88321 164160 88401
rect 164470 88321 164480 88401
rect 164790 88321 164800 88401
rect 165110 88321 165120 88401
rect 165430 88321 165440 88401
rect 165750 88321 165760 88401
rect 166070 88321 166080 88401
rect 166390 88321 166400 88401
rect 166710 88321 166720 88401
rect 167030 88321 167040 88401
rect 167350 88321 167360 88401
rect 167670 88321 167680 88401
rect 167990 88321 168000 88401
rect 168310 88321 168320 88401
rect 168630 88321 168640 88401
rect 168950 88321 168960 88401
rect 169270 88321 169280 88401
rect 169590 88321 169600 88401
rect 169910 88321 169920 88401
rect 170230 88321 170240 88401
rect 170550 88321 170560 88401
rect 170870 88321 170880 88401
rect 30360 88180 30440 88190
rect 30680 88180 30760 88190
rect 31000 88180 31080 88190
rect 31320 88180 31400 88190
rect 31640 88180 31720 88190
rect 31960 88180 32040 88190
rect 32280 88180 32360 88190
rect 32600 88180 32680 88190
rect 32920 88180 33000 88190
rect 33240 88180 33320 88190
rect 33560 88180 33640 88190
rect 33880 88180 33960 88190
rect 34200 88180 34280 88190
rect 34520 88180 34600 88190
rect 34840 88180 34920 88190
rect 35160 88180 35240 88190
rect 35480 88180 35560 88190
rect 35800 88180 35880 88190
rect 36120 88180 36200 88190
rect 36440 88180 36520 88190
rect 36760 88180 36840 88190
rect 37080 88180 37160 88190
rect 37400 88180 37480 88190
rect 37720 88180 37800 88190
rect 40180 88180 40260 88190
rect 40500 88180 40580 88190
rect 40820 88180 40900 88190
rect 41140 88180 41220 88190
rect 42560 88180 42640 88190
rect 42880 88180 42960 88190
rect 43200 88180 43280 88190
rect 43520 88180 43600 88190
rect 18970 88150 19050 88160
rect 19290 88150 19370 88160
rect 19610 88150 19690 88160
rect 19930 88150 20010 88160
rect 20250 88150 20330 88160
rect 20570 88150 20650 88160
rect 20890 88150 20970 88160
rect 21210 88150 21290 88160
rect 21530 88150 21610 88160
rect 21850 88150 21930 88160
rect 22170 88150 22250 88160
rect 22490 88150 22570 88160
rect 22810 88150 22890 88160
rect 23130 88150 23210 88160
rect 23450 88150 23530 88160
rect 23770 88150 23850 88160
rect 24090 88150 24170 88160
rect 24410 88150 24490 88160
rect 24730 88150 24810 88160
rect 25050 88150 25130 88160
rect 25370 88150 25450 88160
rect 25690 88150 25770 88160
rect 26010 88150 26090 88160
rect 26330 88150 26410 88160
rect 19050 88070 19060 88150
rect 19370 88070 19380 88150
rect 19690 88070 19700 88150
rect 20010 88070 20020 88150
rect 20330 88070 20340 88150
rect 20650 88070 20660 88150
rect 20970 88070 20980 88150
rect 21290 88070 21300 88150
rect 21610 88070 21620 88150
rect 21930 88070 21940 88150
rect 22250 88070 22260 88150
rect 22570 88070 22580 88150
rect 22890 88070 22900 88150
rect 23210 88070 23220 88150
rect 23530 88070 23540 88150
rect 23850 88070 23860 88150
rect 24170 88070 24180 88150
rect 24490 88070 24500 88150
rect 24810 88070 24820 88150
rect 25130 88070 25140 88150
rect 25450 88070 25460 88150
rect 25770 88070 25780 88150
rect 26090 88070 26100 88150
rect 26410 88070 26420 88150
rect 30440 88100 30450 88180
rect 30760 88100 30770 88180
rect 31080 88100 31090 88180
rect 31400 88100 31410 88180
rect 31720 88100 31730 88180
rect 32040 88100 32050 88180
rect 32360 88100 32370 88180
rect 32680 88100 32690 88180
rect 33000 88100 33010 88180
rect 33320 88100 33330 88180
rect 33640 88100 33650 88180
rect 33960 88100 33970 88180
rect 34280 88100 34290 88180
rect 34600 88100 34610 88180
rect 34920 88100 34930 88180
rect 35240 88100 35250 88180
rect 35560 88100 35570 88180
rect 35880 88100 35890 88180
rect 36200 88100 36210 88180
rect 36520 88100 36530 88180
rect 36840 88100 36850 88180
rect 37160 88100 37170 88180
rect 37480 88100 37490 88180
rect 37800 88100 37810 88180
rect 40260 88100 40270 88180
rect 40580 88100 40590 88180
rect 40900 88100 40910 88180
rect 41220 88100 41230 88180
rect 42640 88100 42650 88180
rect 42960 88100 42970 88180
rect 43280 88100 43290 88180
rect 43600 88100 43610 88180
rect 146400 88171 146480 88181
rect 146720 88171 146800 88181
rect 147040 88171 147120 88181
rect 147360 88171 147440 88181
rect 148780 88171 148860 88181
rect 149100 88171 149180 88181
rect 149420 88171 149500 88181
rect 149740 88171 149820 88181
rect 152200 88171 152280 88181
rect 152520 88171 152600 88181
rect 152840 88171 152920 88181
rect 153160 88171 153240 88181
rect 153480 88171 153560 88181
rect 153800 88171 153880 88181
rect 154120 88171 154200 88181
rect 154440 88171 154520 88181
rect 154760 88171 154840 88181
rect 155080 88171 155160 88181
rect 155400 88171 155480 88181
rect 155720 88171 155800 88181
rect 156040 88171 156120 88181
rect 156360 88171 156440 88181
rect 156680 88171 156760 88181
rect 157000 88171 157080 88181
rect 157320 88171 157400 88181
rect 157640 88171 157720 88181
rect 157960 88171 158040 88181
rect 158280 88171 158360 88181
rect 158600 88171 158680 88181
rect 158920 88171 159000 88181
rect 159240 88171 159320 88181
rect 159560 88171 159640 88181
rect 146480 88091 146490 88171
rect 146800 88091 146810 88171
rect 147120 88091 147130 88171
rect 147440 88091 147450 88171
rect 148860 88091 148870 88171
rect 149180 88091 149190 88171
rect 149500 88091 149510 88171
rect 149820 88091 149830 88171
rect 152280 88091 152290 88171
rect 152600 88091 152610 88171
rect 152920 88091 152930 88171
rect 153240 88091 153250 88171
rect 153560 88091 153570 88171
rect 153880 88091 153890 88171
rect 154200 88091 154210 88171
rect 154520 88091 154530 88171
rect 154840 88091 154850 88171
rect 155160 88091 155170 88171
rect 155480 88091 155490 88171
rect 155800 88091 155810 88171
rect 156120 88091 156130 88171
rect 156440 88091 156450 88171
rect 156760 88091 156770 88171
rect 157080 88091 157090 88171
rect 157400 88091 157410 88171
rect 157720 88091 157730 88171
rect 158040 88091 158050 88171
rect 158360 88091 158370 88171
rect 158680 88091 158690 88171
rect 159000 88091 159010 88171
rect 159320 88091 159330 88171
rect 159640 88091 159650 88171
rect 163590 88141 163670 88151
rect 163910 88141 163990 88151
rect 164230 88141 164310 88151
rect 164550 88141 164630 88151
rect 164870 88141 164950 88151
rect 165190 88141 165270 88151
rect 165510 88141 165590 88151
rect 165830 88141 165910 88151
rect 166150 88141 166230 88151
rect 166470 88141 166550 88151
rect 166790 88141 166870 88151
rect 167110 88141 167190 88151
rect 167430 88141 167510 88151
rect 167750 88141 167830 88151
rect 168070 88141 168150 88151
rect 168390 88141 168470 88151
rect 168710 88141 168790 88151
rect 169030 88141 169110 88151
rect 169350 88141 169430 88151
rect 169670 88141 169750 88151
rect 169990 88141 170070 88151
rect 170310 88141 170390 88151
rect 170630 88141 170710 88151
rect 170950 88141 171030 88151
rect 163670 88061 163680 88141
rect 163990 88061 164000 88141
rect 164310 88061 164320 88141
rect 164630 88061 164640 88141
rect 164950 88061 164960 88141
rect 165270 88061 165280 88141
rect 165590 88061 165600 88141
rect 165910 88061 165920 88141
rect 166230 88061 166240 88141
rect 166550 88061 166560 88141
rect 166870 88061 166880 88141
rect 167190 88061 167200 88141
rect 167510 88061 167520 88141
rect 167830 88061 167840 88141
rect 168150 88061 168160 88141
rect 168470 88061 168480 88141
rect 168790 88061 168800 88141
rect 169110 88061 169120 88141
rect 169430 88061 169440 88141
rect 169750 88061 169760 88141
rect 170070 88061 170080 88141
rect 170390 88061 170400 88141
rect 170710 88061 170720 88141
rect 171030 88061 171040 88141
rect 30520 88020 30600 88030
rect 30840 88020 30920 88030
rect 31160 88020 31240 88030
rect 31480 88020 31560 88030
rect 31800 88020 31880 88030
rect 32120 88020 32200 88030
rect 32440 88020 32520 88030
rect 32760 88020 32840 88030
rect 33080 88020 33160 88030
rect 33400 88020 33480 88030
rect 33720 88020 33800 88030
rect 34040 88020 34120 88030
rect 34360 88020 34440 88030
rect 34680 88020 34760 88030
rect 35000 88020 35080 88030
rect 35320 88020 35400 88030
rect 35640 88020 35720 88030
rect 35960 88020 36040 88030
rect 36280 88020 36360 88030
rect 36600 88020 36680 88030
rect 36920 88020 37000 88030
rect 37240 88020 37320 88030
rect 37560 88020 37640 88030
rect 40340 88020 40420 88030
rect 40660 88020 40740 88030
rect 40980 88020 41060 88030
rect 42720 88020 42800 88030
rect 43040 88020 43120 88030
rect 43360 88020 43440 88030
rect 19130 87990 19210 88000
rect 19450 87990 19530 88000
rect 19770 87990 19850 88000
rect 20090 87990 20170 88000
rect 20410 87990 20490 88000
rect 20730 87990 20810 88000
rect 21050 87990 21130 88000
rect 21370 87990 21450 88000
rect 21690 87990 21770 88000
rect 22010 87990 22090 88000
rect 22330 87990 22410 88000
rect 22650 87990 22730 88000
rect 22970 87990 23050 88000
rect 23290 87990 23370 88000
rect 23610 87990 23690 88000
rect 23930 87990 24010 88000
rect 24250 87990 24330 88000
rect 24570 87990 24650 88000
rect 24890 87990 24970 88000
rect 25210 87990 25290 88000
rect 25530 87990 25610 88000
rect 25850 87990 25930 88000
rect 26170 87990 26250 88000
rect 19210 87910 19220 87990
rect 19530 87910 19540 87990
rect 19850 87910 19860 87990
rect 20170 87910 20180 87990
rect 20490 87910 20500 87990
rect 20810 87910 20820 87990
rect 21130 87910 21140 87990
rect 21450 87910 21460 87990
rect 21770 87910 21780 87990
rect 22090 87910 22100 87990
rect 22410 87910 22420 87990
rect 22730 87910 22740 87990
rect 23050 87910 23060 87990
rect 23370 87910 23380 87990
rect 23690 87910 23700 87990
rect 24010 87910 24020 87990
rect 24330 87910 24340 87990
rect 24650 87910 24660 87990
rect 24970 87910 24980 87990
rect 25290 87910 25300 87990
rect 25610 87910 25620 87990
rect 25930 87910 25940 87990
rect 26250 87910 26260 87990
rect 30600 87940 30610 88020
rect 30920 87940 30930 88020
rect 31240 87940 31250 88020
rect 31560 87940 31570 88020
rect 31880 87940 31890 88020
rect 32200 87940 32210 88020
rect 32520 87940 32530 88020
rect 32840 87940 32850 88020
rect 33160 87940 33170 88020
rect 33480 87940 33490 88020
rect 33800 87940 33810 88020
rect 34120 87940 34130 88020
rect 34440 87940 34450 88020
rect 34760 87940 34770 88020
rect 35080 87940 35090 88020
rect 35400 87940 35410 88020
rect 35720 87940 35730 88020
rect 36040 87940 36050 88020
rect 36360 87940 36370 88020
rect 36680 87940 36690 88020
rect 37000 87940 37010 88020
rect 37320 87940 37330 88020
rect 37640 87940 37650 88020
rect 40420 87940 40430 88020
rect 40740 87940 40750 88020
rect 41060 87940 41070 88020
rect 42800 87940 42810 88020
rect 43120 87940 43130 88020
rect 43440 87940 43450 88020
rect 146560 88011 146640 88021
rect 146880 88011 146960 88021
rect 147200 88011 147280 88021
rect 148940 88011 149020 88021
rect 149260 88011 149340 88021
rect 149580 88011 149660 88021
rect 152360 88011 152440 88021
rect 152680 88011 152760 88021
rect 153000 88011 153080 88021
rect 153320 88011 153400 88021
rect 153640 88011 153720 88021
rect 153960 88011 154040 88021
rect 154280 88011 154360 88021
rect 154600 88011 154680 88021
rect 154920 88011 155000 88021
rect 155240 88011 155320 88021
rect 155560 88011 155640 88021
rect 155880 88011 155960 88021
rect 156200 88011 156280 88021
rect 156520 88011 156600 88021
rect 156840 88011 156920 88021
rect 157160 88011 157240 88021
rect 157480 88011 157560 88021
rect 157800 88011 157880 88021
rect 158120 88011 158200 88021
rect 158440 88011 158520 88021
rect 158760 88011 158840 88021
rect 159080 88011 159160 88021
rect 159400 88011 159480 88021
rect 146640 87931 146650 88011
rect 146960 87931 146970 88011
rect 147280 87931 147290 88011
rect 149020 87931 149030 88011
rect 149340 87931 149350 88011
rect 149660 87931 149670 88011
rect 152440 87931 152450 88011
rect 152760 87931 152770 88011
rect 153080 87931 153090 88011
rect 153400 87931 153410 88011
rect 153720 87931 153730 88011
rect 154040 87931 154050 88011
rect 154360 87931 154370 88011
rect 154680 87931 154690 88011
rect 155000 87931 155010 88011
rect 155320 87931 155330 88011
rect 155640 87931 155650 88011
rect 155960 87931 155970 88011
rect 156280 87931 156290 88011
rect 156600 87931 156610 88011
rect 156920 87931 156930 88011
rect 157240 87931 157250 88011
rect 157560 87931 157570 88011
rect 157880 87931 157890 88011
rect 158200 87931 158210 88011
rect 158520 87931 158530 88011
rect 158840 87931 158850 88011
rect 159160 87931 159170 88011
rect 159480 87931 159490 88011
rect 163750 87981 163830 87991
rect 164070 87981 164150 87991
rect 164390 87981 164470 87991
rect 164710 87981 164790 87991
rect 165030 87981 165110 87991
rect 165350 87981 165430 87991
rect 165670 87981 165750 87991
rect 165990 87981 166070 87991
rect 166310 87981 166390 87991
rect 166630 87981 166710 87991
rect 166950 87981 167030 87991
rect 167270 87981 167350 87991
rect 167590 87981 167670 87991
rect 167910 87981 167990 87991
rect 168230 87981 168310 87991
rect 168550 87981 168630 87991
rect 168870 87981 168950 87991
rect 169190 87981 169270 87991
rect 169510 87981 169590 87991
rect 169830 87981 169910 87991
rect 170150 87981 170230 87991
rect 170470 87981 170550 87991
rect 170790 87981 170870 87991
rect 163830 87901 163840 87981
rect 164150 87901 164160 87981
rect 164470 87901 164480 87981
rect 164790 87901 164800 87981
rect 165110 87901 165120 87981
rect 165430 87901 165440 87981
rect 165750 87901 165760 87981
rect 166070 87901 166080 87981
rect 166390 87901 166400 87981
rect 166710 87901 166720 87981
rect 167030 87901 167040 87981
rect 167350 87901 167360 87981
rect 167670 87901 167680 87981
rect 167990 87901 168000 87981
rect 168310 87901 168320 87981
rect 168630 87901 168640 87981
rect 168950 87901 168960 87981
rect 169270 87901 169280 87981
rect 169590 87901 169600 87981
rect 169910 87901 169920 87981
rect 170230 87901 170240 87981
rect 170550 87901 170560 87981
rect 170870 87901 170880 87981
rect 30360 87860 30440 87870
rect 30680 87860 30760 87870
rect 31000 87860 31080 87870
rect 31320 87860 31400 87870
rect 31640 87860 31720 87870
rect 31960 87860 32040 87870
rect 32280 87860 32360 87870
rect 32600 87860 32680 87870
rect 32920 87860 33000 87870
rect 33240 87860 33320 87870
rect 33560 87860 33640 87870
rect 33880 87860 33960 87870
rect 34200 87860 34280 87870
rect 34520 87860 34600 87870
rect 34840 87860 34920 87870
rect 35160 87860 35240 87870
rect 35480 87860 35560 87870
rect 35800 87860 35880 87870
rect 36120 87860 36200 87870
rect 36440 87860 36520 87870
rect 36760 87860 36840 87870
rect 37080 87860 37160 87870
rect 37400 87860 37480 87870
rect 37720 87860 37800 87870
rect 40180 87860 40260 87870
rect 40500 87860 40580 87870
rect 40820 87860 40900 87870
rect 41140 87860 41220 87870
rect 42560 87860 42640 87870
rect 42880 87860 42960 87870
rect 43200 87860 43280 87870
rect 43520 87860 43600 87870
rect 18970 87830 19050 87840
rect 19290 87830 19370 87840
rect 19610 87830 19690 87840
rect 19930 87830 20010 87840
rect 20250 87830 20330 87840
rect 20570 87830 20650 87840
rect 20890 87830 20970 87840
rect 21210 87830 21290 87840
rect 21530 87830 21610 87840
rect 21850 87830 21930 87840
rect 22170 87830 22250 87840
rect 22490 87830 22570 87840
rect 22810 87830 22890 87840
rect 23130 87830 23210 87840
rect 23450 87830 23530 87840
rect 23770 87830 23850 87840
rect 24090 87830 24170 87840
rect 24410 87830 24490 87840
rect 24730 87830 24810 87840
rect 25050 87830 25130 87840
rect 25370 87830 25450 87840
rect 25690 87830 25770 87840
rect 26010 87830 26090 87840
rect 26330 87830 26410 87840
rect 19050 87750 19060 87830
rect 19370 87750 19380 87830
rect 19690 87750 19700 87830
rect 20010 87750 20020 87830
rect 20330 87750 20340 87830
rect 20650 87750 20660 87830
rect 20970 87750 20980 87830
rect 21290 87750 21300 87830
rect 21610 87750 21620 87830
rect 21930 87750 21940 87830
rect 22250 87750 22260 87830
rect 22570 87750 22580 87830
rect 22890 87750 22900 87830
rect 23210 87750 23220 87830
rect 23530 87750 23540 87830
rect 23850 87750 23860 87830
rect 24170 87750 24180 87830
rect 24490 87750 24500 87830
rect 24810 87750 24820 87830
rect 25130 87750 25140 87830
rect 25450 87750 25460 87830
rect 25770 87750 25780 87830
rect 26090 87750 26100 87830
rect 26410 87750 26420 87830
rect 30440 87780 30450 87860
rect 30760 87780 30770 87860
rect 31080 87780 31090 87860
rect 31400 87780 31410 87860
rect 31720 87780 31730 87860
rect 32040 87780 32050 87860
rect 32360 87780 32370 87860
rect 32680 87780 32690 87860
rect 33000 87780 33010 87860
rect 33320 87780 33330 87860
rect 33640 87780 33650 87860
rect 33960 87780 33970 87860
rect 34280 87780 34290 87860
rect 34600 87780 34610 87860
rect 34920 87780 34930 87860
rect 35240 87780 35250 87860
rect 35560 87780 35570 87860
rect 35880 87780 35890 87860
rect 36200 87780 36210 87860
rect 36520 87780 36530 87860
rect 36840 87780 36850 87860
rect 37160 87780 37170 87860
rect 37480 87780 37490 87860
rect 37800 87780 37810 87860
rect 40260 87780 40270 87860
rect 40580 87780 40590 87860
rect 40900 87780 40910 87860
rect 41220 87780 41230 87860
rect 42640 87780 42650 87860
rect 42960 87780 42970 87860
rect 43280 87780 43290 87860
rect 43600 87780 43610 87860
rect 146400 87851 146480 87861
rect 146720 87851 146800 87861
rect 147040 87851 147120 87861
rect 147360 87851 147440 87861
rect 148780 87851 148860 87861
rect 149100 87851 149180 87861
rect 149420 87851 149500 87861
rect 149740 87851 149820 87861
rect 152200 87851 152280 87861
rect 152520 87851 152600 87861
rect 152840 87851 152920 87861
rect 153160 87851 153240 87861
rect 153480 87851 153560 87861
rect 153800 87851 153880 87861
rect 154120 87851 154200 87861
rect 154440 87851 154520 87861
rect 154760 87851 154840 87861
rect 155080 87851 155160 87861
rect 155400 87851 155480 87861
rect 155720 87851 155800 87861
rect 156040 87851 156120 87861
rect 156360 87851 156440 87861
rect 156680 87851 156760 87861
rect 157000 87851 157080 87861
rect 157320 87851 157400 87861
rect 157640 87851 157720 87861
rect 157960 87851 158040 87861
rect 158280 87851 158360 87861
rect 158600 87851 158680 87861
rect 158920 87851 159000 87861
rect 159240 87851 159320 87861
rect 159560 87851 159640 87861
rect 146480 87771 146490 87851
rect 146800 87771 146810 87851
rect 147120 87771 147130 87851
rect 147440 87771 147450 87851
rect 148860 87771 148870 87851
rect 149180 87771 149190 87851
rect 149500 87771 149510 87851
rect 149820 87771 149830 87851
rect 152280 87771 152290 87851
rect 152600 87771 152610 87851
rect 152920 87771 152930 87851
rect 153240 87771 153250 87851
rect 153560 87771 153570 87851
rect 153880 87771 153890 87851
rect 154200 87771 154210 87851
rect 154520 87771 154530 87851
rect 154840 87771 154850 87851
rect 155160 87771 155170 87851
rect 155480 87771 155490 87851
rect 155800 87771 155810 87851
rect 156120 87771 156130 87851
rect 156440 87771 156450 87851
rect 156760 87771 156770 87851
rect 157080 87771 157090 87851
rect 157400 87771 157410 87851
rect 157720 87771 157730 87851
rect 158040 87771 158050 87851
rect 158360 87771 158370 87851
rect 158680 87771 158690 87851
rect 159000 87771 159010 87851
rect 159320 87771 159330 87851
rect 159640 87771 159650 87851
rect 163590 87821 163670 87831
rect 163910 87821 163990 87831
rect 164230 87821 164310 87831
rect 164550 87821 164630 87831
rect 164870 87821 164950 87831
rect 165190 87821 165270 87831
rect 165510 87821 165590 87831
rect 165830 87821 165910 87831
rect 166150 87821 166230 87831
rect 166470 87821 166550 87831
rect 166790 87821 166870 87831
rect 167110 87821 167190 87831
rect 167430 87821 167510 87831
rect 167750 87821 167830 87831
rect 168070 87821 168150 87831
rect 168390 87821 168470 87831
rect 168710 87821 168790 87831
rect 169030 87821 169110 87831
rect 169350 87821 169430 87831
rect 169670 87821 169750 87831
rect 169990 87821 170070 87831
rect 170310 87821 170390 87831
rect 170630 87821 170710 87831
rect 170950 87821 171030 87831
rect 163670 87741 163680 87821
rect 163990 87741 164000 87821
rect 164310 87741 164320 87821
rect 164630 87741 164640 87821
rect 164950 87741 164960 87821
rect 165270 87741 165280 87821
rect 165590 87741 165600 87821
rect 165910 87741 165920 87821
rect 166230 87741 166240 87821
rect 166550 87741 166560 87821
rect 166870 87741 166880 87821
rect 167190 87741 167200 87821
rect 167510 87741 167520 87821
rect 167830 87741 167840 87821
rect 168150 87741 168160 87821
rect 168470 87741 168480 87821
rect 168790 87741 168800 87821
rect 169110 87741 169120 87821
rect 169430 87741 169440 87821
rect 169750 87741 169760 87821
rect 170070 87741 170080 87821
rect 170390 87741 170400 87821
rect 170710 87741 170720 87821
rect 171030 87741 171040 87821
rect 30520 87700 30600 87710
rect 30840 87700 30920 87710
rect 31160 87700 31240 87710
rect 31480 87700 31560 87710
rect 31800 87700 31880 87710
rect 32120 87700 32200 87710
rect 32440 87700 32520 87710
rect 32760 87700 32840 87710
rect 33080 87700 33160 87710
rect 33400 87700 33480 87710
rect 33720 87700 33800 87710
rect 34040 87700 34120 87710
rect 34360 87700 34440 87710
rect 34680 87700 34760 87710
rect 35000 87700 35080 87710
rect 35320 87700 35400 87710
rect 35640 87700 35720 87710
rect 35960 87700 36040 87710
rect 36280 87700 36360 87710
rect 36600 87700 36680 87710
rect 36920 87700 37000 87710
rect 37240 87700 37320 87710
rect 37560 87700 37640 87710
rect 40340 87700 40420 87710
rect 40660 87700 40740 87710
rect 40980 87700 41060 87710
rect 42720 87700 42800 87710
rect 43040 87700 43120 87710
rect 43360 87700 43440 87710
rect 19130 87670 19210 87680
rect 19450 87670 19530 87680
rect 19770 87670 19850 87680
rect 20090 87670 20170 87680
rect 20410 87670 20490 87680
rect 20730 87670 20810 87680
rect 21050 87670 21130 87680
rect 21370 87670 21450 87680
rect 21690 87670 21770 87680
rect 22010 87670 22090 87680
rect 22330 87670 22410 87680
rect 22650 87670 22730 87680
rect 22970 87670 23050 87680
rect 23290 87670 23370 87680
rect 23610 87670 23690 87680
rect 23930 87670 24010 87680
rect 24250 87670 24330 87680
rect 24570 87670 24650 87680
rect 24890 87670 24970 87680
rect 25210 87670 25290 87680
rect 25530 87670 25610 87680
rect 25850 87670 25930 87680
rect 26170 87670 26250 87680
rect 19210 87590 19220 87670
rect 19530 87590 19540 87670
rect 19850 87590 19860 87670
rect 20170 87590 20180 87670
rect 20490 87590 20500 87670
rect 20810 87590 20820 87670
rect 21130 87590 21140 87670
rect 21450 87590 21460 87670
rect 21770 87590 21780 87670
rect 22090 87590 22100 87670
rect 22410 87590 22420 87670
rect 22730 87590 22740 87670
rect 23050 87590 23060 87670
rect 23370 87590 23380 87670
rect 23690 87590 23700 87670
rect 24010 87590 24020 87670
rect 24330 87590 24340 87670
rect 24650 87590 24660 87670
rect 24970 87590 24980 87670
rect 25290 87590 25300 87670
rect 25610 87590 25620 87670
rect 25930 87590 25940 87670
rect 26250 87590 26260 87670
rect 30600 87620 30610 87700
rect 30920 87620 30930 87700
rect 31240 87620 31250 87700
rect 31560 87620 31570 87700
rect 31880 87620 31890 87700
rect 32200 87620 32210 87700
rect 32520 87620 32530 87700
rect 32840 87620 32850 87700
rect 33160 87620 33170 87700
rect 33480 87620 33490 87700
rect 33800 87620 33810 87700
rect 34120 87620 34130 87700
rect 34440 87620 34450 87700
rect 34760 87620 34770 87700
rect 35080 87620 35090 87700
rect 35400 87620 35410 87700
rect 35720 87620 35730 87700
rect 36040 87620 36050 87700
rect 36360 87620 36370 87700
rect 36680 87620 36690 87700
rect 37000 87620 37010 87700
rect 37320 87620 37330 87700
rect 37640 87620 37650 87700
rect 40420 87620 40430 87700
rect 40740 87620 40750 87700
rect 41060 87620 41070 87700
rect 42800 87620 42810 87700
rect 43120 87620 43130 87700
rect 43440 87620 43450 87700
rect 146560 87691 146640 87701
rect 146880 87691 146960 87701
rect 147200 87691 147280 87701
rect 148940 87691 149020 87701
rect 149260 87691 149340 87701
rect 149580 87691 149660 87701
rect 152360 87691 152440 87701
rect 152680 87691 152760 87701
rect 153000 87691 153080 87701
rect 153320 87691 153400 87701
rect 153640 87691 153720 87701
rect 153960 87691 154040 87701
rect 154280 87691 154360 87701
rect 154600 87691 154680 87701
rect 154920 87691 155000 87701
rect 155240 87691 155320 87701
rect 155560 87691 155640 87701
rect 155880 87691 155960 87701
rect 156200 87691 156280 87701
rect 156520 87691 156600 87701
rect 156840 87691 156920 87701
rect 157160 87691 157240 87701
rect 157480 87691 157560 87701
rect 157800 87691 157880 87701
rect 158120 87691 158200 87701
rect 158440 87691 158520 87701
rect 158760 87691 158840 87701
rect 159080 87691 159160 87701
rect 159400 87691 159480 87701
rect 146640 87611 146650 87691
rect 146960 87611 146970 87691
rect 147280 87611 147290 87691
rect 149020 87611 149030 87691
rect 149340 87611 149350 87691
rect 149660 87611 149670 87691
rect 152440 87611 152450 87691
rect 152760 87611 152770 87691
rect 153080 87611 153090 87691
rect 153400 87611 153410 87691
rect 153720 87611 153730 87691
rect 154040 87611 154050 87691
rect 154360 87611 154370 87691
rect 154680 87611 154690 87691
rect 155000 87611 155010 87691
rect 155320 87611 155330 87691
rect 155640 87611 155650 87691
rect 155960 87611 155970 87691
rect 156280 87611 156290 87691
rect 156600 87611 156610 87691
rect 156920 87611 156930 87691
rect 157240 87611 157250 87691
rect 157560 87611 157570 87691
rect 157880 87611 157890 87691
rect 158200 87611 158210 87691
rect 158520 87611 158530 87691
rect 158840 87611 158850 87691
rect 159160 87611 159170 87691
rect 159480 87611 159490 87691
rect 163750 87661 163830 87671
rect 164070 87661 164150 87671
rect 164390 87661 164470 87671
rect 164710 87661 164790 87671
rect 165030 87661 165110 87671
rect 165350 87661 165430 87671
rect 165670 87661 165750 87671
rect 165990 87661 166070 87671
rect 166310 87661 166390 87671
rect 166630 87661 166710 87671
rect 166950 87661 167030 87671
rect 167270 87661 167350 87671
rect 167590 87661 167670 87671
rect 167910 87661 167990 87671
rect 168230 87661 168310 87671
rect 168550 87661 168630 87671
rect 168870 87661 168950 87671
rect 169190 87661 169270 87671
rect 169510 87661 169590 87671
rect 169830 87661 169910 87671
rect 170150 87661 170230 87671
rect 170470 87661 170550 87671
rect 170790 87661 170870 87671
rect 163830 87581 163840 87661
rect 164150 87581 164160 87661
rect 164470 87581 164480 87661
rect 164790 87581 164800 87661
rect 165110 87581 165120 87661
rect 165430 87581 165440 87661
rect 165750 87581 165760 87661
rect 166070 87581 166080 87661
rect 166390 87581 166400 87661
rect 166710 87581 166720 87661
rect 167030 87581 167040 87661
rect 167350 87581 167360 87661
rect 167670 87581 167680 87661
rect 167990 87581 168000 87661
rect 168310 87581 168320 87661
rect 168630 87581 168640 87661
rect 168950 87581 168960 87661
rect 169270 87581 169280 87661
rect 169590 87581 169600 87661
rect 169910 87581 169920 87661
rect 170230 87581 170240 87661
rect 170550 87581 170560 87661
rect 170870 87581 170880 87661
rect 18980 87440 19060 87450
rect 19160 87440 19240 87450
rect 19340 87440 19420 87450
rect 19520 87440 19600 87450
rect 19700 87440 19780 87450
rect 19880 87440 19960 87450
rect 20060 87440 20140 87450
rect 20240 87440 20320 87450
rect 20420 87440 20500 87450
rect 20600 87440 20680 87450
rect 20780 87440 20860 87450
rect 20960 87440 21040 87450
rect 21140 87440 21220 87450
rect 21320 87440 21400 87450
rect 21500 87440 21580 87450
rect 21680 87440 21760 87450
rect 21860 87440 21940 87450
rect 22040 87440 22120 87450
rect 22220 87440 22300 87450
rect 22400 87440 22480 87450
rect 22580 87440 22660 87450
rect 22760 87440 22840 87450
rect 22940 87440 23020 87450
rect 23120 87440 23200 87450
rect 23300 87440 23380 87450
rect 23480 87440 23560 87450
rect 23660 87440 23740 87450
rect 23840 87440 23920 87450
rect 24020 87440 24100 87450
rect 24200 87440 24280 87450
rect 24380 87440 24460 87450
rect 24560 87440 24640 87450
rect 24740 87440 24820 87450
rect 24920 87440 25000 87450
rect 25100 87440 25180 87450
rect 25280 87440 25360 87450
rect 25460 87440 25540 87450
rect 25640 87440 25720 87450
rect 25820 87440 25900 87450
rect 26000 87440 26080 87450
rect 26180 87440 26260 87450
rect 26360 87440 26440 87450
rect 26540 87440 26620 87450
rect 146300 87440 146380 87450
rect 146440 87440 146520 87450
rect 146580 87440 146660 87450
rect 146720 87440 146800 87450
rect 146860 87440 146940 87450
rect 147000 87440 147080 87450
rect 147140 87440 147220 87450
rect 147280 87440 147360 87450
rect 147420 87440 147500 87450
rect 147560 87440 147640 87450
rect 148600 87440 148680 87450
rect 148740 87440 148820 87450
rect 148880 87440 148960 87450
rect 149020 87440 149100 87450
rect 149160 87440 149240 87450
rect 149300 87440 149380 87450
rect 149440 87440 149520 87450
rect 149580 87440 149660 87450
rect 149720 87440 149800 87450
rect 149860 87440 149940 87450
rect 152080 87440 152160 87450
rect 152260 87440 152340 87450
rect 152440 87440 152520 87450
rect 152620 87440 152700 87450
rect 152800 87440 152880 87450
rect 152980 87440 153060 87450
rect 153160 87440 153240 87450
rect 153340 87440 153420 87450
rect 153520 87440 153600 87450
rect 153700 87440 153780 87450
rect 153880 87440 153960 87450
rect 154060 87440 154140 87450
rect 154240 87440 154320 87450
rect 154420 87440 154500 87450
rect 154600 87440 154680 87450
rect 154780 87440 154860 87450
rect 154960 87440 155040 87450
rect 155140 87440 155220 87450
rect 155320 87440 155400 87450
rect 155500 87440 155580 87450
rect 155680 87440 155760 87450
rect 155860 87440 155940 87450
rect 156040 87440 156120 87450
rect 156220 87440 156300 87450
rect 156400 87440 156480 87450
rect 156580 87440 156660 87450
rect 156760 87440 156840 87450
rect 156940 87440 157020 87450
rect 157120 87440 157200 87450
rect 157300 87440 157380 87450
rect 157480 87440 157560 87450
rect 157660 87440 157740 87450
rect 157840 87440 157920 87450
rect 158020 87440 158100 87450
rect 158200 87440 158280 87450
rect 158380 87440 158460 87450
rect 158560 87440 158640 87450
rect 158740 87440 158820 87450
rect 158920 87440 159000 87450
rect 159100 87440 159180 87450
rect 159280 87440 159360 87450
rect 159460 87440 159540 87450
rect 159640 87440 159720 87450
rect 163380 87440 163460 87450
rect 163560 87440 163640 87450
rect 163740 87440 163820 87450
rect 163920 87440 164000 87450
rect 164100 87440 164180 87450
rect 164280 87440 164360 87450
rect 164460 87440 164540 87450
rect 164640 87440 164720 87450
rect 164820 87440 164900 87450
rect 165000 87440 165080 87450
rect 165180 87440 165260 87450
rect 165360 87440 165440 87450
rect 165540 87440 165620 87450
rect 165720 87440 165800 87450
rect 165900 87440 165980 87450
rect 166080 87440 166160 87450
rect 166260 87440 166340 87450
rect 166440 87440 166520 87450
rect 166620 87440 166700 87450
rect 166800 87440 166880 87450
rect 166980 87440 167060 87450
rect 167160 87440 167240 87450
rect 167340 87440 167420 87450
rect 167520 87440 167600 87450
rect 167700 87440 167780 87450
rect 167880 87440 167960 87450
rect 168060 87440 168140 87450
rect 168240 87440 168320 87450
rect 168420 87440 168500 87450
rect 168600 87440 168680 87450
rect 168780 87440 168860 87450
rect 168960 87440 169040 87450
rect 169140 87440 169220 87450
rect 169320 87440 169400 87450
rect 169500 87440 169580 87450
rect 169680 87440 169760 87450
rect 169860 87440 169940 87450
rect 170040 87440 170120 87450
rect 170220 87440 170300 87450
rect 170400 87440 170480 87450
rect 170580 87440 170660 87450
rect 170760 87440 170840 87450
rect 170940 87440 171020 87450
rect 19060 87360 19070 87440
rect 19240 87360 19250 87440
rect 19420 87360 19430 87440
rect 19600 87360 19610 87440
rect 19780 87360 19790 87440
rect 19960 87360 19970 87440
rect 20140 87360 20150 87440
rect 20320 87360 20330 87440
rect 20500 87360 20510 87440
rect 20680 87360 20690 87440
rect 20860 87360 20870 87440
rect 21040 87360 21050 87440
rect 21220 87360 21230 87440
rect 21400 87360 21410 87440
rect 21580 87360 21590 87440
rect 21760 87360 21770 87440
rect 21940 87360 21950 87440
rect 22120 87360 22130 87440
rect 22300 87360 22310 87440
rect 22480 87360 22490 87440
rect 22660 87360 22670 87440
rect 22840 87360 22850 87440
rect 23020 87360 23030 87440
rect 23200 87360 23210 87440
rect 23380 87360 23390 87440
rect 23560 87360 23570 87440
rect 23740 87360 23750 87440
rect 23920 87360 23930 87440
rect 24100 87360 24110 87440
rect 24280 87360 24290 87440
rect 24460 87360 24470 87440
rect 24640 87360 24650 87440
rect 24820 87360 24830 87440
rect 25000 87360 25010 87440
rect 25180 87360 25190 87440
rect 25360 87360 25370 87440
rect 25540 87360 25550 87440
rect 25720 87360 25730 87440
rect 25900 87360 25910 87440
rect 26080 87360 26090 87440
rect 26260 87360 26270 87440
rect 26440 87360 26450 87440
rect 26620 87360 26630 87440
rect 146380 87360 146390 87440
rect 146520 87360 146530 87440
rect 146660 87360 146670 87440
rect 146800 87360 146810 87440
rect 146940 87360 146950 87440
rect 147080 87360 147090 87440
rect 147220 87360 147230 87440
rect 147360 87360 147370 87440
rect 147500 87360 147510 87440
rect 147640 87360 147650 87440
rect 148680 87360 148690 87440
rect 148820 87360 148830 87440
rect 148960 87360 148970 87440
rect 149100 87360 149110 87440
rect 149240 87360 149250 87440
rect 149380 87360 149390 87440
rect 149520 87360 149530 87440
rect 149660 87360 149670 87440
rect 149800 87360 149810 87440
rect 149940 87360 149950 87440
rect 152160 87360 152170 87440
rect 152340 87360 152350 87440
rect 152520 87360 152530 87440
rect 152700 87360 152710 87440
rect 152880 87360 152890 87440
rect 153060 87360 153070 87440
rect 153240 87360 153250 87440
rect 153420 87360 153430 87440
rect 153600 87360 153610 87440
rect 153780 87360 153790 87440
rect 153960 87360 153970 87440
rect 154140 87360 154150 87440
rect 154320 87360 154330 87440
rect 154500 87360 154510 87440
rect 154680 87360 154690 87440
rect 154860 87360 154870 87440
rect 155040 87360 155050 87440
rect 155220 87360 155230 87440
rect 155400 87360 155410 87440
rect 155580 87360 155590 87440
rect 155760 87360 155770 87440
rect 155940 87360 155950 87440
rect 156120 87360 156130 87440
rect 156300 87360 156310 87440
rect 156480 87360 156490 87440
rect 156660 87360 156670 87440
rect 156840 87360 156850 87440
rect 157020 87360 157030 87440
rect 157200 87360 157210 87440
rect 157380 87360 157390 87440
rect 157560 87360 157570 87440
rect 157740 87360 157750 87440
rect 157920 87360 157930 87440
rect 158100 87360 158110 87440
rect 158280 87360 158290 87440
rect 158460 87360 158470 87440
rect 158640 87360 158650 87440
rect 158820 87360 158830 87440
rect 159000 87360 159010 87440
rect 159180 87360 159190 87440
rect 159360 87360 159370 87440
rect 159540 87360 159550 87440
rect 159720 87360 159730 87440
rect 163460 87360 163470 87440
rect 163640 87360 163650 87440
rect 163820 87360 163830 87440
rect 164000 87360 164010 87440
rect 164180 87360 164190 87440
rect 164360 87360 164370 87440
rect 164540 87360 164550 87440
rect 164720 87360 164730 87440
rect 164900 87360 164910 87440
rect 165080 87360 165090 87440
rect 165260 87360 165270 87440
rect 165440 87360 165450 87440
rect 165620 87360 165630 87440
rect 165800 87360 165810 87440
rect 165980 87360 165990 87440
rect 166160 87360 166170 87440
rect 166340 87360 166350 87440
rect 166520 87360 166530 87440
rect 166700 87360 166710 87440
rect 166880 87360 166890 87440
rect 167060 87360 167070 87440
rect 167240 87360 167250 87440
rect 167420 87360 167430 87440
rect 167600 87360 167610 87440
rect 167780 87360 167790 87440
rect 167960 87360 167970 87440
rect 168140 87360 168150 87440
rect 168320 87360 168330 87440
rect 168500 87360 168510 87440
rect 168680 87360 168690 87440
rect 168860 87360 168870 87440
rect 169040 87360 169050 87440
rect 169220 87360 169230 87440
rect 169400 87360 169410 87440
rect 169580 87360 169590 87440
rect 169760 87360 169770 87440
rect 169940 87360 169950 87440
rect 170120 87360 170130 87440
rect 170300 87360 170310 87440
rect 170480 87360 170490 87440
rect 170660 87360 170670 87440
rect 170840 87360 170850 87440
rect 171020 87360 171030 87440
rect 161885 87345 161965 87355
rect 162065 87345 162145 87355
rect 162245 87345 162325 87355
rect 162425 87345 162505 87355
rect 162605 87345 162685 87355
rect 18980 87290 19060 87300
rect 19160 87290 19240 87300
rect 19340 87290 19420 87300
rect 19520 87290 19600 87300
rect 19700 87290 19780 87300
rect 19880 87290 19960 87300
rect 20060 87290 20140 87300
rect 20240 87290 20320 87300
rect 20420 87290 20500 87300
rect 20600 87290 20680 87300
rect 20780 87290 20860 87300
rect 20960 87290 21040 87300
rect 21140 87290 21220 87300
rect 21320 87290 21400 87300
rect 21500 87290 21580 87300
rect 21680 87290 21760 87300
rect 21860 87290 21940 87300
rect 22040 87290 22120 87300
rect 22220 87290 22300 87300
rect 22400 87290 22480 87300
rect 22580 87290 22660 87300
rect 22760 87290 22840 87300
rect 22940 87290 23020 87300
rect 23120 87290 23200 87300
rect 23300 87290 23380 87300
rect 23480 87290 23560 87300
rect 23660 87290 23740 87300
rect 23840 87290 23920 87300
rect 24020 87290 24100 87300
rect 24200 87290 24280 87300
rect 24380 87290 24460 87300
rect 24560 87290 24640 87300
rect 24740 87290 24820 87300
rect 24920 87290 25000 87300
rect 25100 87290 25180 87300
rect 25280 87290 25360 87300
rect 25460 87290 25540 87300
rect 25640 87290 25720 87300
rect 25820 87290 25900 87300
rect 26000 87290 26080 87300
rect 26180 87290 26260 87300
rect 26360 87290 26440 87300
rect 26540 87290 26620 87300
rect 152080 87290 152160 87300
rect 152260 87290 152340 87300
rect 152440 87290 152520 87300
rect 152620 87290 152700 87300
rect 152800 87290 152880 87300
rect 152980 87290 153060 87300
rect 153160 87290 153240 87300
rect 153340 87290 153420 87300
rect 153520 87290 153600 87300
rect 153700 87290 153780 87300
rect 153880 87290 153960 87300
rect 154060 87290 154140 87300
rect 154240 87290 154320 87300
rect 154420 87290 154500 87300
rect 154600 87290 154680 87300
rect 154780 87290 154860 87300
rect 154960 87290 155040 87300
rect 155140 87290 155220 87300
rect 155320 87290 155400 87300
rect 155500 87290 155580 87300
rect 155680 87290 155760 87300
rect 155860 87290 155940 87300
rect 156040 87290 156120 87300
rect 156220 87290 156300 87300
rect 156400 87290 156480 87300
rect 156580 87290 156660 87300
rect 156760 87290 156840 87300
rect 156940 87290 157020 87300
rect 157120 87290 157200 87300
rect 157300 87290 157380 87300
rect 157480 87290 157560 87300
rect 157660 87290 157740 87300
rect 157840 87290 157920 87300
rect 158020 87290 158100 87300
rect 158200 87290 158280 87300
rect 158380 87290 158460 87300
rect 158560 87290 158640 87300
rect 158740 87290 158820 87300
rect 158920 87290 159000 87300
rect 159100 87290 159180 87300
rect 159280 87290 159360 87300
rect 159460 87290 159540 87300
rect 159640 87290 159720 87300
rect 19060 87210 19070 87290
rect 19240 87210 19250 87290
rect 19420 87210 19430 87290
rect 19600 87210 19610 87290
rect 19780 87210 19790 87290
rect 19960 87210 19970 87290
rect 20140 87210 20150 87290
rect 20320 87210 20330 87290
rect 20500 87210 20510 87290
rect 20680 87210 20690 87290
rect 20860 87210 20870 87290
rect 21040 87210 21050 87290
rect 21220 87210 21230 87290
rect 21400 87210 21410 87290
rect 21580 87210 21590 87290
rect 21760 87210 21770 87290
rect 21940 87210 21950 87290
rect 22120 87210 22130 87290
rect 22300 87210 22310 87290
rect 22480 87210 22490 87290
rect 22660 87210 22670 87290
rect 22840 87210 22850 87290
rect 23020 87210 23030 87290
rect 23200 87210 23210 87290
rect 23380 87210 23390 87290
rect 23560 87210 23570 87290
rect 23740 87210 23750 87290
rect 23920 87210 23930 87290
rect 24100 87210 24110 87290
rect 24280 87210 24290 87290
rect 24460 87210 24470 87290
rect 24640 87210 24650 87290
rect 24820 87210 24830 87290
rect 25000 87210 25010 87290
rect 25180 87210 25190 87290
rect 25360 87210 25370 87290
rect 25540 87210 25550 87290
rect 25720 87210 25730 87290
rect 25900 87210 25910 87290
rect 26080 87210 26090 87290
rect 26260 87210 26270 87290
rect 26440 87210 26450 87290
rect 26620 87210 26630 87290
rect 152160 87210 152170 87290
rect 152340 87210 152350 87290
rect 152520 87210 152530 87290
rect 152700 87210 152710 87290
rect 152880 87210 152890 87290
rect 153060 87210 153070 87290
rect 153240 87210 153250 87290
rect 153420 87210 153430 87290
rect 153600 87210 153610 87290
rect 153780 87210 153790 87290
rect 153960 87210 153970 87290
rect 154140 87210 154150 87290
rect 154320 87210 154330 87290
rect 154500 87210 154510 87290
rect 154680 87210 154690 87290
rect 154860 87210 154870 87290
rect 155040 87210 155050 87290
rect 155220 87210 155230 87290
rect 155400 87210 155410 87290
rect 155580 87210 155590 87290
rect 155760 87210 155770 87290
rect 155940 87210 155950 87290
rect 156120 87210 156130 87290
rect 156300 87210 156310 87290
rect 156480 87210 156490 87290
rect 156660 87210 156670 87290
rect 156840 87210 156850 87290
rect 157020 87210 157030 87290
rect 157200 87210 157210 87290
rect 157380 87210 157390 87290
rect 157560 87210 157570 87290
rect 157740 87210 157750 87290
rect 157920 87210 157930 87290
rect 158100 87210 158110 87290
rect 158280 87210 158290 87290
rect 158460 87210 158470 87290
rect 158640 87210 158650 87290
rect 158820 87210 158830 87290
rect 159000 87210 159010 87290
rect 159180 87210 159190 87290
rect 159360 87210 159370 87290
rect 159540 87210 159550 87290
rect 159720 87210 159730 87290
rect 161965 87265 161975 87345
rect 162145 87265 162155 87345
rect 162325 87265 162335 87345
rect 162505 87265 162515 87345
rect 162685 87265 162695 87345
rect 163380 87290 163460 87300
rect 163560 87290 163640 87300
rect 163740 87290 163820 87300
rect 163920 87290 164000 87300
rect 164100 87290 164180 87300
rect 164280 87290 164360 87300
rect 164460 87290 164540 87300
rect 164640 87290 164720 87300
rect 164820 87290 164900 87300
rect 165000 87290 165080 87300
rect 165180 87290 165260 87300
rect 165360 87290 165440 87300
rect 165540 87290 165620 87300
rect 165720 87290 165800 87300
rect 165900 87290 165980 87300
rect 166080 87290 166160 87300
rect 166260 87290 166340 87300
rect 166440 87290 166520 87300
rect 166620 87290 166700 87300
rect 166800 87290 166880 87300
rect 166980 87290 167060 87300
rect 167160 87290 167240 87300
rect 167340 87290 167420 87300
rect 167520 87290 167600 87300
rect 167700 87290 167780 87300
rect 167880 87290 167960 87300
rect 168060 87290 168140 87300
rect 168240 87290 168320 87300
rect 168420 87290 168500 87300
rect 168600 87290 168680 87300
rect 168780 87290 168860 87300
rect 168960 87290 169040 87300
rect 169140 87290 169220 87300
rect 169320 87290 169400 87300
rect 169500 87290 169580 87300
rect 169680 87290 169760 87300
rect 169860 87290 169940 87300
rect 170040 87290 170120 87300
rect 170220 87290 170300 87300
rect 170400 87290 170480 87300
rect 170580 87290 170660 87300
rect 170760 87290 170840 87300
rect 170940 87290 171020 87300
rect 163460 87210 163470 87290
rect 163640 87210 163650 87290
rect 163820 87210 163830 87290
rect 164000 87210 164010 87290
rect 164180 87210 164190 87290
rect 164360 87210 164370 87290
rect 164540 87210 164550 87290
rect 164720 87210 164730 87290
rect 164900 87210 164910 87290
rect 165080 87210 165090 87290
rect 165260 87210 165270 87290
rect 165440 87210 165450 87290
rect 165620 87210 165630 87290
rect 165800 87210 165810 87290
rect 165980 87210 165990 87290
rect 166160 87210 166170 87290
rect 166340 87210 166350 87290
rect 166520 87210 166530 87290
rect 166700 87210 166710 87290
rect 166880 87210 166890 87290
rect 167060 87210 167070 87290
rect 167240 87210 167250 87290
rect 167420 87210 167430 87290
rect 167600 87210 167610 87290
rect 167780 87210 167790 87290
rect 167960 87210 167970 87290
rect 168140 87210 168150 87290
rect 168320 87210 168330 87290
rect 168500 87210 168510 87290
rect 168680 87210 168690 87290
rect 168860 87210 168870 87290
rect 169040 87210 169050 87290
rect 169220 87210 169230 87290
rect 169400 87210 169410 87290
rect 169580 87210 169590 87290
rect 169760 87210 169770 87290
rect 169940 87210 169950 87290
rect 170120 87210 170130 87290
rect 170300 87210 170310 87290
rect 170480 87210 170490 87290
rect 170660 87210 170670 87290
rect 170840 87210 170850 87290
rect 171020 87210 171030 87290
rect 146100 87150 146160 87180
rect 147580 87150 147640 87180
rect 148400 87150 148460 87180
rect 149880 87150 149940 87180
rect 161885 87165 161965 87175
rect 162065 87165 162145 87175
rect 162245 87165 162325 87175
rect 162425 87165 162505 87175
rect 162605 87165 162685 87175
rect 146100 87030 146160 87060
rect 146210 87040 146220 87130
rect 19130 86910 19160 86940
rect 19250 86910 19280 86940
rect 26420 86910 26450 86940
rect 26540 86910 26570 86940
rect 146100 86910 146160 86940
rect 19010 86880 19070 86910
rect 19130 86880 19190 86910
rect 19250 86880 19310 86910
rect 26300 86880 26360 86910
rect 26420 86880 26480 86910
rect 26540 86880 26600 86910
rect 19130 86790 19160 86820
rect 19250 86790 19280 86820
rect 26420 86790 26450 86820
rect 26540 86790 26570 86820
rect 146100 86790 146160 86820
rect 19010 86760 19070 86790
rect 19130 86760 19190 86790
rect 19250 86760 19310 86790
rect 26300 86760 26360 86790
rect 26420 86760 26480 86790
rect 26540 86760 26600 86790
rect 146100 86670 146160 86700
rect 146100 86550 146160 86580
rect 146100 86430 146160 86460
rect 146100 86310 146160 86340
rect 146100 86190 146160 86220
rect 36020 86180 36100 86190
rect 36200 86180 36280 86190
rect 36380 86180 36460 86190
rect 36560 86180 36640 86190
rect 36740 86180 36820 86190
rect 36920 86180 37000 86190
rect 37100 86180 37180 86190
rect 37280 86180 37360 86190
rect 37460 86180 37540 86190
rect 37640 86180 37720 86190
rect 37820 86180 37900 86190
rect 38000 86180 38080 86190
rect 38180 86180 38260 86190
rect 38360 86180 38440 86190
rect 38540 86180 38620 86190
rect 38720 86180 38800 86190
rect 38900 86180 38980 86190
rect 39080 86180 39160 86190
rect 39260 86180 39340 86190
rect 39440 86180 39520 86190
rect 39620 86180 39700 86190
rect 39800 86180 39880 86190
rect 39980 86180 40060 86190
rect 40160 86180 40240 86190
rect 40340 86180 40420 86190
rect 40520 86180 40600 86190
rect 40700 86180 40780 86190
rect 40880 86180 40960 86190
rect 41060 86180 41140 86190
rect 41240 86180 41320 86190
rect 41420 86180 41500 86190
rect 41600 86180 41680 86190
rect 36100 86100 36110 86180
rect 36280 86100 36290 86180
rect 36460 86100 36470 86180
rect 36640 86100 36650 86180
rect 36820 86100 36830 86180
rect 37000 86100 37010 86180
rect 37180 86100 37190 86180
rect 37360 86100 37370 86180
rect 37540 86100 37550 86180
rect 37720 86100 37730 86180
rect 37900 86100 37910 86180
rect 38080 86100 38090 86180
rect 38260 86100 38270 86180
rect 38440 86100 38450 86180
rect 38620 86100 38630 86180
rect 38800 86100 38810 86180
rect 38980 86100 38990 86180
rect 39160 86100 39170 86180
rect 39340 86100 39350 86180
rect 39520 86100 39530 86180
rect 39700 86100 39710 86180
rect 39880 86100 39890 86180
rect 40060 86100 40070 86180
rect 40240 86100 40250 86180
rect 40420 86100 40430 86180
rect 40600 86100 40610 86180
rect 40780 86100 40790 86180
rect 40960 86100 40970 86180
rect 41140 86100 41150 86180
rect 41320 86100 41330 86180
rect 41500 86100 41510 86180
rect 41680 86100 41690 86180
rect 146100 86070 146160 86100
rect 146100 85950 146160 85980
rect 36020 85880 36100 85890
rect 36200 85880 36280 85890
rect 36380 85880 36460 85890
rect 36560 85880 36640 85890
rect 36740 85880 36820 85890
rect 36920 85880 37000 85890
rect 37100 85880 37180 85890
rect 37280 85880 37360 85890
rect 37460 85880 37540 85890
rect 37640 85880 37720 85890
rect 37820 85880 37900 85890
rect 38000 85880 38080 85890
rect 38180 85880 38260 85890
rect 38360 85880 38440 85890
rect 38540 85880 38620 85890
rect 38720 85880 38800 85890
rect 38900 85880 38980 85890
rect 39080 85880 39160 85890
rect 39260 85880 39340 85890
rect 39440 85880 39520 85890
rect 39620 85880 39700 85890
rect 39800 85880 39880 85890
rect 39980 85880 40060 85890
rect 40160 85880 40240 85890
rect 40340 85880 40420 85890
rect 40520 85880 40600 85890
rect 40700 85880 40780 85890
rect 40880 85880 40960 85890
rect 41060 85880 41140 85890
rect 41240 85880 41320 85890
rect 41420 85880 41500 85890
rect 41600 85880 41680 85890
rect 36100 85800 36110 85880
rect 36280 85800 36290 85880
rect 36460 85800 36470 85880
rect 36640 85800 36650 85880
rect 36820 85800 36830 85880
rect 37000 85800 37010 85880
rect 37180 85800 37190 85880
rect 37360 85800 37370 85880
rect 37540 85800 37550 85880
rect 37720 85800 37730 85880
rect 37900 85800 37910 85880
rect 38080 85800 38090 85880
rect 38260 85800 38270 85880
rect 38440 85800 38450 85880
rect 38620 85800 38630 85880
rect 38800 85800 38810 85880
rect 38980 85800 38990 85880
rect 39160 85800 39170 85880
rect 39340 85800 39350 85880
rect 39520 85800 39530 85880
rect 39700 85800 39710 85880
rect 39880 85800 39890 85880
rect 40060 85800 40070 85880
rect 40240 85800 40250 85880
rect 40420 85800 40430 85880
rect 40600 85800 40610 85880
rect 40780 85800 40790 85880
rect 40960 85800 40970 85880
rect 41140 85800 41150 85880
rect 41320 85800 41330 85880
rect 41500 85800 41510 85880
rect 41680 85800 41690 85880
rect 46660 85660 47160 85840
rect 146100 85830 146160 85860
rect 146100 85710 146160 85740
rect 146300 85650 146310 87040
rect 146690 87000 146810 87060
rect 146970 87000 147090 87060
rect 147580 87030 147640 87060
rect 148400 87030 148460 87060
rect 148820 87050 149620 87140
rect 148950 87020 149070 87050
rect 149230 87020 149350 87050
rect 149070 87010 149130 87020
rect 149350 87010 149410 87020
rect 149070 87000 149190 87010
rect 149350 87000 149470 87010
rect 146810 86990 146870 87000
rect 146570 86980 146650 86990
rect 146810 86980 146930 86990
rect 146650 86900 146660 86980
rect 146810 86880 146870 86980
rect 146930 86900 146940 86980
rect 147090 86880 147150 87000
rect 146410 86830 147140 86840
rect 146410 86750 146420 86830
rect 147220 86825 147230 86880
rect 147270 86850 147390 86910
rect 146460 86815 147250 86825
rect 146450 86765 146460 86815
rect 146500 86560 146510 86750
rect 146690 86700 146810 86760
rect 146970 86700 147090 86760
rect 147220 86736 147230 86815
rect 147390 86736 147450 86850
rect 147520 86736 147530 86970
rect 147580 86910 147640 86940
rect 148400 86910 148460 86940
rect 148510 86900 148520 86990
rect 147580 86790 147640 86820
rect 148400 86790 148460 86820
rect 148600 86736 148610 86900
rect 148650 86870 148770 86930
rect 149070 86900 149130 87000
rect 149190 86920 149200 87000
rect 149350 86900 149410 87000
rect 149470 86920 149480 87000
rect 148770 86845 148830 86870
rect 149530 86865 149620 87050
rect 148910 86860 149620 86865
rect 148900 86850 149630 86860
rect 148910 86845 149630 86850
rect 148770 86835 149630 86845
rect 148770 86750 148830 86835
rect 149530 86785 149630 86835
rect 148910 86755 149630 86785
rect 148950 86736 149070 86755
rect 149230 86736 149350 86755
rect 149530 86736 149630 86755
rect 149820 86736 149830 87150
rect 152080 87140 152160 87150
rect 152260 87140 152340 87150
rect 152440 87140 152520 87150
rect 152620 87140 152700 87150
rect 152800 87140 152880 87150
rect 152980 87140 153060 87150
rect 153160 87140 153240 87150
rect 153340 87140 153420 87150
rect 153520 87140 153600 87150
rect 153700 87140 153780 87150
rect 153880 87140 153960 87150
rect 154060 87140 154140 87150
rect 154240 87140 154320 87150
rect 154420 87140 154500 87150
rect 154600 87140 154680 87150
rect 154780 87140 154860 87150
rect 154960 87140 155040 87150
rect 155140 87140 155220 87150
rect 155320 87140 155400 87150
rect 155500 87140 155580 87150
rect 155680 87140 155760 87150
rect 155860 87140 155940 87150
rect 156040 87140 156120 87150
rect 156220 87140 156300 87150
rect 156400 87140 156480 87150
rect 156580 87140 156660 87150
rect 156760 87140 156840 87150
rect 156940 87140 157020 87150
rect 157120 87140 157200 87150
rect 157300 87140 157380 87150
rect 157480 87140 157560 87150
rect 157660 87140 157740 87150
rect 157840 87140 157920 87150
rect 158020 87140 158100 87150
rect 158200 87140 158280 87150
rect 158380 87140 158460 87150
rect 158560 87140 158640 87150
rect 158740 87140 158820 87150
rect 158920 87140 159000 87150
rect 159100 87140 159180 87150
rect 159280 87140 159360 87150
rect 159460 87140 159540 87150
rect 159640 87140 159720 87150
rect 152160 87060 152170 87140
rect 152340 87060 152350 87140
rect 152520 87060 152530 87140
rect 152700 87060 152710 87140
rect 152880 87060 152890 87140
rect 153060 87060 153070 87140
rect 153240 87060 153250 87140
rect 153420 87060 153430 87140
rect 153600 87060 153610 87140
rect 153780 87060 153790 87140
rect 153960 87060 153970 87140
rect 154140 87060 154150 87140
rect 154320 87060 154330 87140
rect 154500 87060 154510 87140
rect 154680 87060 154690 87140
rect 154860 87060 154870 87140
rect 155040 87060 155050 87140
rect 155220 87060 155230 87140
rect 155400 87060 155410 87140
rect 155580 87060 155590 87140
rect 155760 87060 155770 87140
rect 155940 87060 155950 87140
rect 156120 87060 156130 87140
rect 156300 87060 156310 87140
rect 156480 87060 156490 87140
rect 156660 87060 156670 87140
rect 156840 87060 156850 87140
rect 157020 87060 157030 87140
rect 157200 87060 157210 87140
rect 157380 87060 157390 87140
rect 157560 87060 157570 87140
rect 157740 87060 157750 87140
rect 157920 87060 157930 87140
rect 158100 87060 158110 87140
rect 158280 87060 158290 87140
rect 158460 87060 158470 87140
rect 158640 87060 158650 87140
rect 158820 87060 158830 87140
rect 159000 87060 159010 87140
rect 159180 87060 159190 87140
rect 159360 87060 159370 87140
rect 159540 87060 159550 87140
rect 159720 87060 159730 87140
rect 161965 87085 161975 87165
rect 162145 87085 162155 87165
rect 162325 87085 162335 87165
rect 162505 87085 162515 87165
rect 162685 87085 162695 87165
rect 163380 87140 163460 87150
rect 163560 87140 163640 87150
rect 163740 87140 163820 87150
rect 163920 87140 164000 87150
rect 164100 87140 164180 87150
rect 164280 87140 164360 87150
rect 164460 87140 164540 87150
rect 164640 87140 164720 87150
rect 164820 87140 164900 87150
rect 165000 87140 165080 87150
rect 165180 87140 165260 87150
rect 165360 87140 165440 87150
rect 165540 87140 165620 87150
rect 165720 87140 165800 87150
rect 165900 87140 165980 87150
rect 166080 87140 166160 87150
rect 166260 87140 166340 87150
rect 166440 87140 166520 87150
rect 166620 87140 166700 87150
rect 166800 87140 166880 87150
rect 166980 87140 167060 87150
rect 167160 87140 167240 87150
rect 167340 87140 167420 87150
rect 167520 87140 167600 87150
rect 167700 87140 167780 87150
rect 167880 87140 167960 87150
rect 168060 87140 168140 87150
rect 168240 87140 168320 87150
rect 168420 87140 168500 87150
rect 168600 87140 168680 87150
rect 168780 87140 168860 87150
rect 168960 87140 169040 87150
rect 169140 87140 169220 87150
rect 169320 87140 169400 87150
rect 169500 87140 169580 87150
rect 169680 87140 169760 87150
rect 169860 87140 169940 87150
rect 170040 87140 170120 87150
rect 170220 87140 170300 87150
rect 170400 87140 170480 87150
rect 170580 87140 170660 87150
rect 170760 87140 170840 87150
rect 170940 87140 171020 87150
rect 163460 87060 163470 87140
rect 163640 87060 163650 87140
rect 163820 87060 163830 87140
rect 164000 87060 164010 87140
rect 164180 87060 164190 87140
rect 164360 87060 164370 87140
rect 164540 87060 164550 87140
rect 164720 87060 164730 87140
rect 164900 87060 164910 87140
rect 165080 87060 165090 87140
rect 165260 87060 165270 87140
rect 165440 87060 165450 87140
rect 165620 87060 165630 87140
rect 165800 87060 165810 87140
rect 165980 87060 165990 87140
rect 166160 87060 166170 87140
rect 166340 87060 166350 87140
rect 166520 87060 166530 87140
rect 166700 87060 166710 87140
rect 166880 87060 166890 87140
rect 167060 87060 167070 87140
rect 167240 87060 167250 87140
rect 167420 87060 167430 87140
rect 167600 87060 167610 87140
rect 167780 87060 167790 87140
rect 167960 87060 167970 87140
rect 168140 87060 168150 87140
rect 168320 87060 168330 87140
rect 168500 87060 168510 87140
rect 168680 87060 168690 87140
rect 168860 87060 168870 87140
rect 169040 87060 169050 87140
rect 169220 87060 169230 87140
rect 169400 87060 169410 87140
rect 169580 87060 169590 87140
rect 169760 87060 169770 87140
rect 169940 87060 169950 87140
rect 170120 87060 170130 87140
rect 170300 87060 170310 87140
rect 170480 87060 170490 87140
rect 170660 87060 170670 87140
rect 170840 87060 170850 87140
rect 171020 87060 171030 87140
rect 149880 87030 149940 87060
rect 149880 86910 149940 86940
rect 152220 86890 152250 86920
rect 152340 86890 152370 86920
rect 159520 86890 159550 86920
rect 159640 86890 159670 86920
rect 152100 86860 152160 86890
rect 152220 86860 152280 86890
rect 152340 86860 152400 86890
rect 159400 86860 159460 86890
rect 159520 86860 159580 86890
rect 159640 86860 159700 86890
rect 149880 86790 149940 86820
rect 152220 86770 152250 86800
rect 152340 86770 152370 86800
rect 159520 86770 159550 86800
rect 159640 86770 159670 86800
rect 163520 86770 163550 86800
rect 163640 86770 163670 86800
rect 170810 86770 170840 86800
rect 170930 86770 170960 86800
rect 152100 86740 152160 86770
rect 152220 86740 152280 86770
rect 152340 86740 152400 86770
rect 152810 86736 158990 86760
rect 159400 86740 159460 86770
rect 159520 86740 159580 86770
rect 159640 86740 159700 86770
rect 163400 86740 163460 86770
rect 163520 86740 163580 86770
rect 163640 86740 163700 86770
rect 170690 86740 170750 86770
rect 170810 86740 170870 86770
rect 170930 86740 170990 86770
rect 164280 86736 164360 86740
rect 164460 86736 164540 86740
rect 164640 86736 164720 86740
rect 164820 86736 164900 86740
rect 165000 86736 165080 86740
rect 165180 86736 165260 86740
rect 165360 86736 165440 86740
rect 165540 86736 165620 86740
rect 165720 86736 165800 86740
rect 165900 86736 165980 86740
rect 166080 86736 166160 86740
rect 166260 86736 166340 86740
rect 166440 86736 166520 86740
rect 166620 86736 166700 86740
rect 166800 86736 166880 86740
rect 166980 86736 167060 86740
rect 167160 86736 167240 86740
rect 167340 86736 167420 86740
rect 167520 86736 167600 86740
rect 167700 86736 167780 86740
rect 167880 86736 167960 86740
rect 168060 86736 168140 86740
rect 168240 86736 168320 86740
rect 168420 86736 168500 86740
rect 168600 86736 168680 86740
rect 168780 86736 168860 86740
rect 168960 86736 169040 86740
rect 169140 86736 169220 86740
rect 169320 86736 169400 86740
rect 169500 86736 169580 86740
rect 169680 86736 169760 86740
rect 169860 86736 169940 86740
rect 170040 86736 170120 86740
rect 146810 86690 146870 86700
rect 146570 86680 146650 86690
rect 146710 86680 146790 86690
rect 146810 86680 146930 86690
rect 146990 86680 147070 86690
rect 146650 86600 146660 86680
rect 146790 86600 146800 86680
rect 146810 86580 146870 86680
rect 146930 86600 146940 86680
rect 147070 86600 147080 86680
rect 147090 86580 147150 86700
rect 146500 86550 147130 86560
rect 146500 86540 146510 86550
rect 146690 86410 146810 86470
rect 146970 86410 147090 86470
rect 146690 86320 146700 86410
rect 146800 86380 146870 86410
rect 146810 86290 146870 86380
rect 146970 86320 146980 86410
rect 147090 86290 147150 86410
rect 146410 86240 147140 86250
rect 146410 86160 146420 86240
rect 146460 86225 147150 86235
rect 146450 86175 146460 86225
rect 146500 85970 146510 86160
rect 146690 86110 146810 86170
rect 146970 86110 147090 86170
rect 146810 86100 146870 86110
rect 146570 86090 146650 86100
rect 146710 86090 146790 86100
rect 146810 86090 146930 86100
rect 146990 86090 147070 86100
rect 146650 86010 146660 86090
rect 146790 86010 146800 86090
rect 146810 85990 146870 86090
rect 146930 86010 146940 86090
rect 147070 86010 147080 86090
rect 147090 85990 147150 86110
rect 146500 85960 147130 85970
rect 146500 85950 146510 85960
rect 146690 85820 146810 85880
rect 146970 85820 147090 85880
rect 146690 85730 146700 85820
rect 146800 85790 146870 85820
rect 146810 85700 146870 85790
rect 146970 85730 146980 85820
rect 147090 85700 147150 85820
rect 146410 85650 147140 85660
rect 146460 85635 147150 85645
rect 146100 85590 146160 85620
rect 146450 85585 146460 85635
rect 146690 85520 146810 85580
rect 146970 85520 147090 85580
rect 146810 85510 146870 85520
rect 146570 85500 146650 85510
rect 146710 85500 146790 85510
rect 146810 85500 146930 85510
rect 146990 85500 147070 85510
rect 36020 85470 36100 85480
rect 36200 85470 36280 85480
rect 36380 85470 36460 85480
rect 36560 85470 36640 85480
rect 36740 85470 36820 85480
rect 36920 85470 37000 85480
rect 37100 85470 37180 85480
rect 37280 85470 37360 85480
rect 37460 85470 37540 85480
rect 37640 85470 37720 85480
rect 37820 85470 37900 85480
rect 38000 85470 38080 85480
rect 38180 85470 38260 85480
rect 38360 85470 38440 85480
rect 38540 85470 38620 85480
rect 38720 85470 38800 85480
rect 38900 85470 38980 85480
rect 39080 85470 39160 85480
rect 39260 85470 39340 85480
rect 39440 85470 39520 85480
rect 39620 85470 39700 85480
rect 39800 85470 39880 85480
rect 39980 85470 40060 85480
rect 40160 85470 40240 85480
rect 40340 85470 40420 85480
rect 40520 85470 40600 85480
rect 40700 85470 40780 85480
rect 40880 85470 40960 85480
rect 41060 85470 41140 85480
rect 41240 85470 41320 85480
rect 146100 85470 146160 85500
rect 36100 85390 36110 85470
rect 36280 85390 36290 85470
rect 36460 85390 36470 85470
rect 36640 85390 36650 85470
rect 36820 85390 36830 85470
rect 37000 85390 37010 85470
rect 37180 85390 37190 85470
rect 37360 85390 37370 85470
rect 37540 85390 37550 85470
rect 37720 85390 37730 85470
rect 37900 85390 37910 85470
rect 38080 85390 38090 85470
rect 38260 85390 38270 85470
rect 38440 85390 38450 85470
rect 38620 85390 38630 85470
rect 38800 85390 38810 85470
rect 38980 85390 38990 85470
rect 39160 85390 39170 85470
rect 39340 85390 39350 85470
rect 39520 85390 39530 85470
rect 39700 85390 39710 85470
rect 39880 85390 39890 85470
rect 40060 85390 40070 85470
rect 40240 85390 40250 85470
rect 40420 85390 40430 85470
rect 40600 85390 40610 85470
rect 40780 85390 40790 85470
rect 40960 85390 40970 85470
rect 41140 85390 41150 85470
rect 41320 85390 41330 85470
rect 146650 85420 146660 85500
rect 146790 85420 146800 85500
rect 146810 85400 146870 85500
rect 146930 85420 146940 85500
rect 147070 85420 147080 85500
rect 147090 85400 147150 85520
rect 146100 85350 146160 85380
rect 146100 85230 146160 85260
rect 36020 85170 36100 85180
rect 36200 85170 36280 85180
rect 36380 85170 36460 85180
rect 36560 85170 36640 85180
rect 36740 85170 36820 85180
rect 36920 85170 37000 85180
rect 37100 85170 37180 85180
rect 37280 85170 37360 85180
rect 37460 85170 37540 85180
rect 37640 85170 37720 85180
rect 37820 85170 37900 85180
rect 38000 85170 38080 85180
rect 38180 85170 38260 85180
rect 38360 85170 38440 85180
rect 38540 85170 38620 85180
rect 38720 85170 38800 85180
rect 38900 85170 38980 85180
rect 39080 85170 39160 85180
rect 39260 85170 39340 85180
rect 39440 85170 39520 85180
rect 39620 85170 39700 85180
rect 39800 85170 39880 85180
rect 39980 85170 40060 85180
rect 40160 85170 40240 85180
rect 40340 85170 40420 85180
rect 40520 85170 40600 85180
rect 40700 85170 40780 85180
rect 40880 85170 40960 85180
rect 41060 85170 41140 85180
rect 41240 85170 41320 85180
rect 36100 85090 36110 85170
rect 36280 85090 36290 85170
rect 36460 85090 36470 85170
rect 36640 85090 36650 85170
rect 36820 85090 36830 85170
rect 37000 85090 37010 85170
rect 37180 85090 37190 85170
rect 37360 85090 37370 85170
rect 37540 85090 37550 85170
rect 37720 85090 37730 85170
rect 37900 85090 37910 85170
rect 38080 85090 38090 85170
rect 38260 85090 38270 85170
rect 38440 85090 38450 85170
rect 38620 85090 38630 85170
rect 38800 85090 38810 85170
rect 38980 85090 38990 85170
rect 39160 85090 39170 85170
rect 39340 85090 39350 85170
rect 39520 85090 39530 85170
rect 39700 85090 39710 85170
rect 39880 85090 39890 85170
rect 40060 85090 40070 85170
rect 40240 85090 40250 85170
rect 40420 85090 40430 85170
rect 40600 85090 40610 85170
rect 40780 85090 40790 85170
rect 40960 85090 40970 85170
rect 41140 85090 41150 85170
rect 41320 85090 41330 85170
rect 146100 85110 146160 85140
rect 36000 85030 41400 85040
rect 146100 84990 146160 85020
rect 146690 84940 146810 85000
rect 146970 84940 147090 85000
rect 146810 84930 146870 84940
rect 146570 84920 146650 84930
rect 146810 84920 146930 84930
rect 146100 84870 146160 84900
rect 36020 84850 36100 84860
rect 36200 84850 36280 84860
rect 36380 84850 36460 84860
rect 36560 84850 36640 84860
rect 36740 84850 36820 84860
rect 36920 84850 37000 84860
rect 37100 84850 37180 84860
rect 37280 84850 37360 84860
rect 37460 84850 37540 84860
rect 37640 84850 37720 84860
rect 37820 84850 37900 84860
rect 38000 84850 38080 84860
rect 38180 84850 38260 84860
rect 38360 84850 38440 84860
rect 38540 84850 38620 84860
rect 38720 84850 38800 84860
rect 38900 84850 38980 84860
rect 39080 84850 39160 84860
rect 39260 84850 39340 84860
rect 39440 84850 39520 84860
rect 39620 84850 39700 84860
rect 39800 84850 39880 84860
rect 39980 84850 40060 84860
rect 40160 84850 40240 84860
rect 40340 84850 40420 84860
rect 40520 84850 40600 84860
rect 40700 84850 40780 84860
rect 40880 84850 40960 84860
rect 41060 84850 41140 84860
rect 41240 84850 41320 84860
rect 36100 84770 36110 84850
rect 36280 84770 36290 84850
rect 36460 84770 36470 84850
rect 36640 84770 36650 84850
rect 36820 84770 36830 84850
rect 37000 84770 37010 84850
rect 37180 84770 37190 84850
rect 37360 84770 37370 84850
rect 37540 84770 37550 84850
rect 37720 84770 37730 84850
rect 37900 84770 37910 84850
rect 38080 84770 38090 84850
rect 38260 84770 38270 84850
rect 38440 84770 38450 84850
rect 38620 84770 38630 84850
rect 38800 84770 38810 84850
rect 38980 84770 38990 84850
rect 39160 84770 39170 84850
rect 39340 84770 39350 84850
rect 39520 84770 39530 84850
rect 39700 84770 39710 84850
rect 39880 84770 39890 84850
rect 40060 84770 40070 84850
rect 40240 84770 40250 84850
rect 40420 84770 40430 84850
rect 40600 84770 40610 84850
rect 40780 84770 40790 84850
rect 40960 84770 40970 84850
rect 41140 84770 41150 84850
rect 41320 84770 41330 84850
rect 146650 84840 146660 84920
rect 146810 84820 146870 84920
rect 146930 84840 146940 84920
rect 147090 84820 147150 84940
rect 146100 84750 146160 84780
rect 146500 84770 147140 84780
rect 146460 84755 147150 84765
rect 36000 84700 36040 84710
rect 36140 84700 36220 84710
rect 36320 84700 36400 84710
rect 36500 84700 36580 84710
rect 36680 84700 36760 84710
rect 36860 84700 36940 84710
rect 37040 84700 37120 84710
rect 37220 84700 37300 84710
rect 37400 84700 37480 84710
rect 37580 84700 37660 84710
rect 37760 84700 37840 84710
rect 146450 84705 146460 84755
rect 36040 84620 36050 84700
rect 36220 84620 36230 84700
rect 36400 84620 36410 84700
rect 36580 84620 36590 84700
rect 36760 84620 36770 84700
rect 36940 84620 36950 84700
rect 37120 84620 37130 84700
rect 37300 84620 37310 84700
rect 37480 84620 37490 84700
rect 37660 84620 37670 84700
rect 37840 84620 37850 84700
rect 40160 84695 40240 84705
rect 40340 84695 40420 84705
rect 40520 84695 40600 84705
rect 40700 84695 40780 84705
rect 40880 84695 40960 84705
rect 41060 84695 41140 84705
rect 41240 84695 41320 84705
rect 40240 84615 40250 84695
rect 40420 84615 40430 84695
rect 40600 84615 40610 84695
rect 40780 84615 40790 84695
rect 40960 84615 40970 84695
rect 41140 84615 41150 84695
rect 41320 84615 41330 84695
rect 146100 84630 146160 84660
rect 146690 84640 146810 84700
rect 146970 84640 147090 84700
rect 146810 84630 146870 84640
rect 146570 84620 146650 84630
rect 146710 84620 146790 84630
rect 146810 84620 146930 84630
rect 146990 84620 147070 84630
rect 146650 84540 146660 84620
rect 146790 84540 146800 84620
rect 36020 84530 36100 84540
rect 36200 84530 36280 84540
rect 36380 84530 36460 84540
rect 36560 84530 36640 84540
rect 36740 84530 36820 84540
rect 36920 84530 37000 84540
rect 37100 84530 37180 84540
rect 37280 84530 37360 84540
rect 37460 84530 37540 84540
rect 37640 84530 37720 84540
rect 37820 84530 37900 84540
rect 38000 84530 38080 84540
rect 38180 84530 38260 84540
rect 38360 84530 38440 84540
rect 38540 84530 38620 84540
rect 38720 84530 38800 84540
rect 38900 84530 38980 84540
rect 39080 84530 39160 84540
rect 39260 84530 39340 84540
rect 39440 84530 39520 84540
rect 39620 84530 39700 84540
rect 39800 84530 39880 84540
rect 39980 84530 40060 84540
rect 40160 84530 40240 84540
rect 40340 84530 40420 84540
rect 40520 84530 40600 84540
rect 40700 84530 40780 84540
rect 40880 84530 40960 84540
rect 41060 84530 41140 84540
rect 41240 84530 41320 84540
rect 36100 84450 36110 84530
rect 36280 84450 36290 84530
rect 36460 84450 36470 84530
rect 36640 84450 36650 84530
rect 36820 84450 36830 84530
rect 37000 84450 37010 84530
rect 37180 84450 37190 84530
rect 37360 84450 37370 84530
rect 37540 84450 37550 84530
rect 37720 84450 37730 84530
rect 37900 84450 37910 84530
rect 38080 84450 38090 84530
rect 38260 84450 38270 84530
rect 38440 84450 38450 84530
rect 38620 84450 38630 84530
rect 38800 84450 38810 84530
rect 38980 84450 38990 84530
rect 39160 84450 39170 84530
rect 39340 84450 39350 84530
rect 39520 84450 39530 84530
rect 39700 84450 39710 84530
rect 39880 84450 39890 84530
rect 40060 84450 40070 84530
rect 40240 84450 40250 84530
rect 40420 84450 40430 84530
rect 40600 84450 40610 84530
rect 40780 84450 40790 84530
rect 40960 84450 40970 84530
rect 41140 84450 41150 84530
rect 41320 84450 41330 84530
rect 146100 84510 146160 84540
rect 146810 84520 146870 84620
rect 146930 84540 146940 84620
rect 147070 84540 147080 84620
rect 147090 84520 147150 84640
rect 146510 84490 147130 84500
rect 146100 84390 146160 84420
rect 146610 84360 146970 84420
rect 36000 84350 41400 84360
rect 146100 84270 146160 84300
rect 146300 84230 146420 84290
rect 146420 84220 146480 84230
rect 36020 84210 36100 84220
rect 36200 84210 36280 84220
rect 36380 84210 36460 84220
rect 36560 84210 36640 84220
rect 36740 84210 36820 84220
rect 36920 84210 37000 84220
rect 37100 84210 37180 84220
rect 37280 84210 37360 84220
rect 37460 84210 37540 84220
rect 37640 84210 37720 84220
rect 37820 84210 37900 84220
rect 38000 84210 38080 84220
rect 38180 84210 38260 84220
rect 38360 84210 38440 84220
rect 38540 84210 38620 84220
rect 38720 84210 38800 84220
rect 38900 84210 38980 84220
rect 39080 84210 39160 84220
rect 39260 84210 39340 84220
rect 39440 84210 39520 84220
rect 39620 84210 39700 84220
rect 39800 84210 39880 84220
rect 39980 84210 40060 84220
rect 40160 84210 40240 84220
rect 40340 84210 40420 84220
rect 40520 84210 40600 84220
rect 40700 84210 40780 84220
rect 40880 84210 40960 84220
rect 41060 84210 41140 84220
rect 41240 84210 41320 84220
rect 146420 84210 147050 84220
rect 36100 84130 36110 84210
rect 36280 84130 36290 84210
rect 36460 84130 36470 84210
rect 36640 84130 36650 84210
rect 36820 84130 36830 84210
rect 37000 84130 37010 84210
rect 37180 84130 37190 84210
rect 37360 84130 37370 84210
rect 37540 84130 37550 84210
rect 37720 84130 37730 84210
rect 37900 84130 37910 84210
rect 38080 84130 38090 84210
rect 38260 84130 38270 84210
rect 38440 84130 38450 84210
rect 38620 84130 38630 84210
rect 38800 84130 38810 84210
rect 38980 84130 38990 84210
rect 39160 84130 39170 84210
rect 39340 84130 39350 84210
rect 39520 84130 39530 84210
rect 39700 84130 39710 84210
rect 39880 84130 39890 84210
rect 40060 84130 40070 84210
rect 40240 84130 40250 84210
rect 40420 84130 40430 84210
rect 40600 84130 40610 84210
rect 40780 84130 40790 84210
rect 40960 84130 40970 84210
rect 41140 84130 41150 84210
rect 41320 84130 41330 84210
rect 146420 84205 146480 84210
rect 146420 84195 147090 84205
rect 146100 84150 146160 84180
rect 146420 84110 146480 84195
rect 146100 84030 146160 84060
rect 146300 83970 146420 84030
rect 146420 83945 146480 83970
rect 146530 83960 146540 84130
rect 146610 84100 146970 84160
rect 147090 84145 147100 84195
rect 146530 83950 147140 83960
rect 36020 83910 36100 83920
rect 36200 83910 36280 83920
rect 36380 83910 36460 83920
rect 36560 83910 36640 83920
rect 36740 83910 36820 83920
rect 36920 83910 37000 83920
rect 37100 83910 37180 83920
rect 37280 83910 37360 83920
rect 37460 83910 37540 83920
rect 37640 83910 37720 83920
rect 37820 83910 37900 83920
rect 38000 83910 38080 83920
rect 38180 83910 38260 83920
rect 38360 83910 38440 83920
rect 38540 83910 38620 83920
rect 38720 83910 38800 83920
rect 38900 83910 38980 83920
rect 39080 83910 39160 83920
rect 39260 83910 39340 83920
rect 39440 83910 39520 83920
rect 39620 83910 39700 83920
rect 39800 83910 39880 83920
rect 39980 83910 40060 83920
rect 40160 83910 40240 83920
rect 40340 83910 40420 83920
rect 40520 83910 40600 83920
rect 40700 83910 40780 83920
rect 40880 83910 40960 83920
rect 41060 83910 41140 83920
rect 41240 83910 41320 83920
rect 146100 83910 146160 83940
rect 146420 83935 147090 83945
rect 36100 83830 36110 83910
rect 36280 83830 36290 83910
rect 36460 83830 36470 83910
rect 36640 83830 36650 83910
rect 36820 83830 36830 83910
rect 37000 83830 37010 83910
rect 37180 83830 37190 83910
rect 37360 83830 37370 83910
rect 37540 83830 37550 83910
rect 37720 83830 37730 83910
rect 37900 83830 37910 83910
rect 38080 83830 38090 83910
rect 38260 83830 38270 83910
rect 38440 83830 38450 83910
rect 38620 83830 38630 83910
rect 38800 83830 38810 83910
rect 38980 83830 38990 83910
rect 39160 83830 39170 83910
rect 39340 83830 39350 83910
rect 39520 83830 39530 83910
rect 39700 83830 39710 83910
rect 39880 83830 39890 83910
rect 40060 83830 40070 83910
rect 40240 83830 40250 83910
rect 40420 83830 40430 83910
rect 40600 83830 40610 83910
rect 40780 83830 40790 83910
rect 40960 83830 40970 83910
rect 41140 83830 41150 83910
rect 41320 83830 41330 83910
rect 146420 83850 146480 83935
rect 146610 83840 146970 83900
rect 147090 83885 147100 83935
rect 146100 83790 146160 83820
rect 36000 83770 41400 83780
rect 146300 83710 146420 83770
rect 146420 83700 146480 83710
rect 146100 83670 146160 83700
rect 146420 83690 147050 83700
rect 146420 83685 146480 83690
rect 146420 83675 147090 83685
rect 36020 83590 36100 83600
rect 36200 83590 36280 83600
rect 36380 83590 36460 83600
rect 36560 83590 36640 83600
rect 36740 83590 36820 83600
rect 36920 83590 37000 83600
rect 37100 83590 37180 83600
rect 37280 83590 37360 83600
rect 37460 83590 37540 83600
rect 37640 83590 37720 83600
rect 37820 83590 37900 83600
rect 38000 83590 38080 83600
rect 38180 83590 38260 83600
rect 38360 83590 38440 83600
rect 38540 83590 38620 83600
rect 38720 83590 38800 83600
rect 38900 83590 38980 83600
rect 39080 83590 39160 83600
rect 39260 83590 39340 83600
rect 39440 83590 39520 83600
rect 39620 83590 39700 83600
rect 39800 83590 39880 83600
rect 39980 83590 40060 83600
rect 40160 83590 40240 83600
rect 40340 83590 40420 83600
rect 40520 83590 40600 83600
rect 40700 83590 40780 83600
rect 40880 83590 40960 83600
rect 41060 83590 41140 83600
rect 41240 83590 41320 83600
rect 146420 83590 146480 83675
rect 36100 83510 36110 83590
rect 36280 83510 36290 83590
rect 36460 83510 36470 83590
rect 36640 83510 36650 83590
rect 36820 83510 36830 83590
rect 37000 83510 37010 83590
rect 37180 83510 37190 83590
rect 37360 83510 37370 83590
rect 37540 83510 37550 83590
rect 37720 83510 37730 83590
rect 37900 83510 37910 83590
rect 38080 83510 38090 83590
rect 38260 83510 38270 83590
rect 38440 83510 38450 83590
rect 38620 83510 38630 83590
rect 38800 83510 38810 83590
rect 38980 83510 38990 83590
rect 39160 83510 39170 83590
rect 39340 83510 39350 83590
rect 39520 83510 39530 83590
rect 39700 83510 39710 83590
rect 39880 83510 39890 83590
rect 40060 83510 40070 83590
rect 40240 83510 40250 83590
rect 40420 83510 40430 83590
rect 40600 83510 40610 83590
rect 40780 83510 40790 83590
rect 40960 83510 40970 83590
rect 41140 83510 41150 83590
rect 41320 83510 41330 83590
rect 146100 83550 146160 83580
rect 36000 83425 36040 83435
rect 36140 83425 36220 83435
rect 36320 83425 36400 83435
rect 36500 83425 36580 83435
rect 36680 83425 36760 83435
rect 36860 83425 36940 83435
rect 37040 83425 37120 83435
rect 37220 83425 37300 83435
rect 37400 83425 37480 83435
rect 37580 83425 37660 83435
rect 37760 83425 37840 83435
rect 40160 83430 40240 83440
rect 40340 83430 40420 83440
rect 40520 83430 40600 83440
rect 40700 83430 40780 83440
rect 40880 83430 40960 83440
rect 41060 83430 41140 83440
rect 41240 83430 41320 83440
rect 146100 83430 146160 83460
rect 146300 83450 146420 83510
rect 36040 83345 36050 83425
rect 36220 83345 36230 83425
rect 36400 83345 36410 83425
rect 36580 83345 36590 83425
rect 36760 83345 36770 83425
rect 36940 83345 36950 83425
rect 37120 83345 37130 83425
rect 37300 83345 37310 83425
rect 37480 83345 37490 83425
rect 37660 83345 37670 83425
rect 37840 83345 37850 83425
rect 40240 83350 40250 83430
rect 40420 83350 40430 83430
rect 40600 83350 40610 83430
rect 40780 83350 40790 83430
rect 40960 83350 40970 83430
rect 41140 83350 41150 83430
rect 41320 83350 41330 83430
rect 146420 83425 146480 83450
rect 146530 83440 146540 83610
rect 146610 83580 146970 83640
rect 147090 83625 147100 83675
rect 146530 83430 147140 83440
rect 146420 83415 147090 83425
rect 146100 83310 146160 83340
rect 146420 83330 146480 83415
rect 146610 83320 146970 83380
rect 147090 83365 147100 83415
rect 36020 83270 36100 83280
rect 36200 83270 36280 83280
rect 36380 83270 36460 83280
rect 36560 83270 36640 83280
rect 36740 83270 36820 83280
rect 36920 83270 37000 83280
rect 37100 83270 37180 83280
rect 37280 83270 37360 83280
rect 37460 83270 37540 83280
rect 37640 83270 37720 83280
rect 37820 83270 37900 83280
rect 38000 83270 38080 83280
rect 38180 83270 38260 83280
rect 38360 83270 38440 83280
rect 38540 83270 38620 83280
rect 38720 83270 38800 83280
rect 38900 83270 38980 83280
rect 39080 83270 39160 83280
rect 39260 83270 39340 83280
rect 39440 83270 39520 83280
rect 39620 83270 39700 83280
rect 39800 83270 39880 83280
rect 39980 83270 40060 83280
rect 40160 83270 40240 83280
rect 40340 83270 40420 83280
rect 40520 83270 40600 83280
rect 40700 83270 40780 83280
rect 40880 83270 40960 83280
rect 41060 83270 41140 83280
rect 41240 83270 41320 83280
rect 36100 83190 36110 83270
rect 36280 83190 36290 83270
rect 36460 83190 36470 83270
rect 36640 83190 36650 83270
rect 36820 83190 36830 83270
rect 37000 83190 37010 83270
rect 37180 83190 37190 83270
rect 37360 83190 37370 83270
rect 37540 83190 37550 83270
rect 37720 83190 37730 83270
rect 37900 83190 37910 83270
rect 38080 83190 38090 83270
rect 38260 83190 38270 83270
rect 38440 83190 38450 83270
rect 38620 83190 38630 83270
rect 38800 83190 38810 83270
rect 38980 83190 38990 83270
rect 39160 83190 39170 83270
rect 39340 83190 39350 83270
rect 39520 83190 39530 83270
rect 39700 83190 39710 83270
rect 39880 83190 39890 83270
rect 40060 83190 40070 83270
rect 40240 83190 40250 83270
rect 40420 83190 40430 83270
rect 40600 83190 40610 83270
rect 40780 83190 40790 83270
rect 40960 83190 40970 83270
rect 41140 83190 41150 83270
rect 41320 83190 41330 83270
rect 146100 83190 146160 83220
rect 36000 83090 41400 83100
rect 146100 83070 146160 83100
rect 36020 82950 36100 82960
rect 36200 82950 36280 82960
rect 36380 82950 36460 82960
rect 36560 82950 36640 82960
rect 36740 82950 36820 82960
rect 36920 82950 37000 82960
rect 37100 82950 37180 82960
rect 37280 82950 37360 82960
rect 37460 82950 37540 82960
rect 37640 82950 37720 82960
rect 37820 82950 37900 82960
rect 38000 82950 38080 82960
rect 38180 82950 38260 82960
rect 38360 82950 38440 82960
rect 38540 82950 38620 82960
rect 38720 82950 38800 82960
rect 38900 82950 38980 82960
rect 39080 82950 39160 82960
rect 39260 82950 39340 82960
rect 39440 82950 39520 82960
rect 39620 82950 39700 82960
rect 39800 82950 39880 82960
rect 39980 82950 40060 82960
rect 40160 82950 40240 82960
rect 40340 82950 40420 82960
rect 40520 82950 40600 82960
rect 40700 82950 40780 82960
rect 40880 82950 40960 82960
rect 41060 82950 41140 82960
rect 41240 82950 41320 82960
rect 146100 82950 146160 82980
rect 36100 82870 36110 82950
rect 36280 82870 36290 82950
rect 36460 82870 36470 82950
rect 36640 82870 36650 82950
rect 36820 82870 36830 82950
rect 37000 82870 37010 82950
rect 37180 82870 37190 82950
rect 37360 82870 37370 82950
rect 37540 82870 37550 82950
rect 37720 82870 37730 82950
rect 37900 82870 37910 82950
rect 38080 82870 38090 82950
rect 38260 82870 38270 82950
rect 38440 82870 38450 82950
rect 38620 82870 38630 82950
rect 38800 82870 38810 82950
rect 38980 82870 38990 82950
rect 39160 82870 39170 82950
rect 39340 82870 39350 82950
rect 39520 82870 39530 82950
rect 39700 82870 39710 82950
rect 39880 82870 39890 82950
rect 40060 82870 40070 82950
rect 40240 82870 40250 82950
rect 40420 82870 40430 82950
rect 40600 82870 40610 82950
rect 40780 82870 40790 82950
rect 40960 82870 40970 82950
rect 41140 82870 41150 82950
rect 41320 82870 41330 82950
rect 146100 82830 146160 82860
rect 146100 82710 146160 82740
rect 36020 82650 36100 82660
rect 36200 82650 36280 82660
rect 36380 82650 36460 82660
rect 36560 82650 36640 82660
rect 36740 82650 36820 82660
rect 36920 82650 37000 82660
rect 37100 82650 37180 82660
rect 37280 82650 37360 82660
rect 37460 82650 37540 82660
rect 37640 82650 37720 82660
rect 37820 82650 37900 82660
rect 38000 82650 38080 82660
rect 38180 82650 38260 82660
rect 38360 82650 38440 82660
rect 38540 82650 38620 82660
rect 38720 82650 38800 82660
rect 38900 82650 38980 82660
rect 39080 82650 39160 82660
rect 39260 82650 39340 82660
rect 39440 82650 39520 82660
rect 39620 82650 39700 82660
rect 39800 82650 39880 82660
rect 39980 82650 40060 82660
rect 40160 82650 40240 82660
rect 40340 82650 40420 82660
rect 40520 82650 40600 82660
rect 40700 82650 40780 82660
rect 40880 82650 40960 82660
rect 41060 82650 41140 82660
rect 41240 82650 41320 82660
rect 36100 82570 36110 82650
rect 36280 82570 36290 82650
rect 36460 82570 36470 82650
rect 36640 82570 36650 82650
rect 36820 82570 36830 82650
rect 37000 82570 37010 82650
rect 37180 82570 37190 82650
rect 37360 82570 37370 82650
rect 37540 82570 37550 82650
rect 37720 82570 37730 82650
rect 37900 82570 37910 82650
rect 38080 82570 38090 82650
rect 38260 82570 38270 82650
rect 38440 82570 38450 82650
rect 38620 82570 38630 82650
rect 38800 82570 38810 82650
rect 38980 82570 38990 82650
rect 39160 82570 39170 82650
rect 39340 82570 39350 82650
rect 39520 82570 39530 82650
rect 39700 82570 39710 82650
rect 39880 82570 39890 82650
rect 40060 82570 40070 82650
rect 40240 82570 40250 82650
rect 40420 82570 40430 82650
rect 40600 82570 40610 82650
rect 40780 82570 40790 82650
rect 40960 82570 40970 82650
rect 41140 82570 41150 82650
rect 41320 82570 41330 82650
rect 146100 82590 146160 82620
rect 36000 82510 41400 82520
rect 146100 82470 146160 82500
rect 146100 82350 146160 82380
rect 36020 82330 36100 82340
rect 36200 82330 36280 82340
rect 36380 82330 36460 82340
rect 36560 82330 36640 82340
rect 36740 82330 36820 82340
rect 36920 82330 37000 82340
rect 37100 82330 37180 82340
rect 37280 82330 37360 82340
rect 37460 82330 37540 82340
rect 37640 82330 37720 82340
rect 37820 82330 37900 82340
rect 38000 82330 38080 82340
rect 38180 82330 38260 82340
rect 38360 82330 38440 82340
rect 38540 82330 38620 82340
rect 38720 82330 38800 82340
rect 38900 82330 38980 82340
rect 39080 82330 39160 82340
rect 39260 82330 39340 82340
rect 39440 82330 39520 82340
rect 39620 82330 39700 82340
rect 39800 82330 39880 82340
rect 39980 82330 40060 82340
rect 40160 82330 40240 82340
rect 40340 82330 40420 82340
rect 40520 82330 40600 82340
rect 40700 82330 40780 82340
rect 40880 82330 40960 82340
rect 41060 82330 41140 82340
rect 41240 82330 41320 82340
rect 36100 82250 36110 82330
rect 36280 82250 36290 82330
rect 36460 82250 36470 82330
rect 36640 82250 36650 82330
rect 36820 82250 36830 82330
rect 37000 82250 37010 82330
rect 37180 82250 37190 82330
rect 37360 82250 37370 82330
rect 37540 82250 37550 82330
rect 37720 82250 37730 82330
rect 37900 82250 37910 82330
rect 38080 82250 38090 82330
rect 38260 82250 38270 82330
rect 38440 82250 38450 82330
rect 38620 82250 38630 82330
rect 38800 82250 38810 82330
rect 38980 82250 38990 82330
rect 39160 82250 39170 82330
rect 39340 82250 39350 82330
rect 39520 82250 39530 82330
rect 39700 82250 39710 82330
rect 39880 82250 39890 82330
rect 40060 82250 40070 82330
rect 40240 82250 40250 82330
rect 40420 82250 40430 82330
rect 40600 82250 40610 82330
rect 40780 82250 40790 82330
rect 40960 82250 40970 82330
rect 41140 82250 41150 82330
rect 41320 82250 41330 82330
rect 146100 82230 146160 82260
rect 36000 82165 36040 82175
rect 36140 82165 36220 82175
rect 36320 82165 36400 82175
rect 36500 82165 36580 82175
rect 36680 82165 36760 82175
rect 36860 82165 36940 82175
rect 37040 82165 37120 82175
rect 37220 82165 37300 82175
rect 37400 82165 37480 82175
rect 37580 82165 37660 82175
rect 37760 82165 37840 82175
rect 40160 82170 40240 82180
rect 40340 82170 40420 82180
rect 40520 82170 40600 82180
rect 40700 82170 40780 82180
rect 40880 82170 40960 82180
rect 41060 82170 41140 82180
rect 41240 82170 41320 82180
rect 36040 82085 36050 82165
rect 36220 82085 36230 82165
rect 36400 82085 36410 82165
rect 36580 82085 36590 82165
rect 36760 82085 36770 82165
rect 36940 82085 36950 82165
rect 37120 82085 37130 82165
rect 37300 82085 37310 82165
rect 37480 82085 37490 82165
rect 37660 82085 37670 82165
rect 37840 82085 37850 82165
rect 40240 82090 40250 82170
rect 40420 82090 40430 82170
rect 40600 82090 40610 82170
rect 40780 82090 40790 82170
rect 40960 82090 40970 82170
rect 41140 82090 41150 82170
rect 41320 82090 41330 82170
rect 146100 82110 146160 82140
rect 36020 82010 36100 82020
rect 36200 82010 36280 82020
rect 36380 82010 36460 82020
rect 36560 82010 36640 82020
rect 36740 82010 36820 82020
rect 36920 82010 37000 82020
rect 37100 82010 37180 82020
rect 37280 82010 37360 82020
rect 37460 82010 37540 82020
rect 37640 82010 37720 82020
rect 37820 82010 37900 82020
rect 38000 82010 38080 82020
rect 38180 82010 38260 82020
rect 38360 82010 38440 82020
rect 38540 82010 38620 82020
rect 38720 82010 38800 82020
rect 38900 82010 38980 82020
rect 39080 82010 39160 82020
rect 39260 82010 39340 82020
rect 39440 82010 39520 82020
rect 39620 82010 39700 82020
rect 39800 82010 39880 82020
rect 39980 82010 40060 82020
rect 40160 82010 40240 82020
rect 40340 82010 40420 82020
rect 40520 82010 40600 82020
rect 40700 82010 40780 82020
rect 40880 82010 40960 82020
rect 41060 82010 41140 82020
rect 41240 82010 41320 82020
rect 36100 81930 36110 82010
rect 36280 81930 36290 82010
rect 36460 81930 36470 82010
rect 36640 81930 36650 82010
rect 36820 81930 36830 82010
rect 37000 81930 37010 82010
rect 37180 81930 37190 82010
rect 37360 81930 37370 82010
rect 37540 81930 37550 82010
rect 37720 81930 37730 82010
rect 37900 81930 37910 82010
rect 38080 81930 38090 82010
rect 38260 81930 38270 82010
rect 38440 81930 38450 82010
rect 38620 81930 38630 82010
rect 38800 81930 38810 82010
rect 38980 81930 38990 82010
rect 39160 81930 39170 82010
rect 39340 81930 39350 82010
rect 39520 81930 39530 82010
rect 39700 81930 39710 82010
rect 39880 81930 39890 82010
rect 40060 81930 40070 82010
rect 40240 81930 40250 82010
rect 40420 81930 40430 82010
rect 40600 81930 40610 82010
rect 40780 81930 40790 82010
rect 40960 81930 40970 82010
rect 41140 81930 41150 82010
rect 41320 81930 41330 82010
rect 146100 81990 146160 82020
rect 36000 81830 41400 81840
rect 46660 81760 47160 81940
rect 146100 81870 146160 81900
rect 146100 81750 146160 81780
rect 36020 81690 36100 81700
rect 36200 81690 36280 81700
rect 36380 81690 36460 81700
rect 36560 81690 36640 81700
rect 36740 81690 36820 81700
rect 36920 81690 37000 81700
rect 37100 81690 37180 81700
rect 37280 81690 37360 81700
rect 37460 81690 37540 81700
rect 37640 81690 37720 81700
rect 37820 81690 37900 81700
rect 38000 81690 38080 81700
rect 38180 81690 38260 81700
rect 38360 81690 38440 81700
rect 38540 81690 38620 81700
rect 38720 81690 38800 81700
rect 38900 81690 38980 81700
rect 39080 81690 39160 81700
rect 39260 81690 39340 81700
rect 39440 81690 39520 81700
rect 39620 81690 39700 81700
rect 39800 81690 39880 81700
rect 39980 81690 40060 81700
rect 40160 81690 40240 81700
rect 40340 81690 40420 81700
rect 40520 81690 40600 81700
rect 40700 81690 40780 81700
rect 40880 81690 40960 81700
rect 41060 81690 41140 81700
rect 41240 81690 41320 81700
rect 36100 81610 36110 81690
rect 36280 81610 36290 81690
rect 36460 81610 36470 81690
rect 36640 81610 36650 81690
rect 36820 81610 36830 81690
rect 37000 81610 37010 81690
rect 37180 81610 37190 81690
rect 37360 81610 37370 81690
rect 37540 81610 37550 81690
rect 37720 81610 37730 81690
rect 37900 81610 37910 81690
rect 38080 81610 38090 81690
rect 38260 81610 38270 81690
rect 38440 81610 38450 81690
rect 38620 81610 38630 81690
rect 38800 81610 38810 81690
rect 38980 81610 38990 81690
rect 39160 81610 39170 81690
rect 39340 81610 39350 81690
rect 39520 81610 39530 81690
rect 39700 81610 39710 81690
rect 39880 81610 39890 81690
rect 40060 81610 40070 81690
rect 40240 81610 40250 81690
rect 40420 81610 40430 81690
rect 40600 81610 40610 81690
rect 40780 81610 40790 81690
rect 40960 81610 40970 81690
rect 41140 81610 41150 81690
rect 41320 81610 41330 81690
rect 146100 81630 146160 81660
rect 146100 81510 146160 81540
rect 36020 81390 36100 81400
rect 36200 81390 36280 81400
rect 36380 81390 36460 81400
rect 36560 81390 36640 81400
rect 36740 81390 36820 81400
rect 36920 81390 37000 81400
rect 37100 81390 37180 81400
rect 37280 81390 37360 81400
rect 37460 81390 37540 81400
rect 37640 81390 37720 81400
rect 37820 81390 37900 81400
rect 38000 81390 38080 81400
rect 38180 81390 38260 81400
rect 38360 81390 38440 81400
rect 38540 81390 38620 81400
rect 38720 81390 38800 81400
rect 38900 81390 38980 81400
rect 39080 81390 39160 81400
rect 39260 81390 39340 81400
rect 39440 81390 39520 81400
rect 39620 81390 39700 81400
rect 39800 81390 39880 81400
rect 39980 81390 40060 81400
rect 40160 81390 40240 81400
rect 40340 81390 40420 81400
rect 40520 81390 40600 81400
rect 40700 81390 40780 81400
rect 40880 81390 40960 81400
rect 41060 81390 41140 81400
rect 41240 81390 41320 81400
rect 146100 81390 146160 81420
rect 36100 81310 36110 81390
rect 36280 81310 36290 81390
rect 36460 81310 36470 81390
rect 36640 81310 36650 81390
rect 36820 81310 36830 81390
rect 37000 81310 37010 81390
rect 37180 81310 37190 81390
rect 37360 81310 37370 81390
rect 37540 81310 37550 81390
rect 37720 81310 37730 81390
rect 37900 81310 37910 81390
rect 38080 81310 38090 81390
rect 38260 81310 38270 81390
rect 38440 81310 38450 81390
rect 38620 81310 38630 81390
rect 38800 81310 38810 81390
rect 38980 81310 38990 81390
rect 39160 81310 39170 81390
rect 39340 81310 39350 81390
rect 39520 81310 39530 81390
rect 39700 81310 39710 81390
rect 39880 81310 39890 81390
rect 40060 81310 40070 81390
rect 40240 81310 40250 81390
rect 40420 81310 40430 81390
rect 40600 81310 40610 81390
rect 40780 81310 40790 81390
rect 40960 81310 40970 81390
rect 41140 81310 41150 81390
rect 41320 81310 41330 81390
rect 146100 81270 146160 81300
rect 36000 81250 41400 81260
rect 146100 81150 146160 81180
rect 36020 81070 36100 81080
rect 36200 81070 36280 81080
rect 36380 81070 36460 81080
rect 36560 81070 36640 81080
rect 36740 81070 36820 81080
rect 36920 81070 37000 81080
rect 37100 81070 37180 81080
rect 37280 81070 37360 81080
rect 37460 81070 37540 81080
rect 37640 81070 37720 81080
rect 37820 81070 37900 81080
rect 38000 81070 38080 81080
rect 38180 81070 38260 81080
rect 38360 81070 38440 81080
rect 38540 81070 38620 81080
rect 38720 81070 38800 81080
rect 38900 81070 38980 81080
rect 39080 81070 39160 81080
rect 39260 81070 39340 81080
rect 39440 81070 39520 81080
rect 39620 81070 39700 81080
rect 39800 81070 39880 81080
rect 39980 81070 40060 81080
rect 40160 81070 40240 81080
rect 40340 81070 40420 81080
rect 40520 81070 40600 81080
rect 40700 81070 40780 81080
rect 40880 81070 40960 81080
rect 41060 81070 41140 81080
rect 41240 81070 41320 81080
rect 36100 80990 36110 81070
rect 36280 80990 36290 81070
rect 36460 80990 36470 81070
rect 36640 80990 36650 81070
rect 36820 80990 36830 81070
rect 37000 80990 37010 81070
rect 37180 80990 37190 81070
rect 37360 80990 37370 81070
rect 37540 80990 37550 81070
rect 37720 80990 37730 81070
rect 37900 80990 37910 81070
rect 38080 80990 38090 81070
rect 38260 80990 38270 81070
rect 38440 80990 38450 81070
rect 38620 80990 38630 81070
rect 38800 80990 38810 81070
rect 38980 80990 38990 81070
rect 39160 80990 39170 81070
rect 39340 80990 39350 81070
rect 39520 80990 39530 81070
rect 39700 80990 39710 81070
rect 39880 80990 39890 81070
rect 40060 80990 40070 81070
rect 40240 80990 40250 81070
rect 40420 80990 40430 81070
rect 40600 80990 40610 81070
rect 40780 80990 40790 81070
rect 40960 80990 40970 81070
rect 41140 80990 41150 81070
rect 41320 80990 41330 81070
rect 146100 81030 146160 81060
rect 40160 80910 40240 80920
rect 40340 80910 40420 80920
rect 40520 80910 40600 80920
rect 40700 80910 40780 80920
rect 40880 80910 40960 80920
rect 41060 80910 41140 80920
rect 41240 80910 41320 80920
rect 146100 80910 146160 80940
rect 36000 80900 36040 80910
rect 36140 80900 36220 80910
rect 36320 80900 36400 80910
rect 36500 80900 36580 80910
rect 36680 80900 36760 80910
rect 36860 80900 36940 80910
rect 37040 80900 37120 80910
rect 37220 80900 37300 80910
rect 37400 80900 37480 80910
rect 37580 80900 37660 80910
rect 37760 80900 37840 80910
rect 36040 80820 36050 80900
rect 36220 80820 36230 80900
rect 36400 80820 36410 80900
rect 36580 80820 36590 80900
rect 36760 80820 36770 80900
rect 36940 80820 36950 80900
rect 37120 80820 37130 80900
rect 37300 80820 37310 80900
rect 37480 80820 37490 80900
rect 37660 80820 37670 80900
rect 37840 80820 37850 80900
rect 40240 80830 40250 80910
rect 40420 80830 40430 80910
rect 40600 80830 40610 80910
rect 40780 80830 40790 80910
rect 40960 80830 40970 80910
rect 41140 80830 41150 80910
rect 41320 80830 41330 80910
rect 146100 80790 146160 80820
rect 36020 80750 36100 80760
rect 36200 80750 36280 80760
rect 36380 80750 36460 80760
rect 36560 80750 36640 80760
rect 36740 80750 36820 80760
rect 36920 80750 37000 80760
rect 37100 80750 37180 80760
rect 37280 80750 37360 80760
rect 37460 80750 37540 80760
rect 37640 80750 37720 80760
rect 37820 80750 37900 80760
rect 38000 80750 38080 80760
rect 38180 80750 38260 80760
rect 38360 80750 38440 80760
rect 38540 80750 38620 80760
rect 38720 80750 38800 80760
rect 38900 80750 38980 80760
rect 39080 80750 39160 80760
rect 39260 80750 39340 80760
rect 39440 80750 39520 80760
rect 39620 80750 39700 80760
rect 39800 80750 39880 80760
rect 39980 80750 40060 80760
rect 40160 80750 40240 80760
rect 40340 80750 40420 80760
rect 40520 80750 40600 80760
rect 40700 80750 40780 80760
rect 40880 80750 40960 80760
rect 41060 80750 41140 80760
rect 41240 80750 41320 80760
rect 36100 80670 36110 80750
rect 36280 80670 36290 80750
rect 36460 80670 36470 80750
rect 36640 80670 36650 80750
rect 36820 80670 36830 80750
rect 37000 80670 37010 80750
rect 37180 80670 37190 80750
rect 37360 80670 37370 80750
rect 37540 80670 37550 80750
rect 37720 80670 37730 80750
rect 37900 80670 37910 80750
rect 38080 80670 38090 80750
rect 38260 80670 38270 80750
rect 38440 80670 38450 80750
rect 38620 80670 38630 80750
rect 38800 80670 38810 80750
rect 38980 80670 38990 80750
rect 39160 80670 39170 80750
rect 39340 80670 39350 80750
rect 39520 80670 39530 80750
rect 39700 80670 39710 80750
rect 39880 80670 39890 80750
rect 40060 80670 40070 80750
rect 40240 80670 40250 80750
rect 40420 80670 40430 80750
rect 40600 80670 40610 80750
rect 40780 80670 40790 80750
rect 40960 80670 40970 80750
rect 41140 80670 41150 80750
rect 41320 80670 41330 80750
rect 146100 80670 146160 80700
rect 36000 80570 41400 80580
rect 146100 80550 146160 80580
rect 36020 80430 36100 80440
rect 36200 80430 36280 80440
rect 36380 80430 36460 80440
rect 36560 80430 36640 80440
rect 36740 80430 36820 80440
rect 36920 80430 37000 80440
rect 37100 80430 37180 80440
rect 37280 80430 37360 80440
rect 37460 80430 37540 80440
rect 37640 80430 37720 80440
rect 37820 80430 37900 80440
rect 38000 80430 38080 80440
rect 38180 80430 38260 80440
rect 38360 80430 38440 80440
rect 38540 80430 38620 80440
rect 38720 80430 38800 80440
rect 38900 80430 38980 80440
rect 39080 80430 39160 80440
rect 39260 80430 39340 80440
rect 39440 80430 39520 80440
rect 39620 80430 39700 80440
rect 39800 80430 39880 80440
rect 39980 80430 40060 80440
rect 40160 80430 40240 80440
rect 40340 80430 40420 80440
rect 40520 80430 40600 80440
rect 40700 80430 40780 80440
rect 40880 80430 40960 80440
rect 41060 80430 41140 80440
rect 41240 80430 41320 80440
rect 146100 80430 146160 80460
rect 36100 80350 36110 80430
rect 36280 80350 36290 80430
rect 36460 80350 36470 80430
rect 36640 80350 36650 80430
rect 36820 80350 36830 80430
rect 37000 80350 37010 80430
rect 37180 80350 37190 80430
rect 37360 80350 37370 80430
rect 37540 80350 37550 80430
rect 37720 80350 37730 80430
rect 37900 80350 37910 80430
rect 38080 80350 38090 80430
rect 38260 80350 38270 80430
rect 38440 80350 38450 80430
rect 38620 80350 38630 80430
rect 38800 80350 38810 80430
rect 38980 80350 38990 80430
rect 39160 80350 39170 80430
rect 39340 80350 39350 80430
rect 39520 80350 39530 80430
rect 39700 80350 39710 80430
rect 39880 80350 39890 80430
rect 40060 80350 40070 80430
rect 40240 80350 40250 80430
rect 40420 80350 40430 80430
rect 40600 80350 40610 80430
rect 40780 80350 40790 80430
rect 40960 80350 40970 80430
rect 41140 80350 41150 80430
rect 41320 80350 41330 80430
rect 146100 80310 146160 80340
rect 146100 80190 146160 80220
rect 36020 80130 36100 80140
rect 36200 80130 36280 80140
rect 36380 80130 36460 80140
rect 36560 80130 36640 80140
rect 36740 80130 36820 80140
rect 36920 80130 37000 80140
rect 37100 80130 37180 80140
rect 37280 80130 37360 80140
rect 37460 80130 37540 80140
rect 37640 80130 37720 80140
rect 37820 80130 37900 80140
rect 38000 80130 38080 80140
rect 38180 80130 38260 80140
rect 38360 80130 38440 80140
rect 38540 80130 38620 80140
rect 38720 80130 38800 80140
rect 38900 80130 38980 80140
rect 39080 80130 39160 80140
rect 39260 80130 39340 80140
rect 39440 80130 39520 80140
rect 39620 80130 39700 80140
rect 39800 80130 39880 80140
rect 39980 80130 40060 80140
rect 40160 80130 40240 80140
rect 40340 80130 40420 80140
rect 40520 80130 40600 80140
rect 40700 80130 40780 80140
rect 40880 80130 40960 80140
rect 41060 80130 41140 80140
rect 41240 80130 41320 80140
rect 36100 80050 36110 80130
rect 36280 80050 36290 80130
rect 36460 80050 36470 80130
rect 36640 80050 36650 80130
rect 36820 80050 36830 80130
rect 37000 80050 37010 80130
rect 37180 80050 37190 80130
rect 37360 80050 37370 80130
rect 37540 80050 37550 80130
rect 37720 80050 37730 80130
rect 37900 80050 37910 80130
rect 38080 80050 38090 80130
rect 38260 80050 38270 80130
rect 38440 80050 38450 80130
rect 38620 80050 38630 80130
rect 38800 80050 38810 80130
rect 38980 80050 38990 80130
rect 39160 80050 39170 80130
rect 39340 80050 39350 80130
rect 39520 80050 39530 80130
rect 39700 80050 39710 80130
rect 39880 80050 39890 80130
rect 40060 80050 40070 80130
rect 40240 80050 40250 80130
rect 40420 80050 40430 80130
rect 40600 80050 40610 80130
rect 40780 80050 40790 80130
rect 40960 80050 40970 80130
rect 41140 80050 41150 80130
rect 41320 80050 41330 80130
rect 146100 80070 146160 80100
rect 36000 79990 41400 80000
rect 146100 79950 146160 79980
rect 146100 79830 146160 79860
rect 36020 79810 36100 79820
rect 36200 79810 36280 79820
rect 36380 79810 36460 79820
rect 36560 79810 36640 79820
rect 36740 79810 36820 79820
rect 36920 79810 37000 79820
rect 37100 79810 37180 79820
rect 37280 79810 37360 79820
rect 37460 79810 37540 79820
rect 37640 79810 37720 79820
rect 37820 79810 37900 79820
rect 38000 79810 38080 79820
rect 38180 79810 38260 79820
rect 38360 79810 38440 79820
rect 38540 79810 38620 79820
rect 38720 79810 38800 79820
rect 38900 79810 38980 79820
rect 39080 79810 39160 79820
rect 39260 79810 39340 79820
rect 39440 79810 39520 79820
rect 39620 79810 39700 79820
rect 39800 79810 39880 79820
rect 39980 79810 40060 79820
rect 40160 79810 40240 79820
rect 40340 79810 40420 79820
rect 40520 79810 40600 79820
rect 40700 79810 40780 79820
rect 40880 79810 40960 79820
rect 41060 79810 41140 79820
rect 41240 79810 41320 79820
rect 36100 79730 36110 79810
rect 36280 79730 36290 79810
rect 36460 79730 36470 79810
rect 36640 79730 36650 79810
rect 36820 79730 36830 79810
rect 37000 79730 37010 79810
rect 37180 79730 37190 79810
rect 37360 79730 37370 79810
rect 37540 79730 37550 79810
rect 37720 79730 37730 79810
rect 37900 79730 37910 79810
rect 38080 79730 38090 79810
rect 38260 79730 38270 79810
rect 38440 79730 38450 79810
rect 38620 79730 38630 79810
rect 38800 79730 38810 79810
rect 38980 79730 38990 79810
rect 39160 79730 39170 79810
rect 39340 79730 39350 79810
rect 39520 79730 39530 79810
rect 39700 79730 39710 79810
rect 39880 79730 39890 79810
rect 40060 79730 40070 79810
rect 40240 79730 40250 79810
rect 40420 79730 40430 79810
rect 40600 79730 40610 79810
rect 40780 79730 40790 79810
rect 40960 79730 40970 79810
rect 41140 79730 41150 79810
rect 41320 79730 41330 79810
rect 146100 79710 146160 79740
rect 36000 79650 36040 79660
rect 36140 79650 36220 79660
rect 36320 79650 36400 79660
rect 36500 79650 36580 79660
rect 36680 79650 36760 79660
rect 36860 79650 36940 79660
rect 37040 79650 37120 79660
rect 37220 79650 37300 79660
rect 37400 79650 37480 79660
rect 37580 79650 37660 79660
rect 37760 79650 37840 79660
rect 36040 79570 36050 79650
rect 36220 79570 36230 79650
rect 36400 79570 36410 79650
rect 36580 79570 36590 79650
rect 36760 79570 36770 79650
rect 36940 79570 36950 79650
rect 37120 79570 37130 79650
rect 37300 79570 37310 79650
rect 37480 79570 37490 79650
rect 37660 79570 37670 79650
rect 37840 79570 37850 79650
rect 40160 79635 40240 79645
rect 40340 79635 40420 79645
rect 40520 79635 40600 79645
rect 40700 79635 40780 79645
rect 40880 79635 40960 79645
rect 41060 79635 41140 79645
rect 41240 79635 41320 79645
rect 40240 79555 40250 79635
rect 40420 79555 40430 79635
rect 40600 79555 40610 79635
rect 40780 79555 40790 79635
rect 40960 79555 40970 79635
rect 41140 79555 41150 79635
rect 41320 79555 41330 79635
rect 146100 79590 146160 79620
rect 36020 79490 36100 79500
rect 36200 79490 36280 79500
rect 36380 79490 36460 79500
rect 36560 79490 36640 79500
rect 36740 79490 36820 79500
rect 36920 79490 37000 79500
rect 37100 79490 37180 79500
rect 37280 79490 37360 79500
rect 37460 79490 37540 79500
rect 37640 79490 37720 79500
rect 37820 79490 37900 79500
rect 38000 79490 38080 79500
rect 38180 79490 38260 79500
rect 38360 79490 38440 79500
rect 38540 79490 38620 79500
rect 38720 79490 38800 79500
rect 38900 79490 38980 79500
rect 39080 79490 39160 79500
rect 39260 79490 39340 79500
rect 39440 79490 39520 79500
rect 39620 79490 39700 79500
rect 39800 79490 39880 79500
rect 39980 79490 40060 79500
rect 40160 79490 40240 79500
rect 40340 79490 40420 79500
rect 40520 79490 40600 79500
rect 40700 79490 40780 79500
rect 40880 79490 40960 79500
rect 41060 79490 41140 79500
rect 41240 79490 41320 79500
rect 36100 79410 36110 79490
rect 36280 79410 36290 79490
rect 36460 79410 36470 79490
rect 36640 79410 36650 79490
rect 36820 79410 36830 79490
rect 37000 79410 37010 79490
rect 37180 79410 37190 79490
rect 37360 79410 37370 79490
rect 37540 79410 37550 79490
rect 37720 79410 37730 79490
rect 37900 79410 37910 79490
rect 38080 79410 38090 79490
rect 38260 79410 38270 79490
rect 38440 79410 38450 79490
rect 38620 79410 38630 79490
rect 38800 79410 38810 79490
rect 38980 79410 38990 79490
rect 39160 79410 39170 79490
rect 39340 79410 39350 79490
rect 39520 79410 39530 79490
rect 39700 79410 39710 79490
rect 39880 79410 39890 79490
rect 40060 79410 40070 79490
rect 40240 79410 40250 79490
rect 40420 79410 40430 79490
rect 40600 79410 40610 79490
rect 40780 79410 40790 79490
rect 40960 79410 40970 79490
rect 41140 79410 41150 79490
rect 41320 79410 41330 79490
rect 146100 79470 146160 79500
rect 146100 79350 146160 79380
rect 36000 79310 41400 79320
rect 146100 79230 146160 79260
rect 36020 79170 36100 79180
rect 36200 79170 36280 79180
rect 36380 79170 36460 79180
rect 36560 79170 36640 79180
rect 36740 79170 36820 79180
rect 36920 79170 37000 79180
rect 37100 79170 37180 79180
rect 37280 79170 37360 79180
rect 37460 79170 37540 79180
rect 37640 79170 37720 79180
rect 37820 79170 37900 79180
rect 38000 79170 38080 79180
rect 38180 79170 38260 79180
rect 38360 79170 38440 79180
rect 38540 79170 38620 79180
rect 38720 79170 38800 79180
rect 38900 79170 38980 79180
rect 39080 79170 39160 79180
rect 39260 79170 39340 79180
rect 39440 79170 39520 79180
rect 39620 79170 39700 79180
rect 39800 79170 39880 79180
rect 39980 79170 40060 79180
rect 40160 79170 40240 79180
rect 40340 79170 40420 79180
rect 40520 79170 40600 79180
rect 40700 79170 40780 79180
rect 40880 79170 40960 79180
rect 41060 79170 41140 79180
rect 41240 79170 41320 79180
rect 36100 79090 36110 79170
rect 36280 79090 36290 79170
rect 36460 79090 36470 79170
rect 36640 79090 36650 79170
rect 36820 79090 36830 79170
rect 37000 79090 37010 79170
rect 37180 79090 37190 79170
rect 37360 79090 37370 79170
rect 37540 79090 37550 79170
rect 37720 79090 37730 79170
rect 37900 79090 37910 79170
rect 38080 79090 38090 79170
rect 38260 79090 38270 79170
rect 38440 79090 38450 79170
rect 38620 79090 38630 79170
rect 38800 79090 38810 79170
rect 38980 79090 38990 79170
rect 39160 79090 39170 79170
rect 39340 79090 39350 79170
rect 39520 79090 39530 79170
rect 39700 79090 39710 79170
rect 39880 79090 39890 79170
rect 40060 79090 40070 79170
rect 40240 79090 40250 79170
rect 40420 79090 40430 79170
rect 40600 79090 40610 79170
rect 40780 79090 40790 79170
rect 40960 79090 40970 79170
rect 41140 79090 41150 79170
rect 41320 79090 41330 79170
rect 146100 79110 146160 79140
rect 146100 78990 146160 79020
rect 36020 78870 36100 78880
rect 36200 78870 36280 78880
rect 36380 78870 36460 78880
rect 36560 78870 36640 78880
rect 36740 78870 36820 78880
rect 36920 78870 37000 78880
rect 37100 78870 37180 78880
rect 37280 78870 37360 78880
rect 37460 78870 37540 78880
rect 37640 78870 37720 78880
rect 37820 78870 37900 78880
rect 38000 78870 38080 78880
rect 38180 78870 38260 78880
rect 38360 78870 38440 78880
rect 38540 78870 38620 78880
rect 38720 78870 38800 78880
rect 38900 78870 38980 78880
rect 39080 78870 39160 78880
rect 39260 78870 39340 78880
rect 39440 78870 39520 78880
rect 39620 78870 39700 78880
rect 39800 78870 39880 78880
rect 39980 78870 40060 78880
rect 40160 78870 40240 78880
rect 40340 78870 40420 78880
rect 40520 78870 40600 78880
rect 40700 78870 40780 78880
rect 40880 78870 40960 78880
rect 41060 78870 41140 78880
rect 41240 78870 41320 78880
rect 146100 78870 146160 78900
rect 36100 78790 36110 78870
rect 36280 78790 36290 78870
rect 36460 78790 36470 78870
rect 36640 78790 36650 78870
rect 36820 78790 36830 78870
rect 37000 78790 37010 78870
rect 37180 78790 37190 78870
rect 37360 78790 37370 78870
rect 37540 78790 37550 78870
rect 37720 78790 37730 78870
rect 37900 78790 37910 78870
rect 38080 78790 38090 78870
rect 38260 78790 38270 78870
rect 38440 78790 38450 78870
rect 38620 78790 38630 78870
rect 38800 78790 38810 78870
rect 38980 78790 38990 78870
rect 39160 78790 39170 78870
rect 39340 78790 39350 78870
rect 39520 78790 39530 78870
rect 39700 78790 39710 78870
rect 39880 78790 39890 78870
rect 40060 78790 40070 78870
rect 40240 78790 40250 78870
rect 40420 78790 40430 78870
rect 40600 78790 40610 78870
rect 40780 78790 40790 78870
rect 40960 78790 40970 78870
rect 41140 78790 41150 78870
rect 41320 78790 41330 78870
rect 146100 78750 146160 78780
rect 36000 78730 41400 78740
rect 146100 78630 146160 78660
rect 36020 78550 36100 78560
rect 36200 78550 36280 78560
rect 36380 78550 36460 78560
rect 36560 78550 36640 78560
rect 36740 78550 36820 78560
rect 36920 78550 37000 78560
rect 37100 78550 37180 78560
rect 37280 78550 37360 78560
rect 37460 78550 37540 78560
rect 37640 78550 37720 78560
rect 37820 78550 37900 78560
rect 38000 78550 38080 78560
rect 38180 78550 38260 78560
rect 38360 78550 38440 78560
rect 38540 78550 38620 78560
rect 38720 78550 38800 78560
rect 38900 78550 38980 78560
rect 39080 78550 39160 78560
rect 39260 78550 39340 78560
rect 39440 78550 39520 78560
rect 39620 78550 39700 78560
rect 39800 78550 39880 78560
rect 39980 78550 40060 78560
rect 40160 78550 40240 78560
rect 40340 78550 40420 78560
rect 40520 78550 40600 78560
rect 40700 78550 40780 78560
rect 40880 78550 40960 78560
rect 41060 78550 41140 78560
rect 41240 78550 41320 78560
rect 36100 78470 36110 78550
rect 36280 78470 36290 78550
rect 36460 78470 36470 78550
rect 36640 78470 36650 78550
rect 36820 78470 36830 78550
rect 37000 78470 37010 78550
rect 37180 78470 37190 78550
rect 37360 78470 37370 78550
rect 37540 78470 37550 78550
rect 37720 78470 37730 78550
rect 37900 78470 37910 78550
rect 38080 78470 38090 78550
rect 38260 78470 38270 78550
rect 38440 78470 38450 78550
rect 38620 78470 38630 78550
rect 38800 78470 38810 78550
rect 38980 78470 38990 78550
rect 39160 78470 39170 78550
rect 39340 78470 39350 78550
rect 39520 78470 39530 78550
rect 39700 78470 39710 78550
rect 39880 78470 39890 78550
rect 40060 78470 40070 78550
rect 40240 78470 40250 78550
rect 40420 78470 40430 78550
rect 40600 78470 40610 78550
rect 40780 78470 40790 78550
rect 40960 78470 40970 78550
rect 41140 78470 41150 78550
rect 41320 78470 41330 78550
rect 146100 78510 146160 78540
rect 36000 78395 36040 78405
rect 36140 78395 36220 78405
rect 36320 78395 36400 78405
rect 36500 78395 36580 78405
rect 36680 78395 36760 78405
rect 36860 78395 36940 78405
rect 37040 78395 37120 78405
rect 37220 78395 37300 78405
rect 37400 78395 37480 78405
rect 37580 78395 37660 78405
rect 37760 78395 37840 78405
rect 36040 78315 36050 78395
rect 36220 78315 36230 78395
rect 36400 78315 36410 78395
rect 36580 78315 36590 78395
rect 36760 78315 36770 78395
rect 36940 78315 36950 78395
rect 37120 78315 37130 78395
rect 37300 78315 37310 78395
rect 37480 78315 37490 78395
rect 37660 78315 37670 78395
rect 37840 78315 37850 78395
rect 146100 78390 146160 78420
rect 40160 78375 40240 78385
rect 40340 78375 40420 78385
rect 40520 78375 40600 78385
rect 40700 78375 40780 78385
rect 40880 78375 40960 78385
rect 41060 78375 41140 78385
rect 41240 78375 41320 78385
rect 40240 78295 40250 78375
rect 40420 78295 40430 78375
rect 40600 78295 40610 78375
rect 40780 78295 40790 78375
rect 40960 78295 40970 78375
rect 41140 78295 41150 78375
rect 41320 78295 41330 78375
rect 146100 78270 146160 78300
rect 36020 78230 36100 78240
rect 36200 78230 36280 78240
rect 36380 78230 36460 78240
rect 36560 78230 36640 78240
rect 36740 78230 36820 78240
rect 36920 78230 37000 78240
rect 37100 78230 37180 78240
rect 37280 78230 37360 78240
rect 37460 78230 37540 78240
rect 37640 78230 37720 78240
rect 37820 78230 37900 78240
rect 38000 78230 38080 78240
rect 38180 78230 38260 78240
rect 38360 78230 38440 78240
rect 38540 78230 38620 78240
rect 38720 78230 38800 78240
rect 38900 78230 38980 78240
rect 39080 78230 39160 78240
rect 39260 78230 39340 78240
rect 39440 78230 39520 78240
rect 39620 78230 39700 78240
rect 39800 78230 39880 78240
rect 39980 78230 40060 78240
rect 40160 78230 40240 78240
rect 40340 78230 40420 78240
rect 40520 78230 40600 78240
rect 40700 78230 40780 78240
rect 40880 78230 40960 78240
rect 41060 78230 41140 78240
rect 41240 78230 41320 78240
rect 36100 78150 36110 78230
rect 36280 78150 36290 78230
rect 36460 78150 36470 78230
rect 36640 78150 36650 78230
rect 36820 78150 36830 78230
rect 37000 78150 37010 78230
rect 37180 78150 37190 78230
rect 37360 78150 37370 78230
rect 37540 78150 37550 78230
rect 37720 78150 37730 78230
rect 37900 78150 37910 78230
rect 38080 78150 38090 78230
rect 38260 78150 38270 78230
rect 38440 78150 38450 78230
rect 38620 78150 38630 78230
rect 38800 78150 38810 78230
rect 38980 78150 38990 78230
rect 39160 78150 39170 78230
rect 39340 78150 39350 78230
rect 39520 78150 39530 78230
rect 39700 78150 39710 78230
rect 39880 78150 39890 78230
rect 40060 78150 40070 78230
rect 40240 78150 40250 78230
rect 40420 78150 40430 78230
rect 40600 78150 40610 78230
rect 40780 78150 40790 78230
rect 40960 78150 40970 78230
rect 41140 78150 41150 78230
rect 41320 78150 41330 78230
rect 46555 78090 46560 78160
rect 146100 78150 146160 78180
rect 36000 78050 41400 78060
rect 36020 77910 36100 77920
rect 36200 77910 36280 77920
rect 36380 77910 36460 77920
rect 36560 77910 36640 77920
rect 36740 77910 36820 77920
rect 36920 77910 37000 77920
rect 37100 77910 37180 77920
rect 37280 77910 37360 77920
rect 37460 77910 37540 77920
rect 37640 77910 37720 77920
rect 37820 77910 37900 77920
rect 38000 77910 38080 77920
rect 38180 77910 38260 77920
rect 38360 77910 38440 77920
rect 38540 77910 38620 77920
rect 38720 77910 38800 77920
rect 38900 77910 38980 77920
rect 39080 77910 39160 77920
rect 39260 77910 39340 77920
rect 39440 77910 39520 77920
rect 39620 77910 39700 77920
rect 39800 77910 39880 77920
rect 39980 77910 40060 77920
rect 40160 77910 40240 77920
rect 40340 77910 40420 77920
rect 40520 77910 40600 77920
rect 40700 77910 40780 77920
rect 40880 77910 40960 77920
rect 41060 77910 41140 77920
rect 41240 77910 41320 77920
rect 36100 77830 36110 77910
rect 36280 77830 36290 77910
rect 36460 77830 36470 77910
rect 36640 77830 36650 77910
rect 36820 77830 36830 77910
rect 37000 77830 37010 77910
rect 37180 77830 37190 77910
rect 37360 77830 37370 77910
rect 37540 77830 37550 77910
rect 37720 77830 37730 77910
rect 37900 77830 37910 77910
rect 38080 77830 38090 77910
rect 38260 77830 38270 77910
rect 38440 77830 38450 77910
rect 38620 77830 38630 77910
rect 38800 77830 38810 77910
rect 38980 77830 38990 77910
rect 39160 77830 39170 77910
rect 39340 77830 39350 77910
rect 39520 77830 39530 77910
rect 39700 77830 39710 77910
rect 39880 77830 39890 77910
rect 40060 77830 40070 77910
rect 40240 77830 40250 77910
rect 40420 77830 40430 77910
rect 40600 77830 40610 77910
rect 40780 77830 40790 77910
rect 40960 77830 40970 77910
rect 41140 77830 41150 77910
rect 41320 77830 41330 77910
rect 46660 77860 47160 78040
rect 146100 78030 146160 78060
rect 146100 77910 146160 77940
rect 146100 77790 146160 77820
rect 146100 77670 146160 77700
rect 36020 77610 36100 77620
rect 36200 77610 36280 77620
rect 36380 77610 36460 77620
rect 36560 77610 36640 77620
rect 36740 77610 36820 77620
rect 36920 77610 37000 77620
rect 37100 77610 37180 77620
rect 37280 77610 37360 77620
rect 37460 77610 37540 77620
rect 37640 77610 37720 77620
rect 37820 77610 37900 77620
rect 38000 77610 38080 77620
rect 38180 77610 38260 77620
rect 38360 77610 38440 77620
rect 38540 77610 38620 77620
rect 38720 77610 38800 77620
rect 38900 77610 38980 77620
rect 39080 77610 39160 77620
rect 39260 77610 39340 77620
rect 39440 77610 39520 77620
rect 39620 77610 39700 77620
rect 39800 77610 39880 77620
rect 39980 77610 40060 77620
rect 40160 77610 40240 77620
rect 40340 77610 40420 77620
rect 40520 77610 40600 77620
rect 40700 77610 40780 77620
rect 40880 77610 40960 77620
rect 41060 77610 41140 77620
rect 41240 77610 41320 77620
rect 36100 77530 36110 77610
rect 36280 77530 36290 77610
rect 36460 77530 36470 77610
rect 36640 77530 36650 77610
rect 36820 77530 36830 77610
rect 37000 77530 37010 77610
rect 37180 77530 37190 77610
rect 37360 77530 37370 77610
rect 37540 77530 37550 77610
rect 37720 77530 37730 77610
rect 37900 77530 37910 77610
rect 38080 77530 38090 77610
rect 38260 77530 38270 77610
rect 38440 77530 38450 77610
rect 38620 77530 38630 77610
rect 38800 77530 38810 77610
rect 38980 77530 38990 77610
rect 39160 77530 39170 77610
rect 39340 77530 39350 77610
rect 39520 77530 39530 77610
rect 39700 77530 39710 77610
rect 39880 77530 39890 77610
rect 40060 77530 40070 77610
rect 40240 77530 40250 77610
rect 40420 77530 40430 77610
rect 40600 77530 40610 77610
rect 40780 77530 40790 77610
rect 40960 77530 40970 77610
rect 41140 77530 41150 77610
rect 41320 77530 41330 77610
rect 146100 77550 146160 77580
rect 146100 77430 146160 77460
rect 146100 77310 146160 77340
rect 36020 77200 36100 77210
rect 36200 77200 36280 77210
rect 36380 77200 36460 77210
rect 36560 77200 36640 77210
rect 36740 77200 36820 77210
rect 36920 77200 37000 77210
rect 37100 77200 37180 77210
rect 37280 77200 37360 77210
rect 37460 77200 37540 77210
rect 37640 77200 37720 77210
rect 37820 77200 37900 77210
rect 38000 77200 38080 77210
rect 38180 77200 38260 77210
rect 38360 77200 38440 77210
rect 38540 77200 38620 77210
rect 38720 77200 38800 77210
rect 38900 77200 38980 77210
rect 39080 77200 39160 77210
rect 39260 77200 39340 77210
rect 39440 77200 39520 77210
rect 39620 77200 39700 77210
rect 39800 77200 39880 77210
rect 39980 77200 40060 77210
rect 40160 77200 40240 77210
rect 40340 77200 40420 77210
rect 40520 77200 40600 77210
rect 40700 77200 40780 77210
rect 40880 77200 40960 77210
rect 41060 77200 41140 77210
rect 41240 77200 41320 77210
rect 41420 77200 41500 77210
rect 41600 77200 41680 77210
rect 36100 77120 36110 77200
rect 36280 77120 36290 77200
rect 36460 77120 36470 77200
rect 36640 77120 36650 77200
rect 36820 77120 36830 77200
rect 37000 77120 37010 77200
rect 37180 77120 37190 77200
rect 37360 77120 37370 77200
rect 37540 77120 37550 77200
rect 37720 77120 37730 77200
rect 37900 77120 37910 77200
rect 38080 77120 38090 77200
rect 38260 77120 38270 77200
rect 38440 77120 38450 77200
rect 38620 77120 38630 77200
rect 38800 77120 38810 77200
rect 38980 77120 38990 77200
rect 39160 77120 39170 77200
rect 39340 77120 39350 77200
rect 39520 77120 39530 77200
rect 39700 77120 39710 77200
rect 39880 77120 39890 77200
rect 40060 77120 40070 77200
rect 40240 77120 40250 77200
rect 40420 77120 40430 77200
rect 40600 77120 40610 77200
rect 40780 77120 40790 77200
rect 40960 77120 40970 77200
rect 41140 77120 41150 77200
rect 41320 77120 41330 77200
rect 41500 77120 41510 77200
rect 41680 77120 41690 77200
rect 146100 77190 146160 77220
rect 146100 77070 146160 77100
rect 146100 76950 146160 76980
rect 36020 76900 36100 76910
rect 36200 76900 36280 76910
rect 36380 76900 36460 76910
rect 36560 76900 36640 76910
rect 36740 76900 36820 76910
rect 36920 76900 37000 76910
rect 37100 76900 37180 76910
rect 37280 76900 37360 76910
rect 37460 76900 37540 76910
rect 37640 76900 37720 76910
rect 37820 76900 37900 76910
rect 38000 76900 38080 76910
rect 38180 76900 38260 76910
rect 38360 76900 38440 76910
rect 38540 76900 38620 76910
rect 38720 76900 38800 76910
rect 38900 76900 38980 76910
rect 39080 76900 39160 76910
rect 39260 76900 39340 76910
rect 39440 76900 39520 76910
rect 39620 76900 39700 76910
rect 39800 76900 39880 76910
rect 39980 76900 40060 76910
rect 40160 76900 40240 76910
rect 40340 76900 40420 76910
rect 40520 76900 40600 76910
rect 40700 76900 40780 76910
rect 40880 76900 40960 76910
rect 41060 76900 41140 76910
rect 41240 76900 41320 76910
rect 41420 76900 41500 76910
rect 41600 76900 41680 76910
rect 36100 76820 36110 76900
rect 36280 76820 36290 76900
rect 36460 76820 36470 76900
rect 36640 76820 36650 76900
rect 36820 76820 36830 76900
rect 37000 76820 37010 76900
rect 37180 76820 37190 76900
rect 37360 76820 37370 76900
rect 37540 76820 37550 76900
rect 37720 76820 37730 76900
rect 37900 76820 37910 76900
rect 38080 76820 38090 76900
rect 38260 76820 38270 76900
rect 38440 76820 38450 76900
rect 38620 76820 38630 76900
rect 38800 76820 38810 76900
rect 38980 76820 38990 76900
rect 39160 76820 39170 76900
rect 39340 76820 39350 76900
rect 39520 76820 39530 76900
rect 39700 76820 39710 76900
rect 39880 76820 39890 76900
rect 40060 76820 40070 76900
rect 40240 76820 40250 76900
rect 40420 76820 40430 76900
rect 40600 76820 40610 76900
rect 40780 76820 40790 76900
rect 40960 76820 40970 76900
rect 41140 76820 41150 76900
rect 41320 76820 41330 76900
rect 41500 76820 41510 76900
rect 41680 76820 41690 76900
rect 146100 76830 146160 76860
rect 146100 76710 146160 76740
rect 146100 76590 146160 76620
rect 146100 76470 146160 76500
rect 146100 76350 146160 76380
rect 19130 76200 19160 76255
rect 19250 76200 19280 76255
rect 26420 76200 26450 76255
rect 26540 76200 26570 76255
rect 146100 76230 146160 76260
rect 147580 76230 147640 76246
rect 148400 76230 148460 76246
rect 149880 76230 149940 76246
rect 152220 76210 152250 76240
rect 152340 76210 152370 76240
rect 159520 76210 159550 76240
rect 159640 76210 159670 76240
rect 163520 76210 163550 76240
rect 163640 76210 163670 76240
rect 170810 76210 170840 76240
rect 170930 76210 170960 76240
rect 152100 76180 152160 76210
rect 152220 76180 152280 76210
rect 152340 76180 152400 76210
rect 159400 76180 159460 76210
rect 159520 76180 159580 76210
rect 159640 76180 159700 76210
rect 163400 76180 163460 76210
rect 163520 76180 163580 76210
rect 163640 76180 163700 76210
rect 170690 76180 170750 76210
rect 170810 76180 170870 76210
rect 170930 76180 170990 76210
rect 146100 76110 146160 76140
rect 147580 76110 147640 76140
rect 148400 76110 148460 76140
rect 149880 76110 149940 76140
rect 152220 76060 152250 76120
rect 152340 76060 152370 76120
rect 159520 76060 159550 76120
rect 159640 76060 159670 76120
rect 163520 76060 163550 76120
rect 163640 76060 163670 76120
rect 170810 76060 170840 76120
rect 170930 76060 170960 76120
rect 146100 75990 146160 76020
rect 147580 75990 147640 76020
rect 148400 75990 148460 76020
rect 149880 75990 149940 76020
rect 18980 75940 19060 75950
rect 19160 75940 19240 75950
rect 19340 75940 19420 75950
rect 19520 75940 19600 75950
rect 19700 75940 19780 75950
rect 19880 75940 19960 75950
rect 20060 75940 20140 75950
rect 20240 75940 20320 75950
rect 20420 75940 20500 75950
rect 20600 75940 20680 75950
rect 20780 75940 20860 75950
rect 20960 75940 21040 75950
rect 21140 75940 21220 75950
rect 21320 75940 21400 75950
rect 21500 75940 21580 75950
rect 21680 75940 21760 75950
rect 21860 75940 21940 75950
rect 22040 75940 22120 75950
rect 22220 75940 22300 75950
rect 22400 75940 22480 75950
rect 22580 75940 22660 75950
rect 22760 75940 22840 75950
rect 22940 75940 23020 75950
rect 23120 75940 23200 75950
rect 23300 75940 23380 75950
rect 23480 75940 23560 75950
rect 23660 75940 23740 75950
rect 23840 75940 23920 75950
rect 24020 75940 24100 75950
rect 24200 75940 24280 75950
rect 24380 75940 24460 75950
rect 24560 75940 24640 75950
rect 24740 75940 24820 75950
rect 24920 75940 25000 75950
rect 25100 75940 25180 75950
rect 25280 75940 25360 75950
rect 25460 75940 25540 75950
rect 25640 75940 25720 75950
rect 25820 75940 25900 75950
rect 26000 75940 26080 75950
rect 26180 75940 26260 75950
rect 26360 75940 26440 75950
rect 26540 75940 26620 75950
rect 19060 75860 19070 75940
rect 19240 75860 19250 75940
rect 19420 75860 19430 75940
rect 19600 75860 19610 75940
rect 19780 75860 19790 75940
rect 19960 75860 19970 75940
rect 20140 75860 20150 75940
rect 20320 75860 20330 75940
rect 20500 75860 20510 75940
rect 20680 75860 20690 75940
rect 20860 75860 20870 75940
rect 21040 75860 21050 75940
rect 21220 75860 21230 75940
rect 21400 75860 21410 75940
rect 21580 75860 21590 75940
rect 21760 75860 21770 75940
rect 21940 75860 21950 75940
rect 22120 75860 22130 75940
rect 22300 75860 22310 75940
rect 22480 75860 22490 75940
rect 22660 75860 22670 75940
rect 22840 75860 22850 75940
rect 23020 75860 23030 75940
rect 23200 75860 23210 75940
rect 23380 75860 23390 75940
rect 23560 75860 23570 75940
rect 23740 75860 23750 75940
rect 23920 75860 23930 75940
rect 24100 75860 24110 75940
rect 24280 75860 24290 75940
rect 24460 75860 24470 75940
rect 24640 75860 24650 75940
rect 24820 75860 24830 75940
rect 25000 75860 25010 75940
rect 25180 75860 25190 75940
rect 25360 75860 25370 75940
rect 25540 75860 25550 75940
rect 25720 75860 25730 75940
rect 25900 75860 25910 75940
rect 26080 75860 26090 75940
rect 26260 75860 26270 75940
rect 26440 75860 26450 75940
rect 26620 75860 26630 75940
rect 146100 75870 146160 75900
rect 147580 75870 147640 75900
rect 148400 75870 148460 75900
rect 149880 75870 149940 75900
rect 18980 75790 19060 75800
rect 19160 75790 19240 75800
rect 19340 75790 19420 75800
rect 19520 75790 19600 75800
rect 19700 75790 19780 75800
rect 19880 75790 19960 75800
rect 20060 75790 20140 75800
rect 20240 75790 20320 75800
rect 20420 75790 20500 75800
rect 20600 75790 20680 75800
rect 20780 75790 20860 75800
rect 20960 75790 21040 75800
rect 21140 75790 21220 75800
rect 21320 75790 21400 75800
rect 21500 75790 21580 75800
rect 21680 75790 21760 75800
rect 21860 75790 21940 75800
rect 22040 75790 22120 75800
rect 22220 75790 22300 75800
rect 22400 75790 22480 75800
rect 22580 75790 22660 75800
rect 22760 75790 22840 75800
rect 22940 75790 23020 75800
rect 23120 75790 23200 75800
rect 23300 75790 23380 75800
rect 23480 75790 23560 75800
rect 23660 75790 23740 75800
rect 23840 75790 23920 75800
rect 24020 75790 24100 75800
rect 24200 75790 24280 75800
rect 24380 75790 24460 75800
rect 24560 75790 24640 75800
rect 24740 75790 24820 75800
rect 24920 75790 25000 75800
rect 25100 75790 25180 75800
rect 25280 75790 25360 75800
rect 25460 75790 25540 75800
rect 25640 75790 25720 75800
rect 25820 75790 25900 75800
rect 26000 75790 26080 75800
rect 26180 75790 26260 75800
rect 26360 75790 26440 75800
rect 26540 75790 26620 75800
rect 152080 75790 152160 75800
rect 152260 75790 152340 75800
rect 152440 75790 152520 75800
rect 152620 75790 152700 75800
rect 152800 75790 152880 75800
rect 152980 75790 153060 75800
rect 153160 75790 153240 75800
rect 153340 75790 153420 75800
rect 153520 75790 153600 75800
rect 153700 75790 153780 75800
rect 153880 75790 153960 75800
rect 154060 75790 154140 75800
rect 154240 75790 154320 75800
rect 154420 75790 154500 75800
rect 154600 75790 154680 75800
rect 154780 75790 154860 75800
rect 154960 75790 155040 75800
rect 155140 75790 155220 75800
rect 155320 75790 155400 75800
rect 155500 75790 155580 75800
rect 155680 75790 155760 75800
rect 155860 75790 155940 75800
rect 156040 75790 156120 75800
rect 156220 75790 156300 75800
rect 156400 75790 156480 75800
rect 156580 75790 156660 75800
rect 156760 75790 156840 75800
rect 156940 75790 157020 75800
rect 157120 75790 157200 75800
rect 157300 75790 157380 75800
rect 157480 75790 157560 75800
rect 157660 75790 157740 75800
rect 157840 75790 157920 75800
rect 158020 75790 158100 75800
rect 158200 75790 158280 75800
rect 158380 75790 158460 75800
rect 158560 75790 158640 75800
rect 158740 75790 158820 75800
rect 158920 75790 159000 75800
rect 159100 75790 159180 75800
rect 159280 75790 159360 75800
rect 159460 75790 159540 75800
rect 159640 75790 159720 75800
rect 163380 75790 163460 75800
rect 163560 75790 163640 75800
rect 163740 75790 163820 75800
rect 163920 75790 164000 75800
rect 164100 75790 164180 75800
rect 164280 75790 164360 75800
rect 164460 75790 164540 75800
rect 164640 75790 164720 75800
rect 164820 75790 164900 75800
rect 165000 75790 165080 75800
rect 165180 75790 165260 75800
rect 165360 75790 165440 75800
rect 165540 75790 165620 75800
rect 165720 75790 165800 75800
rect 165900 75790 165980 75800
rect 166080 75790 166160 75800
rect 166260 75790 166340 75800
rect 166440 75790 166520 75800
rect 166620 75790 166700 75800
rect 166800 75790 166880 75800
rect 166980 75790 167060 75800
rect 167160 75790 167240 75800
rect 167340 75790 167420 75800
rect 167520 75790 167600 75800
rect 167700 75790 167780 75800
rect 167880 75790 167960 75800
rect 168060 75790 168140 75800
rect 168240 75790 168320 75800
rect 168420 75790 168500 75800
rect 168600 75790 168680 75800
rect 168780 75790 168860 75800
rect 168960 75790 169040 75800
rect 169140 75790 169220 75800
rect 169320 75790 169400 75800
rect 169500 75790 169580 75800
rect 169680 75790 169760 75800
rect 169860 75790 169940 75800
rect 170040 75790 170120 75800
rect 170220 75790 170300 75800
rect 170400 75790 170480 75800
rect 170580 75790 170660 75800
rect 170760 75790 170840 75800
rect 170940 75790 171020 75800
rect 19060 75710 19070 75790
rect 19240 75710 19250 75790
rect 19420 75710 19430 75790
rect 19600 75710 19610 75790
rect 19780 75710 19790 75790
rect 19960 75710 19970 75790
rect 20140 75710 20150 75790
rect 20320 75710 20330 75790
rect 20500 75710 20510 75790
rect 20680 75710 20690 75790
rect 20860 75710 20870 75790
rect 21040 75710 21050 75790
rect 21220 75710 21230 75790
rect 21400 75710 21410 75790
rect 21580 75710 21590 75790
rect 21760 75710 21770 75790
rect 21940 75710 21950 75790
rect 22120 75710 22130 75790
rect 22300 75710 22310 75790
rect 22480 75710 22490 75790
rect 22660 75710 22670 75790
rect 22840 75710 22850 75790
rect 23020 75710 23030 75790
rect 23200 75710 23210 75790
rect 23380 75710 23390 75790
rect 23560 75710 23570 75790
rect 23740 75710 23750 75790
rect 23920 75710 23930 75790
rect 24100 75710 24110 75790
rect 24280 75710 24290 75790
rect 24460 75710 24470 75790
rect 24640 75710 24650 75790
rect 24820 75710 24830 75790
rect 25000 75710 25010 75790
rect 25180 75710 25190 75790
rect 25360 75710 25370 75790
rect 25540 75710 25550 75790
rect 25720 75710 25730 75790
rect 25900 75710 25910 75790
rect 26080 75710 26090 75790
rect 26260 75710 26270 75790
rect 26440 75710 26450 75790
rect 26620 75710 26630 75790
rect 152160 75710 152170 75790
rect 152340 75710 152350 75790
rect 152520 75710 152530 75790
rect 152700 75710 152710 75790
rect 152880 75710 152890 75790
rect 153060 75710 153070 75790
rect 153240 75710 153250 75790
rect 153420 75710 153430 75790
rect 153600 75710 153610 75790
rect 153780 75710 153790 75790
rect 153960 75710 153970 75790
rect 154140 75710 154150 75790
rect 154320 75710 154330 75790
rect 154500 75710 154510 75790
rect 154680 75710 154690 75790
rect 154860 75710 154870 75790
rect 155040 75710 155050 75790
rect 155220 75710 155230 75790
rect 155400 75710 155410 75790
rect 155580 75710 155590 75790
rect 155760 75710 155770 75790
rect 155940 75710 155950 75790
rect 156120 75710 156130 75790
rect 156300 75710 156310 75790
rect 156480 75710 156490 75790
rect 156660 75710 156670 75790
rect 156840 75710 156850 75790
rect 157020 75710 157030 75790
rect 157200 75710 157210 75790
rect 157380 75710 157390 75790
rect 157560 75710 157570 75790
rect 157740 75710 157750 75790
rect 157920 75710 157930 75790
rect 158100 75710 158110 75790
rect 158280 75710 158290 75790
rect 158460 75710 158470 75790
rect 158640 75710 158650 75790
rect 158820 75710 158830 75790
rect 159000 75710 159010 75790
rect 159180 75710 159190 75790
rect 159360 75710 159370 75790
rect 159540 75710 159550 75790
rect 159720 75710 159730 75790
rect 160430 75765 160510 75775
rect 160590 75765 160670 75775
rect 160750 75765 160830 75775
rect 160910 75765 160990 75775
rect 161070 75765 161150 75775
rect 160510 75685 160520 75765
rect 160590 75685 160600 75765
rect 160670 75685 160680 75765
rect 160750 75685 160760 75765
rect 160830 75685 160840 75765
rect 160910 75685 160920 75765
rect 160990 75685 161000 75765
rect 161070 75685 161080 75765
rect 161150 75685 161160 75765
rect 163460 75710 163470 75790
rect 163640 75710 163650 75790
rect 163820 75710 163830 75790
rect 164000 75710 164010 75790
rect 164180 75710 164190 75790
rect 164360 75710 164370 75790
rect 164540 75710 164550 75790
rect 164720 75710 164730 75790
rect 164900 75710 164910 75790
rect 165080 75710 165090 75790
rect 165260 75710 165270 75790
rect 165440 75710 165450 75790
rect 165620 75710 165630 75790
rect 165800 75710 165810 75790
rect 165980 75710 165990 75790
rect 166160 75710 166170 75790
rect 166340 75710 166350 75790
rect 166520 75710 166530 75790
rect 166700 75710 166710 75790
rect 166880 75710 166890 75790
rect 167060 75710 167070 75790
rect 167240 75710 167250 75790
rect 167420 75710 167430 75790
rect 167600 75710 167610 75790
rect 167780 75710 167790 75790
rect 167960 75710 167970 75790
rect 168140 75710 168150 75790
rect 168320 75710 168330 75790
rect 168500 75710 168510 75790
rect 168680 75710 168690 75790
rect 168860 75710 168870 75790
rect 169040 75710 169050 75790
rect 169220 75710 169230 75790
rect 169400 75710 169410 75790
rect 169580 75710 169590 75790
rect 169760 75710 169770 75790
rect 169940 75710 169950 75790
rect 170120 75710 170130 75790
rect 170300 75710 170310 75790
rect 170480 75710 170490 75790
rect 170660 75710 170670 75790
rect 170840 75710 170850 75790
rect 171020 75710 171030 75790
rect 18980 75640 19060 75650
rect 19160 75640 19240 75650
rect 19340 75640 19420 75650
rect 19520 75640 19600 75650
rect 19700 75640 19780 75650
rect 19880 75640 19960 75650
rect 20060 75640 20140 75650
rect 20240 75640 20320 75650
rect 20420 75640 20500 75650
rect 20600 75640 20680 75650
rect 20780 75640 20860 75650
rect 20960 75640 21040 75650
rect 21140 75640 21220 75650
rect 21320 75640 21400 75650
rect 21500 75640 21580 75650
rect 21680 75640 21760 75650
rect 21860 75640 21940 75650
rect 22040 75640 22120 75650
rect 22220 75640 22300 75650
rect 22400 75640 22480 75650
rect 22580 75640 22660 75650
rect 22760 75640 22840 75650
rect 22940 75640 23020 75650
rect 23120 75640 23200 75650
rect 23300 75640 23380 75650
rect 23480 75640 23560 75650
rect 23660 75640 23740 75650
rect 23840 75640 23920 75650
rect 24020 75640 24100 75650
rect 24200 75640 24280 75650
rect 24380 75640 24460 75650
rect 24560 75640 24640 75650
rect 24740 75640 24820 75650
rect 24920 75640 25000 75650
rect 25100 75640 25180 75650
rect 25280 75640 25360 75650
rect 25460 75640 25540 75650
rect 25640 75640 25720 75650
rect 25820 75640 25900 75650
rect 26000 75640 26080 75650
rect 26180 75640 26260 75650
rect 26360 75640 26440 75650
rect 26540 75640 26620 75650
rect 146300 75640 146380 75650
rect 146440 75640 146520 75650
rect 146580 75640 146660 75650
rect 146720 75640 146800 75650
rect 146860 75640 146940 75650
rect 147000 75640 147080 75650
rect 147140 75640 147220 75650
rect 147280 75640 147360 75650
rect 147420 75640 147500 75650
rect 147560 75640 147640 75650
rect 148600 75640 148680 75650
rect 148740 75640 148820 75650
rect 148880 75640 148960 75650
rect 149020 75640 149100 75650
rect 149160 75640 149240 75650
rect 149300 75640 149380 75650
rect 149440 75640 149520 75650
rect 149580 75640 149660 75650
rect 149720 75640 149800 75650
rect 149860 75640 149940 75650
rect 152080 75640 152160 75650
rect 152260 75640 152340 75650
rect 152440 75640 152520 75650
rect 152620 75640 152700 75650
rect 152800 75640 152880 75650
rect 152980 75640 153060 75650
rect 153160 75640 153240 75650
rect 153340 75640 153420 75650
rect 153520 75640 153600 75650
rect 153700 75640 153780 75650
rect 153880 75640 153960 75650
rect 154060 75640 154140 75650
rect 154240 75640 154320 75650
rect 154420 75640 154500 75650
rect 154600 75640 154680 75650
rect 154780 75640 154860 75650
rect 154960 75640 155040 75650
rect 155140 75640 155220 75650
rect 155320 75640 155400 75650
rect 155500 75640 155580 75650
rect 155680 75640 155760 75650
rect 155860 75640 155940 75650
rect 156040 75640 156120 75650
rect 156220 75640 156300 75650
rect 156400 75640 156480 75650
rect 156580 75640 156660 75650
rect 156760 75640 156840 75650
rect 156940 75640 157020 75650
rect 157120 75640 157200 75650
rect 157300 75640 157380 75650
rect 157480 75640 157560 75650
rect 157660 75640 157740 75650
rect 157840 75640 157920 75650
rect 158020 75640 158100 75650
rect 158200 75640 158280 75650
rect 158380 75640 158460 75650
rect 158560 75640 158640 75650
rect 158740 75640 158820 75650
rect 158920 75640 159000 75650
rect 159100 75640 159180 75650
rect 159280 75640 159360 75650
rect 159460 75640 159540 75650
rect 159640 75640 159720 75650
rect 163380 75640 163460 75650
rect 163560 75640 163640 75650
rect 163740 75640 163820 75650
rect 163920 75640 164000 75650
rect 164100 75640 164180 75650
rect 164280 75640 164360 75650
rect 164460 75640 164540 75650
rect 164640 75640 164720 75650
rect 164820 75640 164900 75650
rect 165000 75640 165080 75650
rect 165180 75640 165260 75650
rect 165360 75640 165440 75650
rect 165540 75640 165620 75650
rect 165720 75640 165800 75650
rect 165900 75640 165980 75650
rect 166080 75640 166160 75650
rect 166260 75640 166340 75650
rect 166440 75640 166520 75650
rect 166620 75640 166700 75650
rect 166800 75640 166880 75650
rect 166980 75640 167060 75650
rect 167160 75640 167240 75650
rect 167340 75640 167420 75650
rect 167520 75640 167600 75650
rect 167700 75640 167780 75650
rect 167880 75640 167960 75650
rect 168060 75640 168140 75650
rect 168240 75640 168320 75650
rect 168420 75640 168500 75650
rect 168600 75640 168680 75650
rect 168780 75640 168860 75650
rect 168960 75640 169040 75650
rect 169140 75640 169220 75650
rect 169320 75640 169400 75650
rect 169500 75640 169580 75650
rect 169680 75640 169760 75650
rect 169860 75640 169940 75650
rect 170040 75640 170120 75650
rect 170220 75640 170300 75650
rect 170400 75640 170480 75650
rect 170580 75640 170660 75650
rect 170760 75640 170840 75650
rect 170940 75640 171020 75650
rect 19060 75560 19070 75640
rect 19240 75560 19250 75640
rect 19420 75560 19430 75640
rect 19600 75560 19610 75640
rect 19780 75560 19790 75640
rect 19960 75560 19970 75640
rect 20140 75560 20150 75640
rect 20320 75560 20330 75640
rect 20500 75560 20510 75640
rect 20680 75560 20690 75640
rect 20860 75560 20870 75640
rect 21040 75560 21050 75640
rect 21220 75560 21230 75640
rect 21400 75560 21410 75640
rect 21580 75560 21590 75640
rect 21760 75560 21770 75640
rect 21940 75560 21950 75640
rect 22120 75560 22130 75640
rect 22300 75560 22310 75640
rect 22480 75560 22490 75640
rect 22660 75560 22670 75640
rect 22840 75560 22850 75640
rect 23020 75560 23030 75640
rect 23200 75560 23210 75640
rect 23380 75560 23390 75640
rect 23560 75560 23570 75640
rect 23740 75560 23750 75640
rect 23920 75560 23930 75640
rect 24100 75560 24110 75640
rect 24280 75560 24290 75640
rect 24460 75560 24470 75640
rect 24640 75560 24650 75640
rect 24820 75560 24830 75640
rect 25000 75560 25010 75640
rect 25180 75560 25190 75640
rect 25360 75560 25370 75640
rect 25540 75560 25550 75640
rect 25720 75560 25730 75640
rect 25900 75560 25910 75640
rect 26080 75560 26090 75640
rect 26260 75560 26270 75640
rect 26440 75560 26450 75640
rect 26620 75560 26630 75640
rect 146380 75581 146390 75640
rect 146520 75581 146530 75640
rect 146660 75581 146670 75640
rect 146800 75581 146810 75640
rect 146940 75581 146950 75640
rect 147080 75581 147090 75640
rect 147220 75581 147230 75640
rect 147360 75581 147370 75640
rect 147500 75581 147510 75640
rect 147640 75581 147650 75640
rect 148680 75581 148690 75640
rect 148820 75581 148830 75640
rect 148960 75581 148970 75640
rect 149100 75581 149110 75640
rect 149240 75581 149250 75640
rect 149380 75581 149390 75640
rect 149520 75581 149530 75640
rect 149660 75581 149670 75640
rect 149800 75581 149810 75640
rect 149940 75581 149950 75640
rect 152160 75581 152170 75640
rect 152340 75581 152350 75640
rect 152520 75581 152530 75640
rect 152700 75581 152710 75640
rect 152880 75581 152890 75640
rect 153060 75581 153070 75640
rect 153240 75581 153250 75640
rect 153420 75581 153430 75640
rect 153600 75581 153610 75640
rect 153780 75581 153790 75640
rect 153960 75581 153970 75640
rect 154140 75581 154150 75640
rect 154320 75581 154330 75640
rect 154500 75581 154510 75640
rect 154680 75581 154690 75640
rect 154860 75581 154870 75640
rect 155040 75581 155050 75640
rect 155220 75581 155230 75640
rect 155400 75581 155410 75640
rect 155580 75581 155590 75640
rect 155760 75581 155770 75640
rect 155940 75581 155950 75640
rect 156120 75581 156130 75640
rect 156300 75581 156310 75640
rect 156480 75581 156490 75640
rect 156660 75581 156670 75640
rect 156840 75581 156850 75640
rect 157020 75581 157030 75640
rect 157200 75581 157210 75640
rect 157380 75581 157390 75640
rect 157560 75581 157570 75640
rect 157740 75581 157750 75640
rect 157920 75581 157930 75640
rect 158100 75581 158110 75640
rect 158280 75581 158290 75640
rect 158460 75581 158470 75640
rect 158640 75581 158650 75640
rect 158820 75581 158830 75640
rect 159000 75581 159010 75640
rect 159180 75581 159190 75640
rect 159360 75581 159370 75640
rect 159540 75581 159550 75640
rect 159720 75581 159730 75640
rect 163460 75581 163470 75640
rect 163640 75581 163650 75640
rect 163820 75581 163830 75640
rect 164000 75581 164010 75640
rect 164180 75581 164190 75640
rect 164360 75581 164370 75640
rect 164540 75581 164550 75640
rect 164720 75581 164730 75640
rect 164900 75581 164910 75640
rect 165080 75581 165090 75640
rect 165260 75581 165270 75640
rect 165440 75581 165450 75640
rect 165620 75581 165630 75640
rect 165800 75581 165810 75640
rect 165980 75581 165990 75640
rect 166160 75581 166170 75640
rect 166340 75581 166350 75640
rect 166520 75581 166530 75640
rect 166700 75581 166710 75640
rect 166880 75581 166890 75640
rect 167060 75581 167070 75640
rect 167240 75581 167250 75640
rect 167420 75581 167430 75640
rect 167600 75581 167610 75640
rect 167780 75581 167790 75640
rect 167960 75581 167970 75640
rect 168140 75581 168150 75640
rect 168320 75581 168330 75640
rect 168500 75581 168510 75640
rect 168680 75581 168690 75640
rect 168860 75581 168870 75640
rect 169040 75581 169050 75640
rect 169220 75581 169230 75640
rect 169400 75581 169410 75640
rect 169580 75581 169590 75640
rect 169760 75581 169770 75640
rect 169940 75581 169950 75640
rect 170120 75581 170130 75640
rect 170300 75581 170310 75640
rect 170480 75581 170490 75640
rect 170660 75581 170670 75640
rect 170840 75581 170850 75640
rect 171020 75581 171030 75640
rect 146040 75500 147700 75581
rect 148340 75500 150000 75581
rect 152000 75500 159800 75581
rect 163210 75560 171100 75581
rect 163300 75500 171100 75560
rect 30360 75420 30440 75430
rect 30680 75420 30760 75430
rect 31000 75420 31080 75430
rect 31320 75420 31400 75430
rect 31640 75420 31720 75430
rect 31960 75420 32040 75430
rect 32280 75420 32360 75430
rect 32600 75420 32680 75430
rect 32920 75420 33000 75430
rect 33240 75420 33320 75430
rect 33560 75420 33640 75430
rect 33880 75420 33960 75430
rect 34200 75420 34280 75430
rect 34520 75420 34600 75430
rect 34840 75420 34920 75430
rect 35160 75420 35240 75430
rect 35480 75420 35560 75430
rect 35800 75420 35880 75430
rect 36120 75420 36200 75430
rect 36440 75420 36520 75430
rect 36760 75420 36840 75430
rect 37080 75420 37160 75430
rect 37400 75420 37480 75430
rect 37720 75420 37800 75430
rect 40180 75420 40260 75430
rect 40500 75420 40580 75430
rect 40820 75420 40900 75430
rect 41140 75420 41220 75430
rect 42560 75420 42640 75430
rect 42880 75420 42960 75430
rect 43200 75420 43280 75430
rect 43520 75420 43600 75430
rect 18970 75390 19050 75400
rect 19290 75390 19370 75400
rect 19610 75390 19690 75400
rect 19930 75390 20010 75400
rect 20250 75390 20330 75400
rect 20570 75390 20650 75400
rect 20890 75390 20970 75400
rect 21210 75390 21290 75400
rect 21530 75390 21610 75400
rect 21850 75390 21930 75400
rect 22170 75390 22250 75400
rect 22490 75390 22570 75400
rect 22810 75390 22890 75400
rect 23130 75390 23210 75400
rect 23450 75390 23530 75400
rect 23770 75390 23850 75400
rect 24090 75390 24170 75400
rect 24410 75390 24490 75400
rect 24730 75390 24810 75400
rect 25050 75390 25130 75400
rect 25370 75390 25450 75400
rect 25690 75390 25770 75400
rect 26010 75390 26090 75400
rect 26330 75390 26410 75400
rect 19050 75310 19060 75390
rect 19370 75310 19380 75390
rect 19690 75310 19700 75390
rect 20010 75310 20020 75390
rect 20330 75310 20340 75390
rect 20650 75310 20660 75390
rect 20970 75310 20980 75390
rect 21290 75310 21300 75390
rect 21610 75310 21620 75390
rect 21930 75310 21940 75390
rect 22250 75310 22260 75390
rect 22570 75310 22580 75390
rect 22890 75310 22900 75390
rect 23210 75310 23220 75390
rect 23530 75310 23540 75390
rect 23850 75310 23860 75390
rect 24170 75310 24180 75390
rect 24490 75310 24500 75390
rect 24810 75310 24820 75390
rect 25130 75310 25140 75390
rect 25450 75310 25460 75390
rect 25770 75310 25780 75390
rect 26090 75310 26100 75390
rect 26410 75310 26420 75390
rect 30440 75340 30450 75420
rect 30760 75340 30770 75420
rect 31080 75340 31090 75420
rect 31400 75340 31410 75420
rect 31720 75340 31730 75420
rect 32040 75340 32050 75420
rect 32360 75340 32370 75420
rect 32680 75340 32690 75420
rect 33000 75340 33010 75420
rect 33320 75340 33330 75420
rect 33640 75340 33650 75420
rect 33960 75340 33970 75420
rect 34280 75340 34290 75420
rect 34600 75340 34610 75420
rect 34920 75340 34930 75420
rect 35240 75340 35250 75420
rect 35560 75340 35570 75420
rect 35880 75340 35890 75420
rect 36200 75340 36210 75420
rect 36520 75340 36530 75420
rect 36840 75340 36850 75420
rect 37160 75340 37170 75420
rect 37480 75340 37490 75420
rect 37800 75340 37810 75420
rect 40260 75340 40270 75420
rect 40580 75340 40590 75420
rect 40900 75340 40910 75420
rect 41220 75340 41230 75420
rect 42640 75340 42650 75420
rect 42960 75340 42970 75420
rect 43280 75340 43290 75420
rect 43600 75340 43610 75420
rect 146400 75411 146480 75421
rect 146720 75411 146800 75421
rect 147040 75411 147120 75421
rect 147360 75411 147440 75421
rect 148780 75411 148860 75421
rect 149100 75411 149180 75421
rect 149420 75411 149500 75421
rect 149740 75411 149820 75421
rect 152200 75411 152280 75421
rect 152520 75411 152600 75421
rect 152840 75411 152920 75421
rect 153160 75411 153240 75421
rect 153480 75411 153560 75421
rect 153800 75411 153880 75421
rect 154120 75411 154200 75421
rect 154440 75411 154520 75421
rect 154760 75411 154840 75421
rect 155080 75411 155160 75421
rect 155400 75411 155480 75421
rect 155720 75411 155800 75421
rect 156040 75411 156120 75421
rect 156360 75411 156440 75421
rect 156680 75411 156760 75421
rect 157000 75411 157080 75421
rect 157320 75411 157400 75421
rect 157640 75411 157720 75421
rect 157960 75411 158040 75421
rect 158280 75411 158360 75421
rect 158600 75411 158680 75421
rect 158920 75411 159000 75421
rect 159240 75411 159320 75421
rect 159560 75411 159640 75421
rect 146480 75331 146490 75411
rect 146800 75331 146810 75411
rect 147120 75331 147130 75411
rect 147440 75331 147450 75411
rect 148860 75331 148870 75411
rect 149180 75331 149190 75411
rect 149500 75331 149510 75411
rect 149820 75331 149830 75411
rect 152280 75331 152290 75411
rect 152600 75331 152610 75411
rect 152920 75331 152930 75411
rect 153240 75331 153250 75411
rect 153560 75331 153570 75411
rect 153880 75331 153890 75411
rect 154200 75331 154210 75411
rect 154520 75331 154530 75411
rect 154840 75331 154850 75411
rect 155160 75331 155170 75411
rect 155480 75331 155490 75411
rect 155800 75331 155810 75411
rect 156120 75331 156130 75411
rect 156440 75331 156450 75411
rect 156760 75331 156770 75411
rect 157080 75331 157090 75411
rect 157400 75331 157410 75411
rect 157720 75331 157730 75411
rect 158040 75331 158050 75411
rect 158360 75331 158370 75411
rect 158680 75331 158690 75411
rect 159000 75331 159010 75411
rect 159320 75331 159330 75411
rect 159640 75331 159650 75411
rect 163590 75381 163670 75391
rect 163910 75381 163990 75391
rect 164230 75381 164310 75391
rect 164550 75381 164630 75391
rect 164870 75381 164950 75391
rect 165190 75381 165270 75391
rect 165510 75381 165590 75391
rect 165830 75381 165910 75391
rect 166150 75381 166230 75391
rect 166470 75381 166550 75391
rect 166790 75381 166870 75391
rect 167110 75381 167190 75391
rect 167430 75381 167510 75391
rect 167750 75381 167830 75391
rect 168070 75381 168150 75391
rect 168390 75381 168470 75391
rect 168710 75381 168790 75391
rect 169030 75381 169110 75391
rect 169350 75381 169430 75391
rect 169670 75381 169750 75391
rect 169990 75381 170070 75391
rect 170310 75381 170390 75391
rect 170630 75381 170710 75391
rect 170950 75381 171030 75391
rect 163670 75301 163680 75381
rect 163990 75301 164000 75381
rect 164310 75301 164320 75381
rect 164630 75301 164640 75381
rect 164950 75301 164960 75381
rect 165270 75301 165280 75381
rect 165590 75301 165600 75381
rect 165910 75301 165920 75381
rect 166230 75301 166240 75381
rect 166550 75301 166560 75381
rect 166870 75301 166880 75381
rect 167190 75301 167200 75381
rect 167510 75301 167520 75381
rect 167830 75301 167840 75381
rect 168150 75301 168160 75381
rect 168470 75301 168480 75381
rect 168790 75301 168800 75381
rect 169110 75301 169120 75381
rect 169430 75301 169440 75381
rect 169750 75301 169760 75381
rect 170070 75301 170080 75381
rect 170390 75301 170400 75381
rect 170710 75301 170720 75381
rect 171030 75301 171040 75381
rect 30520 75260 30600 75270
rect 30840 75260 30920 75270
rect 31160 75260 31240 75270
rect 31480 75260 31560 75270
rect 31800 75260 31880 75270
rect 32120 75260 32200 75270
rect 32440 75260 32520 75270
rect 32760 75260 32840 75270
rect 33080 75260 33160 75270
rect 33400 75260 33480 75270
rect 33720 75260 33800 75270
rect 34040 75260 34120 75270
rect 34360 75260 34440 75270
rect 34680 75260 34760 75270
rect 35000 75260 35080 75270
rect 35320 75260 35400 75270
rect 35640 75260 35720 75270
rect 35960 75260 36040 75270
rect 36280 75260 36360 75270
rect 36600 75260 36680 75270
rect 36920 75260 37000 75270
rect 37240 75260 37320 75270
rect 37560 75260 37640 75270
rect 40340 75260 40420 75270
rect 40660 75260 40740 75270
rect 40980 75260 41060 75270
rect 42720 75260 42800 75270
rect 43040 75260 43120 75270
rect 43360 75260 43440 75270
rect 19130 75230 19210 75240
rect 19450 75230 19530 75240
rect 19770 75230 19850 75240
rect 20090 75230 20170 75240
rect 20410 75230 20490 75240
rect 20730 75230 20810 75240
rect 21050 75230 21130 75240
rect 21370 75230 21450 75240
rect 21690 75230 21770 75240
rect 22010 75230 22090 75240
rect 22330 75230 22410 75240
rect 22650 75230 22730 75240
rect 22970 75230 23050 75240
rect 23290 75230 23370 75240
rect 23610 75230 23690 75240
rect 23930 75230 24010 75240
rect 24250 75230 24330 75240
rect 24570 75230 24650 75240
rect 24890 75230 24970 75240
rect 25210 75230 25290 75240
rect 25530 75230 25610 75240
rect 25850 75230 25930 75240
rect 26170 75230 26250 75240
rect 19210 75150 19220 75230
rect 19530 75150 19540 75230
rect 19850 75150 19860 75230
rect 20170 75150 20180 75230
rect 20490 75150 20500 75230
rect 20810 75150 20820 75230
rect 21130 75150 21140 75230
rect 21450 75150 21460 75230
rect 21770 75150 21780 75230
rect 22090 75150 22100 75230
rect 22410 75150 22420 75230
rect 22730 75150 22740 75230
rect 23050 75150 23060 75230
rect 23370 75150 23380 75230
rect 23690 75150 23700 75230
rect 24010 75150 24020 75230
rect 24330 75150 24340 75230
rect 24650 75150 24660 75230
rect 24970 75150 24980 75230
rect 25290 75150 25300 75230
rect 25610 75150 25620 75230
rect 25930 75150 25940 75230
rect 26250 75150 26260 75230
rect 30600 75180 30610 75260
rect 30920 75180 30930 75260
rect 31240 75180 31250 75260
rect 31560 75180 31570 75260
rect 31880 75180 31890 75260
rect 32200 75180 32210 75260
rect 32520 75180 32530 75260
rect 32840 75180 32850 75260
rect 33160 75180 33170 75260
rect 33480 75180 33490 75260
rect 33800 75180 33810 75260
rect 34120 75180 34130 75260
rect 34440 75180 34450 75260
rect 34760 75180 34770 75260
rect 35080 75180 35090 75260
rect 35400 75180 35410 75260
rect 35720 75180 35730 75260
rect 36040 75180 36050 75260
rect 36360 75180 36370 75260
rect 36680 75180 36690 75260
rect 37000 75180 37010 75260
rect 37320 75180 37330 75260
rect 37640 75180 37650 75260
rect 40420 75180 40430 75260
rect 40740 75180 40750 75260
rect 41060 75180 41070 75260
rect 42800 75180 42810 75260
rect 43120 75180 43130 75260
rect 43440 75180 43450 75260
rect 146560 75251 146640 75261
rect 146880 75251 146960 75261
rect 147200 75251 147280 75261
rect 148940 75251 149020 75261
rect 149260 75251 149340 75261
rect 149580 75251 149660 75261
rect 152360 75251 152440 75261
rect 152680 75251 152760 75261
rect 153000 75251 153080 75261
rect 153320 75251 153400 75261
rect 153640 75251 153720 75261
rect 153960 75251 154040 75261
rect 154280 75251 154360 75261
rect 154600 75251 154680 75261
rect 154920 75251 155000 75261
rect 155240 75251 155320 75261
rect 155560 75251 155640 75261
rect 155880 75251 155960 75261
rect 156200 75251 156280 75261
rect 156520 75251 156600 75261
rect 156840 75251 156920 75261
rect 157160 75251 157240 75261
rect 157480 75251 157560 75261
rect 157800 75251 157880 75261
rect 158120 75251 158200 75261
rect 158440 75251 158520 75261
rect 158760 75251 158840 75261
rect 159080 75251 159160 75261
rect 159400 75251 159480 75261
rect 146640 75171 146650 75251
rect 146960 75171 146970 75251
rect 147280 75171 147290 75251
rect 149020 75171 149030 75251
rect 149340 75171 149350 75251
rect 149660 75171 149670 75251
rect 152440 75171 152450 75251
rect 152760 75171 152770 75251
rect 153080 75171 153090 75251
rect 153400 75171 153410 75251
rect 153720 75171 153730 75251
rect 154040 75171 154050 75251
rect 154360 75171 154370 75251
rect 154680 75171 154690 75251
rect 155000 75171 155010 75251
rect 155320 75171 155330 75251
rect 155640 75171 155650 75251
rect 155960 75171 155970 75251
rect 156280 75171 156290 75251
rect 156600 75171 156610 75251
rect 156920 75171 156930 75251
rect 157240 75171 157250 75251
rect 157560 75171 157570 75251
rect 157880 75171 157890 75251
rect 158200 75171 158210 75251
rect 158520 75171 158530 75251
rect 158840 75171 158850 75251
rect 159160 75171 159170 75251
rect 159480 75171 159490 75251
rect 163750 75221 163830 75231
rect 164070 75221 164150 75231
rect 164390 75221 164470 75231
rect 164710 75221 164790 75231
rect 165030 75221 165110 75231
rect 165350 75221 165430 75231
rect 165670 75221 165750 75231
rect 165990 75221 166070 75231
rect 166310 75221 166390 75231
rect 166630 75221 166710 75231
rect 166950 75221 167030 75231
rect 167270 75221 167350 75231
rect 167590 75221 167670 75231
rect 167910 75221 167990 75231
rect 168230 75221 168310 75231
rect 168550 75221 168630 75231
rect 168870 75221 168950 75231
rect 169190 75221 169270 75231
rect 169510 75221 169590 75231
rect 169830 75221 169910 75231
rect 170150 75221 170230 75231
rect 170470 75221 170550 75231
rect 170790 75221 170870 75231
rect 163830 75141 163840 75221
rect 164150 75141 164160 75221
rect 164470 75141 164480 75221
rect 164790 75141 164800 75221
rect 165110 75141 165120 75221
rect 165430 75141 165440 75221
rect 165750 75141 165760 75221
rect 166070 75141 166080 75221
rect 166390 75141 166400 75221
rect 166710 75141 166720 75221
rect 167030 75141 167040 75221
rect 167350 75141 167360 75221
rect 167670 75141 167680 75221
rect 167990 75141 168000 75221
rect 168310 75141 168320 75221
rect 168630 75141 168640 75221
rect 168950 75141 168960 75221
rect 169270 75141 169280 75221
rect 169590 75141 169600 75221
rect 169910 75141 169920 75221
rect 170230 75141 170240 75221
rect 170550 75141 170560 75221
rect 170870 75141 170880 75221
rect 30360 75100 30440 75110
rect 30680 75100 30760 75110
rect 31000 75100 31080 75110
rect 31320 75100 31400 75110
rect 31640 75100 31720 75110
rect 31960 75100 32040 75110
rect 32280 75100 32360 75110
rect 32600 75100 32680 75110
rect 32920 75100 33000 75110
rect 33240 75100 33320 75110
rect 33560 75100 33640 75110
rect 33880 75100 33960 75110
rect 34200 75100 34280 75110
rect 34520 75100 34600 75110
rect 34840 75100 34920 75110
rect 35160 75100 35240 75110
rect 35480 75100 35560 75110
rect 35800 75100 35880 75110
rect 36120 75100 36200 75110
rect 36440 75100 36520 75110
rect 36760 75100 36840 75110
rect 37080 75100 37160 75110
rect 37400 75100 37480 75110
rect 37720 75100 37800 75110
rect 40180 75100 40260 75110
rect 40500 75100 40580 75110
rect 40820 75100 40900 75110
rect 41140 75100 41220 75110
rect 42560 75100 42640 75110
rect 42880 75100 42960 75110
rect 43200 75100 43280 75110
rect 43520 75100 43600 75110
rect 18970 75070 19050 75080
rect 19290 75070 19370 75080
rect 19610 75070 19690 75080
rect 19930 75070 20010 75080
rect 20250 75070 20330 75080
rect 20570 75070 20650 75080
rect 20890 75070 20970 75080
rect 21210 75070 21290 75080
rect 21530 75070 21610 75080
rect 21850 75070 21930 75080
rect 22170 75070 22250 75080
rect 22490 75070 22570 75080
rect 22810 75070 22890 75080
rect 23130 75070 23210 75080
rect 23450 75070 23530 75080
rect 23770 75070 23850 75080
rect 24090 75070 24170 75080
rect 24410 75070 24490 75080
rect 24730 75070 24810 75080
rect 25050 75070 25130 75080
rect 25370 75070 25450 75080
rect 25690 75070 25770 75080
rect 26010 75070 26090 75080
rect 26330 75070 26410 75080
rect 19050 74990 19060 75070
rect 19370 74990 19380 75070
rect 19690 74990 19700 75070
rect 20010 74990 20020 75070
rect 20330 74990 20340 75070
rect 20650 74990 20660 75070
rect 20970 74990 20980 75070
rect 21290 74990 21300 75070
rect 21610 74990 21620 75070
rect 21930 74990 21940 75070
rect 22250 74990 22260 75070
rect 22570 74990 22580 75070
rect 22890 74990 22900 75070
rect 23210 74990 23220 75070
rect 23530 74990 23540 75070
rect 23850 74990 23860 75070
rect 24170 74990 24180 75070
rect 24490 74990 24500 75070
rect 24810 74990 24820 75070
rect 25130 74990 25140 75070
rect 25450 74990 25460 75070
rect 25770 74990 25780 75070
rect 26090 74990 26100 75070
rect 26410 74990 26420 75070
rect 30440 75020 30450 75100
rect 30760 75020 30770 75100
rect 31080 75020 31090 75100
rect 31400 75020 31410 75100
rect 31720 75020 31730 75100
rect 32040 75020 32050 75100
rect 32360 75020 32370 75100
rect 32680 75020 32690 75100
rect 33000 75020 33010 75100
rect 33320 75020 33330 75100
rect 33640 75020 33650 75100
rect 33960 75020 33970 75100
rect 34280 75020 34290 75100
rect 34600 75020 34610 75100
rect 34920 75020 34930 75100
rect 35240 75020 35250 75100
rect 35560 75020 35570 75100
rect 35880 75020 35890 75100
rect 36200 75020 36210 75100
rect 36520 75020 36530 75100
rect 36840 75020 36850 75100
rect 37160 75020 37170 75100
rect 37480 75020 37490 75100
rect 37800 75020 37810 75100
rect 40260 75020 40270 75100
rect 40580 75020 40590 75100
rect 40900 75020 40910 75100
rect 41220 75020 41230 75100
rect 42640 75020 42650 75100
rect 42960 75020 42970 75100
rect 43280 75020 43290 75100
rect 43600 75020 43610 75100
rect 146400 75091 146480 75101
rect 146720 75091 146800 75101
rect 147040 75091 147120 75101
rect 147360 75091 147440 75101
rect 148780 75091 148860 75101
rect 149100 75091 149180 75101
rect 149420 75091 149500 75101
rect 149740 75091 149820 75101
rect 152200 75091 152280 75101
rect 152520 75091 152600 75101
rect 152840 75091 152920 75101
rect 153160 75091 153240 75101
rect 153480 75091 153560 75101
rect 153800 75091 153880 75101
rect 154120 75091 154200 75101
rect 154440 75091 154520 75101
rect 154760 75091 154840 75101
rect 155080 75091 155160 75101
rect 155400 75091 155480 75101
rect 155720 75091 155800 75101
rect 156040 75091 156120 75101
rect 156360 75091 156440 75101
rect 156680 75091 156760 75101
rect 157000 75091 157080 75101
rect 157320 75091 157400 75101
rect 157640 75091 157720 75101
rect 157960 75091 158040 75101
rect 158280 75091 158360 75101
rect 158600 75091 158680 75101
rect 158920 75091 159000 75101
rect 159240 75091 159320 75101
rect 159560 75091 159640 75101
rect 146480 75011 146490 75091
rect 146800 75011 146810 75091
rect 147120 75011 147130 75091
rect 147440 75011 147450 75091
rect 148860 75011 148870 75091
rect 149180 75011 149190 75091
rect 149500 75011 149510 75091
rect 149820 75011 149830 75091
rect 152280 75011 152290 75091
rect 152600 75011 152610 75091
rect 152920 75011 152930 75091
rect 153240 75011 153250 75091
rect 153560 75011 153570 75091
rect 153880 75011 153890 75091
rect 154200 75011 154210 75091
rect 154520 75011 154530 75091
rect 154840 75011 154850 75091
rect 155160 75011 155170 75091
rect 155480 75011 155490 75091
rect 155800 75011 155810 75091
rect 156120 75011 156130 75091
rect 156440 75011 156450 75091
rect 156760 75011 156770 75091
rect 157080 75011 157090 75091
rect 157400 75011 157410 75091
rect 157720 75011 157730 75091
rect 158040 75011 158050 75091
rect 158360 75011 158370 75091
rect 158680 75011 158690 75091
rect 159000 75011 159010 75091
rect 159320 75011 159330 75091
rect 159640 75011 159650 75091
rect 163590 75061 163670 75071
rect 163910 75061 163990 75071
rect 164230 75061 164310 75071
rect 164550 75061 164630 75071
rect 164870 75061 164950 75071
rect 165190 75061 165270 75071
rect 165510 75061 165590 75071
rect 165830 75061 165910 75071
rect 166150 75061 166230 75071
rect 166470 75061 166550 75071
rect 166790 75061 166870 75071
rect 167110 75061 167190 75071
rect 167430 75061 167510 75071
rect 167750 75061 167830 75071
rect 168070 75061 168150 75071
rect 168390 75061 168470 75071
rect 168710 75061 168790 75071
rect 169030 75061 169110 75071
rect 169350 75061 169430 75071
rect 169670 75061 169750 75071
rect 169990 75061 170070 75071
rect 170310 75061 170390 75071
rect 170630 75061 170710 75071
rect 170950 75061 171030 75071
rect 163670 74981 163680 75061
rect 163990 74981 164000 75061
rect 164310 74981 164320 75061
rect 164630 74981 164640 75061
rect 164950 74981 164960 75061
rect 165270 74981 165280 75061
rect 165590 74981 165600 75061
rect 165910 74981 165920 75061
rect 166230 74981 166240 75061
rect 166550 74981 166560 75061
rect 166870 74981 166880 75061
rect 167190 74981 167200 75061
rect 167510 74981 167520 75061
rect 167830 74981 167840 75061
rect 168150 74981 168160 75061
rect 168470 74981 168480 75061
rect 168790 74981 168800 75061
rect 169110 74981 169120 75061
rect 169430 74981 169440 75061
rect 169750 74981 169760 75061
rect 170070 74981 170080 75061
rect 170390 74981 170400 75061
rect 170710 74981 170720 75061
rect 171030 74981 171040 75061
rect 30520 74940 30600 74950
rect 30840 74940 30920 74950
rect 31160 74940 31240 74950
rect 31480 74940 31560 74950
rect 31800 74940 31880 74950
rect 32120 74940 32200 74950
rect 32440 74940 32520 74950
rect 32760 74940 32840 74950
rect 33080 74940 33160 74950
rect 33400 74940 33480 74950
rect 33720 74940 33800 74950
rect 34040 74940 34120 74950
rect 34360 74940 34440 74950
rect 34680 74940 34760 74950
rect 35000 74940 35080 74950
rect 35320 74940 35400 74950
rect 35640 74940 35720 74950
rect 35960 74940 36040 74950
rect 36280 74940 36360 74950
rect 36600 74940 36680 74950
rect 36920 74940 37000 74950
rect 37240 74940 37320 74950
rect 37560 74940 37640 74950
rect 40340 74940 40420 74950
rect 40660 74940 40740 74950
rect 40980 74940 41060 74950
rect 42720 74940 42800 74950
rect 43040 74940 43120 74950
rect 43360 74940 43440 74950
rect 19130 74910 19210 74920
rect 19450 74910 19530 74920
rect 19770 74910 19850 74920
rect 20090 74910 20170 74920
rect 20410 74910 20490 74920
rect 20730 74910 20810 74920
rect 21050 74910 21130 74920
rect 21370 74910 21450 74920
rect 21690 74910 21770 74920
rect 22010 74910 22090 74920
rect 22330 74910 22410 74920
rect 22650 74910 22730 74920
rect 22970 74910 23050 74920
rect 23290 74910 23370 74920
rect 23610 74910 23690 74920
rect 23930 74910 24010 74920
rect 24250 74910 24330 74920
rect 24570 74910 24650 74920
rect 24890 74910 24970 74920
rect 25210 74910 25290 74920
rect 25530 74910 25610 74920
rect 25850 74910 25930 74920
rect 26170 74910 26250 74920
rect 19210 74830 19220 74910
rect 19530 74830 19540 74910
rect 19850 74830 19860 74910
rect 20170 74830 20180 74910
rect 20490 74830 20500 74910
rect 20810 74830 20820 74910
rect 21130 74830 21140 74910
rect 21450 74830 21460 74910
rect 21770 74830 21780 74910
rect 22090 74830 22100 74910
rect 22410 74830 22420 74910
rect 22730 74830 22740 74910
rect 23050 74830 23060 74910
rect 23370 74830 23380 74910
rect 23690 74830 23700 74910
rect 24010 74830 24020 74910
rect 24330 74830 24340 74910
rect 24650 74830 24660 74910
rect 24970 74830 24980 74910
rect 25290 74830 25300 74910
rect 25610 74830 25620 74910
rect 25930 74830 25940 74910
rect 26250 74830 26260 74910
rect 30600 74860 30610 74940
rect 30920 74860 30930 74940
rect 31240 74860 31250 74940
rect 31560 74860 31570 74940
rect 31880 74860 31890 74940
rect 32200 74860 32210 74940
rect 32520 74860 32530 74940
rect 32840 74860 32850 74940
rect 33160 74860 33170 74940
rect 33480 74860 33490 74940
rect 33800 74860 33810 74940
rect 34120 74860 34130 74940
rect 34440 74860 34450 74940
rect 34760 74860 34770 74940
rect 35080 74860 35090 74940
rect 35400 74860 35410 74940
rect 35720 74860 35730 74940
rect 36040 74860 36050 74940
rect 36360 74860 36370 74940
rect 36680 74860 36690 74940
rect 37000 74860 37010 74940
rect 37320 74860 37330 74940
rect 37640 74860 37650 74940
rect 40420 74860 40430 74940
rect 40740 74860 40750 74940
rect 41060 74860 41070 74940
rect 42800 74860 42810 74940
rect 43120 74860 43130 74940
rect 43440 74860 43450 74940
rect 146560 74931 146640 74941
rect 146880 74931 146960 74941
rect 147200 74931 147280 74941
rect 148940 74931 149020 74941
rect 149260 74931 149340 74941
rect 149580 74931 149660 74941
rect 152360 74931 152440 74941
rect 152680 74931 152760 74941
rect 153000 74931 153080 74941
rect 153320 74931 153400 74941
rect 153640 74931 153720 74941
rect 153960 74931 154040 74941
rect 154280 74931 154360 74941
rect 154600 74931 154680 74941
rect 154920 74931 155000 74941
rect 155240 74931 155320 74941
rect 155560 74931 155640 74941
rect 155880 74931 155960 74941
rect 156200 74931 156280 74941
rect 156520 74931 156600 74941
rect 156840 74931 156920 74941
rect 157160 74931 157240 74941
rect 157480 74931 157560 74941
rect 157800 74931 157880 74941
rect 158120 74931 158200 74941
rect 158440 74931 158520 74941
rect 158760 74931 158840 74941
rect 159080 74931 159160 74941
rect 159400 74931 159480 74941
rect 146640 74851 146650 74931
rect 146960 74851 146970 74931
rect 147280 74851 147290 74931
rect 149020 74851 149030 74931
rect 149340 74851 149350 74931
rect 149660 74851 149670 74931
rect 152440 74851 152450 74931
rect 152760 74851 152770 74931
rect 153080 74851 153090 74931
rect 153400 74851 153410 74931
rect 153720 74851 153730 74931
rect 154040 74851 154050 74931
rect 154360 74851 154370 74931
rect 154680 74851 154690 74931
rect 155000 74851 155010 74931
rect 155320 74851 155330 74931
rect 155640 74851 155650 74931
rect 155960 74851 155970 74931
rect 156280 74851 156290 74931
rect 156600 74851 156610 74931
rect 156920 74851 156930 74931
rect 157240 74851 157250 74931
rect 157560 74851 157570 74931
rect 157880 74851 157890 74931
rect 158200 74851 158210 74931
rect 158520 74851 158530 74931
rect 158840 74851 158850 74931
rect 159160 74851 159170 74931
rect 159480 74851 159490 74931
rect 163750 74901 163830 74911
rect 164070 74901 164150 74911
rect 164390 74901 164470 74911
rect 164710 74901 164790 74911
rect 165030 74901 165110 74911
rect 165350 74901 165430 74911
rect 165670 74901 165750 74911
rect 165990 74901 166070 74911
rect 166310 74901 166390 74911
rect 166630 74901 166710 74911
rect 166950 74901 167030 74911
rect 167270 74901 167350 74911
rect 167590 74901 167670 74911
rect 167910 74901 167990 74911
rect 168230 74901 168310 74911
rect 168550 74901 168630 74911
rect 168870 74901 168950 74911
rect 169190 74901 169270 74911
rect 169510 74901 169590 74911
rect 169830 74901 169910 74911
rect 170150 74901 170230 74911
rect 170470 74901 170550 74911
rect 170790 74901 170870 74911
rect 163830 74821 163840 74901
rect 164150 74821 164160 74901
rect 164470 74821 164480 74901
rect 164790 74821 164800 74901
rect 165110 74821 165120 74901
rect 165430 74821 165440 74901
rect 165750 74821 165760 74901
rect 166070 74821 166080 74901
rect 166390 74821 166400 74901
rect 166710 74821 166720 74901
rect 167030 74821 167040 74901
rect 167350 74821 167360 74901
rect 167670 74821 167680 74901
rect 167990 74821 168000 74901
rect 168310 74821 168320 74901
rect 168630 74821 168640 74901
rect 168950 74821 168960 74901
rect 169270 74821 169280 74901
rect 169590 74821 169600 74901
rect 169910 74821 169920 74901
rect 170230 74821 170240 74901
rect 170550 74821 170560 74901
rect 170870 74821 170880 74901
rect 30360 74680 30440 74690
rect 30680 74680 30760 74690
rect 31000 74680 31080 74690
rect 31320 74680 31400 74690
rect 31640 74680 31720 74690
rect 31960 74680 32040 74690
rect 32280 74680 32360 74690
rect 32600 74680 32680 74690
rect 32920 74680 33000 74690
rect 33240 74680 33320 74690
rect 33560 74680 33640 74690
rect 33880 74680 33960 74690
rect 34200 74680 34280 74690
rect 34520 74680 34600 74690
rect 34840 74680 34920 74690
rect 35160 74680 35240 74690
rect 35480 74680 35560 74690
rect 35800 74680 35880 74690
rect 36120 74680 36200 74690
rect 36440 74680 36520 74690
rect 36760 74680 36840 74690
rect 37080 74680 37160 74690
rect 37400 74680 37480 74690
rect 37720 74680 37800 74690
rect 40180 74680 40260 74690
rect 40500 74680 40580 74690
rect 40820 74680 40900 74690
rect 41140 74680 41220 74690
rect 42560 74680 42640 74690
rect 42880 74680 42960 74690
rect 43200 74680 43280 74690
rect 43520 74680 43600 74690
rect 18970 74650 19050 74660
rect 19290 74650 19370 74660
rect 19610 74650 19690 74660
rect 19930 74650 20010 74660
rect 20250 74650 20330 74660
rect 20570 74650 20650 74660
rect 20890 74650 20970 74660
rect 21210 74650 21290 74660
rect 21530 74650 21610 74660
rect 21850 74650 21930 74660
rect 22170 74650 22250 74660
rect 22490 74650 22570 74660
rect 22810 74650 22890 74660
rect 23130 74650 23210 74660
rect 23450 74650 23530 74660
rect 23770 74650 23850 74660
rect 24090 74650 24170 74660
rect 24410 74650 24490 74660
rect 24730 74650 24810 74660
rect 25050 74650 25130 74660
rect 25370 74650 25450 74660
rect 25690 74650 25770 74660
rect 26010 74650 26090 74660
rect 26330 74650 26410 74660
rect 19050 74570 19060 74650
rect 19370 74570 19380 74650
rect 19690 74570 19700 74650
rect 20010 74570 20020 74650
rect 20330 74570 20340 74650
rect 20650 74570 20660 74650
rect 20970 74570 20980 74650
rect 21290 74570 21300 74650
rect 21610 74570 21620 74650
rect 21930 74570 21940 74650
rect 22250 74570 22260 74650
rect 22570 74570 22580 74650
rect 22890 74570 22900 74650
rect 23210 74570 23220 74650
rect 23530 74570 23540 74650
rect 23850 74570 23860 74650
rect 24170 74570 24180 74650
rect 24490 74570 24500 74650
rect 24810 74570 24820 74650
rect 25130 74570 25140 74650
rect 25450 74570 25460 74650
rect 25770 74570 25780 74650
rect 26090 74570 26100 74650
rect 26410 74570 26420 74650
rect 30440 74600 30450 74680
rect 30760 74600 30770 74680
rect 31080 74600 31090 74680
rect 31400 74600 31410 74680
rect 31720 74600 31730 74680
rect 32040 74600 32050 74680
rect 32360 74600 32370 74680
rect 32680 74600 32690 74680
rect 33000 74600 33010 74680
rect 33320 74600 33330 74680
rect 33640 74600 33650 74680
rect 33960 74600 33970 74680
rect 34280 74600 34290 74680
rect 34600 74600 34610 74680
rect 34920 74600 34930 74680
rect 35240 74600 35250 74680
rect 35560 74600 35570 74680
rect 35880 74600 35890 74680
rect 36200 74600 36210 74680
rect 36520 74600 36530 74680
rect 36840 74600 36850 74680
rect 37160 74600 37170 74680
rect 37480 74600 37490 74680
rect 37800 74600 37810 74680
rect 40260 74600 40270 74680
rect 40580 74600 40590 74680
rect 40900 74600 40910 74680
rect 41220 74600 41230 74680
rect 42640 74600 42650 74680
rect 42960 74600 42970 74680
rect 43280 74600 43290 74680
rect 43600 74600 43610 74680
rect 146400 74671 146480 74681
rect 146720 74671 146800 74681
rect 147040 74671 147120 74681
rect 147360 74671 147440 74681
rect 148780 74671 148860 74681
rect 149100 74671 149180 74681
rect 149420 74671 149500 74681
rect 149740 74671 149820 74681
rect 152200 74671 152280 74681
rect 152520 74671 152600 74681
rect 152840 74671 152920 74681
rect 153160 74671 153240 74681
rect 153480 74671 153560 74681
rect 153800 74671 153880 74681
rect 154120 74671 154200 74681
rect 154440 74671 154520 74681
rect 154760 74671 154840 74681
rect 155080 74671 155160 74681
rect 155400 74671 155480 74681
rect 155720 74671 155800 74681
rect 156040 74671 156120 74681
rect 156360 74671 156440 74681
rect 156680 74671 156760 74681
rect 157000 74671 157080 74681
rect 157320 74671 157400 74681
rect 157640 74671 157720 74681
rect 157960 74671 158040 74681
rect 158280 74671 158360 74681
rect 158600 74671 158680 74681
rect 158920 74671 159000 74681
rect 159240 74671 159320 74681
rect 159560 74671 159640 74681
rect 146480 74591 146490 74671
rect 146800 74591 146810 74671
rect 147120 74591 147130 74671
rect 147440 74591 147450 74671
rect 148860 74591 148870 74671
rect 149180 74591 149190 74671
rect 149500 74591 149510 74671
rect 149820 74591 149830 74671
rect 152280 74591 152290 74671
rect 152600 74591 152610 74671
rect 152920 74591 152930 74671
rect 153240 74591 153250 74671
rect 153560 74591 153570 74671
rect 153880 74591 153890 74671
rect 154200 74591 154210 74671
rect 154520 74591 154530 74671
rect 154840 74591 154850 74671
rect 155160 74591 155170 74671
rect 155480 74591 155490 74671
rect 155800 74591 155810 74671
rect 156120 74591 156130 74671
rect 156440 74591 156450 74671
rect 156760 74591 156770 74671
rect 157080 74591 157090 74671
rect 157400 74591 157410 74671
rect 157720 74591 157730 74671
rect 158040 74591 158050 74671
rect 158360 74591 158370 74671
rect 158680 74591 158690 74671
rect 159000 74591 159010 74671
rect 159320 74591 159330 74671
rect 159640 74591 159650 74671
rect 163590 74641 163670 74651
rect 163910 74641 163990 74651
rect 164230 74641 164310 74651
rect 164550 74641 164630 74651
rect 164870 74641 164950 74651
rect 165190 74641 165270 74651
rect 165510 74641 165590 74651
rect 165830 74641 165910 74651
rect 166150 74641 166230 74651
rect 166470 74641 166550 74651
rect 166790 74641 166870 74651
rect 167110 74641 167190 74651
rect 167430 74641 167510 74651
rect 167750 74641 167830 74651
rect 168070 74641 168150 74651
rect 168390 74641 168470 74651
rect 168710 74641 168790 74651
rect 169030 74641 169110 74651
rect 169350 74641 169430 74651
rect 169670 74641 169750 74651
rect 169990 74641 170070 74651
rect 170310 74641 170390 74651
rect 170630 74641 170710 74651
rect 170950 74641 171030 74651
rect 163670 74561 163680 74641
rect 163990 74561 164000 74641
rect 164310 74561 164320 74641
rect 164630 74561 164640 74641
rect 164950 74561 164960 74641
rect 165270 74561 165280 74641
rect 165590 74561 165600 74641
rect 165910 74561 165920 74641
rect 166230 74561 166240 74641
rect 166550 74561 166560 74641
rect 166870 74561 166880 74641
rect 167190 74561 167200 74641
rect 167510 74561 167520 74641
rect 167830 74561 167840 74641
rect 168150 74561 168160 74641
rect 168470 74561 168480 74641
rect 168790 74561 168800 74641
rect 169110 74561 169120 74641
rect 169430 74561 169440 74641
rect 169750 74561 169760 74641
rect 170070 74561 170080 74641
rect 170390 74561 170400 74641
rect 170710 74561 170720 74641
rect 171030 74561 171040 74641
rect 30520 74520 30600 74530
rect 30840 74520 30920 74530
rect 31160 74520 31240 74530
rect 31480 74520 31560 74530
rect 31800 74520 31880 74530
rect 32120 74520 32200 74530
rect 32440 74520 32520 74530
rect 32760 74520 32840 74530
rect 33080 74520 33160 74530
rect 33400 74520 33480 74530
rect 33720 74520 33800 74530
rect 34040 74520 34120 74530
rect 34360 74520 34440 74530
rect 34680 74520 34760 74530
rect 35000 74520 35080 74530
rect 35320 74520 35400 74530
rect 35640 74520 35720 74530
rect 35960 74520 36040 74530
rect 36280 74520 36360 74530
rect 36600 74520 36680 74530
rect 36920 74520 37000 74530
rect 37240 74520 37320 74530
rect 37560 74520 37640 74530
rect 40340 74520 40420 74530
rect 40660 74520 40740 74530
rect 40980 74520 41060 74530
rect 42720 74520 42800 74530
rect 43040 74520 43120 74530
rect 43360 74520 43440 74530
rect 19130 74490 19210 74500
rect 19450 74490 19530 74500
rect 19770 74490 19850 74500
rect 20090 74490 20170 74500
rect 20410 74490 20490 74500
rect 20730 74490 20810 74500
rect 21050 74490 21130 74500
rect 21370 74490 21450 74500
rect 21690 74490 21770 74500
rect 22010 74490 22090 74500
rect 22330 74490 22410 74500
rect 22650 74490 22730 74500
rect 22970 74490 23050 74500
rect 23290 74490 23370 74500
rect 23610 74490 23690 74500
rect 23930 74490 24010 74500
rect 24250 74490 24330 74500
rect 24570 74490 24650 74500
rect 24890 74490 24970 74500
rect 25210 74490 25290 74500
rect 25530 74490 25610 74500
rect 25850 74490 25930 74500
rect 26170 74490 26250 74500
rect 19210 74410 19220 74490
rect 19530 74410 19540 74490
rect 19850 74410 19860 74490
rect 20170 74410 20180 74490
rect 20490 74410 20500 74490
rect 20810 74410 20820 74490
rect 21130 74410 21140 74490
rect 21450 74410 21460 74490
rect 21770 74410 21780 74490
rect 22090 74410 22100 74490
rect 22410 74410 22420 74490
rect 22730 74410 22740 74490
rect 23050 74410 23060 74490
rect 23370 74410 23380 74490
rect 23690 74410 23700 74490
rect 24010 74410 24020 74490
rect 24330 74410 24340 74490
rect 24650 74410 24660 74490
rect 24970 74410 24980 74490
rect 25290 74410 25300 74490
rect 25610 74410 25620 74490
rect 25930 74410 25940 74490
rect 26250 74410 26260 74490
rect 30600 74440 30610 74520
rect 30920 74440 30930 74520
rect 31240 74440 31250 74520
rect 31560 74440 31570 74520
rect 31880 74440 31890 74520
rect 32200 74440 32210 74520
rect 32520 74440 32530 74520
rect 32840 74440 32850 74520
rect 33160 74440 33170 74520
rect 33480 74440 33490 74520
rect 33800 74440 33810 74520
rect 34120 74440 34130 74520
rect 34440 74440 34450 74520
rect 34760 74440 34770 74520
rect 35080 74440 35090 74520
rect 35400 74440 35410 74520
rect 35720 74440 35730 74520
rect 36040 74440 36050 74520
rect 36360 74440 36370 74520
rect 36680 74440 36690 74520
rect 37000 74440 37010 74520
rect 37320 74440 37330 74520
rect 37640 74440 37650 74520
rect 40420 74440 40430 74520
rect 40740 74440 40750 74520
rect 41060 74440 41070 74520
rect 42800 74440 42810 74520
rect 43120 74440 43130 74520
rect 43440 74440 43450 74520
rect 146560 74511 146640 74521
rect 146880 74511 146960 74521
rect 147200 74511 147280 74521
rect 148940 74511 149020 74521
rect 149260 74511 149340 74521
rect 149580 74511 149660 74521
rect 152360 74511 152440 74521
rect 152680 74511 152760 74521
rect 153000 74511 153080 74521
rect 153320 74511 153400 74521
rect 153640 74511 153720 74521
rect 153960 74511 154040 74521
rect 154280 74511 154360 74521
rect 154600 74511 154680 74521
rect 154920 74511 155000 74521
rect 155240 74511 155320 74521
rect 155560 74511 155640 74521
rect 155880 74511 155960 74521
rect 156200 74511 156280 74521
rect 156520 74511 156600 74521
rect 156840 74511 156920 74521
rect 157160 74511 157240 74521
rect 157480 74511 157560 74521
rect 157800 74511 157880 74521
rect 158120 74511 158200 74521
rect 158440 74511 158520 74521
rect 158760 74511 158840 74521
rect 159080 74511 159160 74521
rect 159400 74511 159480 74521
rect 146640 74431 146650 74511
rect 146960 74431 146970 74511
rect 147280 74431 147290 74511
rect 149020 74431 149030 74511
rect 149340 74431 149350 74511
rect 149660 74431 149670 74511
rect 152440 74431 152450 74511
rect 152760 74431 152770 74511
rect 153080 74431 153090 74511
rect 153400 74431 153410 74511
rect 153720 74431 153730 74511
rect 154040 74431 154050 74511
rect 154360 74431 154370 74511
rect 154680 74431 154690 74511
rect 155000 74431 155010 74511
rect 155320 74431 155330 74511
rect 155640 74431 155650 74511
rect 155960 74431 155970 74511
rect 156280 74431 156290 74511
rect 156600 74431 156610 74511
rect 156920 74431 156930 74511
rect 157240 74431 157250 74511
rect 157560 74431 157570 74511
rect 157880 74431 157890 74511
rect 158200 74431 158210 74511
rect 158520 74431 158530 74511
rect 158840 74431 158850 74511
rect 159160 74431 159170 74511
rect 159480 74431 159490 74511
rect 163750 74481 163830 74491
rect 164070 74481 164150 74491
rect 164390 74481 164470 74491
rect 164710 74481 164790 74491
rect 165030 74481 165110 74491
rect 165350 74481 165430 74491
rect 165670 74481 165750 74491
rect 165990 74481 166070 74491
rect 166310 74481 166390 74491
rect 166630 74481 166710 74491
rect 166950 74481 167030 74491
rect 167270 74481 167350 74491
rect 167590 74481 167670 74491
rect 167910 74481 167990 74491
rect 168230 74481 168310 74491
rect 168550 74481 168630 74491
rect 168870 74481 168950 74491
rect 169190 74481 169270 74491
rect 169510 74481 169590 74491
rect 169830 74481 169910 74491
rect 170150 74481 170230 74491
rect 170470 74481 170550 74491
rect 170790 74481 170870 74491
rect 163830 74401 163840 74481
rect 164150 74401 164160 74481
rect 164470 74401 164480 74481
rect 164790 74401 164800 74481
rect 165110 74401 165120 74481
rect 165430 74401 165440 74481
rect 165750 74401 165760 74481
rect 166070 74401 166080 74481
rect 166390 74401 166400 74481
rect 166710 74401 166720 74481
rect 167030 74401 167040 74481
rect 167350 74401 167360 74481
rect 167670 74401 167680 74481
rect 167990 74401 168000 74481
rect 168310 74401 168320 74481
rect 168630 74401 168640 74481
rect 168950 74401 168960 74481
rect 169270 74401 169280 74481
rect 169590 74401 169600 74481
rect 169910 74401 169920 74481
rect 170230 74401 170240 74481
rect 170550 74401 170560 74481
rect 170870 74401 170880 74481
rect 30360 74360 30440 74370
rect 30680 74360 30760 74370
rect 31000 74360 31080 74370
rect 31320 74360 31400 74370
rect 31640 74360 31720 74370
rect 31960 74360 32040 74370
rect 32280 74360 32360 74370
rect 32600 74360 32680 74370
rect 32920 74360 33000 74370
rect 33240 74360 33320 74370
rect 33560 74360 33640 74370
rect 33880 74360 33960 74370
rect 34200 74360 34280 74370
rect 34520 74360 34600 74370
rect 34840 74360 34920 74370
rect 35160 74360 35240 74370
rect 35480 74360 35560 74370
rect 35800 74360 35880 74370
rect 36120 74360 36200 74370
rect 36440 74360 36520 74370
rect 36760 74360 36840 74370
rect 37080 74360 37160 74370
rect 37400 74360 37480 74370
rect 37720 74360 37800 74370
rect 40180 74360 40260 74370
rect 40500 74360 40580 74370
rect 40820 74360 40900 74370
rect 41140 74360 41220 74370
rect 42560 74360 42640 74370
rect 42880 74360 42960 74370
rect 43200 74360 43280 74370
rect 43520 74360 43600 74370
rect 18970 74330 19050 74340
rect 19290 74330 19370 74340
rect 19610 74330 19690 74340
rect 19930 74330 20010 74340
rect 20250 74330 20330 74340
rect 20570 74330 20650 74340
rect 20890 74330 20970 74340
rect 21210 74330 21290 74340
rect 21530 74330 21610 74340
rect 21850 74330 21930 74340
rect 22170 74330 22250 74340
rect 22490 74330 22570 74340
rect 22810 74330 22890 74340
rect 23130 74330 23210 74340
rect 23450 74330 23530 74340
rect 23770 74330 23850 74340
rect 24090 74330 24170 74340
rect 24410 74330 24490 74340
rect 24730 74330 24810 74340
rect 25050 74330 25130 74340
rect 25370 74330 25450 74340
rect 25690 74330 25770 74340
rect 26010 74330 26090 74340
rect 26330 74330 26410 74340
rect 19050 74250 19060 74330
rect 19370 74250 19380 74330
rect 19690 74250 19700 74330
rect 20010 74250 20020 74330
rect 20330 74250 20340 74330
rect 20650 74250 20660 74330
rect 20970 74250 20980 74330
rect 21290 74250 21300 74330
rect 21610 74250 21620 74330
rect 21930 74250 21940 74330
rect 22250 74250 22260 74330
rect 22570 74250 22580 74330
rect 22890 74250 22900 74330
rect 23210 74250 23220 74330
rect 23530 74250 23540 74330
rect 23850 74250 23860 74330
rect 24170 74250 24180 74330
rect 24490 74250 24500 74330
rect 24810 74250 24820 74330
rect 25130 74250 25140 74330
rect 25450 74250 25460 74330
rect 25770 74250 25780 74330
rect 26090 74250 26100 74330
rect 26410 74250 26420 74330
rect 30440 74280 30450 74360
rect 30760 74280 30770 74360
rect 31080 74280 31090 74360
rect 31400 74280 31410 74360
rect 31720 74280 31730 74360
rect 32040 74280 32050 74360
rect 32360 74280 32370 74360
rect 32680 74280 32690 74360
rect 33000 74280 33010 74360
rect 33320 74280 33330 74360
rect 33640 74280 33650 74360
rect 33960 74280 33970 74360
rect 34280 74280 34290 74360
rect 34600 74280 34610 74360
rect 34920 74280 34930 74360
rect 35240 74280 35250 74360
rect 35560 74280 35570 74360
rect 35880 74280 35890 74360
rect 36200 74280 36210 74360
rect 36520 74280 36530 74360
rect 36840 74280 36850 74360
rect 37160 74280 37170 74360
rect 37480 74280 37490 74360
rect 37800 74280 37810 74360
rect 40260 74280 40270 74360
rect 40580 74280 40590 74360
rect 40900 74280 40910 74360
rect 41220 74280 41230 74360
rect 42640 74280 42650 74360
rect 42960 74280 42970 74360
rect 43280 74280 43290 74360
rect 43600 74280 43610 74360
rect 146400 74351 146480 74361
rect 146720 74351 146800 74361
rect 147040 74351 147120 74361
rect 147360 74351 147440 74361
rect 148780 74351 148860 74361
rect 149100 74351 149180 74361
rect 149420 74351 149500 74361
rect 149740 74351 149820 74361
rect 152200 74351 152280 74361
rect 152520 74351 152600 74361
rect 152840 74351 152920 74361
rect 153160 74351 153240 74361
rect 153480 74351 153560 74361
rect 153800 74351 153880 74361
rect 154120 74351 154200 74361
rect 154440 74351 154520 74361
rect 154760 74351 154840 74361
rect 155080 74351 155160 74361
rect 155400 74351 155480 74361
rect 155720 74351 155800 74361
rect 156040 74351 156120 74361
rect 156360 74351 156440 74361
rect 156680 74351 156760 74361
rect 157000 74351 157080 74361
rect 157320 74351 157400 74361
rect 157640 74351 157720 74361
rect 157960 74351 158040 74361
rect 158280 74351 158360 74361
rect 158600 74351 158680 74361
rect 158920 74351 159000 74361
rect 159240 74351 159320 74361
rect 159560 74351 159640 74361
rect 146480 74271 146490 74351
rect 146800 74271 146810 74351
rect 147120 74271 147130 74351
rect 147440 74271 147450 74351
rect 148860 74271 148870 74351
rect 149180 74271 149190 74351
rect 149500 74271 149510 74351
rect 149820 74271 149830 74351
rect 152280 74271 152290 74351
rect 152600 74271 152610 74351
rect 152920 74271 152930 74351
rect 153240 74271 153250 74351
rect 153560 74271 153570 74351
rect 153880 74271 153890 74351
rect 154200 74271 154210 74351
rect 154520 74271 154530 74351
rect 154840 74271 154850 74351
rect 155160 74271 155170 74351
rect 155480 74271 155490 74351
rect 155800 74271 155810 74351
rect 156120 74271 156130 74351
rect 156440 74271 156450 74351
rect 156760 74271 156770 74351
rect 157080 74271 157090 74351
rect 157400 74271 157410 74351
rect 157720 74271 157730 74351
rect 158040 74271 158050 74351
rect 158360 74271 158370 74351
rect 158680 74271 158690 74351
rect 159000 74271 159010 74351
rect 159320 74271 159330 74351
rect 159640 74271 159650 74351
rect 163590 74321 163670 74331
rect 163910 74321 163990 74331
rect 164230 74321 164310 74331
rect 164550 74321 164630 74331
rect 164870 74321 164950 74331
rect 165190 74321 165270 74331
rect 165510 74321 165590 74331
rect 165830 74321 165910 74331
rect 166150 74321 166230 74331
rect 166470 74321 166550 74331
rect 166790 74321 166870 74331
rect 167110 74321 167190 74331
rect 167430 74321 167510 74331
rect 167750 74321 167830 74331
rect 168070 74321 168150 74331
rect 168390 74321 168470 74331
rect 168710 74321 168790 74331
rect 169030 74321 169110 74331
rect 169350 74321 169430 74331
rect 169670 74321 169750 74331
rect 169990 74321 170070 74331
rect 170310 74321 170390 74331
rect 170630 74321 170710 74331
rect 170950 74321 171030 74331
rect 163670 74241 163680 74321
rect 163990 74241 164000 74321
rect 164310 74241 164320 74321
rect 164630 74241 164640 74321
rect 164950 74241 164960 74321
rect 165270 74241 165280 74321
rect 165590 74241 165600 74321
rect 165910 74241 165920 74321
rect 166230 74241 166240 74321
rect 166550 74241 166560 74321
rect 166870 74241 166880 74321
rect 167190 74241 167200 74321
rect 167510 74241 167520 74321
rect 167830 74241 167840 74321
rect 168150 74241 168160 74321
rect 168470 74241 168480 74321
rect 168790 74241 168800 74321
rect 169110 74241 169120 74321
rect 169430 74241 169440 74321
rect 169750 74241 169760 74321
rect 170070 74241 170080 74321
rect 170390 74241 170400 74321
rect 170710 74241 170720 74321
rect 171030 74241 171040 74321
rect 30520 74200 30600 74210
rect 30840 74200 30920 74210
rect 31160 74200 31240 74210
rect 31480 74200 31560 74210
rect 31800 74200 31880 74210
rect 32120 74200 32200 74210
rect 32440 74200 32520 74210
rect 32760 74200 32840 74210
rect 33080 74200 33160 74210
rect 33400 74200 33480 74210
rect 33720 74200 33800 74210
rect 34040 74200 34120 74210
rect 34360 74200 34440 74210
rect 34680 74200 34760 74210
rect 35000 74200 35080 74210
rect 35320 74200 35400 74210
rect 35640 74200 35720 74210
rect 35960 74200 36040 74210
rect 36280 74200 36360 74210
rect 36600 74200 36680 74210
rect 36920 74200 37000 74210
rect 37240 74200 37320 74210
rect 37560 74200 37640 74210
rect 40340 74200 40420 74210
rect 40660 74200 40740 74210
rect 40980 74200 41060 74210
rect 42720 74200 42800 74210
rect 43040 74200 43120 74210
rect 43360 74200 43440 74210
rect 19130 74170 19210 74180
rect 19450 74170 19530 74180
rect 19770 74170 19850 74180
rect 20090 74170 20170 74180
rect 20410 74170 20490 74180
rect 20730 74170 20810 74180
rect 21050 74170 21130 74180
rect 21370 74170 21450 74180
rect 21690 74170 21770 74180
rect 22010 74170 22090 74180
rect 22330 74170 22410 74180
rect 22650 74170 22730 74180
rect 22970 74170 23050 74180
rect 23290 74170 23370 74180
rect 23610 74170 23690 74180
rect 23930 74170 24010 74180
rect 24250 74170 24330 74180
rect 24570 74170 24650 74180
rect 24890 74170 24970 74180
rect 25210 74170 25290 74180
rect 25530 74170 25610 74180
rect 25850 74170 25930 74180
rect 26170 74170 26250 74180
rect 19210 74090 19220 74170
rect 19530 74090 19540 74170
rect 19850 74090 19860 74170
rect 20170 74090 20180 74170
rect 20490 74090 20500 74170
rect 20810 74090 20820 74170
rect 21130 74090 21140 74170
rect 21450 74090 21460 74170
rect 21770 74090 21780 74170
rect 22090 74090 22100 74170
rect 22410 74090 22420 74170
rect 22730 74090 22740 74170
rect 23050 74090 23060 74170
rect 23370 74090 23380 74170
rect 23690 74090 23700 74170
rect 24010 74090 24020 74170
rect 24330 74090 24340 74170
rect 24650 74090 24660 74170
rect 24970 74090 24980 74170
rect 25290 74090 25300 74170
rect 25610 74090 25620 74170
rect 25930 74090 25940 74170
rect 26250 74090 26260 74170
rect 30600 74120 30610 74200
rect 30920 74120 30930 74200
rect 31240 74120 31250 74200
rect 31560 74120 31570 74200
rect 31880 74120 31890 74200
rect 32200 74120 32210 74200
rect 32520 74120 32530 74200
rect 32840 74120 32850 74200
rect 33160 74120 33170 74200
rect 33480 74120 33490 74200
rect 33800 74120 33810 74200
rect 34120 74120 34130 74200
rect 34440 74120 34450 74200
rect 34760 74120 34770 74200
rect 35080 74120 35090 74200
rect 35400 74120 35410 74200
rect 35720 74120 35730 74200
rect 36040 74120 36050 74200
rect 36360 74120 36370 74200
rect 36680 74120 36690 74200
rect 37000 74120 37010 74200
rect 37320 74120 37330 74200
rect 37640 74120 37650 74200
rect 40420 74120 40430 74200
rect 40740 74120 40750 74200
rect 41060 74120 41070 74200
rect 42800 74120 42810 74200
rect 43120 74120 43130 74200
rect 43440 74120 43450 74200
rect 146560 74191 146640 74201
rect 146880 74191 146960 74201
rect 147200 74191 147280 74201
rect 148940 74191 149020 74201
rect 149260 74191 149340 74201
rect 149580 74191 149660 74201
rect 152360 74191 152440 74201
rect 152680 74191 152760 74201
rect 153000 74191 153080 74201
rect 153320 74191 153400 74201
rect 153640 74191 153720 74201
rect 153960 74191 154040 74201
rect 154280 74191 154360 74201
rect 154600 74191 154680 74201
rect 154920 74191 155000 74201
rect 155240 74191 155320 74201
rect 155560 74191 155640 74201
rect 155880 74191 155960 74201
rect 156200 74191 156280 74201
rect 156520 74191 156600 74201
rect 156840 74191 156920 74201
rect 157160 74191 157240 74201
rect 157480 74191 157560 74201
rect 157800 74191 157880 74201
rect 158120 74191 158200 74201
rect 158440 74191 158520 74201
rect 158760 74191 158840 74201
rect 159080 74191 159160 74201
rect 159400 74191 159480 74201
rect 46660 73960 47160 74140
rect 146640 74111 146650 74191
rect 146960 74111 146970 74191
rect 147280 74111 147290 74191
rect 149020 74111 149030 74191
rect 149340 74111 149350 74191
rect 149660 74111 149670 74191
rect 152440 74111 152450 74191
rect 152760 74111 152770 74191
rect 153080 74111 153090 74191
rect 153400 74111 153410 74191
rect 153720 74111 153730 74191
rect 154040 74111 154050 74191
rect 154360 74111 154370 74191
rect 154680 74111 154690 74191
rect 155000 74111 155010 74191
rect 155320 74111 155330 74191
rect 155640 74111 155650 74191
rect 155960 74111 155970 74191
rect 156280 74111 156290 74191
rect 156600 74111 156610 74191
rect 156920 74111 156930 74191
rect 157240 74111 157250 74191
rect 157560 74111 157570 74191
rect 157880 74111 157890 74191
rect 158200 74111 158210 74191
rect 158520 74111 158530 74191
rect 158840 74111 158850 74191
rect 159160 74111 159170 74191
rect 159480 74111 159490 74191
rect 163750 74161 163830 74171
rect 164070 74161 164150 74171
rect 164390 74161 164470 74171
rect 164710 74161 164790 74171
rect 165030 74161 165110 74171
rect 165350 74161 165430 74171
rect 165670 74161 165750 74171
rect 165990 74161 166070 74171
rect 166310 74161 166390 74171
rect 166630 74161 166710 74171
rect 166950 74161 167030 74171
rect 167270 74161 167350 74171
rect 167590 74161 167670 74171
rect 167910 74161 167990 74171
rect 168230 74161 168310 74171
rect 168550 74161 168630 74171
rect 168870 74161 168950 74171
rect 169190 74161 169270 74171
rect 169510 74161 169590 74171
rect 169830 74161 169910 74171
rect 170150 74161 170230 74171
rect 170470 74161 170550 74171
rect 170790 74161 170870 74171
rect 163830 74081 163840 74161
rect 164150 74081 164160 74161
rect 164470 74081 164480 74161
rect 164790 74081 164800 74161
rect 165110 74081 165120 74161
rect 165430 74081 165440 74161
rect 165750 74081 165760 74161
rect 166070 74081 166080 74161
rect 166390 74081 166400 74161
rect 166710 74081 166720 74161
rect 167030 74081 167040 74161
rect 167350 74081 167360 74161
rect 167670 74081 167680 74161
rect 167990 74081 168000 74161
rect 168310 74081 168320 74161
rect 168630 74081 168640 74161
rect 168950 74081 168960 74161
rect 169270 74081 169280 74161
rect 169590 74081 169600 74161
rect 169910 74081 169920 74161
rect 170230 74081 170240 74161
rect 170550 74081 170560 74161
rect 170870 74081 170880 74161
rect 18980 73940 19060 73950
rect 19160 73940 19240 73950
rect 19340 73940 19420 73950
rect 19520 73940 19600 73950
rect 19700 73940 19780 73950
rect 19880 73940 19960 73950
rect 20060 73940 20140 73950
rect 20240 73940 20320 73950
rect 20420 73940 20500 73950
rect 20600 73940 20680 73950
rect 20780 73940 20860 73950
rect 20960 73940 21040 73950
rect 21140 73940 21220 73950
rect 21320 73940 21400 73950
rect 21500 73940 21580 73950
rect 21680 73940 21760 73950
rect 21860 73940 21940 73950
rect 22040 73940 22120 73950
rect 22220 73940 22300 73950
rect 22400 73940 22480 73950
rect 22580 73940 22660 73950
rect 22760 73940 22840 73950
rect 22940 73940 23020 73950
rect 23120 73940 23200 73950
rect 23300 73940 23380 73950
rect 23480 73940 23560 73950
rect 23660 73940 23740 73950
rect 23840 73940 23920 73950
rect 24020 73940 24100 73950
rect 24200 73940 24280 73950
rect 24380 73940 24460 73950
rect 24560 73940 24640 73950
rect 24740 73940 24820 73950
rect 24920 73940 25000 73950
rect 25100 73940 25180 73950
rect 25280 73940 25360 73950
rect 25460 73940 25540 73950
rect 25640 73940 25720 73950
rect 25820 73940 25900 73950
rect 26000 73940 26080 73950
rect 26180 73940 26260 73950
rect 26360 73940 26440 73950
rect 26540 73940 26620 73950
rect 30280 73940 30360 73950
rect 30460 73940 30540 73950
rect 30640 73940 30720 73950
rect 30820 73940 30900 73950
rect 31000 73940 31080 73950
rect 31180 73940 31260 73950
rect 31360 73940 31440 73950
rect 31540 73940 31620 73950
rect 31720 73940 31800 73950
rect 31900 73940 31980 73950
rect 32080 73940 32160 73950
rect 32260 73940 32340 73950
rect 32440 73940 32520 73950
rect 32620 73940 32700 73950
rect 32800 73940 32880 73950
rect 32980 73940 33060 73950
rect 33160 73940 33240 73950
rect 33340 73940 33420 73950
rect 33520 73940 33600 73950
rect 33700 73940 33780 73950
rect 33880 73940 33960 73950
rect 34060 73940 34140 73950
rect 34240 73940 34320 73950
rect 34420 73940 34500 73950
rect 34600 73940 34680 73950
rect 34780 73940 34860 73950
rect 34960 73940 35040 73950
rect 35140 73940 35220 73950
rect 35320 73940 35400 73950
rect 35500 73940 35580 73950
rect 35680 73940 35760 73950
rect 35860 73940 35940 73950
rect 36040 73940 36120 73950
rect 36220 73940 36300 73950
rect 36400 73940 36480 73950
rect 36580 73940 36660 73950
rect 36760 73940 36840 73950
rect 36940 73940 37020 73950
rect 37120 73940 37200 73950
rect 37300 73940 37380 73950
rect 37480 73940 37560 73950
rect 37660 73940 37740 73950
rect 37840 73940 37920 73950
rect 40060 73940 40140 73950
rect 40200 73940 40280 73950
rect 40340 73940 40420 73950
rect 40480 73940 40560 73950
rect 40620 73940 40700 73950
rect 40760 73940 40840 73950
rect 40900 73940 40980 73950
rect 41040 73940 41120 73950
rect 41180 73940 41260 73950
rect 41320 73940 41400 73950
rect 42360 73940 42440 73950
rect 42500 73940 42580 73950
rect 42640 73940 42720 73950
rect 42780 73940 42860 73950
rect 42920 73940 43000 73950
rect 43060 73940 43140 73950
rect 43200 73940 43280 73950
rect 43340 73940 43420 73950
rect 43480 73940 43560 73950
rect 43620 73940 43700 73950
rect 146300 73940 146380 73950
rect 146440 73940 146520 73950
rect 146580 73940 146660 73950
rect 146720 73940 146800 73950
rect 146860 73940 146940 73950
rect 147000 73940 147080 73950
rect 147140 73940 147220 73950
rect 147280 73940 147360 73950
rect 147420 73940 147500 73950
rect 147560 73940 147640 73950
rect 148600 73940 148680 73950
rect 148740 73940 148820 73950
rect 148880 73940 148960 73950
rect 149020 73940 149100 73950
rect 149160 73940 149240 73950
rect 149300 73940 149380 73950
rect 149440 73940 149520 73950
rect 149580 73940 149660 73950
rect 149720 73940 149800 73950
rect 149860 73940 149940 73950
rect 152080 73940 152160 73950
rect 152260 73940 152340 73950
rect 152440 73940 152520 73950
rect 152620 73940 152700 73950
rect 152800 73940 152880 73950
rect 152980 73940 153060 73950
rect 153160 73940 153240 73950
rect 153340 73940 153420 73950
rect 153520 73940 153600 73950
rect 153700 73940 153780 73950
rect 153880 73940 153960 73950
rect 154060 73940 154140 73950
rect 154240 73940 154320 73950
rect 154420 73940 154500 73950
rect 154600 73940 154680 73950
rect 154780 73940 154860 73950
rect 154960 73940 155040 73950
rect 155140 73940 155220 73950
rect 155320 73940 155400 73950
rect 155500 73940 155580 73950
rect 155680 73940 155760 73950
rect 155860 73940 155940 73950
rect 156040 73940 156120 73950
rect 156220 73940 156300 73950
rect 156400 73940 156480 73950
rect 156580 73940 156660 73950
rect 156760 73940 156840 73950
rect 156940 73940 157020 73950
rect 157120 73940 157200 73950
rect 157300 73940 157380 73950
rect 157480 73940 157560 73950
rect 157660 73940 157740 73950
rect 157840 73940 157920 73950
rect 158020 73940 158100 73950
rect 158200 73940 158280 73950
rect 158380 73940 158460 73950
rect 158560 73940 158640 73950
rect 158740 73940 158820 73950
rect 158920 73940 159000 73950
rect 159100 73940 159180 73950
rect 159280 73940 159360 73950
rect 159460 73940 159540 73950
rect 159640 73940 159720 73950
rect 163380 73940 163460 73950
rect 163560 73940 163640 73950
rect 163740 73940 163820 73950
rect 163920 73940 164000 73950
rect 164100 73940 164180 73950
rect 164280 73940 164360 73950
rect 164460 73940 164540 73950
rect 164640 73940 164720 73950
rect 164820 73940 164900 73950
rect 165000 73940 165080 73950
rect 165180 73940 165260 73950
rect 165360 73940 165440 73950
rect 165540 73940 165620 73950
rect 165720 73940 165800 73950
rect 165900 73940 165980 73950
rect 166080 73940 166160 73950
rect 166260 73940 166340 73950
rect 166440 73940 166520 73950
rect 166620 73940 166700 73950
rect 166800 73940 166880 73950
rect 166980 73940 167060 73950
rect 167160 73940 167240 73950
rect 167340 73940 167420 73950
rect 167520 73940 167600 73950
rect 167700 73940 167780 73950
rect 167880 73940 167960 73950
rect 168060 73940 168140 73950
rect 168240 73940 168320 73950
rect 168420 73940 168500 73950
rect 168600 73940 168680 73950
rect 168780 73940 168860 73950
rect 168960 73940 169040 73950
rect 169140 73940 169220 73950
rect 169320 73940 169400 73950
rect 169500 73940 169580 73950
rect 169680 73940 169760 73950
rect 169860 73940 169940 73950
rect 170040 73940 170120 73950
rect 170220 73940 170300 73950
rect 170400 73940 170480 73950
rect 170580 73940 170660 73950
rect 170760 73940 170840 73950
rect 170940 73940 171020 73950
rect 19060 73860 19070 73940
rect 19240 73860 19250 73940
rect 19420 73860 19430 73940
rect 19600 73860 19610 73940
rect 19780 73860 19790 73940
rect 19960 73860 19970 73940
rect 20140 73860 20150 73940
rect 20320 73860 20330 73940
rect 20500 73860 20510 73940
rect 20680 73860 20690 73940
rect 20860 73860 20870 73940
rect 21040 73860 21050 73940
rect 21220 73860 21230 73940
rect 21400 73860 21410 73940
rect 21580 73860 21590 73940
rect 21760 73860 21770 73940
rect 21940 73860 21950 73940
rect 22120 73860 22130 73940
rect 22300 73860 22310 73940
rect 22480 73860 22490 73940
rect 22660 73860 22670 73940
rect 22840 73860 22850 73940
rect 23020 73860 23030 73940
rect 23200 73860 23210 73940
rect 23380 73860 23390 73940
rect 23560 73860 23570 73940
rect 23740 73860 23750 73940
rect 23920 73860 23930 73940
rect 24100 73860 24110 73940
rect 24280 73860 24290 73940
rect 24460 73860 24470 73940
rect 24640 73860 24650 73940
rect 24820 73860 24830 73940
rect 25000 73860 25010 73940
rect 25180 73860 25190 73940
rect 25360 73860 25370 73940
rect 25540 73860 25550 73940
rect 25720 73860 25730 73940
rect 25900 73860 25910 73940
rect 26080 73860 26090 73940
rect 26260 73860 26270 73940
rect 26440 73860 26450 73940
rect 26620 73860 26630 73940
rect 30360 73860 30370 73940
rect 30540 73860 30550 73940
rect 30720 73860 30730 73940
rect 30900 73860 30910 73940
rect 31080 73860 31090 73940
rect 31260 73860 31270 73940
rect 31440 73860 31450 73940
rect 31620 73860 31630 73940
rect 31800 73860 31810 73940
rect 31980 73860 31990 73940
rect 32160 73860 32170 73940
rect 32340 73860 32350 73940
rect 32520 73860 32530 73940
rect 32700 73860 32710 73940
rect 32880 73860 32890 73940
rect 33060 73860 33070 73940
rect 33240 73860 33250 73940
rect 33420 73860 33430 73940
rect 33600 73860 33610 73940
rect 33780 73860 33790 73940
rect 33960 73860 33970 73940
rect 34140 73860 34150 73940
rect 34320 73860 34330 73940
rect 34500 73860 34510 73940
rect 34680 73860 34690 73940
rect 34860 73860 34870 73940
rect 35040 73860 35050 73940
rect 35220 73860 35230 73940
rect 35400 73860 35410 73940
rect 35580 73860 35590 73940
rect 35760 73860 35770 73940
rect 35940 73860 35950 73940
rect 36120 73860 36130 73940
rect 36300 73860 36310 73940
rect 36480 73860 36490 73940
rect 36660 73860 36670 73940
rect 36840 73860 36850 73940
rect 37020 73860 37030 73940
rect 37200 73860 37210 73940
rect 37380 73860 37390 73940
rect 37560 73860 37570 73940
rect 37740 73860 37750 73940
rect 37920 73860 37930 73940
rect 40140 73860 40150 73940
rect 40280 73860 40290 73940
rect 40420 73860 40430 73940
rect 40560 73860 40570 73940
rect 40700 73860 40710 73940
rect 40840 73860 40850 73940
rect 40980 73860 40990 73940
rect 41120 73860 41130 73940
rect 41260 73860 41270 73940
rect 41400 73860 41410 73940
rect 42440 73860 42450 73940
rect 42580 73860 42590 73940
rect 42720 73860 42730 73940
rect 42860 73860 42870 73940
rect 43000 73860 43010 73940
rect 43140 73860 43150 73940
rect 43280 73860 43290 73940
rect 43420 73860 43430 73940
rect 43560 73860 43570 73940
rect 43700 73860 43710 73940
rect 146380 73860 146390 73940
rect 146520 73860 146530 73940
rect 146660 73860 146670 73940
rect 146800 73860 146810 73940
rect 146940 73860 146950 73940
rect 147080 73860 147090 73940
rect 147220 73860 147230 73940
rect 147360 73860 147370 73940
rect 147500 73860 147510 73940
rect 147640 73860 147650 73940
rect 148680 73860 148690 73940
rect 148820 73860 148830 73940
rect 148960 73860 148970 73940
rect 149100 73860 149110 73940
rect 149240 73860 149250 73940
rect 149380 73860 149390 73940
rect 149520 73860 149530 73940
rect 149660 73860 149670 73940
rect 149800 73860 149810 73940
rect 149940 73860 149950 73940
rect 152160 73860 152170 73940
rect 152340 73860 152350 73940
rect 152520 73860 152530 73940
rect 152700 73860 152710 73940
rect 152880 73860 152890 73940
rect 153060 73860 153070 73940
rect 153240 73860 153250 73940
rect 153420 73860 153430 73940
rect 153600 73860 153610 73940
rect 153780 73860 153790 73940
rect 153960 73860 153970 73940
rect 154140 73860 154150 73940
rect 154320 73860 154330 73940
rect 154500 73860 154510 73940
rect 154680 73860 154690 73940
rect 154860 73860 154870 73940
rect 155040 73860 155050 73940
rect 155220 73860 155230 73940
rect 155400 73860 155410 73940
rect 155580 73860 155590 73940
rect 155760 73860 155770 73940
rect 155940 73860 155950 73940
rect 156120 73860 156130 73940
rect 156300 73860 156310 73940
rect 156480 73860 156490 73940
rect 156660 73860 156670 73940
rect 156840 73860 156850 73940
rect 157020 73860 157030 73940
rect 157200 73860 157210 73940
rect 157380 73860 157390 73940
rect 157560 73860 157570 73940
rect 157740 73860 157750 73940
rect 157920 73860 157930 73940
rect 158100 73860 158110 73940
rect 158280 73860 158290 73940
rect 158460 73860 158470 73940
rect 158640 73860 158650 73940
rect 158820 73860 158830 73940
rect 159000 73860 159010 73940
rect 159180 73860 159190 73940
rect 159360 73860 159370 73940
rect 159540 73860 159550 73940
rect 159720 73860 159730 73940
rect 163460 73860 163470 73940
rect 163640 73860 163650 73940
rect 163820 73860 163830 73940
rect 164000 73860 164010 73940
rect 164180 73860 164190 73940
rect 164360 73860 164370 73940
rect 164540 73860 164550 73940
rect 164720 73860 164730 73940
rect 164900 73860 164910 73940
rect 165080 73860 165090 73940
rect 165260 73860 165270 73940
rect 165440 73860 165450 73940
rect 165620 73860 165630 73940
rect 165800 73860 165810 73940
rect 165980 73860 165990 73940
rect 166160 73860 166170 73940
rect 166340 73860 166350 73940
rect 166520 73860 166530 73940
rect 166700 73860 166710 73940
rect 166880 73860 166890 73940
rect 167060 73860 167070 73940
rect 167240 73860 167250 73940
rect 167420 73860 167430 73940
rect 167600 73860 167610 73940
rect 167780 73860 167790 73940
rect 167960 73860 167970 73940
rect 168140 73860 168150 73940
rect 168320 73860 168330 73940
rect 168500 73860 168510 73940
rect 168680 73860 168690 73940
rect 168860 73860 168870 73940
rect 169040 73860 169050 73940
rect 169220 73860 169230 73940
rect 169400 73860 169410 73940
rect 169580 73860 169590 73940
rect 169760 73860 169770 73940
rect 169940 73860 169950 73940
rect 170120 73860 170130 73940
rect 170300 73860 170310 73940
rect 170480 73860 170490 73940
rect 170660 73860 170670 73940
rect 170840 73860 170850 73940
rect 171020 73860 171030 73940
rect 161885 73845 161965 73855
rect 162065 73845 162145 73855
rect 162245 73845 162325 73855
rect 162425 73845 162505 73855
rect 162605 73845 162685 73855
rect 28850 73815 28930 73825
rect 29010 73815 29090 73825
rect 29170 73815 29250 73825
rect 29330 73815 29410 73825
rect 29490 73815 29570 73825
rect 18980 73790 19060 73800
rect 19160 73790 19240 73800
rect 19340 73790 19420 73800
rect 19520 73790 19600 73800
rect 19700 73790 19780 73800
rect 19880 73790 19960 73800
rect 20060 73790 20140 73800
rect 20240 73790 20320 73800
rect 20420 73790 20500 73800
rect 20600 73790 20680 73800
rect 20780 73790 20860 73800
rect 20960 73790 21040 73800
rect 21140 73790 21220 73800
rect 21320 73790 21400 73800
rect 21500 73790 21580 73800
rect 21680 73790 21760 73800
rect 21860 73790 21940 73800
rect 22040 73790 22120 73800
rect 22220 73790 22300 73800
rect 22400 73790 22480 73800
rect 22580 73790 22660 73800
rect 22760 73790 22840 73800
rect 22940 73790 23020 73800
rect 23120 73790 23200 73800
rect 23300 73790 23380 73800
rect 23480 73790 23560 73800
rect 23660 73790 23740 73800
rect 23840 73790 23920 73800
rect 24020 73790 24100 73800
rect 24200 73790 24280 73800
rect 24380 73790 24460 73800
rect 24560 73790 24640 73800
rect 24740 73790 24820 73800
rect 24920 73790 25000 73800
rect 25100 73790 25180 73800
rect 25280 73790 25360 73800
rect 25460 73790 25540 73800
rect 25640 73790 25720 73800
rect 25820 73790 25900 73800
rect 26000 73790 26080 73800
rect 26180 73790 26260 73800
rect 26360 73790 26440 73800
rect 26540 73790 26620 73800
rect 19060 73710 19070 73790
rect 19240 73710 19250 73790
rect 19420 73710 19430 73790
rect 19600 73710 19610 73790
rect 19780 73710 19790 73790
rect 19960 73710 19970 73790
rect 20140 73710 20150 73790
rect 20320 73710 20330 73790
rect 20500 73710 20510 73790
rect 20680 73710 20690 73790
rect 20860 73710 20870 73790
rect 21040 73710 21050 73790
rect 21220 73710 21230 73790
rect 21400 73710 21410 73790
rect 21580 73710 21590 73790
rect 21760 73710 21770 73790
rect 21940 73710 21950 73790
rect 22120 73710 22130 73790
rect 22300 73710 22310 73790
rect 22480 73710 22490 73790
rect 22660 73710 22670 73790
rect 22840 73710 22850 73790
rect 23020 73710 23030 73790
rect 23200 73710 23210 73790
rect 23380 73710 23390 73790
rect 23560 73710 23570 73790
rect 23740 73710 23750 73790
rect 23920 73710 23930 73790
rect 24100 73710 24110 73790
rect 24280 73710 24290 73790
rect 24460 73710 24470 73790
rect 24640 73710 24650 73790
rect 24820 73710 24830 73790
rect 25000 73710 25010 73790
rect 25180 73710 25190 73790
rect 25360 73710 25370 73790
rect 25540 73710 25550 73790
rect 25720 73710 25730 73790
rect 25900 73710 25910 73790
rect 26080 73710 26090 73790
rect 26260 73710 26270 73790
rect 26440 73710 26450 73790
rect 26620 73710 26630 73790
rect 28930 73735 28940 73815
rect 29010 73735 29020 73815
rect 29090 73735 29100 73815
rect 29170 73735 29180 73815
rect 29250 73735 29260 73815
rect 29330 73735 29340 73815
rect 29410 73735 29420 73815
rect 29490 73735 29500 73815
rect 29570 73735 29580 73815
rect 30280 73790 30360 73800
rect 30460 73790 30540 73800
rect 30640 73790 30720 73800
rect 30820 73790 30900 73800
rect 31000 73790 31080 73800
rect 31180 73790 31260 73800
rect 31360 73790 31440 73800
rect 31540 73790 31620 73800
rect 31720 73790 31800 73800
rect 31900 73790 31980 73800
rect 32080 73790 32160 73800
rect 32260 73790 32340 73800
rect 32440 73790 32520 73800
rect 32620 73790 32700 73800
rect 32800 73790 32880 73800
rect 32980 73790 33060 73800
rect 33160 73790 33240 73800
rect 33340 73790 33420 73800
rect 33520 73790 33600 73800
rect 33700 73790 33780 73800
rect 33880 73790 33960 73800
rect 34060 73790 34140 73800
rect 34240 73790 34320 73800
rect 34420 73790 34500 73800
rect 34600 73790 34680 73800
rect 34780 73790 34860 73800
rect 34960 73790 35040 73800
rect 35140 73790 35220 73800
rect 35320 73790 35400 73800
rect 35500 73790 35580 73800
rect 35680 73790 35760 73800
rect 35860 73790 35940 73800
rect 36040 73790 36120 73800
rect 36220 73790 36300 73800
rect 36400 73790 36480 73800
rect 36580 73790 36660 73800
rect 36760 73790 36840 73800
rect 36940 73790 37020 73800
rect 37120 73790 37200 73800
rect 37300 73790 37380 73800
rect 37480 73790 37560 73800
rect 37660 73790 37740 73800
rect 37840 73790 37920 73800
rect 152080 73790 152160 73800
rect 152260 73790 152340 73800
rect 152440 73790 152520 73800
rect 152620 73790 152700 73800
rect 152800 73790 152880 73800
rect 152980 73790 153060 73800
rect 153160 73790 153240 73800
rect 153340 73790 153420 73800
rect 153520 73790 153600 73800
rect 153700 73790 153780 73800
rect 153880 73790 153960 73800
rect 154060 73790 154140 73800
rect 154240 73790 154320 73800
rect 154420 73790 154500 73800
rect 154600 73790 154680 73800
rect 154780 73790 154860 73800
rect 154960 73790 155040 73800
rect 155140 73790 155220 73800
rect 155320 73790 155400 73800
rect 155500 73790 155580 73800
rect 155680 73790 155760 73800
rect 155860 73790 155940 73800
rect 156040 73790 156120 73800
rect 156220 73790 156300 73800
rect 156400 73790 156480 73800
rect 156580 73790 156660 73800
rect 156760 73790 156840 73800
rect 156940 73790 157020 73800
rect 157120 73790 157200 73800
rect 157300 73790 157380 73800
rect 157480 73790 157560 73800
rect 157660 73790 157740 73800
rect 157840 73790 157920 73800
rect 158020 73790 158100 73800
rect 158200 73790 158280 73800
rect 158380 73790 158460 73800
rect 158560 73790 158640 73800
rect 158740 73790 158820 73800
rect 158920 73790 159000 73800
rect 159100 73790 159180 73800
rect 159280 73790 159360 73800
rect 159460 73790 159540 73800
rect 159640 73790 159720 73800
rect 30360 73710 30370 73790
rect 30540 73710 30550 73790
rect 30720 73710 30730 73790
rect 30900 73710 30910 73790
rect 31080 73710 31090 73790
rect 31260 73710 31270 73790
rect 31440 73710 31450 73790
rect 31620 73710 31630 73790
rect 31800 73710 31810 73790
rect 31980 73710 31990 73790
rect 32160 73710 32170 73790
rect 32340 73710 32350 73790
rect 32520 73710 32530 73790
rect 32700 73710 32710 73790
rect 32880 73710 32890 73790
rect 33060 73710 33070 73790
rect 33240 73710 33250 73790
rect 33420 73710 33430 73790
rect 33600 73710 33610 73790
rect 33780 73710 33790 73790
rect 33960 73710 33970 73790
rect 34140 73710 34150 73790
rect 34320 73710 34330 73790
rect 34500 73710 34510 73790
rect 34680 73710 34690 73790
rect 34860 73710 34870 73790
rect 35040 73710 35050 73790
rect 35220 73710 35230 73790
rect 35400 73710 35410 73790
rect 35580 73710 35590 73790
rect 35760 73710 35770 73790
rect 35940 73710 35950 73790
rect 36120 73710 36130 73790
rect 36300 73710 36310 73790
rect 36480 73710 36490 73790
rect 36660 73710 36670 73790
rect 36840 73710 36850 73790
rect 37020 73710 37030 73790
rect 37200 73710 37210 73790
rect 37380 73710 37390 73790
rect 37560 73710 37570 73790
rect 37740 73710 37750 73790
rect 37920 73710 37930 73790
rect 40060 73690 40120 73720
rect 41540 73690 41600 73720
rect 42360 73690 42420 73720
rect 43840 73690 43900 73720
rect 152160 73710 152170 73790
rect 152340 73710 152350 73790
rect 152520 73710 152530 73790
rect 152700 73710 152710 73790
rect 152880 73710 152890 73790
rect 153060 73710 153070 73790
rect 153240 73710 153250 73790
rect 153420 73710 153430 73790
rect 153600 73710 153610 73790
rect 153780 73710 153790 73790
rect 153960 73710 153970 73790
rect 154140 73710 154150 73790
rect 154320 73710 154330 73790
rect 154500 73710 154510 73790
rect 154680 73710 154690 73790
rect 154860 73710 154870 73790
rect 155040 73710 155050 73790
rect 155220 73710 155230 73790
rect 155400 73710 155410 73790
rect 155580 73710 155590 73790
rect 155760 73710 155770 73790
rect 155940 73710 155950 73790
rect 156120 73710 156130 73790
rect 156300 73710 156310 73790
rect 156480 73710 156490 73790
rect 156660 73710 156670 73790
rect 156840 73710 156850 73790
rect 157020 73710 157030 73790
rect 157200 73710 157210 73790
rect 157380 73710 157390 73790
rect 157560 73710 157570 73790
rect 157740 73710 157750 73790
rect 157920 73710 157930 73790
rect 158100 73710 158110 73790
rect 158280 73710 158290 73790
rect 158460 73710 158470 73790
rect 158640 73710 158650 73790
rect 158820 73710 158830 73790
rect 159000 73710 159010 73790
rect 159180 73710 159190 73790
rect 159360 73710 159370 73790
rect 159540 73710 159550 73790
rect 159720 73710 159730 73790
rect 161965 73765 161975 73845
rect 162145 73765 162155 73845
rect 162325 73765 162335 73845
rect 162505 73765 162515 73845
rect 162685 73765 162695 73845
rect 163380 73790 163460 73800
rect 163560 73790 163640 73800
rect 163740 73790 163820 73800
rect 163920 73790 164000 73800
rect 164100 73790 164180 73800
rect 164280 73790 164360 73800
rect 164460 73790 164540 73800
rect 164640 73790 164720 73800
rect 164820 73790 164900 73800
rect 165000 73790 165080 73800
rect 165180 73790 165260 73800
rect 165360 73790 165440 73800
rect 165540 73790 165620 73800
rect 165720 73790 165800 73800
rect 165900 73790 165980 73800
rect 166080 73790 166160 73800
rect 166260 73790 166340 73800
rect 166440 73790 166520 73800
rect 166620 73790 166700 73800
rect 166800 73790 166880 73800
rect 166980 73790 167060 73800
rect 167160 73790 167240 73800
rect 167340 73790 167420 73800
rect 167520 73790 167600 73800
rect 167700 73790 167780 73800
rect 167880 73790 167960 73800
rect 168060 73790 168140 73800
rect 168240 73790 168320 73800
rect 168420 73790 168500 73800
rect 168600 73790 168680 73800
rect 168780 73790 168860 73800
rect 168960 73790 169040 73800
rect 169140 73790 169220 73800
rect 169320 73790 169400 73800
rect 169500 73790 169580 73800
rect 169680 73790 169760 73800
rect 169860 73790 169940 73800
rect 170040 73790 170120 73800
rect 170220 73790 170300 73800
rect 170400 73790 170480 73800
rect 170580 73790 170660 73800
rect 170760 73790 170840 73800
rect 170940 73790 171020 73800
rect 163460 73710 163470 73790
rect 163640 73710 163650 73790
rect 163820 73710 163830 73790
rect 164000 73710 164010 73790
rect 164180 73710 164190 73790
rect 164360 73710 164370 73790
rect 164540 73710 164550 73790
rect 164720 73710 164730 73790
rect 164900 73710 164910 73790
rect 165080 73710 165090 73790
rect 165260 73710 165270 73790
rect 165440 73710 165450 73790
rect 165620 73710 165630 73790
rect 165800 73710 165810 73790
rect 165980 73710 165990 73790
rect 166160 73710 166170 73790
rect 166340 73710 166350 73790
rect 166520 73710 166530 73790
rect 166700 73710 166710 73790
rect 166880 73710 166890 73790
rect 167060 73710 167070 73790
rect 167240 73710 167250 73790
rect 167420 73710 167430 73790
rect 167600 73710 167610 73790
rect 167780 73710 167790 73790
rect 167960 73710 167970 73790
rect 168140 73710 168150 73790
rect 168320 73710 168330 73790
rect 168500 73710 168510 73790
rect 168680 73710 168690 73790
rect 168860 73710 168870 73790
rect 169040 73710 169050 73790
rect 169220 73710 169230 73790
rect 169400 73710 169410 73790
rect 169580 73710 169590 73790
rect 169760 73710 169770 73790
rect 169940 73710 169950 73790
rect 170120 73710 170130 73790
rect 170300 73710 170310 73790
rect 170480 73710 170490 73790
rect 170660 73710 170670 73790
rect 170840 73710 170850 73790
rect 171020 73710 171030 73790
rect 146100 73650 146160 73680
rect 147580 73650 147640 73680
rect 148400 73650 148460 73680
rect 149880 73650 149940 73680
rect 161885 73665 161965 73675
rect 162065 73665 162145 73675
rect 162245 73665 162325 73675
rect 162425 73665 162505 73675
rect 162605 73665 162685 73675
rect 40060 73570 40120 73600
rect 41540 73570 41600 73600
rect 42360 73570 42420 73600
rect 43840 73570 43900 73600
rect 146100 73530 146160 73560
rect 146210 73540 146220 73630
rect 40060 73450 40120 73480
rect 41540 73450 41600 73480
rect 42360 73450 42420 73480
rect 43840 73450 43900 73480
rect 19130 73410 19160 73440
rect 19250 73410 19280 73440
rect 26420 73410 26450 73440
rect 26540 73410 26570 73440
rect 30420 73410 30450 73440
rect 30540 73410 30570 73440
rect 37720 73410 37750 73440
rect 37840 73410 37870 73440
rect 146100 73410 146160 73440
rect 19010 73380 19070 73410
rect 19130 73380 19190 73410
rect 19250 73380 19310 73410
rect 26300 73380 26360 73410
rect 26420 73380 26480 73410
rect 26540 73380 26600 73410
rect 30300 73380 30360 73410
rect 30420 73380 30480 73410
rect 30540 73380 30600 73410
rect 37600 73380 37660 73410
rect 37720 73380 37780 73410
rect 37840 73380 37900 73410
rect 40060 73330 40120 73360
rect 41540 73330 41600 73360
rect 42360 73330 42420 73360
rect 43840 73330 43900 73360
rect 19130 73290 19160 73320
rect 19250 73290 19280 73320
rect 26420 73290 26450 73320
rect 26540 73290 26570 73320
rect 30420 73290 30450 73320
rect 30540 73290 30570 73320
rect 37720 73290 37750 73320
rect 37840 73290 37870 73320
rect 146100 73290 146160 73320
rect 19010 73260 19070 73290
rect 19130 73260 19190 73290
rect 19250 73260 19310 73290
rect 26300 73260 26360 73290
rect 26420 73260 26480 73290
rect 26540 73260 26600 73290
rect 30300 73260 30360 73290
rect 30420 73260 30480 73290
rect 30540 73260 30600 73290
rect 37600 73260 37660 73290
rect 37720 73260 37780 73290
rect 37840 73260 37900 73290
rect 31010 73245 37190 73260
rect 36000 73170 37190 73245
rect 40060 73210 40120 73240
rect 41540 73210 41600 73240
rect 42360 73210 42420 73240
rect 43840 73210 43900 73240
rect 37720 73170 37750 73200
rect 37840 73170 37870 73200
rect 146100 73170 146160 73200
rect 36120 73150 36130 73170
rect 36300 73150 36310 73170
rect 36480 73150 36490 73170
rect 36660 73150 36670 73170
rect 36840 73150 36850 73170
rect 37020 73150 37030 73170
rect 36040 73080 36120 73090
rect 36220 73080 36300 73090
rect 36400 73080 36480 73090
rect 36580 73080 36660 73090
rect 36760 73080 36840 73090
rect 36940 73080 37020 73090
rect 36120 73000 36130 73080
rect 36300 73000 36310 73080
rect 36480 73000 36490 73080
rect 36660 73000 36670 73080
rect 36840 73000 36850 73080
rect 37020 73000 37030 73080
rect 37100 72940 37190 73170
rect 37600 73140 37660 73170
rect 37720 73140 37780 73170
rect 37840 73140 37900 73170
rect 40060 73090 40120 73120
rect 41540 73090 41600 73120
rect 42360 73090 42420 73120
rect 43840 73090 43900 73120
rect 37720 73050 37750 73080
rect 37840 73050 37870 73080
rect 146100 73050 146160 73080
rect 37600 73020 37660 73050
rect 37720 73020 37780 73050
rect 37840 73020 37900 73050
rect 40060 72970 40120 73000
rect 41540 72970 41600 73000
rect 42360 72970 42420 73000
rect 43840 72970 43900 73000
rect 36000 72910 37190 72940
rect 37720 72930 37750 72960
rect 37840 72930 37870 72960
rect 146100 72930 146160 72960
rect 36120 72850 36130 72910
rect 36300 72850 36310 72910
rect 36480 72850 36490 72910
rect 36660 72850 36670 72910
rect 36840 72850 36850 72910
rect 37020 72850 37030 72910
rect 37100 72840 37190 72910
rect 37600 72900 37660 72930
rect 37720 72900 37780 72930
rect 37840 72900 37900 72930
rect 40060 72850 40120 72880
rect 41540 72850 41600 72880
rect 42360 72850 42420 72880
rect 43840 72850 43900 72880
rect 36000 72810 37190 72840
rect 37720 72810 37750 72840
rect 37840 72810 37870 72840
rect 146100 72810 146160 72840
rect 37100 72800 37190 72810
rect 36000 72790 37190 72800
rect 36040 72610 36120 72620
rect 36220 72610 36300 72620
rect 36400 72610 36480 72620
rect 36580 72610 36660 72620
rect 36760 72610 36840 72620
rect 36940 72610 37020 72620
rect 36120 72530 36130 72610
rect 36300 72530 36310 72610
rect 36480 72530 36490 72610
rect 36660 72530 36670 72610
rect 36840 72530 36850 72610
rect 37020 72530 37030 72610
rect 36040 72290 36120 72300
rect 36220 72290 36300 72300
rect 36400 72290 36480 72300
rect 36580 72290 36660 72300
rect 36760 72290 36840 72300
rect 36940 72290 37020 72300
rect 36120 72210 36130 72290
rect 36300 72210 36310 72290
rect 36480 72210 36490 72290
rect 36660 72210 36670 72290
rect 36840 72210 36850 72290
rect 37020 72210 37030 72290
rect 37100 72120 37190 72790
rect 37600 72780 37660 72810
rect 37720 72780 37780 72810
rect 37840 72780 37900 72810
rect 40060 72730 40120 72760
rect 41540 72730 41600 72760
rect 42360 72730 42420 72760
rect 43840 72730 43900 72760
rect 37720 72690 37750 72720
rect 37840 72690 37870 72720
rect 146100 72690 146160 72720
rect 37600 72660 37660 72690
rect 37720 72660 37780 72690
rect 37840 72660 37900 72690
rect 40060 72610 40120 72640
rect 41540 72610 41600 72640
rect 42360 72610 42420 72640
rect 43840 72610 43900 72640
rect 37720 72570 37750 72600
rect 37840 72570 37870 72600
rect 146100 72570 146160 72600
rect 37600 72540 37660 72570
rect 37720 72540 37780 72570
rect 37840 72540 37900 72570
rect 40060 72490 40120 72520
rect 41540 72490 41600 72520
rect 42360 72490 42420 72520
rect 43840 72490 43900 72520
rect 37720 72450 37750 72480
rect 37840 72450 37870 72480
rect 146100 72450 146160 72480
rect 37600 72420 37660 72450
rect 37720 72420 37780 72450
rect 37840 72420 37900 72450
rect 40060 72370 40120 72400
rect 41540 72370 41600 72400
rect 42360 72370 42420 72400
rect 43840 72370 43900 72400
rect 37720 72330 37750 72360
rect 37840 72330 37870 72360
rect 146100 72330 146160 72360
rect 37600 72300 37660 72330
rect 37720 72300 37780 72330
rect 37840 72300 37900 72330
rect 40060 72250 40120 72280
rect 41540 72250 41600 72280
rect 42360 72250 42420 72280
rect 43840 72250 43900 72280
rect 37720 72210 37750 72240
rect 37840 72210 37870 72240
rect 146100 72210 146160 72240
rect 37600 72180 37660 72210
rect 37720 72180 37780 72210
rect 37840 72180 37900 72210
rect 40060 72130 40120 72160
rect 41540 72130 41600 72160
rect 42360 72130 42420 72160
rect 43840 72130 43900 72160
rect 146300 72150 146310 73540
rect 146690 73500 146810 73560
rect 146970 73500 147090 73560
rect 147580 73530 147640 73560
rect 148400 73530 148460 73560
rect 148820 73550 149620 73640
rect 148950 73520 149070 73550
rect 149230 73520 149350 73550
rect 149070 73510 149130 73520
rect 149350 73510 149410 73520
rect 149070 73500 149190 73510
rect 149350 73500 149470 73510
rect 146810 73490 146870 73500
rect 146570 73480 146650 73490
rect 146810 73480 146930 73490
rect 146650 73400 146660 73480
rect 146810 73380 146870 73480
rect 146930 73400 146940 73480
rect 147090 73380 147150 73500
rect 146410 73330 147140 73340
rect 146410 73250 146420 73330
rect 147220 73325 147230 73380
rect 147270 73350 147390 73410
rect 146460 73315 147250 73325
rect 146450 73265 146460 73315
rect 146500 73060 146510 73250
rect 146690 73200 146810 73260
rect 146970 73200 147090 73260
rect 147220 73236 147230 73315
rect 147390 73236 147450 73350
rect 147520 73236 147530 73470
rect 147580 73410 147640 73440
rect 148400 73410 148460 73440
rect 148510 73400 148520 73490
rect 147580 73290 147640 73320
rect 148400 73290 148460 73320
rect 148600 73236 148610 73400
rect 148650 73370 148770 73430
rect 149070 73400 149130 73500
rect 149190 73420 149200 73500
rect 149350 73400 149410 73500
rect 149470 73420 149480 73500
rect 148770 73345 148830 73370
rect 149530 73365 149620 73550
rect 148910 73360 149620 73365
rect 148900 73350 149630 73360
rect 148910 73345 149630 73350
rect 148770 73335 149630 73345
rect 148770 73250 148830 73335
rect 149530 73285 149630 73335
rect 148910 73255 149630 73285
rect 148950 73236 149070 73255
rect 149230 73236 149350 73255
rect 149530 73236 149630 73255
rect 149820 73236 149830 73650
rect 152080 73640 152160 73650
rect 152260 73640 152340 73650
rect 152440 73640 152520 73650
rect 152620 73640 152700 73650
rect 152800 73640 152880 73650
rect 152980 73640 153060 73650
rect 153160 73640 153240 73650
rect 153340 73640 153420 73650
rect 153520 73640 153600 73650
rect 153700 73640 153780 73650
rect 153880 73640 153960 73650
rect 154060 73640 154140 73650
rect 154240 73640 154320 73650
rect 154420 73640 154500 73650
rect 154600 73640 154680 73650
rect 154780 73640 154860 73650
rect 154960 73640 155040 73650
rect 155140 73640 155220 73650
rect 155320 73640 155400 73650
rect 155500 73640 155580 73650
rect 155680 73640 155760 73650
rect 155860 73640 155940 73650
rect 156040 73640 156120 73650
rect 156220 73640 156300 73650
rect 156400 73640 156480 73650
rect 156580 73640 156660 73650
rect 156760 73640 156840 73650
rect 156940 73640 157020 73650
rect 157120 73640 157200 73650
rect 157300 73640 157380 73650
rect 157480 73640 157560 73650
rect 157660 73640 157740 73650
rect 157840 73640 157920 73650
rect 158020 73640 158100 73650
rect 158200 73640 158280 73650
rect 158380 73640 158460 73650
rect 158560 73640 158640 73650
rect 158740 73640 158820 73650
rect 158920 73640 159000 73650
rect 159100 73640 159180 73650
rect 159280 73640 159360 73650
rect 159460 73640 159540 73650
rect 159640 73640 159720 73650
rect 152160 73560 152170 73640
rect 152340 73560 152350 73640
rect 152520 73560 152530 73640
rect 152700 73560 152710 73640
rect 152880 73560 152890 73640
rect 153060 73560 153070 73640
rect 153240 73560 153250 73640
rect 153420 73560 153430 73640
rect 153600 73560 153610 73640
rect 153780 73560 153790 73640
rect 153960 73560 153970 73640
rect 154140 73560 154150 73640
rect 154320 73560 154330 73640
rect 154500 73560 154510 73640
rect 154680 73560 154690 73640
rect 154860 73560 154870 73640
rect 155040 73560 155050 73640
rect 155220 73560 155230 73640
rect 155400 73560 155410 73640
rect 155580 73560 155590 73640
rect 155760 73560 155770 73640
rect 155940 73560 155950 73640
rect 156120 73560 156130 73640
rect 156300 73560 156310 73640
rect 156480 73560 156490 73640
rect 156660 73560 156670 73640
rect 156840 73560 156850 73640
rect 157020 73560 157030 73640
rect 157200 73560 157210 73640
rect 157380 73560 157390 73640
rect 157560 73560 157570 73640
rect 157740 73560 157750 73640
rect 157920 73560 157930 73640
rect 158100 73560 158110 73640
rect 158280 73560 158290 73640
rect 158460 73560 158470 73640
rect 158640 73560 158650 73640
rect 158820 73560 158830 73640
rect 159000 73560 159010 73640
rect 159180 73560 159190 73640
rect 159360 73560 159370 73640
rect 159540 73560 159550 73640
rect 159720 73560 159730 73640
rect 161965 73585 161975 73665
rect 162145 73585 162155 73665
rect 162325 73585 162335 73665
rect 162505 73585 162515 73665
rect 162685 73585 162695 73665
rect 163380 73640 163460 73650
rect 163560 73640 163640 73650
rect 163740 73640 163820 73650
rect 163920 73640 164000 73650
rect 164100 73640 164180 73650
rect 164280 73640 164360 73650
rect 164460 73640 164540 73650
rect 164640 73640 164720 73650
rect 164820 73640 164900 73650
rect 165000 73640 165080 73650
rect 165180 73640 165260 73650
rect 165360 73640 165440 73650
rect 165540 73640 165620 73650
rect 165720 73640 165800 73650
rect 165900 73640 165980 73650
rect 166080 73640 166160 73650
rect 166260 73640 166340 73650
rect 166440 73640 166520 73650
rect 166620 73640 166700 73650
rect 166800 73640 166880 73650
rect 166980 73640 167060 73650
rect 167160 73640 167240 73650
rect 167340 73640 167420 73650
rect 167520 73640 167600 73650
rect 167700 73640 167780 73650
rect 167880 73640 167960 73650
rect 168060 73640 168140 73650
rect 168240 73640 168320 73650
rect 168420 73640 168500 73650
rect 168600 73640 168680 73650
rect 168780 73640 168860 73650
rect 168960 73640 169040 73650
rect 169140 73640 169220 73650
rect 169320 73640 169400 73650
rect 169500 73640 169580 73650
rect 169680 73640 169760 73650
rect 169860 73640 169940 73650
rect 170040 73640 170120 73650
rect 170220 73640 170300 73650
rect 170400 73640 170480 73650
rect 170580 73640 170660 73650
rect 170760 73640 170840 73650
rect 170940 73640 171020 73650
rect 163460 73560 163470 73640
rect 163640 73560 163650 73640
rect 163820 73560 163830 73640
rect 164000 73560 164010 73640
rect 164180 73560 164190 73640
rect 164360 73560 164370 73640
rect 164540 73560 164550 73640
rect 164720 73560 164730 73640
rect 164900 73560 164910 73640
rect 165080 73560 165090 73640
rect 165260 73560 165270 73640
rect 165440 73560 165450 73640
rect 165620 73560 165630 73640
rect 165800 73560 165810 73640
rect 165980 73560 165990 73640
rect 166160 73560 166170 73640
rect 166340 73560 166350 73640
rect 166520 73560 166530 73640
rect 166700 73560 166710 73640
rect 166880 73560 166890 73640
rect 167060 73560 167070 73640
rect 167240 73560 167250 73640
rect 167420 73560 167430 73640
rect 167600 73560 167610 73640
rect 167780 73560 167790 73640
rect 167960 73560 167970 73640
rect 168140 73560 168150 73640
rect 168320 73560 168330 73640
rect 168500 73560 168510 73640
rect 168680 73560 168690 73640
rect 168860 73560 168870 73640
rect 169040 73560 169050 73640
rect 169220 73560 169230 73640
rect 169400 73560 169410 73640
rect 169580 73560 169590 73640
rect 169760 73560 169770 73640
rect 169940 73560 169950 73640
rect 170120 73560 170130 73640
rect 170300 73560 170310 73640
rect 170480 73560 170490 73640
rect 170660 73560 170670 73640
rect 170840 73560 170850 73640
rect 171020 73560 171030 73640
rect 149880 73530 149940 73560
rect 149880 73410 149940 73440
rect 152220 73390 152250 73420
rect 152340 73390 152370 73420
rect 159520 73390 159550 73420
rect 159640 73390 159670 73420
rect 152100 73360 152160 73390
rect 152220 73360 152280 73390
rect 152340 73360 152400 73390
rect 159400 73360 159460 73390
rect 159520 73360 159580 73390
rect 159640 73360 159700 73390
rect 149880 73290 149940 73320
rect 152220 73270 152250 73300
rect 152340 73270 152370 73300
rect 159520 73270 159550 73300
rect 159640 73270 159670 73300
rect 163520 73270 163550 73300
rect 163640 73270 163670 73300
rect 170810 73270 170840 73300
rect 170930 73270 170960 73300
rect 152100 73240 152160 73270
rect 152220 73240 152280 73270
rect 152340 73240 152400 73270
rect 152810 73236 158990 73260
rect 159400 73240 159460 73270
rect 159520 73240 159580 73270
rect 159640 73240 159700 73270
rect 163400 73240 163460 73270
rect 163520 73240 163580 73270
rect 163640 73240 163700 73270
rect 170690 73240 170750 73270
rect 170810 73240 170870 73270
rect 170930 73240 170990 73270
rect 164280 73236 164360 73240
rect 164460 73236 164540 73240
rect 164640 73236 164720 73240
rect 164820 73236 164900 73240
rect 165000 73236 165080 73240
rect 165180 73236 165260 73240
rect 165360 73236 165440 73240
rect 165540 73236 165620 73240
rect 165720 73236 165800 73240
rect 165900 73236 165980 73240
rect 166080 73236 166160 73240
rect 166260 73236 166340 73240
rect 166440 73236 166520 73240
rect 166620 73236 166700 73240
rect 166800 73236 166880 73240
rect 166980 73236 167060 73240
rect 167160 73236 167240 73240
rect 167340 73236 167420 73240
rect 167520 73236 167600 73240
rect 167700 73236 167780 73240
rect 167880 73236 167960 73240
rect 168060 73236 168140 73240
rect 168240 73236 168320 73240
rect 168420 73236 168500 73240
rect 168600 73236 168680 73240
rect 168780 73236 168860 73240
rect 168960 73236 169040 73240
rect 169140 73236 169220 73240
rect 169320 73236 169400 73240
rect 169500 73236 169580 73240
rect 169680 73236 169760 73240
rect 169860 73236 169940 73240
rect 170040 73236 170120 73240
rect 146810 73190 146870 73200
rect 146570 73180 146650 73190
rect 146710 73180 146790 73190
rect 146810 73180 146930 73190
rect 146990 73180 147070 73190
rect 146650 73100 146660 73180
rect 146790 73100 146800 73180
rect 146810 73080 146870 73180
rect 146930 73100 146940 73180
rect 147070 73100 147080 73180
rect 147090 73080 147150 73200
rect 146500 73050 147130 73060
rect 146500 73040 146510 73050
rect 146690 72910 146810 72970
rect 146970 72910 147090 72970
rect 146690 72820 146700 72910
rect 146800 72880 146870 72910
rect 146810 72790 146870 72880
rect 146970 72820 146980 72910
rect 147090 72790 147150 72910
rect 146410 72740 147140 72750
rect 146410 72660 146420 72740
rect 146460 72725 147150 72735
rect 146450 72675 146460 72725
rect 146500 72470 146510 72660
rect 146690 72610 146810 72670
rect 146970 72610 147090 72670
rect 146810 72600 146870 72610
rect 146570 72590 146650 72600
rect 146710 72590 146790 72600
rect 146810 72590 146930 72600
rect 146990 72590 147070 72600
rect 146650 72510 146660 72590
rect 146790 72510 146800 72590
rect 146810 72490 146870 72590
rect 146930 72510 146940 72590
rect 147070 72510 147080 72590
rect 147090 72490 147150 72610
rect 146500 72460 147130 72470
rect 146500 72450 146510 72460
rect 146690 72320 146810 72380
rect 146970 72320 147090 72380
rect 146690 72230 146700 72320
rect 146800 72290 146870 72320
rect 146810 72200 146870 72290
rect 146970 72230 146980 72320
rect 147090 72200 147150 72320
rect 146410 72150 147140 72160
rect 146460 72135 147150 72145
rect 36000 72110 37190 72120
rect 37100 72010 37190 72110
rect 37720 72090 37750 72120
rect 37840 72090 37870 72120
rect 146100 72090 146160 72120
rect 37600 72060 37660 72090
rect 37720 72060 37780 72090
rect 37840 72060 37900 72090
rect 146450 72085 146460 72135
rect 40060 72010 40120 72040
rect 41540 72010 41600 72040
rect 42360 72010 42420 72040
rect 43840 72010 43900 72040
rect 146690 72020 146810 72080
rect 146970 72020 147090 72080
rect 146810 72010 146870 72020
rect 36000 71980 37190 72010
rect 146570 72000 146650 72010
rect 146710 72000 146790 72010
rect 146810 72000 146930 72010
rect 146990 72000 147070 72010
rect 36040 71970 36120 71980
rect 36220 71970 36300 71980
rect 36400 71970 36480 71980
rect 36580 71970 36660 71980
rect 36760 71970 36840 71980
rect 36940 71970 37020 71980
rect 36120 71910 36130 71970
rect 36300 71910 36310 71970
rect 36480 71910 36490 71970
rect 36660 71910 36670 71970
rect 36840 71910 36850 71970
rect 37020 71910 37030 71970
rect 37100 71910 37190 71980
rect 37720 71970 37750 72000
rect 37840 71970 37870 72000
rect 146100 71970 146160 72000
rect 37600 71940 37660 71970
rect 37720 71940 37780 71970
rect 37840 71940 37900 71970
rect 146650 71920 146660 72000
rect 146790 71920 146800 72000
rect 36000 71880 37190 71910
rect 40060 71890 40120 71920
rect 41540 71890 41600 71920
rect 42360 71890 42420 71920
rect 43840 71890 43900 71920
rect 146810 71900 146870 72000
rect 146930 71920 146940 72000
rect 147070 71920 147080 72000
rect 147090 71900 147150 72020
rect 36040 71820 36120 71830
rect 36220 71820 36300 71830
rect 36400 71820 36480 71830
rect 36580 71820 36660 71830
rect 36760 71820 36840 71830
rect 36940 71820 37020 71830
rect 36120 71740 36130 71820
rect 36300 71740 36310 71820
rect 36480 71740 36490 71820
rect 36660 71740 36670 71820
rect 36840 71740 36850 71820
rect 37020 71740 37030 71820
rect 37100 71680 37190 71880
rect 37720 71850 37750 71880
rect 37840 71850 37870 71880
rect 146100 71850 146160 71880
rect 37600 71820 37660 71850
rect 37720 71820 37780 71850
rect 37840 71820 37900 71850
rect 40060 71770 40120 71800
rect 41540 71770 41600 71800
rect 42360 71770 42420 71800
rect 43840 71770 43900 71800
rect 37720 71730 37750 71760
rect 37840 71730 37870 71760
rect 146100 71730 146160 71760
rect 37600 71700 37660 71730
rect 37720 71700 37780 71730
rect 37840 71700 37900 71730
rect 36000 71650 37190 71680
rect 40060 71650 40120 71680
rect 41540 71650 41600 71680
rect 42360 71650 42420 71680
rect 43840 71650 43900 71680
rect 36120 71590 36130 71650
rect 36300 71590 36310 71650
rect 36480 71590 36490 71650
rect 36660 71590 36670 71650
rect 36840 71590 36850 71650
rect 37020 71590 37030 71650
rect 37100 71580 37190 71650
rect 37720 71610 37750 71640
rect 37840 71610 37870 71640
rect 146100 71610 146160 71640
rect 37600 71580 37660 71610
rect 37720 71580 37780 71610
rect 37840 71580 37900 71610
rect 36000 71550 37190 71580
rect 37100 71540 37190 71550
rect 36000 71530 37190 71540
rect 40060 71530 40120 71560
rect 41540 71530 41600 71560
rect 42360 71530 42420 71560
rect 43840 71530 43900 71560
rect 36040 71350 36120 71360
rect 36220 71350 36300 71360
rect 36400 71350 36480 71360
rect 36580 71350 36660 71360
rect 36760 71350 36840 71360
rect 36940 71350 37020 71360
rect 36120 71270 36130 71350
rect 36300 71270 36310 71350
rect 36480 71270 36490 71350
rect 36660 71270 36670 71350
rect 36840 71270 36850 71350
rect 37020 71270 37030 71350
rect 36040 71030 36120 71040
rect 36220 71030 36300 71040
rect 36400 71030 36480 71040
rect 36580 71030 36660 71040
rect 36760 71030 36840 71040
rect 36940 71030 37020 71040
rect 36120 70950 36130 71030
rect 36300 70950 36310 71030
rect 36480 70950 36490 71030
rect 36660 70950 36670 71030
rect 36840 70950 36850 71030
rect 37020 70950 37030 71030
rect 37100 70860 37190 71530
rect 37720 71490 37750 71520
rect 37840 71490 37870 71520
rect 146100 71490 146160 71520
rect 37600 71460 37660 71490
rect 37720 71460 37780 71490
rect 37840 71460 37900 71490
rect 146690 71440 146810 71500
rect 146970 71440 147090 71500
rect 40060 71410 40120 71440
rect 41540 71410 41600 71440
rect 42360 71410 42420 71440
rect 43840 71410 43900 71440
rect 146810 71430 146870 71440
rect 146570 71420 146650 71430
rect 146810 71420 146930 71430
rect 37720 71370 37750 71400
rect 37840 71370 37870 71400
rect 146100 71370 146160 71400
rect 37600 71340 37660 71370
rect 37720 71340 37780 71370
rect 37840 71340 37900 71370
rect 146650 71340 146660 71420
rect 146810 71320 146870 71420
rect 146930 71340 146940 71420
rect 147090 71320 147150 71440
rect 40060 71290 40120 71320
rect 41540 71290 41600 71320
rect 42360 71290 42420 71320
rect 43840 71290 43900 71320
rect 37720 71250 37750 71280
rect 37840 71250 37870 71280
rect 146100 71250 146160 71280
rect 146500 71270 147140 71280
rect 146460 71255 147150 71265
rect 37600 71220 37660 71250
rect 37720 71220 37780 71250
rect 37840 71220 37900 71250
rect 146450 71205 146460 71255
rect 40060 71170 40120 71200
rect 41540 71170 41600 71200
rect 42360 71170 42420 71200
rect 43840 71170 43900 71200
rect 37720 71130 37750 71160
rect 37840 71130 37870 71160
rect 146100 71130 146160 71160
rect 146690 71140 146810 71200
rect 146970 71140 147090 71200
rect 146810 71130 146870 71140
rect 37600 71100 37660 71130
rect 37720 71100 37780 71130
rect 37840 71100 37900 71130
rect 146570 71120 146650 71130
rect 146710 71120 146790 71130
rect 146810 71120 146930 71130
rect 146990 71120 147070 71130
rect 40060 71050 40120 71080
rect 41540 71050 41600 71080
rect 42360 71050 42420 71080
rect 43840 71050 43900 71080
rect 146650 71040 146660 71120
rect 146790 71040 146800 71120
rect 37720 71010 37750 71040
rect 37840 71010 37870 71040
rect 146100 71010 146160 71040
rect 146810 71020 146870 71120
rect 146930 71040 146940 71120
rect 147070 71040 147080 71120
rect 147090 71020 147150 71140
rect 37600 70980 37660 71010
rect 37720 70980 37780 71010
rect 37840 70980 37900 71010
rect 146510 70990 147130 71000
rect 40060 70930 40120 70960
rect 41540 70930 41600 70960
rect 42360 70930 42420 70960
rect 43840 70930 43900 70960
rect 37720 70890 37750 70920
rect 37840 70890 37870 70920
rect 146100 70890 146160 70920
rect 37600 70860 37660 70890
rect 37720 70860 37780 70890
rect 37840 70860 37900 70890
rect 146610 70860 146970 70920
rect 36000 70850 37190 70860
rect 37100 70750 37190 70850
rect 40060 70810 40120 70840
rect 41540 70810 41600 70840
rect 42360 70810 42420 70840
rect 43840 70810 43900 70840
rect 37720 70770 37750 70800
rect 37840 70770 37870 70800
rect 146100 70770 146160 70800
rect 36000 70720 37190 70750
rect 37600 70740 37660 70770
rect 37720 70740 37780 70770
rect 37840 70740 37900 70770
rect 146300 70730 146420 70790
rect 146420 70720 146480 70730
rect 36040 70710 36120 70720
rect 36220 70710 36300 70720
rect 36400 70710 36480 70720
rect 36580 70710 36660 70720
rect 36760 70710 36840 70720
rect 36940 70710 37020 70720
rect 36120 70650 36130 70710
rect 36300 70650 36310 70710
rect 36480 70650 36490 70710
rect 36660 70650 36670 70710
rect 36840 70650 36850 70710
rect 37020 70650 37030 70710
rect 37100 70650 37190 70720
rect 40060 70690 40120 70720
rect 41540 70690 41600 70720
rect 42360 70690 42420 70720
rect 43840 70690 43900 70720
rect 146420 70710 147050 70720
rect 146420 70705 146480 70710
rect 146420 70695 147090 70705
rect 37720 70650 37750 70680
rect 37840 70650 37870 70680
rect 146100 70650 146160 70680
rect 36000 70620 37190 70650
rect 37600 70620 37660 70650
rect 37720 70620 37780 70650
rect 37840 70620 37900 70650
rect 36040 70560 36120 70570
rect 36220 70560 36300 70570
rect 36400 70560 36480 70570
rect 36580 70560 36660 70570
rect 36760 70560 36840 70570
rect 36940 70560 37020 70570
rect 36120 70480 36130 70560
rect 36300 70480 36310 70560
rect 36480 70480 36490 70560
rect 36660 70480 36670 70560
rect 36840 70480 36850 70560
rect 37020 70480 37030 70560
rect 37100 70420 37190 70620
rect 146420 70610 146480 70695
rect 40060 70570 40120 70600
rect 41540 70570 41600 70600
rect 42360 70570 42420 70600
rect 43840 70570 43900 70600
rect 37720 70530 37750 70560
rect 37840 70530 37870 70560
rect 146100 70530 146160 70560
rect 37600 70500 37660 70530
rect 37720 70500 37780 70530
rect 37840 70500 37900 70530
rect 40060 70450 40120 70480
rect 41540 70450 41600 70480
rect 42360 70450 42420 70480
rect 43840 70450 43900 70480
rect 146300 70470 146420 70530
rect 146420 70445 146480 70470
rect 146530 70460 146540 70630
rect 146610 70600 146970 70660
rect 147090 70645 147100 70695
rect 146530 70450 147140 70460
rect 36000 70390 37190 70420
rect 37720 70410 37750 70440
rect 37840 70410 37870 70440
rect 146100 70410 146160 70440
rect 146420 70435 147090 70445
rect 36120 70330 36130 70390
rect 36300 70330 36310 70390
rect 36480 70330 36490 70390
rect 36660 70330 36670 70390
rect 36840 70330 36850 70390
rect 37020 70330 37030 70390
rect 37100 70320 37190 70390
rect 37600 70380 37660 70410
rect 37720 70380 37780 70410
rect 37840 70380 37900 70410
rect 40060 70330 40120 70360
rect 41540 70330 41600 70360
rect 42360 70330 42420 70360
rect 43840 70330 43900 70360
rect 146420 70350 146480 70435
rect 146610 70340 146970 70400
rect 147090 70385 147100 70435
rect 36000 70290 37190 70320
rect 37720 70290 37750 70320
rect 37840 70290 37870 70320
rect 146100 70290 146160 70320
rect 37100 70280 37190 70290
rect 36000 70270 37190 70280
rect 36040 70090 36120 70100
rect 36220 70090 36300 70100
rect 36400 70090 36480 70100
rect 36580 70090 36660 70100
rect 36760 70090 36840 70100
rect 36940 70090 37020 70100
rect 36120 70010 36130 70090
rect 36300 70010 36310 70090
rect 36480 70010 36490 70090
rect 36660 70010 36670 70090
rect 36840 70010 36850 70090
rect 37020 70010 37030 70090
rect 36040 69770 36120 69780
rect 36220 69770 36300 69780
rect 36400 69770 36480 69780
rect 36580 69770 36660 69780
rect 36760 69770 36840 69780
rect 36940 69770 37020 69780
rect 36120 69690 36130 69770
rect 36300 69690 36310 69770
rect 36480 69690 36490 69770
rect 36660 69690 36670 69770
rect 36840 69690 36850 69770
rect 37020 69690 37030 69770
rect 37100 69600 37190 70270
rect 37600 70260 37660 70290
rect 37720 70260 37780 70290
rect 37840 70260 37900 70290
rect 40060 70210 40120 70240
rect 41540 70210 41600 70240
rect 42360 70210 42420 70240
rect 43840 70210 43900 70240
rect 37720 70170 37750 70200
rect 37840 70170 37870 70200
rect 37600 70140 37660 70170
rect 37720 70140 37780 70170
rect 37840 70140 37900 70170
rect 40060 70090 40120 70120
rect 41540 70090 41600 70120
rect 42360 70090 42420 70120
rect 43840 70090 43900 70120
rect 37720 70050 37750 70080
rect 37840 70050 37870 70080
rect 146300 70210 146420 70270
rect 146420 70200 146480 70210
rect 146100 70170 146160 70200
rect 146420 70190 147050 70200
rect 146420 70185 146480 70190
rect 146420 70175 147090 70185
rect 146420 70090 146480 70175
rect 146100 70050 146160 70080
rect 37600 70020 37660 70050
rect 37720 70020 37780 70050
rect 37840 70020 37900 70050
rect 40060 69970 40120 70000
rect 41540 69970 41600 70000
rect 42360 69970 42420 70000
rect 43840 69970 43900 70000
rect 37720 69930 37750 69960
rect 37840 69930 37870 69960
rect 146100 69930 146160 69960
rect 146300 69950 146420 70010
rect 37600 69900 37660 69930
rect 37720 69900 37780 69930
rect 37840 69900 37900 69930
rect 146420 69925 146480 69950
rect 146530 69940 146540 70110
rect 146610 70080 146970 70140
rect 147090 70125 147100 70175
rect 146530 69930 147140 69940
rect 146420 69915 147090 69925
rect 40060 69850 40120 69880
rect 41540 69850 41600 69880
rect 42360 69850 42420 69880
rect 43840 69850 43900 69880
rect 37720 69810 37750 69840
rect 37840 69810 37870 69840
rect 146100 69810 146160 69840
rect 146420 69830 146480 69915
rect 146610 69820 146970 69880
rect 147090 69865 147100 69915
rect 37600 69780 37660 69810
rect 37720 69780 37780 69810
rect 37840 69780 37900 69810
rect 40060 69730 40120 69760
rect 41540 69730 41600 69760
rect 42360 69730 42420 69760
rect 43840 69730 43900 69760
rect 37720 69690 37750 69720
rect 37840 69690 37870 69720
rect 146100 69690 146160 69720
rect 37600 69660 37660 69690
rect 37720 69660 37780 69690
rect 37840 69660 37900 69690
rect 40060 69610 40120 69640
rect 41540 69610 41600 69640
rect 42360 69610 42420 69640
rect 43840 69610 43900 69640
rect 36000 69590 37190 69600
rect 37100 69490 37190 69590
rect 37720 69570 37750 69600
rect 37840 69570 37870 69600
rect 146100 69570 146160 69600
rect 37600 69540 37660 69570
rect 37720 69540 37780 69570
rect 37840 69540 37900 69570
rect 40060 69490 40120 69520
rect 41540 69490 41600 69520
rect 42360 69490 42420 69520
rect 43840 69490 43900 69520
rect 36000 69460 37190 69490
rect 36040 69450 36120 69460
rect 36220 69450 36300 69460
rect 36400 69450 36480 69460
rect 36580 69450 36660 69460
rect 36760 69450 36840 69460
rect 36940 69450 37020 69460
rect 36120 69390 36130 69450
rect 36300 69390 36310 69450
rect 36480 69390 36490 69450
rect 36660 69390 36670 69450
rect 36840 69390 36850 69450
rect 37020 69390 37030 69450
rect 37100 69390 37190 69460
rect 37720 69450 37750 69480
rect 37840 69450 37870 69480
rect 146100 69450 146160 69480
rect 37600 69420 37660 69450
rect 37720 69420 37780 69450
rect 37840 69420 37900 69450
rect 36000 69360 37190 69390
rect 40060 69370 40120 69400
rect 41540 69370 41600 69400
rect 42360 69370 42420 69400
rect 43840 69370 43900 69400
rect 36040 69300 36120 69310
rect 36220 69300 36300 69310
rect 36400 69300 36480 69310
rect 36580 69300 36660 69310
rect 36760 69300 36840 69310
rect 36940 69300 37020 69310
rect 36120 69220 36130 69300
rect 36300 69220 36310 69300
rect 36480 69220 36490 69300
rect 36660 69220 36670 69300
rect 36840 69220 36850 69300
rect 37020 69220 37030 69300
rect 37100 69160 37190 69360
rect 37720 69330 37750 69360
rect 37840 69330 37870 69360
rect 146100 69330 146160 69360
rect 37600 69300 37660 69330
rect 37720 69300 37780 69330
rect 37840 69300 37900 69330
rect 40060 69250 40120 69280
rect 41540 69250 41600 69280
rect 42360 69250 42420 69280
rect 43840 69250 43900 69280
rect 37720 69210 37750 69240
rect 37840 69210 37870 69240
rect 146100 69210 146160 69240
rect 37600 69180 37660 69210
rect 37720 69180 37780 69210
rect 37840 69180 37900 69210
rect 36000 69130 37190 69160
rect 40060 69130 40120 69160
rect 41540 69130 41600 69160
rect 42360 69130 42420 69160
rect 43840 69130 43900 69160
rect 36120 69070 36130 69130
rect 36300 69070 36310 69130
rect 36480 69070 36490 69130
rect 36660 69070 36670 69130
rect 36840 69070 36850 69130
rect 37020 69070 37030 69130
rect 37100 69060 37190 69130
rect 37720 69090 37750 69120
rect 37840 69090 37870 69120
rect 146100 69090 146160 69120
rect 37600 69060 37660 69090
rect 37720 69060 37780 69090
rect 37840 69060 37900 69090
rect 36000 69030 37190 69060
rect 37100 69020 37190 69030
rect 36000 69010 37190 69020
rect 40060 69010 40120 69040
rect 41540 69010 41600 69040
rect 42360 69010 42420 69040
rect 43840 69010 43900 69040
rect 36040 68830 36120 68840
rect 36220 68830 36300 68840
rect 36400 68830 36480 68840
rect 36580 68830 36660 68840
rect 36760 68830 36840 68840
rect 36940 68830 37020 68840
rect 36120 68750 36130 68830
rect 36300 68750 36310 68830
rect 36480 68750 36490 68830
rect 36660 68750 36670 68830
rect 36840 68750 36850 68830
rect 37020 68750 37030 68830
rect 36040 68510 36120 68520
rect 36220 68510 36300 68520
rect 36400 68510 36480 68520
rect 36580 68510 36660 68520
rect 36760 68510 36840 68520
rect 36940 68510 37020 68520
rect 36120 68430 36130 68510
rect 36300 68430 36310 68510
rect 36480 68430 36490 68510
rect 36660 68430 36670 68510
rect 36840 68430 36850 68510
rect 37020 68430 37030 68510
rect 37100 68340 37190 69010
rect 37720 68970 37750 69000
rect 37840 68970 37870 69000
rect 146100 68970 146160 69000
rect 37600 68940 37660 68970
rect 37720 68940 37780 68970
rect 37840 68940 37900 68970
rect 40060 68890 40120 68920
rect 41540 68890 41600 68920
rect 42360 68890 42420 68920
rect 43840 68890 43900 68920
rect 37720 68850 37750 68880
rect 37840 68850 37870 68880
rect 146100 68850 146160 68880
rect 37600 68820 37660 68850
rect 37720 68820 37780 68850
rect 37840 68820 37900 68850
rect 40060 68770 40120 68800
rect 41540 68770 41600 68800
rect 42360 68770 42420 68800
rect 43840 68770 43900 68800
rect 37720 68730 37750 68760
rect 37840 68730 37870 68760
rect 146100 68730 146160 68760
rect 37600 68700 37660 68730
rect 37720 68700 37780 68730
rect 37840 68700 37900 68730
rect 40060 68650 40120 68680
rect 41540 68650 41600 68680
rect 42360 68650 42420 68680
rect 43840 68650 43900 68680
rect 37720 68610 37750 68640
rect 37840 68610 37870 68640
rect 146100 68610 146160 68640
rect 37600 68580 37660 68610
rect 37720 68580 37780 68610
rect 37840 68580 37900 68610
rect 40060 68530 40120 68560
rect 41540 68530 41600 68560
rect 42360 68530 42420 68560
rect 43840 68530 43900 68560
rect 37720 68490 37750 68520
rect 37840 68490 37870 68520
rect 146100 68490 146160 68520
rect 37600 68460 37660 68490
rect 37720 68460 37780 68490
rect 37840 68460 37900 68490
rect 40060 68410 40120 68440
rect 41540 68410 41600 68440
rect 42360 68410 42420 68440
rect 43840 68410 43900 68440
rect 37720 68370 37750 68400
rect 37840 68370 37870 68400
rect 146100 68370 146160 68400
rect 37600 68340 37660 68370
rect 37720 68340 37780 68370
rect 37840 68340 37900 68370
rect 36000 68330 37190 68340
rect 37100 68230 37190 68330
rect 40060 68290 40120 68320
rect 41540 68290 41600 68320
rect 42360 68290 42420 68320
rect 43840 68290 43900 68320
rect 37720 68250 37750 68280
rect 37840 68250 37870 68280
rect 146100 68250 146160 68280
rect 36000 68200 37190 68230
rect 37600 68220 37660 68250
rect 37720 68220 37780 68250
rect 37840 68220 37900 68250
rect 40685 68210 40925 68240
rect 36040 68190 36120 68200
rect 36220 68190 36300 68200
rect 36400 68190 36480 68200
rect 36580 68190 36660 68200
rect 36760 68190 36840 68200
rect 36940 68190 37020 68200
rect 36120 68130 36130 68190
rect 36300 68130 36310 68190
rect 36480 68130 36490 68190
rect 36660 68130 36670 68190
rect 36840 68130 36850 68190
rect 37020 68130 37030 68190
rect 37100 68130 37190 68200
rect 40060 68170 40120 68200
rect 37720 68130 37750 68160
rect 37840 68130 37870 68160
rect 40685 68150 40715 68210
rect 40775 68150 40865 68210
rect 40895 68150 40925 68210
rect 41540 68170 41600 68200
rect 42360 68170 42420 68200
rect 43840 68170 43900 68200
rect 36000 68100 37190 68130
rect 37600 68100 37660 68130
rect 37720 68100 37780 68130
rect 37840 68100 37900 68130
rect 40685 68120 40925 68150
rect 146100 68130 146160 68160
rect 36040 68040 36120 68050
rect 36220 68040 36300 68050
rect 36400 68040 36480 68050
rect 36580 68040 36660 68050
rect 36760 68040 36840 68050
rect 36940 68040 37020 68050
rect 36120 67960 36130 68040
rect 36300 67960 36310 68040
rect 36480 67960 36490 68040
rect 36660 67960 36670 68040
rect 36840 67960 36850 68040
rect 37020 67960 37030 68040
rect 37100 67900 37190 68100
rect 40060 68050 40120 68080
rect 41540 68050 41600 68080
rect 42360 68050 42420 68080
rect 43840 68050 43900 68080
rect 37720 68010 37750 68040
rect 37840 68010 37870 68040
rect 146100 68010 146160 68040
rect 37600 67980 37660 68010
rect 37720 67980 37780 68010
rect 37840 67980 37900 68010
rect 40060 67930 40120 67960
rect 41540 67930 41600 67960
rect 42360 67930 42420 67960
rect 43840 67930 43900 67960
rect 36000 67870 37190 67900
rect 37720 67890 37750 67920
rect 37840 67890 37870 67920
rect 146100 67890 146160 67920
rect 36120 67810 36130 67870
rect 36300 67810 36310 67870
rect 36480 67810 36490 67870
rect 36660 67810 36670 67870
rect 36840 67810 36850 67870
rect 37020 67810 37030 67870
rect 37100 67800 37190 67870
rect 37600 67860 37660 67890
rect 37720 67860 37780 67890
rect 37840 67860 37900 67890
rect 40060 67810 40120 67840
rect 41540 67810 41600 67840
rect 42360 67810 42420 67840
rect 43840 67810 43900 67840
rect 36000 67770 37190 67800
rect 37720 67770 37750 67800
rect 37840 67770 37870 67800
rect 146100 67770 146160 67800
rect 37100 67760 37190 67770
rect 36000 67750 37190 67760
rect 36040 67570 36120 67580
rect 36220 67570 36300 67580
rect 36400 67570 36480 67580
rect 36580 67570 36660 67580
rect 36760 67570 36840 67580
rect 36940 67570 37020 67580
rect 36120 67490 36130 67570
rect 36300 67490 36310 67570
rect 36480 67490 36490 67570
rect 36660 67490 36670 67570
rect 36840 67490 36850 67570
rect 37020 67490 37030 67570
rect 36040 67250 36120 67260
rect 36220 67250 36300 67260
rect 36400 67250 36480 67260
rect 36580 67250 36660 67260
rect 36760 67250 36840 67260
rect 36940 67250 37020 67260
rect 36120 67170 36130 67250
rect 36300 67170 36310 67250
rect 36480 67170 36490 67250
rect 36660 67170 36670 67250
rect 36840 67170 36850 67250
rect 37020 67170 37030 67250
rect 37100 67080 37190 67750
rect 37600 67740 37660 67770
rect 37720 67740 37780 67770
rect 37840 67740 37900 67770
rect 40060 67690 40120 67720
rect 41540 67690 41600 67720
rect 42360 67690 42420 67720
rect 43840 67690 43900 67720
rect 37720 67650 37750 67680
rect 37840 67650 37870 67680
rect 146100 67650 146160 67680
rect 37600 67620 37660 67650
rect 37720 67620 37780 67650
rect 37840 67620 37900 67650
rect 40060 67570 40120 67600
rect 41540 67570 41600 67600
rect 42360 67570 42420 67600
rect 43840 67570 43900 67600
rect 37720 67530 37750 67560
rect 37840 67530 37870 67560
rect 146100 67530 146160 67560
rect 37600 67500 37660 67530
rect 37720 67500 37780 67530
rect 37840 67500 37900 67530
rect 40678 67504 40758 67514
rect 40838 67504 40918 67514
rect 40060 67450 40120 67480
rect 37720 67410 37750 67440
rect 37840 67410 37870 67440
rect 40758 67434 40768 67504
rect 40678 67424 40768 67434
rect 40838 67434 40848 67504
rect 40918 67434 40928 67504
rect 41540 67450 41600 67480
rect 42360 67450 42420 67480
rect 43840 67450 43900 67480
rect 40838 67424 40928 67434
rect 146100 67410 146160 67440
rect 37600 67380 37660 67410
rect 37720 67380 37780 67410
rect 37840 67380 37900 67410
rect 40060 67330 40120 67360
rect 40678 67344 40758 67354
rect 40838 67344 40918 67354
rect 37720 67290 37750 67320
rect 37840 67290 37870 67320
rect 37600 67260 37660 67290
rect 37720 67260 37780 67290
rect 37840 67260 37900 67290
rect 40758 67264 40768 67344
rect 40838 67264 40848 67344
rect 40918 67264 40928 67344
rect 41540 67330 41600 67360
rect 42360 67330 42420 67360
rect 43840 67330 43900 67360
rect 146100 67290 146160 67320
rect 40060 67210 40120 67240
rect 41540 67210 41600 67240
rect 42360 67210 42420 67240
rect 43840 67210 43900 67240
rect 37720 67170 37750 67200
rect 37840 67170 37870 67200
rect 146100 67170 146160 67200
rect 37600 67140 37660 67170
rect 37720 67140 37780 67170
rect 37840 67140 37900 67170
rect 40060 67090 40120 67120
rect 41540 67090 41600 67120
rect 42360 67090 42420 67120
rect 43840 67090 43900 67120
rect 36000 67070 37190 67080
rect 37100 66970 37190 67070
rect 37720 67050 37750 67080
rect 37840 67050 37870 67080
rect 146100 67050 146160 67080
rect 37600 67020 37660 67050
rect 37720 67020 37780 67050
rect 37840 67020 37900 67050
rect 40060 66970 40120 67000
rect 41540 66970 41600 67000
rect 42360 66970 42420 67000
rect 43840 66970 43900 67000
rect 36000 66940 37190 66970
rect 36040 66930 36120 66940
rect 36220 66930 36300 66940
rect 36400 66930 36480 66940
rect 36580 66930 36660 66940
rect 36760 66930 36840 66940
rect 36940 66930 37020 66940
rect 36120 66870 36130 66930
rect 36300 66870 36310 66930
rect 36480 66870 36490 66930
rect 36660 66870 36670 66930
rect 36840 66870 36850 66930
rect 37020 66870 37030 66930
rect 37100 66870 37190 66940
rect 37720 66930 37750 66960
rect 37840 66930 37870 66960
rect 146100 66930 146160 66960
rect 37600 66900 37660 66930
rect 37720 66900 37780 66930
rect 37840 66900 37900 66930
rect 36000 66840 37190 66870
rect 40060 66850 40120 66880
rect 41540 66850 41600 66880
rect 42360 66850 42420 66880
rect 43840 66850 43900 66880
rect 36040 66780 36120 66790
rect 36220 66780 36300 66790
rect 36400 66780 36480 66790
rect 36580 66780 36660 66790
rect 36760 66780 36840 66790
rect 36940 66780 37020 66790
rect 36120 66700 36130 66780
rect 36300 66700 36310 66780
rect 36480 66700 36490 66780
rect 36660 66700 36670 66780
rect 36840 66700 36850 66780
rect 37020 66700 37030 66780
rect 37100 66640 37190 66840
rect 37720 66810 37750 66840
rect 37840 66810 37870 66840
rect 146100 66810 146160 66840
rect 37600 66780 37660 66810
rect 37720 66780 37780 66810
rect 37840 66780 37900 66810
rect 40060 66730 40120 66760
rect 41540 66730 41600 66760
rect 42360 66730 42420 66760
rect 43840 66730 43900 66760
rect 37720 66690 37750 66720
rect 37840 66690 37870 66720
rect 146100 66690 146160 66720
rect 37600 66660 37660 66690
rect 37720 66660 37780 66690
rect 37840 66660 37900 66690
rect 36000 66610 37190 66640
rect 40060 66610 40120 66640
rect 41540 66610 41600 66640
rect 42360 66610 42420 66640
rect 43840 66610 43900 66640
rect 36120 66550 36130 66610
rect 36300 66550 36310 66610
rect 36480 66550 36490 66610
rect 36660 66550 36670 66610
rect 36840 66550 36850 66610
rect 37020 66550 37030 66610
rect 37100 66540 37190 66610
rect 37720 66570 37750 66600
rect 37840 66570 37870 66600
rect 146100 66570 146160 66600
rect 37600 66540 37660 66570
rect 37720 66540 37780 66570
rect 37840 66540 37900 66570
rect 36000 66510 37190 66540
rect 37100 66500 37190 66510
rect 36000 66490 37190 66500
rect 40060 66490 40120 66520
rect 41540 66490 41600 66520
rect 42360 66490 42420 66520
rect 43840 66490 43900 66520
rect 36040 66310 36120 66320
rect 36220 66310 36300 66320
rect 36400 66310 36480 66320
rect 36580 66310 36660 66320
rect 36760 66310 36840 66320
rect 36940 66310 37020 66320
rect 36120 66230 36130 66310
rect 36300 66230 36310 66310
rect 36480 66230 36490 66310
rect 36660 66230 36670 66310
rect 36840 66230 36850 66310
rect 37020 66230 37030 66310
rect 36040 65990 36120 66000
rect 36220 65990 36300 66000
rect 36400 65990 36480 66000
rect 36580 65990 36660 66000
rect 36760 65990 36840 66000
rect 36940 65990 37020 66000
rect 36120 65910 36130 65990
rect 36300 65910 36310 65990
rect 36480 65910 36490 65990
rect 36660 65910 36670 65990
rect 36840 65910 36850 65990
rect 37020 65910 37030 65990
rect 37100 65820 37190 66490
rect 37720 66450 37750 66480
rect 37840 66450 37870 66480
rect 42595 66475 42675 66485
rect 37600 66420 37660 66450
rect 37720 66420 37780 66450
rect 37840 66420 37900 66450
rect 42675 66405 42685 66475
rect 146100 66450 146160 66480
rect 40060 66370 40120 66400
rect 41540 66370 41600 66400
rect 42360 66370 42420 66400
rect 42595 66395 42685 66405
rect 43840 66370 43900 66400
rect 37720 66330 37750 66360
rect 37840 66330 37870 66360
rect 37600 66300 37660 66330
rect 37720 66300 37780 66330
rect 37840 66300 37900 66330
rect 42595 66315 42675 66325
rect 40060 66250 40120 66280
rect 41540 66250 41600 66280
rect 42360 66250 42420 66280
rect 37720 66210 37750 66240
rect 37840 66210 37870 66240
rect 42675 66235 42685 66315
rect 43030 66300 43390 66360
rect 43840 66250 43900 66280
rect 38595 66215 38675 66225
rect 38775 66215 38855 66225
rect 38955 66215 39035 66225
rect 39135 66215 39215 66225
rect 39315 66215 39395 66225
rect 37600 66180 37660 66210
rect 37720 66180 37780 66210
rect 37840 66180 37900 66210
rect 38675 66135 38685 66215
rect 38855 66135 38865 66215
rect 39035 66135 39045 66215
rect 39215 66135 39225 66215
rect 39395 66135 39405 66215
rect 43580 66170 43700 66230
rect 40060 66130 40120 66160
rect 41540 66130 41600 66160
rect 42360 66130 42420 66160
rect 42950 66150 43560 66160
rect 43550 66145 43560 66150
rect 42910 66135 43560 66145
rect 37720 66090 37750 66120
rect 37840 66090 37870 66120
rect 37600 66060 37660 66090
rect 37720 66060 37780 66090
rect 37840 66060 37900 66090
rect 42900 66085 42910 66135
rect 38595 66035 38675 66045
rect 38775 66035 38855 66045
rect 38955 66035 39035 66045
rect 39135 66035 39215 66045
rect 39315 66035 39395 66045
rect 43030 66040 43390 66100
rect 37720 65970 37750 66000
rect 37840 65970 37870 66000
rect 37600 65940 37660 65970
rect 37720 65940 37780 65970
rect 37840 65940 37900 65970
rect 38675 65955 38685 66035
rect 38855 65955 38865 66035
rect 39035 65955 39045 66035
rect 39215 65955 39225 66035
rect 39395 65955 39405 66035
rect 40060 66010 40120 66040
rect 41540 66010 41600 66040
rect 42360 66010 42420 66040
rect 42682 65960 42822 66030
rect 40060 65890 40120 65920
rect 40678 65899 40758 65909
rect 40838 65899 40918 65909
rect 37720 65850 37750 65880
rect 37840 65850 37870 65880
rect 38595 65855 38675 65865
rect 38775 65855 38855 65865
rect 38955 65855 39035 65865
rect 39135 65855 39215 65865
rect 39315 65855 39395 65865
rect 37600 65820 37660 65850
rect 37720 65820 37780 65850
rect 37840 65820 37900 65850
rect 36000 65810 37190 65820
rect 37100 65710 37190 65810
rect 38675 65775 38685 65855
rect 38855 65775 38865 65855
rect 39035 65775 39045 65855
rect 39215 65775 39225 65855
rect 39395 65775 39405 65855
rect 40758 65819 40768 65899
rect 40838 65819 40848 65899
rect 40918 65819 40928 65899
rect 41540 65890 41600 65920
rect 42360 65890 42420 65920
rect 42822 65900 42892 65960
rect 42822 65890 43470 65900
rect 43550 65890 43560 66135
rect 43700 66050 43760 66170
rect 146100 66330 146160 66360
rect 146100 66210 146160 66240
rect 43840 66130 43900 66160
rect 146100 66090 146160 66120
rect 43840 66010 43900 66040
rect 146100 65970 146160 66000
rect 43580 65910 43700 65970
rect 42822 65820 42892 65890
rect 42910 65875 43560 65885
rect 42900 65825 42910 65875
rect 40060 65770 40120 65800
rect 37720 65730 37750 65760
rect 37840 65730 37870 65760
rect 40685 65750 40925 65780
rect 41540 65770 41600 65800
rect 42360 65770 42420 65800
rect 42682 65760 42822 65820
rect 43030 65780 43390 65840
rect 43700 65790 43760 65910
rect 43840 65890 43900 65920
rect 146100 65850 146160 65880
rect 43840 65770 43900 65800
rect 36000 65680 37190 65710
rect 37600 65700 37660 65730
rect 37720 65700 37780 65730
rect 37840 65700 37900 65730
rect 40685 65690 40715 65750
rect 40775 65690 40865 65750
rect 40895 65690 40925 65750
rect 36040 65670 36120 65680
rect 36220 65670 36300 65680
rect 36400 65670 36480 65680
rect 36580 65670 36660 65680
rect 36760 65670 36840 65680
rect 36940 65670 37020 65680
rect 36120 65610 36130 65670
rect 36300 65610 36310 65670
rect 36480 65610 36490 65670
rect 36660 65610 36670 65670
rect 36840 65610 36850 65670
rect 37020 65610 37030 65670
rect 37100 65610 37190 65680
rect 38595 65675 38675 65685
rect 38775 65675 38855 65685
rect 38955 65675 39035 65685
rect 39135 65675 39215 65685
rect 39315 65675 39395 65685
rect 37720 65610 37750 65640
rect 37840 65610 37870 65640
rect 36000 65580 37190 65610
rect 37600 65580 37660 65610
rect 37720 65580 37780 65610
rect 37840 65580 37900 65610
rect 38675 65595 38685 65675
rect 38855 65595 38865 65675
rect 39035 65595 39045 65675
rect 39215 65595 39225 65675
rect 39395 65595 39405 65675
rect 40060 65650 40120 65680
rect 40685 65660 40925 65690
rect 41540 65650 41600 65680
rect 42360 65650 42420 65680
rect 40678 65629 40758 65639
rect 40838 65629 40918 65639
rect 36040 65520 36120 65530
rect 36220 65520 36300 65530
rect 36400 65520 36480 65530
rect 36580 65520 36660 65530
rect 36760 65520 36840 65530
rect 36940 65520 37020 65530
rect 36120 65440 36130 65520
rect 36300 65440 36310 65520
rect 36480 65440 36490 65520
rect 36660 65440 36670 65520
rect 36840 65440 36850 65520
rect 37020 65440 37030 65520
rect 37100 65380 37190 65580
rect 40060 65530 40120 65560
rect 40758 65549 40768 65629
rect 40838 65549 40848 65629
rect 40918 65549 40928 65629
rect 42822 65620 42892 65760
rect 146100 65730 146160 65760
rect 43580 65650 43700 65710
rect 43840 65650 43900 65680
rect 42950 65630 43560 65640
rect 43550 65625 43560 65630
rect 42682 65560 42822 65620
rect 42910 65615 43560 65625
rect 42900 65565 42910 65615
rect 41540 65530 41600 65560
rect 42360 65530 42420 65560
rect 37720 65490 37750 65520
rect 37840 65490 37870 65520
rect 38595 65495 38675 65505
rect 38775 65495 38855 65505
rect 38955 65495 39035 65505
rect 39135 65495 39215 65505
rect 39315 65495 39395 65505
rect 37600 65460 37660 65490
rect 37720 65460 37780 65490
rect 37840 65460 37900 65490
rect 38675 65415 38685 65495
rect 38855 65415 38865 65495
rect 39035 65415 39045 65495
rect 39215 65415 39225 65495
rect 39395 65415 39405 65495
rect 40060 65410 40120 65440
rect 41540 65410 41600 65440
rect 42360 65410 42420 65440
rect 42822 65420 42892 65560
rect 43030 65520 43390 65580
rect 36000 65350 37190 65380
rect 37720 65370 37750 65400
rect 37840 65370 37870 65400
rect 36120 65290 36130 65350
rect 36300 65290 36310 65350
rect 36480 65290 36490 65350
rect 36660 65290 36670 65350
rect 36840 65290 36850 65350
rect 37020 65290 37030 65350
rect 37100 65280 37190 65350
rect 37600 65340 37660 65370
rect 37720 65340 37780 65370
rect 37840 65340 37900 65370
rect 40170 65320 40180 65410
rect 40060 65290 40120 65320
rect 36000 65250 37190 65280
rect 37720 65250 37750 65280
rect 37840 65250 37870 65280
rect 37100 65240 37190 65250
rect 36000 65230 37190 65240
rect 36040 65050 36120 65060
rect 36220 65050 36300 65060
rect 36400 65050 36480 65060
rect 36580 65050 36660 65060
rect 36760 65050 36840 65060
rect 36940 65050 37020 65060
rect 36120 64970 36130 65050
rect 36300 64970 36310 65050
rect 36480 64970 36490 65050
rect 36660 64970 36670 65050
rect 36840 64970 36850 65050
rect 37020 64970 37030 65050
rect 36040 64730 36120 64740
rect 36220 64730 36300 64740
rect 36400 64730 36480 64740
rect 36580 64730 36660 64740
rect 36760 64730 36840 64740
rect 36940 64730 37020 64740
rect 36120 64650 36130 64730
rect 36300 64650 36310 64730
rect 36480 64650 36490 64730
rect 36660 64650 36670 64730
rect 36840 64650 36850 64730
rect 37020 64650 37030 64730
rect 37100 64560 37190 65230
rect 37600 65220 37660 65250
rect 37720 65220 37780 65250
rect 37840 65220 37900 65250
rect 40060 65170 40120 65200
rect 37720 65130 37750 65160
rect 37840 65130 37870 65160
rect 37600 65100 37660 65130
rect 37720 65100 37780 65130
rect 37840 65100 37900 65130
rect 40060 65050 40120 65080
rect 37720 65010 37750 65040
rect 37840 65010 37870 65040
rect 37600 64980 37660 65010
rect 37720 64980 37780 65010
rect 37840 64980 37900 65010
rect 40060 64930 40120 64960
rect 37720 64890 37750 64920
rect 37840 64890 37870 64920
rect 37600 64860 37660 64890
rect 37720 64860 37780 64890
rect 37840 64860 37900 64890
rect 40060 64810 40120 64840
rect 37720 64770 37750 64800
rect 37840 64770 37870 64800
rect 37600 64740 37660 64770
rect 37720 64740 37780 64770
rect 37840 64740 37900 64770
rect 40060 64690 40120 64720
rect 37720 64650 37750 64680
rect 37840 64650 37870 64680
rect 37600 64620 37660 64650
rect 37720 64620 37780 64650
rect 37840 64620 37900 64650
rect 40060 64570 40120 64600
rect 36000 64550 37190 64560
rect 37100 64450 37190 64550
rect 37720 64530 37750 64560
rect 37840 64530 37870 64560
rect 40260 64530 40270 65320
rect 40380 65310 41180 65400
rect 40650 65280 40770 65310
rect 40930 65280 41050 65310
rect 41090 65280 41180 65310
rect 40650 65190 40660 65280
rect 40760 65250 40830 65280
rect 40770 65160 40830 65250
rect 40930 65190 40940 65280
rect 41050 65160 41180 65280
rect 41260 65240 41340 65250
rect 41340 65190 41350 65240
rect 41090 65125 41180 65160
rect 41230 65130 41350 65190
rect 40470 65120 41180 65125
rect 40370 65110 41180 65120
rect 40370 65030 40380 65110
rect 40470 65105 41180 65110
rect 40420 65095 41210 65105
rect 41090 65045 41180 65095
rect 40470 65030 41180 65045
rect 40460 65015 41180 65030
rect 40460 64825 40470 65015
rect 40650 64980 40770 65015
rect 40930 64980 41050 65015
rect 41090 64980 41180 65015
rect 41350 65010 41410 65130
rect 40770 64970 40830 64980
rect 40530 64960 40610 64970
rect 40670 64960 40750 64970
rect 40770 64960 40890 64970
rect 40950 64960 41030 64970
rect 40610 64880 40620 64960
rect 40750 64880 40760 64960
rect 40770 64860 40830 64960
rect 40890 64880 40900 64960
rect 41030 64880 41040 64960
rect 41050 64860 41180 64980
rect 41260 64960 41340 64970
rect 41340 64890 41350 64960
rect 41090 64825 41180 64860
rect 41230 64830 41350 64890
rect 40460 64810 41180 64825
rect 40470 64805 41180 64810
rect 40420 64795 41210 64805
rect 41090 64745 41180 64795
rect 40470 64715 41180 64745
rect 40650 64680 40770 64715
rect 40930 64680 41050 64715
rect 41090 64680 41180 64715
rect 41350 64710 41410 64830
rect 41480 64680 41490 65390
rect 42860 65370 43470 65380
rect 43550 65370 43560 65615
rect 43700 65530 43760 65650
rect 146100 65610 146160 65640
rect 43840 65530 43900 65560
rect 146100 65490 146160 65520
rect 43580 65390 43700 65450
rect 43840 65410 43900 65440
rect 42910 65355 43560 65365
rect 41540 65290 41600 65320
rect 42360 65290 42420 65320
rect 42900 65305 42910 65355
rect 43030 65260 43390 65320
rect 43700 65270 43760 65390
rect 146100 65370 146160 65400
rect 43840 65290 43900 65320
rect 146100 65250 146160 65280
rect 41540 65170 41600 65200
rect 42360 65170 42420 65200
rect 42470 65160 42480 65250
rect 43840 65170 43900 65200
rect 41540 65050 41600 65080
rect 42360 65050 42420 65080
rect 41540 64930 41600 64960
rect 42360 64930 42420 64960
rect 41540 64810 41600 64840
rect 42360 64810 42420 64840
rect 41540 64690 41600 64720
rect 42360 64690 42420 64720
rect 42560 64680 42570 65160
rect 146100 65130 146160 65160
rect 42960 65120 43460 65130
rect 42620 65100 42700 65110
rect 42700 65030 42710 65100
rect 42620 65020 42710 65030
rect 42770 65020 42780 65110
rect 43840 65050 43900 65080
rect 42620 64940 42700 64950
rect 42700 64890 42710 64940
rect 42610 64830 42730 64890
rect 42730 64805 42790 64830
rect 42860 64820 42870 65020
rect 42910 64980 43030 65040
rect 43190 64980 43310 65040
rect 146100 65010 146160 65040
rect 43030 64970 43090 64980
rect 43310 64970 43370 64980
rect 42930 64960 43010 64970
rect 43030 64960 43150 64970
rect 43210 64960 43290 64970
rect 43310 64960 43430 64970
rect 43010 64880 43020 64960
rect 43030 64860 43090 64960
rect 43150 64880 43160 64960
rect 43290 64880 43300 64960
rect 43310 64860 43370 64960
rect 43430 64880 43440 64960
rect 43840 64930 43900 64960
rect 146100 64890 146160 64920
rect 42860 64810 43500 64820
rect 43840 64810 43900 64840
rect 42730 64795 43540 64805
rect 42730 64710 42790 64795
rect 43540 64745 43550 64795
rect 146100 64770 146160 64800
rect 42860 64680 42870 64730
rect 42910 64680 43030 64740
rect 43190 64680 43310 64740
rect 43840 64690 43900 64720
rect 40770 64670 40830 64680
rect 40530 64660 40610 64670
rect 40770 64660 40890 64670
rect 40610 64580 40620 64660
rect 40770 64560 40830 64660
rect 40890 64580 40900 64660
rect 41050 64560 41180 64680
rect 43030 64670 43090 64680
rect 43310 64670 43370 64680
rect 43030 64660 43150 64670
rect 43310 64660 43430 64670
rect 41540 64570 41600 64600
rect 42360 64570 42420 64600
rect 43030 64560 43090 64660
rect 43150 64580 43160 64660
rect 43310 64560 43370 64660
rect 43430 64580 43440 64660
rect 146100 64650 146160 64680
rect 43840 64570 43900 64600
rect 41090 64550 41180 64560
rect 40470 64530 41180 64550
rect 146100 64530 146160 64560
rect 37600 64500 37660 64530
rect 37720 64500 37780 64530
rect 37840 64500 37900 64530
rect 40060 64450 40120 64480
rect 36000 64420 37190 64450
rect 40170 64440 40180 64530
rect 40260 64520 41100 64530
rect 36040 64410 36120 64420
rect 36220 64410 36300 64420
rect 36400 64410 36480 64420
rect 36580 64410 36660 64420
rect 36760 64410 36840 64420
rect 36940 64410 37020 64420
rect 36120 64350 36130 64410
rect 36300 64350 36310 64410
rect 36480 64350 36490 64410
rect 36660 64350 36670 64410
rect 36840 64350 36850 64410
rect 37020 64350 37030 64410
rect 37100 64350 37190 64420
rect 37720 64410 37750 64440
rect 37840 64410 37870 64440
rect 37600 64380 37660 64410
rect 37720 64380 37780 64410
rect 37840 64380 37900 64410
rect 36000 64320 37190 64350
rect 40060 64330 40120 64360
rect 36040 64260 36120 64270
rect 36220 64260 36300 64270
rect 36400 64260 36480 64270
rect 36580 64260 36660 64270
rect 36760 64260 36840 64270
rect 36940 64260 37020 64270
rect 36120 64180 36130 64260
rect 36300 64180 36310 64260
rect 36480 64180 36490 64260
rect 36660 64180 36670 64260
rect 36840 64180 36850 64260
rect 37020 64180 37030 64260
rect 37100 64120 37190 64320
rect 37720 64290 37750 64320
rect 37840 64290 37870 64320
rect 37600 64260 37660 64290
rect 37720 64260 37780 64290
rect 37840 64260 37900 64290
rect 40060 64210 40120 64240
rect 37720 64170 37750 64200
rect 37840 64170 37870 64200
rect 37600 64140 37660 64170
rect 37720 64140 37780 64170
rect 37840 64140 37900 64170
rect 36000 64090 37190 64120
rect 40060 64090 40120 64120
rect 36120 64030 36130 64090
rect 36300 64030 36310 64090
rect 36480 64030 36490 64090
rect 36660 64030 36670 64090
rect 36840 64030 36850 64090
rect 37020 64030 37030 64090
rect 37100 64020 37190 64090
rect 37720 64050 37750 64080
rect 37840 64050 37870 64080
rect 37600 64020 37660 64050
rect 37720 64020 37780 64050
rect 37840 64020 37900 64050
rect 36000 63990 37190 64020
rect 37100 63980 37190 63990
rect 36000 63970 37190 63980
rect 40060 63970 40120 64000
rect 36040 63790 36120 63800
rect 36220 63790 36300 63800
rect 36400 63790 36480 63800
rect 36580 63790 36660 63800
rect 36760 63790 36840 63800
rect 36940 63790 37020 63800
rect 36120 63710 36130 63790
rect 36300 63710 36310 63790
rect 36480 63710 36490 63790
rect 36660 63710 36670 63790
rect 36840 63710 36850 63790
rect 37020 63710 37030 63790
rect 36040 63470 36120 63480
rect 36220 63470 36300 63480
rect 36400 63470 36480 63480
rect 36580 63470 36660 63480
rect 36760 63470 36840 63480
rect 36940 63470 37020 63480
rect 36120 63390 36130 63470
rect 36300 63390 36310 63470
rect 36480 63390 36490 63470
rect 36660 63390 36670 63470
rect 36840 63390 36850 63470
rect 37020 63390 37030 63470
rect 37100 63300 37190 63970
rect 37720 63930 37750 63960
rect 37840 63930 37870 63960
rect 37600 63900 37660 63930
rect 37720 63900 37780 63930
rect 37840 63900 37900 63930
rect 40060 63850 40120 63880
rect 37720 63810 37750 63840
rect 37840 63810 37870 63840
rect 37600 63780 37660 63810
rect 37720 63780 37780 63810
rect 37840 63780 37900 63810
rect 40060 63730 40120 63760
rect 37720 63690 37750 63720
rect 37840 63690 37870 63720
rect 37600 63660 37660 63690
rect 37720 63660 37780 63690
rect 37840 63660 37900 63690
rect 40060 63610 40120 63640
rect 37720 63570 37750 63600
rect 37840 63570 37870 63600
rect 37600 63540 37660 63570
rect 37720 63540 37780 63570
rect 37840 63540 37900 63570
rect 40060 63490 40120 63520
rect 37720 63450 37750 63480
rect 37840 63450 37870 63480
rect 37600 63420 37660 63450
rect 37720 63420 37780 63450
rect 37840 63420 37900 63450
rect 40060 63370 40120 63400
rect 37720 63330 37750 63360
rect 37840 63330 37870 63360
rect 37600 63300 37660 63330
rect 37720 63300 37780 63330
rect 37840 63300 37900 63330
rect 36000 63290 37190 63300
rect 37100 63190 37190 63290
rect 40060 63250 40120 63280
rect 37720 63210 37750 63240
rect 37840 63210 37870 63240
rect 36000 63160 37190 63190
rect 37600 63180 37660 63210
rect 37720 63180 37780 63210
rect 37840 63180 37900 63210
rect 36040 63150 36120 63160
rect 36220 63150 36300 63160
rect 36400 63150 36480 63160
rect 36580 63150 36660 63160
rect 36760 63150 36840 63160
rect 36940 63150 37020 63160
rect 36120 63090 36130 63150
rect 36300 63090 36310 63150
rect 36480 63090 36490 63150
rect 36660 63090 36670 63150
rect 36840 63090 36850 63150
rect 37020 63090 37030 63150
rect 37100 63090 37190 63160
rect 40060 63130 40120 63160
rect 37720 63090 37750 63120
rect 37840 63090 37870 63120
rect 36000 63060 37190 63090
rect 37600 63060 37660 63090
rect 37720 63060 37780 63090
rect 37840 63060 37900 63090
rect 36040 63000 36120 63010
rect 36220 63000 36300 63010
rect 36400 63000 36480 63010
rect 36580 63000 36660 63010
rect 36760 63000 36840 63010
rect 36940 63000 37020 63010
rect 36120 62920 36130 63000
rect 36300 62920 36310 63000
rect 36480 62920 36490 63000
rect 36660 62920 36670 63000
rect 36840 62920 36850 63000
rect 37020 62920 37030 63000
rect 36040 62850 36120 62860
rect 36220 62850 36300 62860
rect 36400 62850 36480 62860
rect 36580 62850 36660 62860
rect 36760 62850 36840 62860
rect 36940 62850 37020 62860
rect 36120 62770 36130 62850
rect 36300 62770 36310 62850
rect 36480 62770 36490 62850
rect 36660 62770 36670 62850
rect 36840 62770 36850 62850
rect 37020 62770 37030 62850
rect 37100 62830 37190 63060
rect 40060 63010 40120 63040
rect 37720 62970 37750 63000
rect 37840 62970 37870 63000
rect 37600 62940 37660 62970
rect 37720 62940 37780 62970
rect 37840 62940 37900 62970
rect 40060 62890 40120 62920
rect 37720 62850 37750 62880
rect 37840 62850 37870 62880
rect 37600 62820 37660 62850
rect 37720 62820 37780 62850
rect 37840 62820 37900 62850
rect 40060 62770 40120 62800
rect 19130 62700 19160 62755
rect 19250 62700 19280 62755
rect 26420 62700 26450 62755
rect 26540 62700 26570 62755
rect 30420 62730 30450 62755
rect 30540 62730 30570 62755
rect 37720 62730 37750 62760
rect 37840 62730 37870 62760
rect 30300 62700 30360 62730
rect 30420 62700 30480 62730
rect 30540 62700 30600 62730
rect 37600 62700 37660 62730
rect 37720 62700 37780 62730
rect 37840 62700 37900 62730
rect 40060 62650 40120 62680
rect 30420 62580 30450 62640
rect 30540 62580 30570 62640
rect 37720 62580 37750 62640
rect 37840 62580 37870 62640
rect 40060 62530 40120 62560
rect 18980 62440 19060 62450
rect 19160 62440 19240 62450
rect 19340 62440 19420 62450
rect 19520 62440 19600 62450
rect 19700 62440 19780 62450
rect 19880 62440 19960 62450
rect 20060 62440 20140 62450
rect 20240 62440 20320 62450
rect 20420 62440 20500 62450
rect 20600 62440 20680 62450
rect 20780 62440 20860 62450
rect 20960 62440 21040 62450
rect 21140 62440 21220 62450
rect 21320 62440 21400 62450
rect 21500 62440 21580 62450
rect 21680 62440 21760 62450
rect 21860 62440 21940 62450
rect 22040 62440 22120 62450
rect 22220 62440 22300 62450
rect 22400 62440 22480 62450
rect 22580 62440 22660 62450
rect 22760 62440 22840 62450
rect 22940 62440 23020 62450
rect 23120 62440 23200 62450
rect 23300 62440 23380 62450
rect 23480 62440 23560 62450
rect 23660 62440 23740 62450
rect 23840 62440 23920 62450
rect 24020 62440 24100 62450
rect 24200 62440 24280 62450
rect 24380 62440 24460 62450
rect 24560 62440 24640 62450
rect 24740 62440 24820 62450
rect 24920 62440 25000 62450
rect 25100 62440 25180 62450
rect 25280 62440 25360 62450
rect 25460 62440 25540 62450
rect 25640 62440 25720 62450
rect 25820 62440 25900 62450
rect 26000 62440 26080 62450
rect 26180 62440 26260 62450
rect 26360 62440 26440 62450
rect 26540 62440 26620 62450
rect 30280 62440 30360 62450
rect 30460 62440 30540 62450
rect 30640 62440 30720 62450
rect 30820 62440 30900 62450
rect 31000 62440 31080 62450
rect 31180 62440 31260 62450
rect 31360 62440 31440 62450
rect 31540 62440 31620 62450
rect 31720 62440 31800 62450
rect 31900 62440 31980 62450
rect 32080 62440 32160 62450
rect 32260 62440 32340 62450
rect 32440 62440 32520 62450
rect 32620 62440 32700 62450
rect 32800 62440 32880 62450
rect 32980 62440 33060 62450
rect 33160 62440 33240 62450
rect 33340 62440 33420 62450
rect 33520 62440 33600 62450
rect 33700 62440 33780 62450
rect 33880 62440 33960 62450
rect 34060 62440 34140 62450
rect 34240 62440 34320 62450
rect 34420 62440 34500 62450
rect 34600 62440 34680 62450
rect 34780 62440 34860 62450
rect 34960 62440 35040 62450
rect 35140 62440 35220 62450
rect 35320 62440 35400 62450
rect 35500 62440 35580 62450
rect 35680 62440 35760 62450
rect 35860 62440 35940 62450
rect 36040 62440 36120 62450
rect 36220 62440 36300 62450
rect 36400 62440 36480 62450
rect 36580 62440 36660 62450
rect 36760 62440 36840 62450
rect 36940 62440 37020 62450
rect 37120 62440 37200 62450
rect 37300 62440 37380 62450
rect 37480 62440 37560 62450
rect 37660 62440 37740 62450
rect 37840 62440 37920 62450
rect 40260 62440 40270 64440
rect 40380 64430 41180 64520
rect 41540 64450 41600 64480
rect 42360 64450 42420 64480
rect 43840 64450 43900 64480
rect 40650 64400 40770 64430
rect 40930 64400 41050 64430
rect 41090 64400 41180 64430
rect 146100 64410 146160 64440
rect 40650 64310 40660 64400
rect 40760 64370 40830 64400
rect 40770 64280 40830 64370
rect 40930 64310 40940 64400
rect 41050 64280 41180 64400
rect 41090 64245 41180 64280
rect 41230 64250 41350 64310
rect 40470 64240 41180 64245
rect 40370 64230 41180 64240
rect 40370 64150 40380 64230
rect 40470 64225 41180 64230
rect 40420 64215 41210 64225
rect 41090 64165 41180 64215
rect 40470 64150 41180 64165
rect 40460 64135 41180 64150
rect 40460 63945 40470 64135
rect 40650 64100 40770 64135
rect 40930 64100 41050 64135
rect 41090 64100 41180 64135
rect 41350 64130 41410 64250
rect 40770 64090 40830 64100
rect 40530 64080 40610 64090
rect 40670 64080 40750 64090
rect 40770 64080 40890 64090
rect 40950 64080 41030 64090
rect 40610 64000 40620 64080
rect 40750 64000 40760 64080
rect 40770 63980 40830 64080
rect 40890 64000 40900 64080
rect 41030 64000 41040 64080
rect 41050 63980 41180 64100
rect 41260 64080 41340 64090
rect 41340 64010 41350 64080
rect 41090 63945 41180 63980
rect 41230 63950 41350 64010
rect 40460 63930 41180 63945
rect 40470 63925 41180 63930
rect 40420 63915 41210 63925
rect 41090 63865 41180 63915
rect 40470 63835 41180 63865
rect 40650 63800 40770 63835
rect 40930 63800 41050 63835
rect 41090 63800 41180 63835
rect 41350 63830 41410 63950
rect 40650 63710 40660 63800
rect 40760 63770 40830 63800
rect 40770 63680 40830 63770
rect 40930 63710 40940 63800
rect 41050 63680 41180 63800
rect 41260 63780 41340 63790
rect 41340 63710 41350 63780
rect 41090 63645 41180 63680
rect 41230 63650 41350 63710
rect 40370 63630 40460 63640
rect 40370 63550 40380 63630
rect 40470 63625 41180 63645
rect 40420 63615 41210 63625
rect 41090 63565 41180 63615
rect 40470 63550 41180 63565
rect 40460 63535 41180 63550
rect 40460 63345 40470 63535
rect 40650 63500 40770 63535
rect 40930 63500 41050 63535
rect 41090 63500 41180 63535
rect 41350 63530 41410 63650
rect 40770 63490 40830 63500
rect 40530 63480 40610 63490
rect 40670 63480 40750 63490
rect 40770 63480 40890 63490
rect 40950 63480 41030 63490
rect 40610 63400 40620 63480
rect 40750 63400 40760 63480
rect 40770 63380 40830 63480
rect 40890 63400 40900 63480
rect 41030 63400 41040 63480
rect 41050 63380 41180 63500
rect 41260 63480 41340 63490
rect 41340 63410 41350 63480
rect 41090 63345 41180 63380
rect 41230 63350 41350 63410
rect 40460 63330 41180 63345
rect 40470 63325 41180 63330
rect 40420 63315 41210 63325
rect 41090 63265 41180 63315
rect 40470 63235 41180 63265
rect 40650 63200 40770 63235
rect 40930 63200 41050 63235
rect 41090 63200 41180 63235
rect 41350 63230 41410 63350
rect 40650 63110 40660 63200
rect 40760 63170 40830 63200
rect 40770 63080 40830 63170
rect 40930 63110 40940 63200
rect 41050 63080 41180 63200
rect 41260 63180 41340 63190
rect 41340 63110 41350 63180
rect 41090 63045 41180 63080
rect 41230 63050 41350 63110
rect 40370 63030 40460 63040
rect 40370 62950 40380 63030
rect 40470 63025 41180 63045
rect 40420 63015 41210 63025
rect 41090 62965 41180 63015
rect 40470 62950 41180 62965
rect 40460 62935 41180 62950
rect 40460 62745 40470 62935
rect 40650 62900 40770 62935
rect 40930 62900 41050 62935
rect 41090 62900 41180 62935
rect 41350 62930 41410 63050
rect 40770 62890 40830 62900
rect 40530 62880 40610 62890
rect 40670 62880 40750 62890
rect 40770 62880 40890 62890
rect 40950 62880 41030 62890
rect 40610 62800 40620 62880
rect 40750 62800 40760 62880
rect 40770 62780 40830 62880
rect 40890 62800 40900 62880
rect 41030 62800 41040 62880
rect 41050 62780 41180 62900
rect 41260 62870 41340 62880
rect 41340 62810 41350 62870
rect 41090 62745 41180 62780
rect 41230 62750 41350 62810
rect 40460 62730 41180 62745
rect 40470 62725 41180 62730
rect 40420 62715 41210 62725
rect 41090 62665 41180 62715
rect 40470 62635 41180 62665
rect 40650 62600 40770 62635
rect 40930 62600 41050 62635
rect 41090 62600 41180 62635
rect 41350 62630 41410 62750
rect 41480 62600 41490 64370
rect 41540 64330 41600 64360
rect 42360 64330 42420 64360
rect 43840 64330 43900 64360
rect 146100 64290 146160 64320
rect 41540 64210 41600 64240
rect 42360 64210 42420 64240
rect 43840 64210 43900 64240
rect 146100 64170 146160 64200
rect 41540 64090 41600 64120
rect 42360 64090 42420 64120
rect 42910 64100 43030 64160
rect 43190 64100 43310 64160
rect 43030 64090 43090 64100
rect 43310 64090 43370 64100
rect 43840 64090 43900 64120
rect 42930 64080 43010 64090
rect 43030 64080 43150 64090
rect 43210 64080 43290 64090
rect 43310 64080 43430 64090
rect 41540 63970 41600 64000
rect 42360 63970 42420 64000
rect 42470 63980 42480 64070
rect 41540 63850 41600 63880
rect 42360 63850 42420 63880
rect 41540 63730 41600 63760
rect 42360 63730 42420 63760
rect 41540 63610 41600 63640
rect 42360 63610 42420 63640
rect 41540 63490 41600 63520
rect 42360 63490 42420 63520
rect 41540 63370 41600 63400
rect 42360 63370 42420 63400
rect 41540 63250 41600 63280
rect 42360 63250 42420 63280
rect 41540 63130 41600 63160
rect 42360 63130 42420 63160
rect 41540 63010 41600 63040
rect 42360 63010 42420 63040
rect 41540 62890 41600 62920
rect 42360 62890 42420 62920
rect 41540 62770 41600 62800
rect 42360 62770 42420 62800
rect 41540 62650 41600 62680
rect 42360 62650 42420 62680
rect 42560 62620 42570 63980
rect 42610 63950 42730 64010
rect 42730 63925 42790 63950
rect 42860 63940 42870 64070
rect 43010 64000 43020 64080
rect 43030 63980 43090 64080
rect 43150 64000 43160 64080
rect 43290 64000 43300 64080
rect 43310 63980 43370 64080
rect 43430 64000 43440 64080
rect 146100 64050 146160 64080
rect 43840 63970 43900 64000
rect 42860 63930 43500 63940
rect 42730 63915 43540 63925
rect 42730 63830 42790 63915
rect 43540 63865 43550 63915
rect 42620 63740 42700 63750
rect 42700 63660 42710 63740
rect 42860 63660 42870 63850
rect 42910 63800 43030 63860
rect 43190 63800 43310 63860
rect 43020 63770 43090 63800
rect 43030 63680 43090 63770
rect 43190 63710 43200 63800
rect 43300 63770 43370 63800
rect 43310 63680 43370 63770
rect 42860 63650 43490 63660
rect 42860 63640 42870 63650
rect 42620 63560 42700 63570
rect 42700 63480 42710 63560
rect 42770 63550 42780 63640
rect 42610 63360 42730 63420
rect 42730 63335 42790 63360
rect 42860 63350 42870 63550
rect 42910 63510 43030 63570
rect 43190 63510 43310 63570
rect 43030 63500 43090 63510
rect 43310 63500 43370 63510
rect 42930 63490 43010 63500
rect 43030 63490 43150 63500
rect 43210 63490 43290 63500
rect 43310 63490 43430 63500
rect 43010 63410 43020 63490
rect 43030 63390 43090 63490
rect 43150 63410 43160 63490
rect 43290 63410 43300 63490
rect 43310 63390 43370 63490
rect 43430 63410 43440 63490
rect 42860 63340 43500 63350
rect 43580 63340 43590 63640
rect 42730 63325 43540 63335
rect 42730 63240 42790 63325
rect 43540 63275 43550 63325
rect 42620 63140 42700 63150
rect 42700 63060 42710 63140
rect 42860 63070 42870 63260
rect 42910 63210 43030 63270
rect 43190 63210 43310 63270
rect 43020 63180 43090 63210
rect 43030 63090 43090 63180
rect 43190 63120 43200 63210
rect 43300 63180 43370 63210
rect 43310 63090 43370 63180
rect 42860 63060 43490 63070
rect 42860 63050 42870 63060
rect 42620 62960 42700 62970
rect 42770 62960 42780 63050
rect 42700 62880 42710 62960
rect 42610 62770 42730 62830
rect 42730 62745 42790 62770
rect 42860 62760 42870 62960
rect 42910 62920 43030 62980
rect 43190 62920 43310 62980
rect 43030 62910 43090 62920
rect 43310 62910 43370 62920
rect 42930 62900 43010 62910
rect 43030 62900 43150 62910
rect 43210 62900 43290 62910
rect 43310 62900 43430 62910
rect 43010 62820 43020 62900
rect 43030 62800 43090 62900
rect 43150 62820 43160 62900
rect 43290 62820 43300 62900
rect 43310 62800 43370 62900
rect 43430 62820 43440 62900
rect 42860 62750 43500 62760
rect 43580 62750 43590 63050
rect 42730 62735 43540 62745
rect 42730 62650 42790 62735
rect 43540 62685 43550 62735
rect 42860 62620 42870 62670
rect 42910 62620 43030 62680
rect 43190 62620 43310 62680
rect 43030 62610 43090 62620
rect 43310 62610 43370 62620
rect 43030 62600 43150 62610
rect 43310 62600 43430 62610
rect 40770 62590 40830 62600
rect 40530 62580 40610 62590
rect 40770 62580 40890 62590
rect 40610 62500 40620 62580
rect 40770 62480 40830 62580
rect 40890 62500 40900 62580
rect 41050 62480 41180 62600
rect 41540 62530 41600 62560
rect 42360 62530 42420 62560
rect 43030 62500 43090 62600
rect 43150 62520 43160 62600
rect 43310 62500 43370 62600
rect 43430 62520 43440 62600
rect 41090 62450 41180 62480
rect 43780 62460 43790 63940
rect 146100 63930 146160 63960
rect 43840 63850 43900 63880
rect 146100 63810 146160 63840
rect 43840 63730 43900 63760
rect 146100 63690 146160 63720
rect 43840 63610 43900 63640
rect 146100 63570 146160 63600
rect 43840 63490 43900 63520
rect 146100 63450 146160 63480
rect 43840 63370 43900 63400
rect 146100 63330 146160 63360
rect 43840 63250 43900 63280
rect 146100 63210 146160 63240
rect 43840 63130 43900 63160
rect 146100 63090 146160 63120
rect 43840 63010 43900 63040
rect 146100 62970 146160 63000
rect 43840 62890 43900 62920
rect 146100 62850 146160 62880
rect 43840 62770 43900 62800
rect 146100 62730 146160 62760
rect 147580 62730 147640 62746
rect 148400 62730 148460 62746
rect 149880 62730 149940 62746
rect 152220 62710 152250 62740
rect 152340 62710 152370 62740
rect 159520 62710 159550 62740
rect 159640 62710 159670 62740
rect 163520 62710 163550 62740
rect 163640 62710 163670 62740
rect 170810 62710 170840 62740
rect 170930 62710 170960 62740
rect 152100 62680 152160 62710
rect 152220 62680 152280 62710
rect 152340 62680 152400 62710
rect 159400 62680 159460 62710
rect 159520 62680 159580 62710
rect 159640 62680 159700 62710
rect 163400 62680 163460 62710
rect 163520 62680 163580 62710
rect 163640 62680 163700 62710
rect 170690 62680 170750 62710
rect 170810 62680 170870 62710
rect 170930 62680 170990 62710
rect 43840 62650 43900 62680
rect 146100 62610 146160 62640
rect 147580 62610 147640 62640
rect 148400 62610 148460 62640
rect 149880 62610 149940 62640
rect 152220 62560 152250 62620
rect 152340 62560 152370 62620
rect 159520 62560 159550 62620
rect 159640 62560 159670 62620
rect 163520 62560 163550 62620
rect 163640 62560 163670 62620
rect 170810 62560 170840 62620
rect 170930 62560 170960 62620
rect 43840 62530 43900 62560
rect 146100 62490 146160 62520
rect 147580 62490 147640 62520
rect 148400 62490 148460 62520
rect 149880 62490 149940 62520
rect 19060 62360 19070 62440
rect 19240 62360 19250 62440
rect 19420 62360 19430 62440
rect 19600 62360 19610 62440
rect 19780 62360 19790 62440
rect 19960 62360 19970 62440
rect 20140 62360 20150 62440
rect 20320 62360 20330 62440
rect 20500 62360 20510 62440
rect 20680 62360 20690 62440
rect 20860 62360 20870 62440
rect 21040 62360 21050 62440
rect 21220 62360 21230 62440
rect 21400 62360 21410 62440
rect 21580 62360 21590 62440
rect 21760 62360 21770 62440
rect 21940 62360 21950 62440
rect 22120 62360 22130 62440
rect 22300 62360 22310 62440
rect 22480 62360 22490 62440
rect 22660 62360 22670 62440
rect 22840 62360 22850 62440
rect 23020 62360 23030 62440
rect 23200 62360 23210 62440
rect 23380 62360 23390 62440
rect 23560 62360 23570 62440
rect 23740 62360 23750 62440
rect 23920 62360 23930 62440
rect 24100 62360 24110 62440
rect 24280 62360 24290 62440
rect 24460 62360 24470 62440
rect 24640 62360 24650 62440
rect 24820 62360 24830 62440
rect 25000 62360 25010 62440
rect 25180 62360 25190 62440
rect 25360 62360 25370 62440
rect 25540 62360 25550 62440
rect 25720 62360 25730 62440
rect 25900 62360 25910 62440
rect 26080 62360 26090 62440
rect 26260 62360 26270 62440
rect 26440 62360 26450 62440
rect 26620 62360 26630 62440
rect 27315 62415 27395 62425
rect 27495 62415 27575 62425
rect 27675 62415 27755 62425
rect 27855 62415 27935 62425
rect 28035 62415 28115 62425
rect 27395 62335 27405 62415
rect 27575 62335 27585 62415
rect 27755 62335 27765 62415
rect 27935 62335 27945 62415
rect 28115 62335 28125 62415
rect 30360 62360 30370 62440
rect 30540 62360 30550 62440
rect 30720 62360 30730 62440
rect 30900 62360 30910 62440
rect 31080 62360 31090 62440
rect 31260 62360 31270 62440
rect 31440 62360 31450 62440
rect 31620 62360 31630 62440
rect 31800 62360 31810 62440
rect 31980 62360 31990 62440
rect 32160 62360 32170 62440
rect 32340 62360 32350 62440
rect 32520 62360 32530 62440
rect 32700 62360 32710 62440
rect 32880 62360 32890 62440
rect 33060 62360 33070 62440
rect 33240 62360 33250 62440
rect 33420 62360 33430 62440
rect 33600 62360 33610 62440
rect 33780 62360 33790 62440
rect 33960 62360 33970 62440
rect 34140 62360 34150 62440
rect 34320 62360 34330 62440
rect 34500 62360 34510 62440
rect 34680 62360 34690 62440
rect 34860 62360 34870 62440
rect 35040 62360 35050 62440
rect 35220 62360 35230 62440
rect 35400 62360 35410 62440
rect 35580 62360 35590 62440
rect 35760 62360 35770 62440
rect 35940 62360 35950 62440
rect 36120 62360 36130 62440
rect 36300 62360 36310 62440
rect 36480 62360 36490 62440
rect 36660 62360 36670 62440
rect 36840 62360 36850 62440
rect 37020 62360 37030 62440
rect 37200 62360 37210 62440
rect 37380 62360 37390 62440
rect 37560 62360 37570 62440
rect 37740 62360 37750 62440
rect 37920 62360 37930 62440
rect 40060 62410 40120 62440
rect 41540 62410 41600 62440
rect 42360 62410 42420 62440
rect 43840 62410 43900 62440
rect 18980 62290 19060 62300
rect 19160 62290 19240 62300
rect 19340 62290 19420 62300
rect 19520 62290 19600 62300
rect 19700 62290 19780 62300
rect 19880 62290 19960 62300
rect 20060 62290 20140 62300
rect 20240 62290 20320 62300
rect 20420 62290 20500 62300
rect 20600 62290 20680 62300
rect 20780 62290 20860 62300
rect 20960 62290 21040 62300
rect 21140 62290 21220 62300
rect 21320 62290 21400 62300
rect 21500 62290 21580 62300
rect 21680 62290 21760 62300
rect 21860 62290 21940 62300
rect 22040 62290 22120 62300
rect 22220 62290 22300 62300
rect 22400 62290 22480 62300
rect 22580 62290 22660 62300
rect 22760 62290 22840 62300
rect 22940 62290 23020 62300
rect 23120 62290 23200 62300
rect 23300 62290 23380 62300
rect 23480 62290 23560 62300
rect 23660 62290 23740 62300
rect 23840 62290 23920 62300
rect 24020 62290 24100 62300
rect 24200 62290 24280 62300
rect 24380 62290 24460 62300
rect 24560 62290 24640 62300
rect 24740 62290 24820 62300
rect 24920 62290 25000 62300
rect 25100 62290 25180 62300
rect 25280 62290 25360 62300
rect 25460 62290 25540 62300
rect 25640 62290 25720 62300
rect 25820 62290 25900 62300
rect 26000 62290 26080 62300
rect 26180 62290 26260 62300
rect 26360 62290 26440 62300
rect 26540 62290 26620 62300
rect 30280 62290 30360 62300
rect 30460 62290 30540 62300
rect 30640 62290 30720 62300
rect 30820 62290 30900 62300
rect 31000 62290 31080 62300
rect 31180 62290 31260 62300
rect 31360 62290 31440 62300
rect 31540 62290 31620 62300
rect 31720 62290 31800 62300
rect 31900 62290 31980 62300
rect 32080 62290 32160 62300
rect 32260 62290 32340 62300
rect 32440 62290 32520 62300
rect 32620 62290 32700 62300
rect 32800 62290 32880 62300
rect 32980 62290 33060 62300
rect 33160 62290 33240 62300
rect 33340 62290 33420 62300
rect 33520 62290 33600 62300
rect 33700 62290 33780 62300
rect 33880 62290 33960 62300
rect 34060 62290 34140 62300
rect 34240 62290 34320 62300
rect 34420 62290 34500 62300
rect 34600 62290 34680 62300
rect 34780 62290 34860 62300
rect 34960 62290 35040 62300
rect 35140 62290 35220 62300
rect 35320 62290 35400 62300
rect 35500 62290 35580 62300
rect 35680 62290 35760 62300
rect 35860 62290 35940 62300
rect 36040 62290 36120 62300
rect 36220 62290 36300 62300
rect 36400 62290 36480 62300
rect 36580 62290 36660 62300
rect 36760 62290 36840 62300
rect 36940 62290 37020 62300
rect 37120 62290 37200 62300
rect 37300 62290 37380 62300
rect 37480 62290 37560 62300
rect 37660 62290 37740 62300
rect 37840 62290 37920 62300
rect 19060 62210 19070 62290
rect 19240 62210 19250 62290
rect 19420 62210 19430 62290
rect 19600 62210 19610 62290
rect 19780 62210 19790 62290
rect 19960 62210 19970 62290
rect 20140 62210 20150 62290
rect 20320 62210 20330 62290
rect 20500 62210 20510 62290
rect 20680 62210 20690 62290
rect 20860 62210 20870 62290
rect 21040 62210 21050 62290
rect 21220 62210 21230 62290
rect 21400 62210 21410 62290
rect 21580 62210 21590 62290
rect 21760 62210 21770 62290
rect 21940 62210 21950 62290
rect 22120 62210 22130 62290
rect 22300 62210 22310 62290
rect 22480 62210 22490 62290
rect 22660 62210 22670 62290
rect 22840 62210 22850 62290
rect 23020 62210 23030 62290
rect 23200 62210 23210 62290
rect 23380 62210 23390 62290
rect 23560 62210 23570 62290
rect 23740 62210 23750 62290
rect 23920 62210 23930 62290
rect 24100 62210 24110 62290
rect 24280 62210 24290 62290
rect 24460 62210 24470 62290
rect 24640 62210 24650 62290
rect 24820 62210 24830 62290
rect 25000 62210 25010 62290
rect 25180 62210 25190 62290
rect 25360 62210 25370 62290
rect 25540 62210 25550 62290
rect 25720 62210 25730 62290
rect 25900 62210 25910 62290
rect 26080 62210 26090 62290
rect 26260 62210 26270 62290
rect 26440 62210 26450 62290
rect 26620 62210 26630 62290
rect 27315 62235 27395 62245
rect 27495 62235 27575 62245
rect 27675 62235 27755 62245
rect 27855 62235 27935 62245
rect 28035 62235 28115 62245
rect 27395 62155 27405 62235
rect 27575 62155 27585 62235
rect 27755 62155 27765 62235
rect 27935 62155 27945 62235
rect 28115 62155 28125 62235
rect 30360 62210 30370 62290
rect 30540 62210 30550 62290
rect 30720 62210 30730 62290
rect 30900 62210 30910 62290
rect 31080 62210 31090 62290
rect 31260 62210 31270 62290
rect 31440 62210 31450 62290
rect 31620 62210 31630 62290
rect 31800 62210 31810 62290
rect 31980 62210 31990 62290
rect 32160 62210 32170 62290
rect 32340 62210 32350 62290
rect 32520 62210 32530 62290
rect 32700 62210 32710 62290
rect 32880 62210 32890 62290
rect 33060 62210 33070 62290
rect 33240 62210 33250 62290
rect 33420 62210 33430 62290
rect 33600 62210 33610 62290
rect 33780 62210 33790 62290
rect 33960 62210 33970 62290
rect 34140 62210 34150 62290
rect 34320 62210 34330 62290
rect 34500 62210 34510 62290
rect 34680 62210 34690 62290
rect 34860 62210 34870 62290
rect 35040 62210 35050 62290
rect 35220 62210 35230 62290
rect 35400 62210 35410 62290
rect 35580 62210 35590 62290
rect 35760 62210 35770 62290
rect 35940 62210 35950 62290
rect 36120 62210 36130 62290
rect 36300 62210 36310 62290
rect 36480 62210 36490 62290
rect 36660 62210 36670 62290
rect 36840 62210 36850 62290
rect 37020 62210 37030 62290
rect 37200 62210 37210 62290
rect 37380 62210 37390 62290
rect 37560 62210 37570 62290
rect 37740 62210 37750 62290
rect 37920 62210 37930 62290
rect 146100 62370 146160 62400
rect 147580 62370 147640 62400
rect 148400 62370 148460 62400
rect 149880 62370 149940 62400
rect 152080 62290 152160 62300
rect 152260 62290 152340 62300
rect 152440 62290 152520 62300
rect 152620 62290 152700 62300
rect 152800 62290 152880 62300
rect 152980 62290 153060 62300
rect 153160 62290 153240 62300
rect 153340 62290 153420 62300
rect 153520 62290 153600 62300
rect 153700 62290 153780 62300
rect 153880 62290 153960 62300
rect 154060 62290 154140 62300
rect 154240 62290 154320 62300
rect 154420 62290 154500 62300
rect 154600 62290 154680 62300
rect 154780 62290 154860 62300
rect 154960 62290 155040 62300
rect 155140 62290 155220 62300
rect 155320 62290 155400 62300
rect 155500 62290 155580 62300
rect 155680 62290 155760 62300
rect 155860 62290 155940 62300
rect 156040 62290 156120 62300
rect 156220 62290 156300 62300
rect 156400 62290 156480 62300
rect 156580 62290 156660 62300
rect 156760 62290 156840 62300
rect 156940 62290 157020 62300
rect 157120 62290 157200 62300
rect 157300 62290 157380 62300
rect 157480 62290 157560 62300
rect 157660 62290 157740 62300
rect 157840 62290 157920 62300
rect 158020 62290 158100 62300
rect 158200 62290 158280 62300
rect 158380 62290 158460 62300
rect 158560 62290 158640 62300
rect 158740 62290 158820 62300
rect 158920 62290 159000 62300
rect 159100 62290 159180 62300
rect 159280 62290 159360 62300
rect 159460 62290 159540 62300
rect 159640 62290 159720 62300
rect 163380 62290 163460 62300
rect 163560 62290 163640 62300
rect 163740 62290 163820 62300
rect 163920 62290 164000 62300
rect 164100 62290 164180 62300
rect 164280 62290 164360 62300
rect 164460 62290 164540 62300
rect 164640 62290 164720 62300
rect 164820 62290 164900 62300
rect 165000 62290 165080 62300
rect 165180 62290 165260 62300
rect 165360 62290 165440 62300
rect 165540 62290 165620 62300
rect 165720 62290 165800 62300
rect 165900 62290 165980 62300
rect 166080 62290 166160 62300
rect 166260 62290 166340 62300
rect 166440 62290 166520 62300
rect 166620 62290 166700 62300
rect 166800 62290 166880 62300
rect 166980 62290 167060 62300
rect 167160 62290 167240 62300
rect 167340 62290 167420 62300
rect 167520 62290 167600 62300
rect 167700 62290 167780 62300
rect 167880 62290 167960 62300
rect 168060 62290 168140 62300
rect 168240 62290 168320 62300
rect 168420 62290 168500 62300
rect 168600 62290 168680 62300
rect 168780 62290 168860 62300
rect 168960 62290 169040 62300
rect 169140 62290 169220 62300
rect 169320 62290 169400 62300
rect 169500 62290 169580 62300
rect 169680 62290 169760 62300
rect 169860 62290 169940 62300
rect 170040 62290 170120 62300
rect 170220 62290 170300 62300
rect 170400 62290 170480 62300
rect 170580 62290 170660 62300
rect 170760 62290 170840 62300
rect 170940 62290 171020 62300
rect 152160 62210 152170 62290
rect 152340 62210 152350 62290
rect 152520 62210 152530 62290
rect 152700 62210 152710 62290
rect 152880 62210 152890 62290
rect 153060 62210 153070 62290
rect 153240 62210 153250 62290
rect 153420 62210 153430 62290
rect 153600 62210 153610 62290
rect 153780 62210 153790 62290
rect 153960 62210 153970 62290
rect 154140 62210 154150 62290
rect 154320 62210 154330 62290
rect 154500 62210 154510 62290
rect 154680 62210 154690 62290
rect 154860 62210 154870 62290
rect 155040 62210 155050 62290
rect 155220 62210 155230 62290
rect 155400 62210 155410 62290
rect 155580 62210 155590 62290
rect 155760 62210 155770 62290
rect 155940 62210 155950 62290
rect 156120 62210 156130 62290
rect 156300 62210 156310 62290
rect 156480 62210 156490 62290
rect 156660 62210 156670 62290
rect 156840 62210 156850 62290
rect 157020 62210 157030 62290
rect 157200 62210 157210 62290
rect 157380 62210 157390 62290
rect 157560 62210 157570 62290
rect 157740 62210 157750 62290
rect 157920 62210 157930 62290
rect 158100 62210 158110 62290
rect 158280 62210 158290 62290
rect 158460 62210 158470 62290
rect 158640 62210 158650 62290
rect 158820 62210 158830 62290
rect 159000 62210 159010 62290
rect 159180 62210 159190 62290
rect 159360 62210 159370 62290
rect 159540 62210 159550 62290
rect 159720 62210 159730 62290
rect 160430 62265 160510 62275
rect 160590 62265 160670 62275
rect 160750 62265 160830 62275
rect 160910 62265 160990 62275
rect 161070 62265 161150 62275
rect 160510 62185 160520 62265
rect 160590 62185 160600 62265
rect 160670 62185 160680 62265
rect 160750 62185 160760 62265
rect 160830 62185 160840 62265
rect 160910 62185 160920 62265
rect 160990 62185 161000 62265
rect 161070 62185 161080 62265
rect 161150 62185 161160 62265
rect 163460 62210 163470 62290
rect 163640 62210 163650 62290
rect 163820 62210 163830 62290
rect 164000 62210 164010 62290
rect 164180 62210 164190 62290
rect 164360 62210 164370 62290
rect 164540 62210 164550 62290
rect 164720 62210 164730 62290
rect 164900 62210 164910 62290
rect 165080 62210 165090 62290
rect 165260 62210 165270 62290
rect 165440 62210 165450 62290
rect 165620 62210 165630 62290
rect 165800 62210 165810 62290
rect 165980 62210 165990 62290
rect 166160 62210 166170 62290
rect 166340 62210 166350 62290
rect 166520 62210 166530 62290
rect 166700 62210 166710 62290
rect 166880 62210 166890 62290
rect 167060 62210 167070 62290
rect 167240 62210 167250 62290
rect 167420 62210 167430 62290
rect 167600 62210 167610 62290
rect 167780 62210 167790 62290
rect 167960 62210 167970 62290
rect 168140 62210 168150 62290
rect 168320 62210 168330 62290
rect 168500 62210 168510 62290
rect 168680 62210 168690 62290
rect 168860 62210 168870 62290
rect 169040 62210 169050 62290
rect 169220 62210 169230 62290
rect 169400 62210 169410 62290
rect 169580 62210 169590 62290
rect 169760 62210 169770 62290
rect 169940 62210 169950 62290
rect 170120 62210 170130 62290
rect 170300 62210 170310 62290
rect 170480 62210 170490 62290
rect 170660 62210 170670 62290
rect 170840 62210 170850 62290
rect 171020 62210 171030 62290
rect 18980 62140 19060 62150
rect 19160 62140 19240 62150
rect 19340 62140 19420 62150
rect 19520 62140 19600 62150
rect 19700 62140 19780 62150
rect 19880 62140 19960 62150
rect 20060 62140 20140 62150
rect 20240 62140 20320 62150
rect 20420 62140 20500 62150
rect 20600 62140 20680 62150
rect 20780 62140 20860 62150
rect 20960 62140 21040 62150
rect 21140 62140 21220 62150
rect 21320 62140 21400 62150
rect 21500 62140 21580 62150
rect 21680 62140 21760 62150
rect 21860 62140 21940 62150
rect 22040 62140 22120 62150
rect 22220 62140 22300 62150
rect 22400 62140 22480 62150
rect 22580 62140 22660 62150
rect 22760 62140 22840 62150
rect 22940 62140 23020 62150
rect 23120 62140 23200 62150
rect 23300 62140 23380 62150
rect 23480 62140 23560 62150
rect 23660 62140 23740 62150
rect 23840 62140 23920 62150
rect 24020 62140 24100 62150
rect 24200 62140 24280 62150
rect 24380 62140 24460 62150
rect 24560 62140 24640 62150
rect 24740 62140 24820 62150
rect 24920 62140 25000 62150
rect 25100 62140 25180 62150
rect 25280 62140 25360 62150
rect 25460 62140 25540 62150
rect 25640 62140 25720 62150
rect 25820 62140 25900 62150
rect 26000 62140 26080 62150
rect 26180 62140 26260 62150
rect 26360 62140 26440 62150
rect 26540 62140 26620 62150
rect 30280 62140 30360 62150
rect 30460 62140 30540 62150
rect 30640 62140 30720 62150
rect 30820 62140 30900 62150
rect 31000 62140 31080 62150
rect 31180 62140 31260 62150
rect 31360 62140 31440 62150
rect 31540 62140 31620 62150
rect 31720 62140 31800 62150
rect 31900 62140 31980 62150
rect 32080 62140 32160 62150
rect 32260 62140 32340 62150
rect 32440 62140 32520 62150
rect 32620 62140 32700 62150
rect 32800 62140 32880 62150
rect 32980 62140 33060 62150
rect 33160 62140 33240 62150
rect 33340 62140 33420 62150
rect 33520 62140 33600 62150
rect 33700 62140 33780 62150
rect 33880 62140 33960 62150
rect 34060 62140 34140 62150
rect 34240 62140 34320 62150
rect 34420 62140 34500 62150
rect 34600 62140 34680 62150
rect 34780 62140 34860 62150
rect 34960 62140 35040 62150
rect 35140 62140 35220 62150
rect 35320 62140 35400 62150
rect 35500 62140 35580 62150
rect 35680 62140 35760 62150
rect 35860 62140 35940 62150
rect 36040 62140 36120 62150
rect 36220 62140 36300 62150
rect 36400 62140 36480 62150
rect 36580 62140 36660 62150
rect 36760 62140 36840 62150
rect 36940 62140 37020 62150
rect 37120 62140 37200 62150
rect 37300 62140 37380 62150
rect 37480 62140 37560 62150
rect 37660 62140 37740 62150
rect 37840 62140 37920 62150
rect 40060 62140 40140 62150
rect 40200 62140 40280 62150
rect 40340 62140 40420 62150
rect 40480 62140 40560 62150
rect 40620 62140 40700 62150
rect 40760 62140 40840 62150
rect 40900 62140 40980 62150
rect 41040 62140 41120 62150
rect 41180 62140 41260 62150
rect 41320 62140 41400 62150
rect 42360 62140 42440 62150
rect 42500 62140 42580 62150
rect 42640 62140 42720 62150
rect 42780 62140 42860 62150
rect 42920 62140 43000 62150
rect 43060 62140 43140 62150
rect 43200 62140 43280 62150
rect 43340 62140 43420 62150
rect 43480 62140 43560 62150
rect 43620 62140 43700 62150
rect 146300 62140 146380 62150
rect 146440 62140 146520 62150
rect 146580 62140 146660 62150
rect 146720 62140 146800 62150
rect 146860 62140 146940 62150
rect 147000 62140 147080 62150
rect 147140 62140 147220 62150
rect 147280 62140 147360 62150
rect 147420 62140 147500 62150
rect 147560 62140 147640 62150
rect 148600 62140 148680 62150
rect 148740 62140 148820 62150
rect 148880 62140 148960 62150
rect 149020 62140 149100 62150
rect 149160 62140 149240 62150
rect 149300 62140 149380 62150
rect 149440 62140 149520 62150
rect 149580 62140 149660 62150
rect 149720 62140 149800 62150
rect 149860 62140 149940 62150
rect 152080 62140 152160 62150
rect 152260 62140 152340 62150
rect 152440 62140 152520 62150
rect 152620 62140 152700 62150
rect 152800 62140 152880 62150
rect 152980 62140 153060 62150
rect 153160 62140 153240 62150
rect 153340 62140 153420 62150
rect 153520 62140 153600 62150
rect 153700 62140 153780 62150
rect 153880 62140 153960 62150
rect 154060 62140 154140 62150
rect 154240 62140 154320 62150
rect 154420 62140 154500 62150
rect 154600 62140 154680 62150
rect 154780 62140 154860 62150
rect 154960 62140 155040 62150
rect 155140 62140 155220 62150
rect 155320 62140 155400 62150
rect 155500 62140 155580 62150
rect 155680 62140 155760 62150
rect 155860 62140 155940 62150
rect 156040 62140 156120 62150
rect 156220 62140 156300 62150
rect 156400 62140 156480 62150
rect 156580 62140 156660 62150
rect 156760 62140 156840 62150
rect 156940 62140 157020 62150
rect 157120 62140 157200 62150
rect 157300 62140 157380 62150
rect 157480 62140 157560 62150
rect 157660 62140 157740 62150
rect 157840 62140 157920 62150
rect 158020 62140 158100 62150
rect 158200 62140 158280 62150
rect 158380 62140 158460 62150
rect 158560 62140 158640 62150
rect 158740 62140 158820 62150
rect 158920 62140 159000 62150
rect 159100 62140 159180 62150
rect 159280 62140 159360 62150
rect 159460 62140 159540 62150
rect 159640 62140 159720 62150
rect 163380 62140 163460 62150
rect 163560 62140 163640 62150
rect 163740 62140 163820 62150
rect 163920 62140 164000 62150
rect 164100 62140 164180 62150
rect 164280 62140 164360 62150
rect 164460 62140 164540 62150
rect 164640 62140 164720 62150
rect 164820 62140 164900 62150
rect 165000 62140 165080 62150
rect 165180 62140 165260 62150
rect 165360 62140 165440 62150
rect 165540 62140 165620 62150
rect 165720 62140 165800 62150
rect 165900 62140 165980 62150
rect 166080 62140 166160 62150
rect 166260 62140 166340 62150
rect 166440 62140 166520 62150
rect 166620 62140 166700 62150
rect 166800 62140 166880 62150
rect 166980 62140 167060 62150
rect 167160 62140 167240 62150
rect 167340 62140 167420 62150
rect 167520 62140 167600 62150
rect 167700 62140 167780 62150
rect 167880 62140 167960 62150
rect 168060 62140 168140 62150
rect 168240 62140 168320 62150
rect 168420 62140 168500 62150
rect 168600 62140 168680 62150
rect 168780 62140 168860 62150
rect 168960 62140 169040 62150
rect 169140 62140 169220 62150
rect 169320 62140 169400 62150
rect 169500 62140 169580 62150
rect 169680 62140 169760 62150
rect 169860 62140 169940 62150
rect 170040 62140 170120 62150
rect 170220 62140 170300 62150
rect 170400 62140 170480 62150
rect 170580 62140 170660 62150
rect 170760 62140 170840 62150
rect 170940 62140 171020 62150
rect 19060 62060 19070 62140
rect 19240 62060 19250 62140
rect 19420 62060 19430 62140
rect 19600 62060 19610 62140
rect 19780 62060 19790 62140
rect 19960 62060 19970 62140
rect 20140 62060 20150 62140
rect 20320 62060 20330 62140
rect 20500 62060 20510 62140
rect 20680 62060 20690 62140
rect 20860 62060 20870 62140
rect 21040 62060 21050 62140
rect 21220 62060 21230 62140
rect 21400 62060 21410 62140
rect 21580 62060 21590 62140
rect 21760 62060 21770 62140
rect 21940 62060 21950 62140
rect 22120 62060 22130 62140
rect 22300 62060 22310 62140
rect 22480 62060 22490 62140
rect 22660 62060 22670 62140
rect 22840 62060 22850 62140
rect 23020 62060 23030 62140
rect 23200 62060 23210 62140
rect 23380 62060 23390 62140
rect 23560 62060 23570 62140
rect 23740 62060 23750 62140
rect 23920 62060 23930 62140
rect 24100 62060 24110 62140
rect 24280 62060 24290 62140
rect 24460 62060 24470 62140
rect 24640 62060 24650 62140
rect 24820 62060 24830 62140
rect 25000 62060 25010 62140
rect 25180 62060 25190 62140
rect 25360 62060 25370 62140
rect 25540 62060 25550 62140
rect 25720 62060 25730 62140
rect 25900 62060 25910 62140
rect 26080 62060 26090 62140
rect 26260 62060 26270 62140
rect 26440 62060 26450 62140
rect 26620 62060 26630 62140
rect 30360 62060 30370 62140
rect 30540 62060 30550 62140
rect 30720 62060 30730 62140
rect 30900 62060 30910 62140
rect 31080 62060 31090 62140
rect 31260 62060 31270 62140
rect 31440 62060 31450 62140
rect 31620 62060 31630 62140
rect 31800 62060 31810 62140
rect 31980 62060 31990 62140
rect 32160 62060 32170 62140
rect 32340 62060 32350 62140
rect 32520 62060 32530 62140
rect 32700 62060 32710 62140
rect 32880 62060 32890 62140
rect 33060 62060 33070 62140
rect 33240 62060 33250 62140
rect 33420 62060 33430 62140
rect 33600 62060 33610 62140
rect 33780 62060 33790 62140
rect 33960 62060 33970 62140
rect 34140 62060 34150 62140
rect 34320 62060 34330 62140
rect 34500 62060 34510 62140
rect 34680 62060 34690 62140
rect 34860 62060 34870 62140
rect 35040 62060 35050 62140
rect 35220 62060 35230 62140
rect 35400 62060 35410 62140
rect 35580 62060 35590 62140
rect 35760 62060 35770 62140
rect 35940 62060 35950 62140
rect 36120 62060 36130 62140
rect 36300 62060 36310 62140
rect 36480 62060 36490 62140
rect 36660 62060 36670 62140
rect 36840 62060 36850 62140
rect 37020 62060 37030 62140
rect 37200 62060 37210 62140
rect 37380 62060 37390 62140
rect 37560 62060 37570 62140
rect 37740 62060 37750 62140
rect 37920 62060 37930 62140
rect 40140 62060 40150 62140
rect 40280 62060 40290 62140
rect 40420 62060 40430 62140
rect 40560 62060 40570 62140
rect 40700 62060 40710 62140
rect 40840 62060 40850 62140
rect 40980 62060 40990 62140
rect 41120 62060 41130 62140
rect 41260 62060 41270 62140
rect 41400 62060 41410 62140
rect 42440 62060 42450 62140
rect 42580 62060 42590 62140
rect 42720 62060 42730 62140
rect 42860 62060 42870 62140
rect 43000 62060 43010 62140
rect 43140 62060 43150 62140
rect 43280 62060 43290 62140
rect 43420 62060 43430 62140
rect 43560 62060 43570 62140
rect 43700 62060 43710 62140
rect 146380 62081 146390 62140
rect 146520 62081 146530 62140
rect 146660 62081 146670 62140
rect 146800 62081 146810 62140
rect 146940 62081 146950 62140
rect 147080 62081 147090 62140
rect 147220 62081 147230 62140
rect 147360 62081 147370 62140
rect 147500 62081 147510 62140
rect 147640 62081 147650 62140
rect 148680 62081 148690 62140
rect 148820 62081 148830 62140
rect 148960 62081 148970 62140
rect 149100 62081 149110 62140
rect 149240 62081 149250 62140
rect 149380 62081 149390 62140
rect 149520 62081 149530 62140
rect 149660 62081 149670 62140
rect 149800 62081 149810 62140
rect 149940 62081 149950 62140
rect 152160 62081 152170 62140
rect 152340 62081 152350 62140
rect 152520 62081 152530 62140
rect 152700 62081 152710 62140
rect 152880 62081 152890 62140
rect 153060 62081 153070 62140
rect 153240 62081 153250 62140
rect 153420 62081 153430 62140
rect 153600 62081 153610 62140
rect 153780 62081 153790 62140
rect 153960 62081 153970 62140
rect 154140 62081 154150 62140
rect 154320 62081 154330 62140
rect 154500 62081 154510 62140
rect 154680 62081 154690 62140
rect 154860 62081 154870 62140
rect 155040 62081 155050 62140
rect 155220 62081 155230 62140
rect 155400 62081 155410 62140
rect 155580 62081 155590 62140
rect 155760 62081 155770 62140
rect 155940 62081 155950 62140
rect 156120 62081 156130 62140
rect 156300 62081 156310 62140
rect 156480 62081 156490 62140
rect 156660 62081 156670 62140
rect 156840 62081 156850 62140
rect 157020 62081 157030 62140
rect 157200 62081 157210 62140
rect 157380 62081 157390 62140
rect 157560 62081 157570 62140
rect 157740 62081 157750 62140
rect 157920 62081 157930 62140
rect 158100 62081 158110 62140
rect 158280 62081 158290 62140
rect 158460 62081 158470 62140
rect 158640 62081 158650 62140
rect 158820 62081 158830 62140
rect 159000 62081 159010 62140
rect 159180 62081 159190 62140
rect 159360 62081 159370 62140
rect 159540 62081 159550 62140
rect 159720 62081 159730 62140
rect 163460 62081 163470 62140
rect 163640 62081 163650 62140
rect 163820 62081 163830 62140
rect 164000 62081 164010 62140
rect 164180 62081 164190 62140
rect 164360 62081 164370 62140
rect 164540 62081 164550 62140
rect 164720 62081 164730 62140
rect 164900 62081 164910 62140
rect 165080 62081 165090 62140
rect 165260 62081 165270 62140
rect 165440 62081 165450 62140
rect 165620 62081 165630 62140
rect 165800 62081 165810 62140
rect 165980 62081 165990 62140
rect 166160 62081 166170 62140
rect 166340 62081 166350 62140
rect 166520 62081 166530 62140
rect 166700 62081 166710 62140
rect 166880 62081 166890 62140
rect 167060 62081 167070 62140
rect 167240 62081 167250 62140
rect 167420 62081 167430 62140
rect 167600 62081 167610 62140
rect 167780 62081 167790 62140
rect 167960 62081 167970 62140
rect 168140 62081 168150 62140
rect 168320 62081 168330 62140
rect 168500 62081 168510 62140
rect 168680 62081 168690 62140
rect 168860 62081 168870 62140
rect 169040 62081 169050 62140
rect 169220 62081 169230 62140
rect 169400 62081 169410 62140
rect 169580 62081 169590 62140
rect 169760 62081 169770 62140
rect 169940 62081 169950 62140
rect 170120 62081 170130 62140
rect 170300 62081 170310 62140
rect 170480 62081 170490 62140
rect 170660 62081 170670 62140
rect 170840 62081 170850 62140
rect 171020 62081 171030 62140
rect 146040 62000 147700 62081
rect 148340 62000 150000 62081
rect 152000 62000 159800 62081
rect 163210 62060 171100 62081
rect 163300 62000 171100 62060
rect 30360 61920 30440 61930
rect 30680 61920 30760 61930
rect 31000 61920 31080 61930
rect 31320 61920 31400 61930
rect 31640 61920 31720 61930
rect 31960 61920 32040 61930
rect 32280 61920 32360 61930
rect 32600 61920 32680 61930
rect 32920 61920 33000 61930
rect 33240 61920 33320 61930
rect 33560 61920 33640 61930
rect 33880 61920 33960 61930
rect 34200 61920 34280 61930
rect 34520 61920 34600 61930
rect 34840 61920 34920 61930
rect 35160 61920 35240 61930
rect 35480 61920 35560 61930
rect 35800 61920 35880 61930
rect 36120 61920 36200 61930
rect 36440 61920 36520 61930
rect 36760 61920 36840 61930
rect 37080 61920 37160 61930
rect 37400 61920 37480 61930
rect 37720 61920 37800 61930
rect 40180 61920 40260 61930
rect 40500 61920 40580 61930
rect 40820 61920 40900 61930
rect 41140 61920 41220 61930
rect 42560 61920 42640 61930
rect 42880 61920 42960 61930
rect 43200 61920 43280 61930
rect 43520 61920 43600 61930
rect 18970 61890 19050 61900
rect 19290 61890 19370 61900
rect 19610 61890 19690 61900
rect 19930 61890 20010 61900
rect 20250 61890 20330 61900
rect 20570 61890 20650 61900
rect 20890 61890 20970 61900
rect 21210 61890 21290 61900
rect 21530 61890 21610 61900
rect 21850 61890 21930 61900
rect 22170 61890 22250 61900
rect 22490 61890 22570 61900
rect 22810 61890 22890 61900
rect 23130 61890 23210 61900
rect 23450 61890 23530 61900
rect 23770 61890 23850 61900
rect 24090 61890 24170 61900
rect 24410 61890 24490 61900
rect 24730 61890 24810 61900
rect 25050 61890 25130 61900
rect 25370 61890 25450 61900
rect 25690 61890 25770 61900
rect 26010 61890 26090 61900
rect 26330 61890 26410 61900
rect 19050 61810 19060 61890
rect 19370 61810 19380 61890
rect 19690 61810 19700 61890
rect 20010 61810 20020 61890
rect 20330 61810 20340 61890
rect 20650 61810 20660 61890
rect 20970 61810 20980 61890
rect 21290 61810 21300 61890
rect 21610 61810 21620 61890
rect 21930 61810 21940 61890
rect 22250 61810 22260 61890
rect 22570 61810 22580 61890
rect 22890 61810 22900 61890
rect 23210 61810 23220 61890
rect 23530 61810 23540 61890
rect 23850 61810 23860 61890
rect 24170 61810 24180 61890
rect 24490 61810 24500 61890
rect 24810 61810 24820 61890
rect 25130 61810 25140 61890
rect 25450 61810 25460 61890
rect 25770 61810 25780 61890
rect 26090 61810 26100 61890
rect 26410 61810 26420 61890
rect 30440 61840 30450 61920
rect 30760 61840 30770 61920
rect 31080 61840 31090 61920
rect 31400 61840 31410 61920
rect 31720 61840 31730 61920
rect 32040 61840 32050 61920
rect 32360 61840 32370 61920
rect 32680 61840 32690 61920
rect 33000 61840 33010 61920
rect 33320 61840 33330 61920
rect 33640 61840 33650 61920
rect 33960 61840 33970 61920
rect 34280 61840 34290 61920
rect 34600 61840 34610 61920
rect 34920 61840 34930 61920
rect 35240 61840 35250 61920
rect 35560 61840 35570 61920
rect 35880 61840 35890 61920
rect 36200 61840 36210 61920
rect 36520 61840 36530 61920
rect 36840 61840 36850 61920
rect 37160 61840 37170 61920
rect 37480 61840 37490 61920
rect 37800 61840 37810 61920
rect 40260 61840 40270 61920
rect 40580 61840 40590 61920
rect 40900 61840 40910 61920
rect 41220 61840 41230 61920
rect 42640 61840 42650 61920
rect 42960 61840 42970 61920
rect 43280 61840 43290 61920
rect 43600 61840 43610 61920
rect 146400 61911 146480 61921
rect 146720 61911 146800 61921
rect 147040 61911 147120 61921
rect 147360 61911 147440 61921
rect 148780 61911 148860 61921
rect 149100 61911 149180 61921
rect 149420 61911 149500 61921
rect 149740 61911 149820 61921
rect 152200 61911 152280 61921
rect 152520 61911 152600 61921
rect 152840 61911 152920 61921
rect 153160 61911 153240 61921
rect 153480 61911 153560 61921
rect 153800 61911 153880 61921
rect 154120 61911 154200 61921
rect 154440 61911 154520 61921
rect 154760 61911 154840 61921
rect 155080 61911 155160 61921
rect 155400 61911 155480 61921
rect 155720 61911 155800 61921
rect 156040 61911 156120 61921
rect 156360 61911 156440 61921
rect 156680 61911 156760 61921
rect 157000 61911 157080 61921
rect 157320 61911 157400 61921
rect 157640 61911 157720 61921
rect 157960 61911 158040 61921
rect 158280 61911 158360 61921
rect 158600 61911 158680 61921
rect 158920 61911 159000 61921
rect 159240 61911 159320 61921
rect 159560 61911 159640 61921
rect 146480 61831 146490 61911
rect 146800 61831 146810 61911
rect 147120 61831 147130 61911
rect 147440 61831 147450 61911
rect 148860 61831 148870 61911
rect 149180 61831 149190 61911
rect 149500 61831 149510 61911
rect 149820 61831 149830 61911
rect 152280 61831 152290 61911
rect 152600 61831 152610 61911
rect 152920 61831 152930 61911
rect 153240 61831 153250 61911
rect 153560 61831 153570 61911
rect 153880 61831 153890 61911
rect 154200 61831 154210 61911
rect 154520 61831 154530 61911
rect 154840 61831 154850 61911
rect 155160 61831 155170 61911
rect 155480 61831 155490 61911
rect 155800 61831 155810 61911
rect 156120 61831 156130 61911
rect 156440 61831 156450 61911
rect 156760 61831 156770 61911
rect 157080 61831 157090 61911
rect 157400 61831 157410 61911
rect 157720 61831 157730 61911
rect 158040 61831 158050 61911
rect 158360 61831 158370 61911
rect 158680 61831 158690 61911
rect 159000 61831 159010 61911
rect 159320 61831 159330 61911
rect 159640 61831 159650 61911
rect 163590 61881 163670 61891
rect 163910 61881 163990 61891
rect 164230 61881 164310 61891
rect 164550 61881 164630 61891
rect 164870 61881 164950 61891
rect 165190 61881 165270 61891
rect 165510 61881 165590 61891
rect 165830 61881 165910 61891
rect 166150 61881 166230 61891
rect 166470 61881 166550 61891
rect 166790 61881 166870 61891
rect 167110 61881 167190 61891
rect 167430 61881 167510 61891
rect 167750 61881 167830 61891
rect 168070 61881 168150 61891
rect 168390 61881 168470 61891
rect 168710 61881 168790 61891
rect 169030 61881 169110 61891
rect 169350 61881 169430 61891
rect 169670 61881 169750 61891
rect 169990 61881 170070 61891
rect 170310 61881 170390 61891
rect 170630 61881 170710 61891
rect 170950 61881 171030 61891
rect 163670 61801 163680 61881
rect 163990 61801 164000 61881
rect 164310 61801 164320 61881
rect 164630 61801 164640 61881
rect 164950 61801 164960 61881
rect 165270 61801 165280 61881
rect 165590 61801 165600 61881
rect 165910 61801 165920 61881
rect 166230 61801 166240 61881
rect 166550 61801 166560 61881
rect 166870 61801 166880 61881
rect 167190 61801 167200 61881
rect 167510 61801 167520 61881
rect 167830 61801 167840 61881
rect 168150 61801 168160 61881
rect 168470 61801 168480 61881
rect 168790 61801 168800 61881
rect 169110 61801 169120 61881
rect 169430 61801 169440 61881
rect 169750 61801 169760 61881
rect 170070 61801 170080 61881
rect 170390 61801 170400 61881
rect 170710 61801 170720 61881
rect 171030 61801 171040 61881
rect 30520 61760 30600 61770
rect 30840 61760 30920 61770
rect 31160 61760 31240 61770
rect 31480 61760 31560 61770
rect 31800 61760 31880 61770
rect 32120 61760 32200 61770
rect 32440 61760 32520 61770
rect 32760 61760 32840 61770
rect 33080 61760 33160 61770
rect 33400 61760 33480 61770
rect 33720 61760 33800 61770
rect 34040 61760 34120 61770
rect 34360 61760 34440 61770
rect 34680 61760 34760 61770
rect 35000 61760 35080 61770
rect 35320 61760 35400 61770
rect 35640 61760 35720 61770
rect 35960 61760 36040 61770
rect 36280 61760 36360 61770
rect 36600 61760 36680 61770
rect 36920 61760 37000 61770
rect 37240 61760 37320 61770
rect 37560 61760 37640 61770
rect 40340 61760 40420 61770
rect 40660 61760 40740 61770
rect 40980 61760 41060 61770
rect 42720 61760 42800 61770
rect 43040 61760 43120 61770
rect 43360 61760 43440 61770
rect 19130 61730 19210 61740
rect 19450 61730 19530 61740
rect 19770 61730 19850 61740
rect 20090 61730 20170 61740
rect 20410 61730 20490 61740
rect 20730 61730 20810 61740
rect 21050 61730 21130 61740
rect 21370 61730 21450 61740
rect 21690 61730 21770 61740
rect 22010 61730 22090 61740
rect 22330 61730 22410 61740
rect 22650 61730 22730 61740
rect 22970 61730 23050 61740
rect 23290 61730 23370 61740
rect 23610 61730 23690 61740
rect 23930 61730 24010 61740
rect 24250 61730 24330 61740
rect 24570 61730 24650 61740
rect 24890 61730 24970 61740
rect 25210 61730 25290 61740
rect 25530 61730 25610 61740
rect 25850 61730 25930 61740
rect 26170 61730 26250 61740
rect 19210 61650 19220 61730
rect 19530 61650 19540 61730
rect 19850 61650 19860 61730
rect 20170 61650 20180 61730
rect 20490 61650 20500 61730
rect 20810 61650 20820 61730
rect 21130 61650 21140 61730
rect 21450 61650 21460 61730
rect 21770 61650 21780 61730
rect 22090 61650 22100 61730
rect 22410 61650 22420 61730
rect 22730 61650 22740 61730
rect 23050 61650 23060 61730
rect 23370 61650 23380 61730
rect 23690 61650 23700 61730
rect 24010 61650 24020 61730
rect 24330 61650 24340 61730
rect 24650 61650 24660 61730
rect 24970 61650 24980 61730
rect 25290 61650 25300 61730
rect 25610 61650 25620 61730
rect 25930 61650 25940 61730
rect 26250 61650 26260 61730
rect 30600 61680 30610 61760
rect 30920 61680 30930 61760
rect 31240 61680 31250 61760
rect 31560 61680 31570 61760
rect 31880 61680 31890 61760
rect 32200 61680 32210 61760
rect 32520 61680 32530 61760
rect 32840 61680 32850 61760
rect 33160 61680 33170 61760
rect 33480 61680 33490 61760
rect 33800 61680 33810 61760
rect 34120 61680 34130 61760
rect 34440 61680 34450 61760
rect 34760 61680 34770 61760
rect 35080 61680 35090 61760
rect 35400 61680 35410 61760
rect 35720 61680 35730 61760
rect 36040 61680 36050 61760
rect 36360 61680 36370 61760
rect 36680 61680 36690 61760
rect 37000 61680 37010 61760
rect 37320 61680 37330 61760
rect 37640 61680 37650 61760
rect 40420 61680 40430 61760
rect 40740 61680 40750 61760
rect 41060 61680 41070 61760
rect 42800 61680 42810 61760
rect 43120 61680 43130 61760
rect 43440 61680 43450 61760
rect 146560 61751 146640 61761
rect 146880 61751 146960 61761
rect 147200 61751 147280 61761
rect 148940 61751 149020 61761
rect 149260 61751 149340 61761
rect 149580 61751 149660 61761
rect 152360 61751 152440 61761
rect 152680 61751 152760 61761
rect 153000 61751 153080 61761
rect 153320 61751 153400 61761
rect 153640 61751 153720 61761
rect 153960 61751 154040 61761
rect 154280 61751 154360 61761
rect 154600 61751 154680 61761
rect 154920 61751 155000 61761
rect 155240 61751 155320 61761
rect 155560 61751 155640 61761
rect 155880 61751 155960 61761
rect 156200 61751 156280 61761
rect 156520 61751 156600 61761
rect 156840 61751 156920 61761
rect 157160 61751 157240 61761
rect 157480 61751 157560 61761
rect 157800 61751 157880 61761
rect 158120 61751 158200 61761
rect 158440 61751 158520 61761
rect 158760 61751 158840 61761
rect 159080 61751 159160 61761
rect 159400 61751 159480 61761
rect 146640 61671 146650 61751
rect 146960 61671 146970 61751
rect 147280 61671 147290 61751
rect 149020 61671 149030 61751
rect 149340 61671 149350 61751
rect 149660 61671 149670 61751
rect 152440 61671 152450 61751
rect 152760 61671 152770 61751
rect 153080 61671 153090 61751
rect 153400 61671 153410 61751
rect 153720 61671 153730 61751
rect 154040 61671 154050 61751
rect 154360 61671 154370 61751
rect 154680 61671 154690 61751
rect 155000 61671 155010 61751
rect 155320 61671 155330 61751
rect 155640 61671 155650 61751
rect 155960 61671 155970 61751
rect 156280 61671 156290 61751
rect 156600 61671 156610 61751
rect 156920 61671 156930 61751
rect 157240 61671 157250 61751
rect 157560 61671 157570 61751
rect 157880 61671 157890 61751
rect 158200 61671 158210 61751
rect 158520 61671 158530 61751
rect 158840 61671 158850 61751
rect 159160 61671 159170 61751
rect 159480 61671 159490 61751
rect 163750 61721 163830 61731
rect 164070 61721 164150 61731
rect 164390 61721 164470 61731
rect 164710 61721 164790 61731
rect 165030 61721 165110 61731
rect 165350 61721 165430 61731
rect 165670 61721 165750 61731
rect 165990 61721 166070 61731
rect 166310 61721 166390 61731
rect 166630 61721 166710 61731
rect 166950 61721 167030 61731
rect 167270 61721 167350 61731
rect 167590 61721 167670 61731
rect 167910 61721 167990 61731
rect 168230 61721 168310 61731
rect 168550 61721 168630 61731
rect 168870 61721 168950 61731
rect 169190 61721 169270 61731
rect 169510 61721 169590 61731
rect 169830 61721 169910 61731
rect 170150 61721 170230 61731
rect 170470 61721 170550 61731
rect 170790 61721 170870 61731
rect 163830 61641 163840 61721
rect 164150 61641 164160 61721
rect 164470 61641 164480 61721
rect 164790 61641 164800 61721
rect 165110 61641 165120 61721
rect 165430 61641 165440 61721
rect 165750 61641 165760 61721
rect 166070 61641 166080 61721
rect 166390 61641 166400 61721
rect 166710 61641 166720 61721
rect 167030 61641 167040 61721
rect 167350 61641 167360 61721
rect 167670 61641 167680 61721
rect 167990 61641 168000 61721
rect 168310 61641 168320 61721
rect 168630 61641 168640 61721
rect 168950 61641 168960 61721
rect 169270 61641 169280 61721
rect 169590 61641 169600 61721
rect 169910 61641 169920 61721
rect 170230 61641 170240 61721
rect 170550 61641 170560 61721
rect 170870 61641 170880 61721
rect 30360 61600 30440 61610
rect 30680 61600 30760 61610
rect 31000 61600 31080 61610
rect 31320 61600 31400 61610
rect 31640 61600 31720 61610
rect 31960 61600 32040 61610
rect 32280 61600 32360 61610
rect 32600 61600 32680 61610
rect 32920 61600 33000 61610
rect 33240 61600 33320 61610
rect 33560 61600 33640 61610
rect 33880 61600 33960 61610
rect 34200 61600 34280 61610
rect 34520 61600 34600 61610
rect 34840 61600 34920 61610
rect 35160 61600 35240 61610
rect 35480 61600 35560 61610
rect 35800 61600 35880 61610
rect 36120 61600 36200 61610
rect 36440 61600 36520 61610
rect 36760 61600 36840 61610
rect 37080 61600 37160 61610
rect 37400 61600 37480 61610
rect 37720 61600 37800 61610
rect 40180 61600 40260 61610
rect 40500 61600 40580 61610
rect 40820 61600 40900 61610
rect 41140 61600 41220 61610
rect 42560 61600 42640 61610
rect 42880 61600 42960 61610
rect 43200 61600 43280 61610
rect 43520 61600 43600 61610
rect 18970 61570 19050 61580
rect 19290 61570 19370 61580
rect 19610 61570 19690 61580
rect 19930 61570 20010 61580
rect 20250 61570 20330 61580
rect 20570 61570 20650 61580
rect 20890 61570 20970 61580
rect 21210 61570 21290 61580
rect 21530 61570 21610 61580
rect 21850 61570 21930 61580
rect 22170 61570 22250 61580
rect 22490 61570 22570 61580
rect 22810 61570 22890 61580
rect 23130 61570 23210 61580
rect 23450 61570 23530 61580
rect 23770 61570 23850 61580
rect 24090 61570 24170 61580
rect 24410 61570 24490 61580
rect 24730 61570 24810 61580
rect 25050 61570 25130 61580
rect 25370 61570 25450 61580
rect 25690 61570 25770 61580
rect 26010 61570 26090 61580
rect 26330 61570 26410 61580
rect 19050 61490 19060 61570
rect 19370 61490 19380 61570
rect 19690 61490 19700 61570
rect 20010 61490 20020 61570
rect 20330 61490 20340 61570
rect 20650 61490 20660 61570
rect 20970 61490 20980 61570
rect 21290 61490 21300 61570
rect 21610 61490 21620 61570
rect 21930 61490 21940 61570
rect 22250 61490 22260 61570
rect 22570 61490 22580 61570
rect 22890 61490 22900 61570
rect 23210 61490 23220 61570
rect 23530 61490 23540 61570
rect 23850 61490 23860 61570
rect 24170 61490 24180 61570
rect 24490 61490 24500 61570
rect 24810 61490 24820 61570
rect 25130 61490 25140 61570
rect 25450 61490 25460 61570
rect 25770 61490 25780 61570
rect 26090 61490 26100 61570
rect 26410 61490 26420 61570
rect 30440 61520 30450 61600
rect 30760 61520 30770 61600
rect 31080 61520 31090 61600
rect 31400 61520 31410 61600
rect 31720 61520 31730 61600
rect 32040 61520 32050 61600
rect 32360 61520 32370 61600
rect 32680 61520 32690 61600
rect 33000 61520 33010 61600
rect 33320 61520 33330 61600
rect 33640 61520 33650 61600
rect 33960 61520 33970 61600
rect 34280 61520 34290 61600
rect 34600 61520 34610 61600
rect 34920 61520 34930 61600
rect 35240 61520 35250 61600
rect 35560 61520 35570 61600
rect 35880 61520 35890 61600
rect 36200 61520 36210 61600
rect 36520 61520 36530 61600
rect 36840 61520 36850 61600
rect 37160 61520 37170 61600
rect 37480 61520 37490 61600
rect 37800 61520 37810 61600
rect 40260 61520 40270 61600
rect 40580 61520 40590 61600
rect 40900 61520 40910 61600
rect 41220 61520 41230 61600
rect 42640 61520 42650 61600
rect 42960 61520 42970 61600
rect 43280 61520 43290 61600
rect 43600 61520 43610 61600
rect 146400 61591 146480 61601
rect 146720 61591 146800 61601
rect 147040 61591 147120 61601
rect 147360 61591 147440 61601
rect 148780 61591 148860 61601
rect 149100 61591 149180 61601
rect 149420 61591 149500 61601
rect 149740 61591 149820 61601
rect 152200 61591 152280 61601
rect 152520 61591 152600 61601
rect 152840 61591 152920 61601
rect 153160 61591 153240 61601
rect 153480 61591 153560 61601
rect 153800 61591 153880 61601
rect 154120 61591 154200 61601
rect 154440 61591 154520 61601
rect 154760 61591 154840 61601
rect 155080 61591 155160 61601
rect 155400 61591 155480 61601
rect 155720 61591 155800 61601
rect 156040 61591 156120 61601
rect 156360 61591 156440 61601
rect 156680 61591 156760 61601
rect 157000 61591 157080 61601
rect 157320 61591 157400 61601
rect 157640 61591 157720 61601
rect 157960 61591 158040 61601
rect 158280 61591 158360 61601
rect 158600 61591 158680 61601
rect 158920 61591 159000 61601
rect 159240 61591 159320 61601
rect 159560 61591 159640 61601
rect 146480 61511 146490 61591
rect 146800 61511 146810 61591
rect 147120 61511 147130 61591
rect 147440 61511 147450 61591
rect 148860 61511 148870 61591
rect 149180 61511 149190 61591
rect 149500 61511 149510 61591
rect 149820 61511 149830 61591
rect 152280 61511 152290 61591
rect 152600 61511 152610 61591
rect 152920 61511 152930 61591
rect 153240 61511 153250 61591
rect 153560 61511 153570 61591
rect 153880 61511 153890 61591
rect 154200 61511 154210 61591
rect 154520 61511 154530 61591
rect 154840 61511 154850 61591
rect 155160 61511 155170 61591
rect 155480 61511 155490 61591
rect 155800 61511 155810 61591
rect 156120 61511 156130 61591
rect 156440 61511 156450 61591
rect 156760 61511 156770 61591
rect 157080 61511 157090 61591
rect 157400 61511 157410 61591
rect 157720 61511 157730 61591
rect 158040 61511 158050 61591
rect 158360 61511 158370 61591
rect 158680 61511 158690 61591
rect 159000 61511 159010 61591
rect 159320 61511 159330 61591
rect 159640 61511 159650 61591
rect 163590 61561 163670 61571
rect 163910 61561 163990 61571
rect 164230 61561 164310 61571
rect 164550 61561 164630 61571
rect 164870 61561 164950 61571
rect 165190 61561 165270 61571
rect 165510 61561 165590 61571
rect 165830 61561 165910 61571
rect 166150 61561 166230 61571
rect 166470 61561 166550 61571
rect 166790 61561 166870 61571
rect 167110 61561 167190 61571
rect 167430 61561 167510 61571
rect 167750 61561 167830 61571
rect 168070 61561 168150 61571
rect 168390 61561 168470 61571
rect 168710 61561 168790 61571
rect 169030 61561 169110 61571
rect 169350 61561 169430 61571
rect 169670 61561 169750 61571
rect 169990 61561 170070 61571
rect 170310 61561 170390 61571
rect 170630 61561 170710 61571
rect 170950 61561 171030 61571
rect 163670 61481 163680 61561
rect 163990 61481 164000 61561
rect 164310 61481 164320 61561
rect 164630 61481 164640 61561
rect 164950 61481 164960 61561
rect 165270 61481 165280 61561
rect 165590 61481 165600 61561
rect 165910 61481 165920 61561
rect 166230 61481 166240 61561
rect 166550 61481 166560 61561
rect 166870 61481 166880 61561
rect 167190 61481 167200 61561
rect 167510 61481 167520 61561
rect 167830 61481 167840 61561
rect 168150 61481 168160 61561
rect 168470 61481 168480 61561
rect 168790 61481 168800 61561
rect 169110 61481 169120 61561
rect 169430 61481 169440 61561
rect 169750 61481 169760 61561
rect 170070 61481 170080 61561
rect 170390 61481 170400 61561
rect 170710 61481 170720 61561
rect 171030 61481 171040 61561
rect 30520 61440 30600 61450
rect 30840 61440 30920 61450
rect 31160 61440 31240 61450
rect 31480 61440 31560 61450
rect 31800 61440 31880 61450
rect 32120 61440 32200 61450
rect 32440 61440 32520 61450
rect 32760 61440 32840 61450
rect 33080 61440 33160 61450
rect 33400 61440 33480 61450
rect 33720 61440 33800 61450
rect 34040 61440 34120 61450
rect 34360 61440 34440 61450
rect 34680 61440 34760 61450
rect 35000 61440 35080 61450
rect 35320 61440 35400 61450
rect 35640 61440 35720 61450
rect 35960 61440 36040 61450
rect 36280 61440 36360 61450
rect 36600 61440 36680 61450
rect 36920 61440 37000 61450
rect 37240 61440 37320 61450
rect 37560 61440 37640 61450
rect 40340 61440 40420 61450
rect 40660 61440 40740 61450
rect 40980 61440 41060 61450
rect 42720 61440 42800 61450
rect 43040 61440 43120 61450
rect 43360 61440 43440 61450
rect 19130 61410 19210 61420
rect 19450 61410 19530 61420
rect 19770 61410 19850 61420
rect 20090 61410 20170 61420
rect 20410 61410 20490 61420
rect 20730 61410 20810 61420
rect 21050 61410 21130 61420
rect 21370 61410 21450 61420
rect 21690 61410 21770 61420
rect 22010 61410 22090 61420
rect 22330 61410 22410 61420
rect 22650 61410 22730 61420
rect 22970 61410 23050 61420
rect 23290 61410 23370 61420
rect 23610 61410 23690 61420
rect 23930 61410 24010 61420
rect 24250 61410 24330 61420
rect 24570 61410 24650 61420
rect 24890 61410 24970 61420
rect 25210 61410 25290 61420
rect 25530 61410 25610 61420
rect 25850 61410 25930 61420
rect 26170 61410 26250 61420
rect 19210 61330 19220 61410
rect 19530 61330 19540 61410
rect 19850 61330 19860 61410
rect 20170 61330 20180 61410
rect 20490 61330 20500 61410
rect 20810 61330 20820 61410
rect 21130 61330 21140 61410
rect 21450 61330 21460 61410
rect 21770 61330 21780 61410
rect 22090 61330 22100 61410
rect 22410 61330 22420 61410
rect 22730 61330 22740 61410
rect 23050 61330 23060 61410
rect 23370 61330 23380 61410
rect 23690 61330 23700 61410
rect 24010 61330 24020 61410
rect 24330 61330 24340 61410
rect 24650 61330 24660 61410
rect 24970 61330 24980 61410
rect 25290 61330 25300 61410
rect 25610 61330 25620 61410
rect 25930 61330 25940 61410
rect 26250 61330 26260 61410
rect 30600 61360 30610 61440
rect 30920 61360 30930 61440
rect 31240 61360 31250 61440
rect 31560 61360 31570 61440
rect 31880 61360 31890 61440
rect 32200 61360 32210 61440
rect 32520 61360 32530 61440
rect 32840 61360 32850 61440
rect 33160 61360 33170 61440
rect 33480 61360 33490 61440
rect 33800 61360 33810 61440
rect 34120 61360 34130 61440
rect 34440 61360 34450 61440
rect 34760 61360 34770 61440
rect 35080 61360 35090 61440
rect 35400 61360 35410 61440
rect 35720 61360 35730 61440
rect 36040 61360 36050 61440
rect 36360 61360 36370 61440
rect 36680 61360 36690 61440
rect 37000 61360 37010 61440
rect 37320 61360 37330 61440
rect 37640 61360 37650 61440
rect 40420 61360 40430 61440
rect 40740 61360 40750 61440
rect 41060 61360 41070 61440
rect 42800 61360 42810 61440
rect 43120 61360 43130 61440
rect 43440 61360 43450 61440
rect 146560 61431 146640 61441
rect 146880 61431 146960 61441
rect 147200 61431 147280 61441
rect 148940 61431 149020 61441
rect 149260 61431 149340 61441
rect 149580 61431 149660 61441
rect 152360 61431 152440 61441
rect 152680 61431 152760 61441
rect 153000 61431 153080 61441
rect 153320 61431 153400 61441
rect 153640 61431 153720 61441
rect 153960 61431 154040 61441
rect 154280 61431 154360 61441
rect 154600 61431 154680 61441
rect 154920 61431 155000 61441
rect 155240 61431 155320 61441
rect 155560 61431 155640 61441
rect 155880 61431 155960 61441
rect 156200 61431 156280 61441
rect 156520 61431 156600 61441
rect 156840 61431 156920 61441
rect 157160 61431 157240 61441
rect 157480 61431 157560 61441
rect 157800 61431 157880 61441
rect 158120 61431 158200 61441
rect 158440 61431 158520 61441
rect 158760 61431 158840 61441
rect 159080 61431 159160 61441
rect 159400 61431 159480 61441
rect 146640 61351 146650 61431
rect 146960 61351 146970 61431
rect 147280 61351 147290 61431
rect 149020 61351 149030 61431
rect 149340 61351 149350 61431
rect 149660 61351 149670 61431
rect 152440 61351 152450 61431
rect 152760 61351 152770 61431
rect 153080 61351 153090 61431
rect 153400 61351 153410 61431
rect 153720 61351 153730 61431
rect 154040 61351 154050 61431
rect 154360 61351 154370 61431
rect 154680 61351 154690 61431
rect 155000 61351 155010 61431
rect 155320 61351 155330 61431
rect 155640 61351 155650 61431
rect 155960 61351 155970 61431
rect 156280 61351 156290 61431
rect 156600 61351 156610 61431
rect 156920 61351 156930 61431
rect 157240 61351 157250 61431
rect 157560 61351 157570 61431
rect 157880 61351 157890 61431
rect 158200 61351 158210 61431
rect 158520 61351 158530 61431
rect 158840 61351 158850 61431
rect 159160 61351 159170 61431
rect 159480 61351 159490 61431
rect 163750 61401 163830 61411
rect 164070 61401 164150 61411
rect 164390 61401 164470 61411
rect 164710 61401 164790 61411
rect 165030 61401 165110 61411
rect 165350 61401 165430 61411
rect 165670 61401 165750 61411
rect 165990 61401 166070 61411
rect 166310 61401 166390 61411
rect 166630 61401 166710 61411
rect 166950 61401 167030 61411
rect 167270 61401 167350 61411
rect 167590 61401 167670 61411
rect 167910 61401 167990 61411
rect 168230 61401 168310 61411
rect 168550 61401 168630 61411
rect 168870 61401 168950 61411
rect 169190 61401 169270 61411
rect 169510 61401 169590 61411
rect 169830 61401 169910 61411
rect 170150 61401 170230 61411
rect 170470 61401 170550 61411
rect 170790 61401 170870 61411
rect 163830 61321 163840 61401
rect 164150 61321 164160 61401
rect 164470 61321 164480 61401
rect 164790 61321 164800 61401
rect 165110 61321 165120 61401
rect 165430 61321 165440 61401
rect 165750 61321 165760 61401
rect 166070 61321 166080 61401
rect 166390 61321 166400 61401
rect 166710 61321 166720 61401
rect 167030 61321 167040 61401
rect 167350 61321 167360 61401
rect 167670 61321 167680 61401
rect 167990 61321 168000 61401
rect 168310 61321 168320 61401
rect 168630 61321 168640 61401
rect 168950 61321 168960 61401
rect 169270 61321 169280 61401
rect 169590 61321 169600 61401
rect 169910 61321 169920 61401
rect 170230 61321 170240 61401
rect 170550 61321 170560 61401
rect 170870 61321 170880 61401
rect 30360 61180 30440 61190
rect 30680 61180 30760 61190
rect 31000 61180 31080 61190
rect 31320 61180 31400 61190
rect 31640 61180 31720 61190
rect 31960 61180 32040 61190
rect 32280 61180 32360 61190
rect 32600 61180 32680 61190
rect 32920 61180 33000 61190
rect 33240 61180 33320 61190
rect 33560 61180 33640 61190
rect 33880 61180 33960 61190
rect 34200 61180 34280 61190
rect 34520 61180 34600 61190
rect 34840 61180 34920 61190
rect 35160 61180 35240 61190
rect 35480 61180 35560 61190
rect 35800 61180 35880 61190
rect 36120 61180 36200 61190
rect 36440 61180 36520 61190
rect 36760 61180 36840 61190
rect 37080 61180 37160 61190
rect 37400 61180 37480 61190
rect 37720 61180 37800 61190
rect 40180 61180 40260 61190
rect 40500 61180 40580 61190
rect 40820 61180 40900 61190
rect 41140 61180 41220 61190
rect 42560 61180 42640 61190
rect 42880 61180 42960 61190
rect 43200 61180 43280 61190
rect 43520 61180 43600 61190
rect 18970 61150 19050 61160
rect 19290 61150 19370 61160
rect 19610 61150 19690 61160
rect 19930 61150 20010 61160
rect 20250 61150 20330 61160
rect 20570 61150 20650 61160
rect 20890 61150 20970 61160
rect 21210 61150 21290 61160
rect 21530 61150 21610 61160
rect 21850 61150 21930 61160
rect 22170 61150 22250 61160
rect 22490 61150 22570 61160
rect 22810 61150 22890 61160
rect 23130 61150 23210 61160
rect 23450 61150 23530 61160
rect 23770 61150 23850 61160
rect 24090 61150 24170 61160
rect 24410 61150 24490 61160
rect 24730 61150 24810 61160
rect 25050 61150 25130 61160
rect 25370 61150 25450 61160
rect 25690 61150 25770 61160
rect 26010 61150 26090 61160
rect 26330 61150 26410 61160
rect 19050 61070 19060 61150
rect 19370 61070 19380 61150
rect 19690 61070 19700 61150
rect 20010 61070 20020 61150
rect 20330 61070 20340 61150
rect 20650 61070 20660 61150
rect 20970 61070 20980 61150
rect 21290 61070 21300 61150
rect 21610 61070 21620 61150
rect 21930 61070 21940 61150
rect 22250 61070 22260 61150
rect 22570 61070 22580 61150
rect 22890 61070 22900 61150
rect 23210 61070 23220 61150
rect 23530 61070 23540 61150
rect 23850 61070 23860 61150
rect 24170 61070 24180 61150
rect 24490 61070 24500 61150
rect 24810 61070 24820 61150
rect 25130 61070 25140 61150
rect 25450 61070 25460 61150
rect 25770 61070 25780 61150
rect 26090 61070 26100 61150
rect 26410 61070 26420 61150
rect 30440 61100 30450 61180
rect 30760 61100 30770 61180
rect 31080 61100 31090 61180
rect 31400 61100 31410 61180
rect 31720 61100 31730 61180
rect 32040 61100 32050 61180
rect 32360 61100 32370 61180
rect 32680 61100 32690 61180
rect 33000 61100 33010 61180
rect 33320 61100 33330 61180
rect 33640 61100 33650 61180
rect 33960 61100 33970 61180
rect 34280 61100 34290 61180
rect 34600 61100 34610 61180
rect 34920 61100 34930 61180
rect 35240 61100 35250 61180
rect 35560 61100 35570 61180
rect 35880 61100 35890 61180
rect 36200 61100 36210 61180
rect 36520 61100 36530 61180
rect 36840 61100 36850 61180
rect 37160 61100 37170 61180
rect 37480 61100 37490 61180
rect 37800 61100 37810 61180
rect 40260 61100 40270 61180
rect 40580 61100 40590 61180
rect 40900 61100 40910 61180
rect 41220 61100 41230 61180
rect 42640 61100 42650 61180
rect 42960 61100 42970 61180
rect 43280 61100 43290 61180
rect 43600 61100 43610 61180
rect 146400 61171 146480 61181
rect 146720 61171 146800 61181
rect 147040 61171 147120 61181
rect 147360 61171 147440 61181
rect 148780 61171 148860 61181
rect 149100 61171 149180 61181
rect 149420 61171 149500 61181
rect 149740 61171 149820 61181
rect 152200 61171 152280 61181
rect 152520 61171 152600 61181
rect 152840 61171 152920 61181
rect 153160 61171 153240 61181
rect 153480 61171 153560 61181
rect 153800 61171 153880 61181
rect 154120 61171 154200 61181
rect 154440 61171 154520 61181
rect 154760 61171 154840 61181
rect 155080 61171 155160 61181
rect 155400 61171 155480 61181
rect 155720 61171 155800 61181
rect 156040 61171 156120 61181
rect 156360 61171 156440 61181
rect 156680 61171 156760 61181
rect 157000 61171 157080 61181
rect 157320 61171 157400 61181
rect 157640 61171 157720 61181
rect 157960 61171 158040 61181
rect 158280 61171 158360 61181
rect 158600 61171 158680 61181
rect 158920 61171 159000 61181
rect 159240 61171 159320 61181
rect 159560 61171 159640 61181
rect 146480 61091 146490 61171
rect 146800 61091 146810 61171
rect 147120 61091 147130 61171
rect 147440 61091 147450 61171
rect 148860 61091 148870 61171
rect 149180 61091 149190 61171
rect 149500 61091 149510 61171
rect 149820 61091 149830 61171
rect 152280 61091 152290 61171
rect 152600 61091 152610 61171
rect 152920 61091 152930 61171
rect 153240 61091 153250 61171
rect 153560 61091 153570 61171
rect 153880 61091 153890 61171
rect 154200 61091 154210 61171
rect 154520 61091 154530 61171
rect 154840 61091 154850 61171
rect 155160 61091 155170 61171
rect 155480 61091 155490 61171
rect 155800 61091 155810 61171
rect 156120 61091 156130 61171
rect 156440 61091 156450 61171
rect 156760 61091 156770 61171
rect 157080 61091 157090 61171
rect 157400 61091 157410 61171
rect 157720 61091 157730 61171
rect 158040 61091 158050 61171
rect 158360 61091 158370 61171
rect 158680 61091 158690 61171
rect 159000 61091 159010 61171
rect 159320 61091 159330 61171
rect 159640 61091 159650 61171
rect 163590 61141 163670 61151
rect 163910 61141 163990 61151
rect 164230 61141 164310 61151
rect 164550 61141 164630 61151
rect 164870 61141 164950 61151
rect 165190 61141 165270 61151
rect 165510 61141 165590 61151
rect 165830 61141 165910 61151
rect 166150 61141 166230 61151
rect 166470 61141 166550 61151
rect 166790 61141 166870 61151
rect 167110 61141 167190 61151
rect 167430 61141 167510 61151
rect 167750 61141 167830 61151
rect 168070 61141 168150 61151
rect 168390 61141 168470 61151
rect 168710 61141 168790 61151
rect 169030 61141 169110 61151
rect 169350 61141 169430 61151
rect 169670 61141 169750 61151
rect 169990 61141 170070 61151
rect 170310 61141 170390 61151
rect 170630 61141 170710 61151
rect 170950 61141 171030 61151
rect 163670 61061 163680 61141
rect 163990 61061 164000 61141
rect 164310 61061 164320 61141
rect 164630 61061 164640 61141
rect 164950 61061 164960 61141
rect 165270 61061 165280 61141
rect 165590 61061 165600 61141
rect 165910 61061 165920 61141
rect 166230 61061 166240 61141
rect 166550 61061 166560 61141
rect 166870 61061 166880 61141
rect 167190 61061 167200 61141
rect 167510 61061 167520 61141
rect 167830 61061 167840 61141
rect 168150 61061 168160 61141
rect 168470 61061 168480 61141
rect 168790 61061 168800 61141
rect 169110 61061 169120 61141
rect 169430 61061 169440 61141
rect 169750 61061 169760 61141
rect 170070 61061 170080 61141
rect 170390 61061 170400 61141
rect 170710 61061 170720 61141
rect 171030 61061 171040 61141
rect 30520 61020 30600 61030
rect 30840 61020 30920 61030
rect 31160 61020 31240 61030
rect 31480 61020 31560 61030
rect 31800 61020 31880 61030
rect 32120 61020 32200 61030
rect 32440 61020 32520 61030
rect 32760 61020 32840 61030
rect 33080 61020 33160 61030
rect 33400 61020 33480 61030
rect 33720 61020 33800 61030
rect 34040 61020 34120 61030
rect 34360 61020 34440 61030
rect 34680 61020 34760 61030
rect 35000 61020 35080 61030
rect 35320 61020 35400 61030
rect 35640 61020 35720 61030
rect 35960 61020 36040 61030
rect 36280 61020 36360 61030
rect 36600 61020 36680 61030
rect 36920 61020 37000 61030
rect 37240 61020 37320 61030
rect 37560 61020 37640 61030
rect 40340 61020 40420 61030
rect 40660 61020 40740 61030
rect 40980 61020 41060 61030
rect 42720 61020 42800 61030
rect 43040 61020 43120 61030
rect 43360 61020 43440 61030
rect 19130 60990 19210 61000
rect 19450 60990 19530 61000
rect 19770 60990 19850 61000
rect 20090 60990 20170 61000
rect 20410 60990 20490 61000
rect 20730 60990 20810 61000
rect 21050 60990 21130 61000
rect 21370 60990 21450 61000
rect 21690 60990 21770 61000
rect 22010 60990 22090 61000
rect 22330 60990 22410 61000
rect 22650 60990 22730 61000
rect 22970 60990 23050 61000
rect 23290 60990 23370 61000
rect 23610 60990 23690 61000
rect 23930 60990 24010 61000
rect 24250 60990 24330 61000
rect 24570 60990 24650 61000
rect 24890 60990 24970 61000
rect 25210 60990 25290 61000
rect 25530 60990 25610 61000
rect 25850 60990 25930 61000
rect 26170 60990 26250 61000
rect 19210 60910 19220 60990
rect 19530 60910 19540 60990
rect 19850 60910 19860 60990
rect 20170 60910 20180 60990
rect 20490 60910 20500 60990
rect 20810 60910 20820 60990
rect 21130 60910 21140 60990
rect 21450 60910 21460 60990
rect 21770 60910 21780 60990
rect 22090 60910 22100 60990
rect 22410 60910 22420 60990
rect 22730 60910 22740 60990
rect 23050 60910 23060 60990
rect 23370 60910 23380 60990
rect 23690 60910 23700 60990
rect 24010 60910 24020 60990
rect 24330 60910 24340 60990
rect 24650 60910 24660 60990
rect 24970 60910 24980 60990
rect 25290 60910 25300 60990
rect 25610 60910 25620 60990
rect 25930 60910 25940 60990
rect 26250 60910 26260 60990
rect 30600 60940 30610 61020
rect 30920 60940 30930 61020
rect 31240 60940 31250 61020
rect 31560 60940 31570 61020
rect 31880 60940 31890 61020
rect 32200 60940 32210 61020
rect 32520 60940 32530 61020
rect 32840 60940 32850 61020
rect 33160 60940 33170 61020
rect 33480 60940 33490 61020
rect 33800 60940 33810 61020
rect 34120 60940 34130 61020
rect 34440 60940 34450 61020
rect 34760 60940 34770 61020
rect 35080 60940 35090 61020
rect 35400 60940 35410 61020
rect 35720 60940 35730 61020
rect 36040 60940 36050 61020
rect 36360 60940 36370 61020
rect 36680 60940 36690 61020
rect 37000 60940 37010 61020
rect 37320 60940 37330 61020
rect 37640 60940 37650 61020
rect 40420 60940 40430 61020
rect 40740 60940 40750 61020
rect 41060 60940 41070 61020
rect 42800 60940 42810 61020
rect 43120 60940 43130 61020
rect 43440 60940 43450 61020
rect 146560 61011 146640 61021
rect 146880 61011 146960 61021
rect 147200 61011 147280 61021
rect 148940 61011 149020 61021
rect 149260 61011 149340 61021
rect 149580 61011 149660 61021
rect 152360 61011 152440 61021
rect 152680 61011 152760 61021
rect 153000 61011 153080 61021
rect 153320 61011 153400 61021
rect 153640 61011 153720 61021
rect 153960 61011 154040 61021
rect 154280 61011 154360 61021
rect 154600 61011 154680 61021
rect 154920 61011 155000 61021
rect 155240 61011 155320 61021
rect 155560 61011 155640 61021
rect 155880 61011 155960 61021
rect 156200 61011 156280 61021
rect 156520 61011 156600 61021
rect 156840 61011 156920 61021
rect 157160 61011 157240 61021
rect 157480 61011 157560 61021
rect 157800 61011 157880 61021
rect 158120 61011 158200 61021
rect 158440 61011 158520 61021
rect 158760 61011 158840 61021
rect 159080 61011 159160 61021
rect 159400 61011 159480 61021
rect 146640 60931 146650 61011
rect 146960 60931 146970 61011
rect 147280 60931 147290 61011
rect 149020 60931 149030 61011
rect 149340 60931 149350 61011
rect 149660 60931 149670 61011
rect 152440 60931 152450 61011
rect 152760 60931 152770 61011
rect 153080 60931 153090 61011
rect 153400 60931 153410 61011
rect 153720 60931 153730 61011
rect 154040 60931 154050 61011
rect 154360 60931 154370 61011
rect 154680 60931 154690 61011
rect 155000 60931 155010 61011
rect 155320 60931 155330 61011
rect 155640 60931 155650 61011
rect 155960 60931 155970 61011
rect 156280 60931 156290 61011
rect 156600 60931 156610 61011
rect 156920 60931 156930 61011
rect 157240 60931 157250 61011
rect 157560 60931 157570 61011
rect 157880 60931 157890 61011
rect 158200 60931 158210 61011
rect 158520 60931 158530 61011
rect 158840 60931 158850 61011
rect 159160 60931 159170 61011
rect 159480 60931 159490 61011
rect 163750 60981 163830 60991
rect 164070 60981 164150 60991
rect 164390 60981 164470 60991
rect 164710 60981 164790 60991
rect 165030 60981 165110 60991
rect 165350 60981 165430 60991
rect 165670 60981 165750 60991
rect 165990 60981 166070 60991
rect 166310 60981 166390 60991
rect 166630 60981 166710 60991
rect 166950 60981 167030 60991
rect 167270 60981 167350 60991
rect 167590 60981 167670 60991
rect 167910 60981 167990 60991
rect 168230 60981 168310 60991
rect 168550 60981 168630 60991
rect 168870 60981 168950 60991
rect 169190 60981 169270 60991
rect 169510 60981 169590 60991
rect 169830 60981 169910 60991
rect 170150 60981 170230 60991
rect 170470 60981 170550 60991
rect 170790 60981 170870 60991
rect 163830 60901 163840 60981
rect 164150 60901 164160 60981
rect 164470 60901 164480 60981
rect 164790 60901 164800 60981
rect 165110 60901 165120 60981
rect 165430 60901 165440 60981
rect 165750 60901 165760 60981
rect 166070 60901 166080 60981
rect 166390 60901 166400 60981
rect 166710 60901 166720 60981
rect 167030 60901 167040 60981
rect 167350 60901 167360 60981
rect 167670 60901 167680 60981
rect 167990 60901 168000 60981
rect 168310 60901 168320 60981
rect 168630 60901 168640 60981
rect 168950 60901 168960 60981
rect 169270 60901 169280 60981
rect 169590 60901 169600 60981
rect 169910 60901 169920 60981
rect 170230 60901 170240 60981
rect 170550 60901 170560 60981
rect 170870 60901 170880 60981
rect 30360 60860 30440 60870
rect 30680 60860 30760 60870
rect 31000 60860 31080 60870
rect 31320 60860 31400 60870
rect 31640 60860 31720 60870
rect 31960 60860 32040 60870
rect 32280 60860 32360 60870
rect 32600 60860 32680 60870
rect 32920 60860 33000 60870
rect 33240 60860 33320 60870
rect 33560 60860 33640 60870
rect 33880 60860 33960 60870
rect 34200 60860 34280 60870
rect 34520 60860 34600 60870
rect 34840 60860 34920 60870
rect 35160 60860 35240 60870
rect 35480 60860 35560 60870
rect 35800 60860 35880 60870
rect 36120 60860 36200 60870
rect 36440 60860 36520 60870
rect 36760 60860 36840 60870
rect 37080 60860 37160 60870
rect 37400 60860 37480 60870
rect 37720 60860 37800 60870
rect 40180 60860 40260 60870
rect 40500 60860 40580 60870
rect 40820 60860 40900 60870
rect 41140 60860 41220 60870
rect 42560 60860 42640 60870
rect 42880 60860 42960 60870
rect 43200 60860 43280 60870
rect 43520 60860 43600 60870
rect 18970 60830 19050 60840
rect 19290 60830 19370 60840
rect 19610 60830 19690 60840
rect 19930 60830 20010 60840
rect 20250 60830 20330 60840
rect 20570 60830 20650 60840
rect 20890 60830 20970 60840
rect 21210 60830 21290 60840
rect 21530 60830 21610 60840
rect 21850 60830 21930 60840
rect 22170 60830 22250 60840
rect 22490 60830 22570 60840
rect 22810 60830 22890 60840
rect 23130 60830 23210 60840
rect 23450 60830 23530 60840
rect 23770 60830 23850 60840
rect 24090 60830 24170 60840
rect 24410 60830 24490 60840
rect 24730 60830 24810 60840
rect 25050 60830 25130 60840
rect 25370 60830 25450 60840
rect 25690 60830 25770 60840
rect 26010 60830 26090 60840
rect 26330 60830 26410 60840
rect 19050 60750 19060 60830
rect 19370 60750 19380 60830
rect 19690 60750 19700 60830
rect 20010 60750 20020 60830
rect 20330 60750 20340 60830
rect 20650 60750 20660 60830
rect 20970 60750 20980 60830
rect 21290 60750 21300 60830
rect 21610 60750 21620 60830
rect 21930 60750 21940 60830
rect 22250 60750 22260 60830
rect 22570 60750 22580 60830
rect 22890 60750 22900 60830
rect 23210 60750 23220 60830
rect 23530 60750 23540 60830
rect 23850 60750 23860 60830
rect 24170 60750 24180 60830
rect 24490 60750 24500 60830
rect 24810 60750 24820 60830
rect 25130 60750 25140 60830
rect 25450 60750 25460 60830
rect 25770 60750 25780 60830
rect 26090 60750 26100 60830
rect 26410 60750 26420 60830
rect 30440 60780 30450 60860
rect 30760 60780 30770 60860
rect 31080 60780 31090 60860
rect 31400 60780 31410 60860
rect 31720 60780 31730 60860
rect 32040 60780 32050 60860
rect 32360 60780 32370 60860
rect 32680 60780 32690 60860
rect 33000 60780 33010 60860
rect 33320 60780 33330 60860
rect 33640 60780 33650 60860
rect 33960 60780 33970 60860
rect 34280 60780 34290 60860
rect 34600 60780 34610 60860
rect 34920 60780 34930 60860
rect 35240 60780 35250 60860
rect 35560 60780 35570 60860
rect 35880 60780 35890 60860
rect 36200 60780 36210 60860
rect 36520 60780 36530 60860
rect 36840 60780 36850 60860
rect 37160 60780 37170 60860
rect 37480 60780 37490 60860
rect 37800 60780 37810 60860
rect 40260 60780 40270 60860
rect 40580 60780 40590 60860
rect 40900 60780 40910 60860
rect 41220 60780 41230 60860
rect 42640 60780 42650 60860
rect 42960 60780 42970 60860
rect 43280 60780 43290 60860
rect 43600 60780 43610 60860
rect 146400 60851 146480 60861
rect 146720 60851 146800 60861
rect 147040 60851 147120 60861
rect 147360 60851 147440 60861
rect 148780 60851 148860 60861
rect 149100 60851 149180 60861
rect 149420 60851 149500 60861
rect 149740 60851 149820 60861
rect 152200 60851 152280 60861
rect 152520 60851 152600 60861
rect 152840 60851 152920 60861
rect 153160 60851 153240 60861
rect 153480 60851 153560 60861
rect 153800 60851 153880 60861
rect 154120 60851 154200 60861
rect 154440 60851 154520 60861
rect 154760 60851 154840 60861
rect 155080 60851 155160 60861
rect 155400 60851 155480 60861
rect 155720 60851 155800 60861
rect 156040 60851 156120 60861
rect 156360 60851 156440 60861
rect 156680 60851 156760 60861
rect 157000 60851 157080 60861
rect 157320 60851 157400 60861
rect 157640 60851 157720 60861
rect 157960 60851 158040 60861
rect 158280 60851 158360 60861
rect 158600 60851 158680 60861
rect 158920 60851 159000 60861
rect 159240 60851 159320 60861
rect 159560 60851 159640 60861
rect 146480 60771 146490 60851
rect 146800 60771 146810 60851
rect 147120 60771 147130 60851
rect 147440 60771 147450 60851
rect 148860 60771 148870 60851
rect 149180 60771 149190 60851
rect 149500 60771 149510 60851
rect 149820 60771 149830 60851
rect 152280 60771 152290 60851
rect 152600 60771 152610 60851
rect 152920 60771 152930 60851
rect 153240 60771 153250 60851
rect 153560 60771 153570 60851
rect 153880 60771 153890 60851
rect 154200 60771 154210 60851
rect 154520 60771 154530 60851
rect 154840 60771 154850 60851
rect 155160 60771 155170 60851
rect 155480 60771 155490 60851
rect 155800 60771 155810 60851
rect 156120 60771 156130 60851
rect 156440 60771 156450 60851
rect 156760 60771 156770 60851
rect 157080 60771 157090 60851
rect 157400 60771 157410 60851
rect 157720 60771 157730 60851
rect 158040 60771 158050 60851
rect 158360 60771 158370 60851
rect 158680 60771 158690 60851
rect 159000 60771 159010 60851
rect 159320 60771 159330 60851
rect 159640 60771 159650 60851
rect 163590 60821 163670 60831
rect 163910 60821 163990 60831
rect 164230 60821 164310 60831
rect 164550 60821 164630 60831
rect 164870 60821 164950 60831
rect 165190 60821 165270 60831
rect 165510 60821 165590 60831
rect 165830 60821 165910 60831
rect 166150 60821 166230 60831
rect 166470 60821 166550 60831
rect 166790 60821 166870 60831
rect 167110 60821 167190 60831
rect 167430 60821 167510 60831
rect 167750 60821 167830 60831
rect 168070 60821 168150 60831
rect 168390 60821 168470 60831
rect 168710 60821 168790 60831
rect 169030 60821 169110 60831
rect 169350 60821 169430 60831
rect 169670 60821 169750 60831
rect 169990 60821 170070 60831
rect 170310 60821 170390 60831
rect 170630 60821 170710 60831
rect 170950 60821 171030 60831
rect 163670 60741 163680 60821
rect 163990 60741 164000 60821
rect 164310 60741 164320 60821
rect 164630 60741 164640 60821
rect 164950 60741 164960 60821
rect 165270 60741 165280 60821
rect 165590 60741 165600 60821
rect 165910 60741 165920 60821
rect 166230 60741 166240 60821
rect 166550 60741 166560 60821
rect 166870 60741 166880 60821
rect 167190 60741 167200 60821
rect 167510 60741 167520 60821
rect 167830 60741 167840 60821
rect 168150 60741 168160 60821
rect 168470 60741 168480 60821
rect 168790 60741 168800 60821
rect 169110 60741 169120 60821
rect 169430 60741 169440 60821
rect 169750 60741 169760 60821
rect 170070 60741 170080 60821
rect 170390 60741 170400 60821
rect 170710 60741 170720 60821
rect 171030 60741 171040 60821
rect 30520 60700 30600 60710
rect 30840 60700 30920 60710
rect 31160 60700 31240 60710
rect 31480 60700 31560 60710
rect 31800 60700 31880 60710
rect 32120 60700 32200 60710
rect 32440 60700 32520 60710
rect 32760 60700 32840 60710
rect 33080 60700 33160 60710
rect 33400 60700 33480 60710
rect 33720 60700 33800 60710
rect 34040 60700 34120 60710
rect 34360 60700 34440 60710
rect 34680 60700 34760 60710
rect 35000 60700 35080 60710
rect 35320 60700 35400 60710
rect 35640 60700 35720 60710
rect 35960 60700 36040 60710
rect 36280 60700 36360 60710
rect 36600 60700 36680 60710
rect 36920 60700 37000 60710
rect 37240 60700 37320 60710
rect 37560 60700 37640 60710
rect 40340 60700 40420 60710
rect 40660 60700 40740 60710
rect 40980 60700 41060 60710
rect 42720 60700 42800 60710
rect 43040 60700 43120 60710
rect 43360 60700 43440 60710
rect 19130 60670 19210 60680
rect 19450 60670 19530 60680
rect 19770 60670 19850 60680
rect 20090 60670 20170 60680
rect 20410 60670 20490 60680
rect 20730 60670 20810 60680
rect 21050 60670 21130 60680
rect 21370 60670 21450 60680
rect 21690 60670 21770 60680
rect 22010 60670 22090 60680
rect 22330 60670 22410 60680
rect 22650 60670 22730 60680
rect 22970 60670 23050 60680
rect 23290 60670 23370 60680
rect 23610 60670 23690 60680
rect 23930 60670 24010 60680
rect 24250 60670 24330 60680
rect 24570 60670 24650 60680
rect 24890 60670 24970 60680
rect 25210 60670 25290 60680
rect 25530 60670 25610 60680
rect 25850 60670 25930 60680
rect 26170 60670 26250 60680
rect 19210 60590 19220 60670
rect 19530 60590 19540 60670
rect 19850 60590 19860 60670
rect 20170 60590 20180 60670
rect 20490 60590 20500 60670
rect 20810 60590 20820 60670
rect 21130 60590 21140 60670
rect 21450 60590 21460 60670
rect 21770 60590 21780 60670
rect 22090 60590 22100 60670
rect 22410 60590 22420 60670
rect 22730 60590 22740 60670
rect 23050 60590 23060 60670
rect 23370 60590 23380 60670
rect 23690 60590 23700 60670
rect 24010 60590 24020 60670
rect 24330 60590 24340 60670
rect 24650 60590 24660 60670
rect 24970 60590 24980 60670
rect 25290 60590 25300 60670
rect 25610 60590 25620 60670
rect 25930 60590 25940 60670
rect 26250 60590 26260 60670
rect 30600 60620 30610 60700
rect 30920 60620 30930 60700
rect 31240 60620 31250 60700
rect 31560 60620 31570 60700
rect 31880 60620 31890 60700
rect 32200 60620 32210 60700
rect 32520 60620 32530 60700
rect 32840 60620 32850 60700
rect 33160 60620 33170 60700
rect 33480 60620 33490 60700
rect 33800 60620 33810 60700
rect 34120 60620 34130 60700
rect 34440 60620 34450 60700
rect 34760 60620 34770 60700
rect 35080 60620 35090 60700
rect 35400 60620 35410 60700
rect 35720 60620 35730 60700
rect 36040 60620 36050 60700
rect 36360 60620 36370 60700
rect 36680 60620 36690 60700
rect 37000 60620 37010 60700
rect 37320 60620 37330 60700
rect 37640 60620 37650 60700
rect 40420 60620 40430 60700
rect 40740 60620 40750 60700
rect 41060 60620 41070 60700
rect 42800 60620 42810 60700
rect 43120 60620 43130 60700
rect 43440 60620 43450 60700
rect 146560 60691 146640 60701
rect 146880 60691 146960 60701
rect 147200 60691 147280 60701
rect 148940 60691 149020 60701
rect 149260 60691 149340 60701
rect 149580 60691 149660 60701
rect 152360 60691 152440 60701
rect 152680 60691 152760 60701
rect 153000 60691 153080 60701
rect 153320 60691 153400 60701
rect 153640 60691 153720 60701
rect 153960 60691 154040 60701
rect 154280 60691 154360 60701
rect 154600 60691 154680 60701
rect 154920 60691 155000 60701
rect 155240 60691 155320 60701
rect 155560 60691 155640 60701
rect 155880 60691 155960 60701
rect 156200 60691 156280 60701
rect 156520 60691 156600 60701
rect 156840 60691 156920 60701
rect 157160 60691 157240 60701
rect 157480 60691 157560 60701
rect 157800 60691 157880 60701
rect 158120 60691 158200 60701
rect 158440 60691 158520 60701
rect 158760 60691 158840 60701
rect 159080 60691 159160 60701
rect 159400 60691 159480 60701
rect 146640 60611 146650 60691
rect 146960 60611 146970 60691
rect 147280 60611 147290 60691
rect 149020 60611 149030 60691
rect 149340 60611 149350 60691
rect 149660 60611 149670 60691
rect 152440 60611 152450 60691
rect 152760 60611 152770 60691
rect 153080 60611 153090 60691
rect 153400 60611 153410 60691
rect 153720 60611 153730 60691
rect 154040 60611 154050 60691
rect 154360 60611 154370 60691
rect 154680 60611 154690 60691
rect 155000 60611 155010 60691
rect 155320 60611 155330 60691
rect 155640 60611 155650 60691
rect 155960 60611 155970 60691
rect 156280 60611 156290 60691
rect 156600 60611 156610 60691
rect 156920 60611 156930 60691
rect 157240 60611 157250 60691
rect 157560 60611 157570 60691
rect 157880 60611 157890 60691
rect 158200 60611 158210 60691
rect 158520 60611 158530 60691
rect 158840 60611 158850 60691
rect 159160 60611 159170 60691
rect 159480 60611 159490 60691
rect 163750 60661 163830 60671
rect 164070 60661 164150 60671
rect 164390 60661 164470 60671
rect 164710 60661 164790 60671
rect 165030 60661 165110 60671
rect 165350 60661 165430 60671
rect 165670 60661 165750 60671
rect 165990 60661 166070 60671
rect 166310 60661 166390 60671
rect 166630 60661 166710 60671
rect 166950 60661 167030 60671
rect 167270 60661 167350 60671
rect 167590 60661 167670 60671
rect 167910 60661 167990 60671
rect 168230 60661 168310 60671
rect 168550 60661 168630 60671
rect 168870 60661 168950 60671
rect 169190 60661 169270 60671
rect 169510 60661 169590 60671
rect 169830 60661 169910 60671
rect 170150 60661 170230 60671
rect 170470 60661 170550 60671
rect 170790 60661 170870 60671
rect 163830 60581 163840 60661
rect 164150 60581 164160 60661
rect 164470 60581 164480 60661
rect 164790 60581 164800 60661
rect 165110 60581 165120 60661
rect 165430 60581 165440 60661
rect 165750 60581 165760 60661
rect 166070 60581 166080 60661
rect 166390 60581 166400 60661
rect 166710 60581 166720 60661
rect 167030 60581 167040 60661
rect 167350 60581 167360 60661
rect 167670 60581 167680 60661
rect 167990 60581 168000 60661
rect 168310 60581 168320 60661
rect 168630 60581 168640 60661
rect 168950 60581 168960 60661
rect 169270 60581 169280 60661
rect 169590 60581 169600 60661
rect 169910 60581 169920 60661
rect 170230 60581 170240 60661
rect 170550 60581 170560 60661
rect 170870 60581 170880 60661
rect 18980 60440 19060 60450
rect 19160 60440 19240 60450
rect 19340 60440 19420 60450
rect 19520 60440 19600 60450
rect 19700 60440 19780 60450
rect 19880 60440 19960 60450
rect 20060 60440 20140 60450
rect 20240 60440 20320 60450
rect 20420 60440 20500 60450
rect 20600 60440 20680 60450
rect 20780 60440 20860 60450
rect 20960 60440 21040 60450
rect 21140 60440 21220 60450
rect 21320 60440 21400 60450
rect 21500 60440 21580 60450
rect 21680 60440 21760 60450
rect 21860 60440 21940 60450
rect 22040 60440 22120 60450
rect 22220 60440 22300 60450
rect 22400 60440 22480 60450
rect 22580 60440 22660 60450
rect 22760 60440 22840 60450
rect 22940 60440 23020 60450
rect 23120 60440 23200 60450
rect 23300 60440 23380 60450
rect 23480 60440 23560 60450
rect 23660 60440 23740 60450
rect 23840 60440 23920 60450
rect 24020 60440 24100 60450
rect 24200 60440 24280 60450
rect 24380 60440 24460 60450
rect 24560 60440 24640 60450
rect 24740 60440 24820 60450
rect 24920 60440 25000 60450
rect 25100 60440 25180 60450
rect 25280 60440 25360 60450
rect 25460 60440 25540 60450
rect 25640 60440 25720 60450
rect 25820 60440 25900 60450
rect 26000 60440 26080 60450
rect 26180 60440 26260 60450
rect 26360 60440 26440 60450
rect 26540 60440 26620 60450
rect 30280 60440 30360 60450
rect 30460 60440 30540 60450
rect 30640 60440 30720 60450
rect 30820 60440 30900 60450
rect 31000 60440 31080 60450
rect 31180 60440 31260 60450
rect 31360 60440 31440 60450
rect 31540 60440 31620 60450
rect 31720 60440 31800 60450
rect 31900 60440 31980 60450
rect 32080 60440 32160 60450
rect 32260 60440 32340 60450
rect 32440 60440 32520 60450
rect 32620 60440 32700 60450
rect 32800 60440 32880 60450
rect 32980 60440 33060 60450
rect 33160 60440 33240 60450
rect 33340 60440 33420 60450
rect 33520 60440 33600 60450
rect 33700 60440 33780 60450
rect 33880 60440 33960 60450
rect 34060 60440 34140 60450
rect 34240 60440 34320 60450
rect 34420 60440 34500 60450
rect 34600 60440 34680 60450
rect 34780 60440 34860 60450
rect 34960 60440 35040 60450
rect 35140 60440 35220 60450
rect 35320 60440 35400 60450
rect 35500 60440 35580 60450
rect 35680 60440 35760 60450
rect 35860 60440 35940 60450
rect 36040 60440 36120 60450
rect 36220 60440 36300 60450
rect 36400 60440 36480 60450
rect 36580 60440 36660 60450
rect 36760 60440 36840 60450
rect 36940 60440 37020 60450
rect 37120 60440 37200 60450
rect 37300 60440 37380 60450
rect 37480 60440 37560 60450
rect 37660 60440 37740 60450
rect 37840 60440 37920 60450
rect 40060 60440 40140 60450
rect 40200 60440 40280 60450
rect 40340 60440 40420 60450
rect 40480 60440 40560 60450
rect 40620 60440 40700 60450
rect 40760 60440 40840 60450
rect 40900 60440 40980 60450
rect 41040 60440 41120 60450
rect 41180 60440 41260 60450
rect 41320 60440 41400 60450
rect 42360 60440 42440 60450
rect 42500 60440 42580 60450
rect 42640 60440 42720 60450
rect 42780 60440 42860 60450
rect 42920 60440 43000 60450
rect 43060 60440 43140 60450
rect 43200 60440 43280 60450
rect 43340 60440 43420 60450
rect 43480 60440 43560 60450
rect 43620 60440 43700 60450
rect 146300 60440 146380 60450
rect 146440 60440 146520 60450
rect 146580 60440 146660 60450
rect 146720 60440 146800 60450
rect 146860 60440 146940 60450
rect 147000 60440 147080 60450
rect 147140 60440 147220 60450
rect 147280 60440 147360 60450
rect 147420 60440 147500 60450
rect 147560 60440 147640 60450
rect 148600 60440 148680 60450
rect 148740 60440 148820 60450
rect 148880 60440 148960 60450
rect 149020 60440 149100 60450
rect 149160 60440 149240 60450
rect 149300 60440 149380 60450
rect 149440 60440 149520 60450
rect 149580 60440 149660 60450
rect 149720 60440 149800 60450
rect 149860 60440 149940 60450
rect 152080 60440 152160 60450
rect 152260 60440 152340 60450
rect 152440 60440 152520 60450
rect 152620 60440 152700 60450
rect 152800 60440 152880 60450
rect 152980 60440 153060 60450
rect 153160 60440 153240 60450
rect 153340 60440 153420 60450
rect 153520 60440 153600 60450
rect 153700 60440 153780 60450
rect 153880 60440 153960 60450
rect 154060 60440 154140 60450
rect 154240 60440 154320 60450
rect 154420 60440 154500 60450
rect 154600 60440 154680 60450
rect 154780 60440 154860 60450
rect 154960 60440 155040 60450
rect 155140 60440 155220 60450
rect 155320 60440 155400 60450
rect 155500 60440 155580 60450
rect 155680 60440 155760 60450
rect 155860 60440 155940 60450
rect 156040 60440 156120 60450
rect 156220 60440 156300 60450
rect 156400 60440 156480 60450
rect 156580 60440 156660 60450
rect 156760 60440 156840 60450
rect 156940 60440 157020 60450
rect 157120 60440 157200 60450
rect 157300 60440 157380 60450
rect 157480 60440 157560 60450
rect 157660 60440 157740 60450
rect 157840 60440 157920 60450
rect 158020 60440 158100 60450
rect 158200 60440 158280 60450
rect 158380 60440 158460 60450
rect 158560 60440 158640 60450
rect 158740 60440 158820 60450
rect 158920 60440 159000 60450
rect 159100 60440 159180 60450
rect 159280 60440 159360 60450
rect 159460 60440 159540 60450
rect 159640 60440 159720 60450
rect 163380 60440 163460 60450
rect 163560 60440 163640 60450
rect 163740 60440 163820 60450
rect 163920 60440 164000 60450
rect 164100 60440 164180 60450
rect 164280 60440 164360 60450
rect 164460 60440 164540 60450
rect 164640 60440 164720 60450
rect 164820 60440 164900 60450
rect 165000 60440 165080 60450
rect 165180 60440 165260 60450
rect 165360 60440 165440 60450
rect 165540 60440 165620 60450
rect 165720 60440 165800 60450
rect 165900 60440 165980 60450
rect 166080 60440 166160 60450
rect 166260 60440 166340 60450
rect 166440 60440 166520 60450
rect 166620 60440 166700 60450
rect 166800 60440 166880 60450
rect 166980 60440 167060 60450
rect 167160 60440 167240 60450
rect 167340 60440 167420 60450
rect 167520 60440 167600 60450
rect 167700 60440 167780 60450
rect 167880 60440 167960 60450
rect 168060 60440 168140 60450
rect 168240 60440 168320 60450
rect 168420 60440 168500 60450
rect 168600 60440 168680 60450
rect 168780 60440 168860 60450
rect 168960 60440 169040 60450
rect 169140 60440 169220 60450
rect 169320 60440 169400 60450
rect 169500 60440 169580 60450
rect 169680 60440 169760 60450
rect 169860 60440 169940 60450
rect 170040 60440 170120 60450
rect 170220 60440 170300 60450
rect 170400 60440 170480 60450
rect 170580 60440 170660 60450
rect 170760 60440 170840 60450
rect 170940 60440 171020 60450
rect 19060 60360 19070 60440
rect 19240 60360 19250 60440
rect 19420 60360 19430 60440
rect 19600 60360 19610 60440
rect 19780 60360 19790 60440
rect 19960 60360 19970 60440
rect 20140 60360 20150 60440
rect 20320 60360 20330 60440
rect 20500 60360 20510 60440
rect 20680 60360 20690 60440
rect 20860 60360 20870 60440
rect 21040 60360 21050 60440
rect 21220 60360 21230 60440
rect 21400 60360 21410 60440
rect 21580 60360 21590 60440
rect 21760 60360 21770 60440
rect 21940 60360 21950 60440
rect 22120 60360 22130 60440
rect 22300 60360 22310 60440
rect 22480 60360 22490 60440
rect 22660 60360 22670 60440
rect 22840 60360 22850 60440
rect 23020 60360 23030 60440
rect 23200 60360 23210 60440
rect 23380 60360 23390 60440
rect 23560 60360 23570 60440
rect 23740 60360 23750 60440
rect 23920 60360 23930 60440
rect 24100 60360 24110 60440
rect 24280 60360 24290 60440
rect 24460 60360 24470 60440
rect 24640 60360 24650 60440
rect 24820 60360 24830 60440
rect 25000 60360 25010 60440
rect 25180 60360 25190 60440
rect 25360 60360 25370 60440
rect 25540 60360 25550 60440
rect 25720 60360 25730 60440
rect 25900 60360 25910 60440
rect 26080 60360 26090 60440
rect 26260 60360 26270 60440
rect 26440 60360 26450 60440
rect 26620 60360 26630 60440
rect 30360 60360 30370 60440
rect 30540 60360 30550 60440
rect 30720 60360 30730 60440
rect 30900 60360 30910 60440
rect 31080 60360 31090 60440
rect 31260 60360 31270 60440
rect 31440 60360 31450 60440
rect 31620 60360 31630 60440
rect 31800 60360 31810 60440
rect 31980 60360 31990 60440
rect 32160 60360 32170 60440
rect 32340 60360 32350 60440
rect 32520 60360 32530 60440
rect 32700 60360 32710 60440
rect 32880 60360 32890 60440
rect 33060 60360 33070 60440
rect 33240 60360 33250 60440
rect 33420 60360 33430 60440
rect 33600 60360 33610 60440
rect 33780 60360 33790 60440
rect 33960 60360 33970 60440
rect 34140 60360 34150 60440
rect 34320 60360 34330 60440
rect 34500 60360 34510 60440
rect 34680 60360 34690 60440
rect 34860 60360 34870 60440
rect 35040 60360 35050 60440
rect 35220 60360 35230 60440
rect 35400 60360 35410 60440
rect 35580 60360 35590 60440
rect 35760 60360 35770 60440
rect 35940 60360 35950 60440
rect 36120 60360 36130 60440
rect 36300 60360 36310 60440
rect 36480 60360 36490 60440
rect 36660 60360 36670 60440
rect 36840 60360 36850 60440
rect 37020 60360 37030 60440
rect 37200 60360 37210 60440
rect 37380 60360 37390 60440
rect 37560 60360 37570 60440
rect 37740 60360 37750 60440
rect 37920 60360 37930 60440
rect 40140 60360 40150 60440
rect 40280 60360 40290 60440
rect 40420 60360 40430 60440
rect 40560 60360 40570 60440
rect 40700 60360 40710 60440
rect 40840 60360 40850 60440
rect 40980 60360 40990 60440
rect 41120 60360 41130 60440
rect 41260 60360 41270 60440
rect 41400 60360 41410 60440
rect 42440 60360 42450 60440
rect 42580 60360 42590 60440
rect 42720 60360 42730 60440
rect 42860 60360 42870 60440
rect 43000 60360 43010 60440
rect 43140 60360 43150 60440
rect 43280 60360 43290 60440
rect 43420 60360 43430 60440
rect 43560 60360 43570 60440
rect 43700 60360 43710 60440
rect 146380 60360 146390 60440
rect 146520 60360 146530 60440
rect 146660 60360 146670 60440
rect 146800 60360 146810 60440
rect 146940 60360 146950 60440
rect 147080 60360 147090 60440
rect 147220 60360 147230 60440
rect 147360 60360 147370 60440
rect 147500 60360 147510 60440
rect 147640 60360 147650 60440
rect 148680 60360 148690 60440
rect 148820 60360 148830 60440
rect 148960 60360 148970 60440
rect 149100 60360 149110 60440
rect 149240 60360 149250 60440
rect 149380 60360 149390 60440
rect 149520 60360 149530 60440
rect 149660 60360 149670 60440
rect 149800 60360 149810 60440
rect 149940 60360 149950 60440
rect 152160 60360 152170 60440
rect 152340 60360 152350 60440
rect 152520 60360 152530 60440
rect 152700 60360 152710 60440
rect 152880 60360 152890 60440
rect 153060 60360 153070 60440
rect 153240 60360 153250 60440
rect 153420 60360 153430 60440
rect 153600 60360 153610 60440
rect 153780 60360 153790 60440
rect 153960 60360 153970 60440
rect 154140 60360 154150 60440
rect 154320 60360 154330 60440
rect 154500 60360 154510 60440
rect 154680 60360 154690 60440
rect 154860 60360 154870 60440
rect 155040 60360 155050 60440
rect 155220 60360 155230 60440
rect 155400 60360 155410 60440
rect 155580 60360 155590 60440
rect 155760 60360 155770 60440
rect 155940 60360 155950 60440
rect 156120 60360 156130 60440
rect 156300 60360 156310 60440
rect 156480 60360 156490 60440
rect 156660 60360 156670 60440
rect 156840 60360 156850 60440
rect 157020 60360 157030 60440
rect 157200 60360 157210 60440
rect 157380 60360 157390 60440
rect 157560 60360 157570 60440
rect 157740 60360 157750 60440
rect 157920 60360 157930 60440
rect 158100 60360 158110 60440
rect 158280 60360 158290 60440
rect 158460 60360 158470 60440
rect 158640 60360 158650 60440
rect 158820 60360 158830 60440
rect 159000 60360 159010 60440
rect 159180 60360 159190 60440
rect 159360 60360 159370 60440
rect 159540 60360 159550 60440
rect 159720 60360 159730 60440
rect 163460 60360 163470 60440
rect 163640 60360 163650 60440
rect 163820 60360 163830 60440
rect 164000 60360 164010 60440
rect 164180 60360 164190 60440
rect 164360 60360 164370 60440
rect 164540 60360 164550 60440
rect 164720 60360 164730 60440
rect 164900 60360 164910 60440
rect 165080 60360 165090 60440
rect 165260 60360 165270 60440
rect 165440 60360 165450 60440
rect 165620 60360 165630 60440
rect 165800 60360 165810 60440
rect 165980 60360 165990 60440
rect 166160 60360 166170 60440
rect 166340 60360 166350 60440
rect 166520 60360 166530 60440
rect 166700 60360 166710 60440
rect 166880 60360 166890 60440
rect 167060 60360 167070 60440
rect 167240 60360 167250 60440
rect 167420 60360 167430 60440
rect 167600 60360 167610 60440
rect 167780 60360 167790 60440
rect 167960 60360 167970 60440
rect 168140 60360 168150 60440
rect 168320 60360 168330 60440
rect 168500 60360 168510 60440
rect 168680 60360 168690 60440
rect 168860 60360 168870 60440
rect 169040 60360 169050 60440
rect 169220 60360 169230 60440
rect 169400 60360 169410 60440
rect 169580 60360 169590 60440
rect 169760 60360 169770 60440
rect 169940 60360 169950 60440
rect 170120 60360 170130 60440
rect 170300 60360 170310 60440
rect 170480 60360 170490 60440
rect 170660 60360 170670 60440
rect 170840 60360 170850 60440
rect 171020 60360 171030 60440
rect 161885 60345 161965 60355
rect 162065 60345 162145 60355
rect 162245 60345 162325 60355
rect 162425 60345 162505 60355
rect 162605 60345 162685 60355
rect 28850 60315 28930 60325
rect 29010 60315 29090 60325
rect 29170 60315 29250 60325
rect 29330 60315 29410 60325
rect 29490 60315 29570 60325
rect 18980 60290 19060 60300
rect 19160 60290 19240 60300
rect 19340 60290 19420 60300
rect 19520 60290 19600 60300
rect 19700 60290 19780 60300
rect 19880 60290 19960 60300
rect 20060 60290 20140 60300
rect 20240 60290 20320 60300
rect 20420 60290 20500 60300
rect 20600 60290 20680 60300
rect 20780 60290 20860 60300
rect 20960 60290 21040 60300
rect 21140 60290 21220 60300
rect 21320 60290 21400 60300
rect 21500 60290 21580 60300
rect 21680 60290 21760 60300
rect 21860 60290 21940 60300
rect 22040 60290 22120 60300
rect 22220 60290 22300 60300
rect 22400 60290 22480 60300
rect 22580 60290 22660 60300
rect 22760 60290 22840 60300
rect 22940 60290 23020 60300
rect 23120 60290 23200 60300
rect 23300 60290 23380 60300
rect 23480 60290 23560 60300
rect 23660 60290 23740 60300
rect 23840 60290 23920 60300
rect 24020 60290 24100 60300
rect 24200 60290 24280 60300
rect 24380 60290 24460 60300
rect 24560 60290 24640 60300
rect 24740 60290 24820 60300
rect 24920 60290 25000 60300
rect 25100 60290 25180 60300
rect 25280 60290 25360 60300
rect 25460 60290 25540 60300
rect 25640 60290 25720 60300
rect 25820 60290 25900 60300
rect 26000 60290 26080 60300
rect 26180 60290 26260 60300
rect 26360 60290 26440 60300
rect 26540 60290 26620 60300
rect 19060 60210 19070 60290
rect 19240 60210 19250 60290
rect 19420 60210 19430 60290
rect 19600 60210 19610 60290
rect 19780 60210 19790 60290
rect 19960 60210 19970 60290
rect 20140 60210 20150 60290
rect 20320 60210 20330 60290
rect 20500 60210 20510 60290
rect 20680 60210 20690 60290
rect 20860 60210 20870 60290
rect 21040 60210 21050 60290
rect 21220 60210 21230 60290
rect 21400 60210 21410 60290
rect 21580 60210 21590 60290
rect 21760 60210 21770 60290
rect 21940 60210 21950 60290
rect 22120 60210 22130 60290
rect 22300 60210 22310 60290
rect 22480 60210 22490 60290
rect 22660 60210 22670 60290
rect 22840 60210 22850 60290
rect 23020 60210 23030 60290
rect 23200 60210 23210 60290
rect 23380 60210 23390 60290
rect 23560 60210 23570 60290
rect 23740 60210 23750 60290
rect 23920 60210 23930 60290
rect 24100 60210 24110 60290
rect 24280 60210 24290 60290
rect 24460 60210 24470 60290
rect 24640 60210 24650 60290
rect 24820 60210 24830 60290
rect 25000 60210 25010 60290
rect 25180 60210 25190 60290
rect 25360 60210 25370 60290
rect 25540 60210 25550 60290
rect 25720 60210 25730 60290
rect 25900 60210 25910 60290
rect 26080 60210 26090 60290
rect 26260 60210 26270 60290
rect 26440 60210 26450 60290
rect 26620 60210 26630 60290
rect 28930 60235 28940 60315
rect 29010 60235 29020 60315
rect 29090 60235 29100 60315
rect 29170 60235 29180 60315
rect 29250 60235 29260 60315
rect 29330 60235 29340 60315
rect 29410 60235 29420 60315
rect 29490 60235 29500 60315
rect 29570 60235 29580 60315
rect 30280 60290 30360 60300
rect 30460 60290 30540 60300
rect 30640 60290 30720 60300
rect 30820 60290 30900 60300
rect 31000 60290 31080 60300
rect 31180 60290 31260 60300
rect 31360 60290 31440 60300
rect 31540 60290 31620 60300
rect 31720 60290 31800 60300
rect 31900 60290 31980 60300
rect 32080 60290 32160 60300
rect 32260 60290 32340 60300
rect 32440 60290 32520 60300
rect 32620 60290 32700 60300
rect 32800 60290 32880 60300
rect 32980 60290 33060 60300
rect 33160 60290 33240 60300
rect 33340 60290 33420 60300
rect 33520 60290 33600 60300
rect 33700 60290 33780 60300
rect 33880 60290 33960 60300
rect 34060 60290 34140 60300
rect 34240 60290 34320 60300
rect 34420 60290 34500 60300
rect 34600 60290 34680 60300
rect 34780 60290 34860 60300
rect 34960 60290 35040 60300
rect 35140 60290 35220 60300
rect 35320 60290 35400 60300
rect 35500 60290 35580 60300
rect 35680 60290 35760 60300
rect 35860 60290 35940 60300
rect 36040 60290 36120 60300
rect 36220 60290 36300 60300
rect 36400 60290 36480 60300
rect 36580 60290 36660 60300
rect 36760 60290 36840 60300
rect 36940 60290 37020 60300
rect 37120 60290 37200 60300
rect 37300 60290 37380 60300
rect 37480 60290 37560 60300
rect 37660 60290 37740 60300
rect 37840 60290 37920 60300
rect 152080 60290 152160 60300
rect 152260 60290 152340 60300
rect 152440 60290 152520 60300
rect 152620 60290 152700 60300
rect 152800 60290 152880 60300
rect 152980 60290 153060 60300
rect 153160 60290 153240 60300
rect 153340 60290 153420 60300
rect 153520 60290 153600 60300
rect 153700 60290 153780 60300
rect 153880 60290 153960 60300
rect 154060 60290 154140 60300
rect 154240 60290 154320 60300
rect 154420 60290 154500 60300
rect 154600 60290 154680 60300
rect 154780 60290 154860 60300
rect 154960 60290 155040 60300
rect 155140 60290 155220 60300
rect 155320 60290 155400 60300
rect 155500 60290 155580 60300
rect 155680 60290 155760 60300
rect 155860 60290 155940 60300
rect 156040 60290 156120 60300
rect 156220 60290 156300 60300
rect 156400 60290 156480 60300
rect 156580 60290 156660 60300
rect 156760 60290 156840 60300
rect 156940 60290 157020 60300
rect 157120 60290 157200 60300
rect 157300 60290 157380 60300
rect 157480 60290 157560 60300
rect 157660 60290 157740 60300
rect 157840 60290 157920 60300
rect 158020 60290 158100 60300
rect 158200 60290 158280 60300
rect 158380 60290 158460 60300
rect 158560 60290 158640 60300
rect 158740 60290 158820 60300
rect 158920 60290 159000 60300
rect 159100 60290 159180 60300
rect 159280 60290 159360 60300
rect 159460 60290 159540 60300
rect 159640 60290 159720 60300
rect 30360 60210 30370 60290
rect 30540 60210 30550 60290
rect 30720 60210 30730 60290
rect 30900 60210 30910 60290
rect 31080 60210 31090 60290
rect 31260 60210 31270 60290
rect 31440 60210 31450 60290
rect 31620 60210 31630 60290
rect 31800 60210 31810 60290
rect 31980 60210 31990 60290
rect 32160 60210 32170 60290
rect 32340 60210 32350 60290
rect 32520 60210 32530 60290
rect 32700 60210 32710 60290
rect 32880 60210 32890 60290
rect 33060 60210 33070 60290
rect 33240 60210 33250 60290
rect 33420 60210 33430 60290
rect 33600 60210 33610 60290
rect 33780 60210 33790 60290
rect 33960 60210 33970 60290
rect 34140 60210 34150 60290
rect 34320 60210 34330 60290
rect 34500 60210 34510 60290
rect 34680 60210 34690 60290
rect 34860 60210 34870 60290
rect 35040 60210 35050 60290
rect 35220 60210 35230 60290
rect 35400 60210 35410 60290
rect 35580 60210 35590 60290
rect 35760 60210 35770 60290
rect 35940 60210 35950 60290
rect 36120 60210 36130 60290
rect 36300 60210 36310 60290
rect 36480 60210 36490 60290
rect 36660 60210 36670 60290
rect 36840 60210 36850 60290
rect 37020 60210 37030 60290
rect 37200 60210 37210 60290
rect 37380 60210 37390 60290
rect 37560 60210 37570 60290
rect 37740 60210 37750 60290
rect 37920 60210 37930 60290
rect 40060 60190 40120 60220
rect 41540 60190 41600 60220
rect 42360 60190 42420 60220
rect 43840 60190 43900 60220
rect 152160 60210 152170 60290
rect 152340 60210 152350 60290
rect 152520 60210 152530 60290
rect 152700 60210 152710 60290
rect 152880 60210 152890 60290
rect 153060 60210 153070 60290
rect 153240 60210 153250 60290
rect 153420 60210 153430 60290
rect 153600 60210 153610 60290
rect 153780 60210 153790 60290
rect 153960 60210 153970 60290
rect 154140 60210 154150 60290
rect 154320 60210 154330 60290
rect 154500 60210 154510 60290
rect 154680 60210 154690 60290
rect 154860 60210 154870 60290
rect 155040 60210 155050 60290
rect 155220 60210 155230 60290
rect 155400 60210 155410 60290
rect 155580 60210 155590 60290
rect 155760 60210 155770 60290
rect 155940 60210 155950 60290
rect 156120 60210 156130 60290
rect 156300 60210 156310 60290
rect 156480 60210 156490 60290
rect 156660 60210 156670 60290
rect 156840 60210 156850 60290
rect 157020 60210 157030 60290
rect 157200 60210 157210 60290
rect 157380 60210 157390 60290
rect 157560 60210 157570 60290
rect 157740 60210 157750 60290
rect 157920 60210 157930 60290
rect 158100 60210 158110 60290
rect 158280 60210 158290 60290
rect 158460 60210 158470 60290
rect 158640 60210 158650 60290
rect 158820 60210 158830 60290
rect 159000 60210 159010 60290
rect 159180 60210 159190 60290
rect 159360 60210 159370 60290
rect 159540 60210 159550 60290
rect 159720 60210 159730 60290
rect 161965 60265 161975 60345
rect 162145 60265 162155 60345
rect 162325 60265 162335 60345
rect 162505 60265 162515 60345
rect 162685 60265 162695 60345
rect 163380 60290 163460 60300
rect 163560 60290 163640 60300
rect 163740 60290 163820 60300
rect 163920 60290 164000 60300
rect 164100 60290 164180 60300
rect 164280 60290 164360 60300
rect 164460 60290 164540 60300
rect 164640 60290 164720 60300
rect 164820 60290 164900 60300
rect 165000 60290 165080 60300
rect 165180 60290 165260 60300
rect 165360 60290 165440 60300
rect 165540 60290 165620 60300
rect 165720 60290 165800 60300
rect 165900 60290 165980 60300
rect 166080 60290 166160 60300
rect 166260 60290 166340 60300
rect 166440 60290 166520 60300
rect 166620 60290 166700 60300
rect 166800 60290 166880 60300
rect 166980 60290 167060 60300
rect 167160 60290 167240 60300
rect 167340 60290 167420 60300
rect 167520 60290 167600 60300
rect 167700 60290 167780 60300
rect 167880 60290 167960 60300
rect 168060 60290 168140 60300
rect 168240 60290 168320 60300
rect 168420 60290 168500 60300
rect 168600 60290 168680 60300
rect 168780 60290 168860 60300
rect 168960 60290 169040 60300
rect 169140 60290 169220 60300
rect 169320 60290 169400 60300
rect 169500 60290 169580 60300
rect 169680 60290 169760 60300
rect 169860 60290 169940 60300
rect 170040 60290 170120 60300
rect 170220 60290 170300 60300
rect 170400 60290 170480 60300
rect 170580 60290 170660 60300
rect 170760 60290 170840 60300
rect 170940 60290 171020 60300
rect 163460 60210 163470 60290
rect 163640 60210 163650 60290
rect 163820 60210 163830 60290
rect 164000 60210 164010 60290
rect 164180 60210 164190 60290
rect 164360 60210 164370 60290
rect 164540 60210 164550 60290
rect 164720 60210 164730 60290
rect 164900 60210 164910 60290
rect 165080 60210 165090 60290
rect 165260 60210 165270 60290
rect 165440 60210 165450 60290
rect 165620 60210 165630 60290
rect 165800 60210 165810 60290
rect 165980 60210 165990 60290
rect 166160 60210 166170 60290
rect 166340 60210 166350 60290
rect 166520 60210 166530 60290
rect 166700 60210 166710 60290
rect 166880 60210 166890 60290
rect 167060 60210 167070 60290
rect 167240 60210 167250 60290
rect 167420 60210 167430 60290
rect 167600 60210 167610 60290
rect 167780 60210 167790 60290
rect 167960 60210 167970 60290
rect 168140 60210 168150 60290
rect 168320 60210 168330 60290
rect 168500 60210 168510 60290
rect 168680 60210 168690 60290
rect 168860 60210 168870 60290
rect 169040 60210 169050 60290
rect 169220 60210 169230 60290
rect 169400 60210 169410 60290
rect 169580 60210 169590 60290
rect 169760 60210 169770 60290
rect 169940 60210 169950 60290
rect 170120 60210 170130 60290
rect 170300 60210 170310 60290
rect 170480 60210 170490 60290
rect 170660 60210 170670 60290
rect 170840 60210 170850 60290
rect 171020 60210 171030 60290
rect 146100 60150 146160 60180
rect 147580 60150 147640 60180
rect 148400 60150 148460 60180
rect 149880 60150 149940 60180
rect 161885 60165 161965 60175
rect 162065 60165 162145 60175
rect 162245 60165 162325 60175
rect 162425 60165 162505 60175
rect 162605 60165 162685 60175
rect 40060 60070 40120 60100
rect 41540 60070 41600 60100
rect 42360 60070 42420 60100
rect 43840 60070 43900 60100
rect 146100 60030 146160 60060
rect 146210 60040 146220 60130
rect 40060 59950 40120 59980
rect 41540 59950 41600 59980
rect 42360 59950 42420 59980
rect 43840 59950 43900 59980
rect 19130 59910 19160 59940
rect 19250 59910 19280 59940
rect 26420 59910 26450 59940
rect 26540 59910 26570 59940
rect 30420 59910 30450 59940
rect 30540 59910 30570 59940
rect 37720 59910 37750 59940
rect 37840 59910 37870 59940
rect 146100 59910 146160 59940
rect 19010 59880 19070 59910
rect 19130 59880 19190 59910
rect 19250 59880 19310 59910
rect 26300 59880 26360 59910
rect 26420 59880 26480 59910
rect 26540 59880 26600 59910
rect 30300 59880 30360 59910
rect 30420 59880 30480 59910
rect 30540 59880 30600 59910
rect 37600 59880 37660 59910
rect 37720 59880 37780 59910
rect 37840 59880 37900 59910
rect 40060 59830 40120 59860
rect 41540 59830 41600 59860
rect 42360 59830 42420 59860
rect 43840 59830 43900 59860
rect 19130 59790 19160 59820
rect 19250 59790 19280 59820
rect 26420 59790 26450 59820
rect 26540 59790 26570 59820
rect 30420 59790 30450 59820
rect 30540 59790 30570 59820
rect 37720 59790 37750 59820
rect 37840 59790 37870 59820
rect 146100 59790 146160 59820
rect 19010 59760 19070 59790
rect 19130 59760 19190 59790
rect 19250 59760 19310 59790
rect 26300 59760 26360 59790
rect 26420 59760 26480 59790
rect 26540 59760 26600 59790
rect 30300 59760 30360 59790
rect 30420 59760 30480 59790
rect 30540 59760 30600 59790
rect 37600 59760 37660 59790
rect 37720 59760 37780 59790
rect 37840 59760 37900 59790
rect 19880 59730 19960 59740
rect 20060 59730 20140 59740
rect 20240 59730 20320 59740
rect 20420 59730 20500 59740
rect 20600 59730 20680 59740
rect 20780 59730 20860 59740
rect 20960 59730 21040 59740
rect 21140 59730 21220 59740
rect 21320 59730 21400 59740
rect 21500 59730 21580 59740
rect 21680 59730 21760 59740
rect 21860 59730 21940 59740
rect 22040 59730 22120 59740
rect 22220 59730 22300 59740
rect 22400 59730 22480 59740
rect 22580 59730 22660 59740
rect 22760 59730 22840 59740
rect 22940 59730 23020 59740
rect 23120 59730 23200 59740
rect 23300 59730 23380 59740
rect 23480 59730 23560 59740
rect 23660 59730 23740 59740
rect 23840 59730 23920 59740
rect 24020 59730 24100 59740
rect 24200 59730 24280 59740
rect 24380 59730 24460 59740
rect 24560 59730 24640 59740
rect 24740 59730 24820 59740
rect 24920 59730 25000 59740
rect 25100 59730 25180 59740
rect 25280 59730 25360 59740
rect 25460 59730 25540 59740
rect 25640 59730 25720 59740
rect 19130 59670 19160 59700
rect 19250 59670 19280 59700
rect 19010 59640 19070 59670
rect 19130 59640 19190 59670
rect 19250 59640 19310 59670
rect 19960 59650 19970 59730
rect 20140 59650 20150 59730
rect 20320 59650 20330 59730
rect 20500 59650 20510 59730
rect 20680 59650 20690 59730
rect 20860 59650 20870 59730
rect 21040 59650 21050 59730
rect 21220 59650 21230 59730
rect 21400 59650 21410 59730
rect 21580 59650 21590 59730
rect 21760 59650 21770 59730
rect 21940 59650 21950 59730
rect 22120 59650 22130 59730
rect 22300 59650 22310 59730
rect 22480 59650 22490 59730
rect 22660 59650 22670 59730
rect 22840 59650 22850 59730
rect 23020 59650 23030 59730
rect 23200 59650 23210 59730
rect 23380 59650 23390 59730
rect 23560 59650 23570 59730
rect 23740 59650 23750 59730
rect 23920 59650 23930 59730
rect 24100 59650 24110 59730
rect 24280 59650 24290 59730
rect 24460 59650 24470 59730
rect 24640 59650 24650 59730
rect 24820 59650 24830 59730
rect 25000 59650 25010 59730
rect 25180 59650 25190 59730
rect 25360 59650 25370 59730
rect 25540 59650 25550 59730
rect 25720 59650 25730 59730
rect 26420 59670 26450 59700
rect 26540 59670 26570 59700
rect 30420 59670 30450 59700
rect 30540 59670 30570 59700
rect 31010 59670 37190 59760
rect 40060 59710 40120 59740
rect 41540 59710 41600 59740
rect 42360 59710 42420 59740
rect 43840 59710 43900 59740
rect 37720 59670 37750 59700
rect 37840 59670 37870 59700
rect 146100 59670 146160 59700
rect 26300 59640 26360 59670
rect 26420 59640 26480 59670
rect 26540 59640 26600 59670
rect 30300 59640 30360 59670
rect 30420 59640 30480 59670
rect 30540 59640 30600 59670
rect 31260 59650 31270 59670
rect 31440 59650 31450 59670
rect 31620 59650 31630 59670
rect 31800 59650 31810 59670
rect 31980 59650 31990 59670
rect 32160 59650 32170 59670
rect 32340 59650 32350 59670
rect 32520 59650 32530 59670
rect 32700 59650 32710 59670
rect 32880 59650 32890 59670
rect 33060 59650 33070 59670
rect 33240 59650 33250 59670
rect 33420 59650 33430 59670
rect 33600 59650 33610 59670
rect 33780 59650 33790 59670
rect 33960 59650 33970 59670
rect 34140 59650 34150 59670
rect 34320 59650 34330 59670
rect 34500 59650 34510 59670
rect 34680 59650 34690 59670
rect 34860 59650 34870 59670
rect 35040 59650 35050 59670
rect 35220 59650 35230 59670
rect 35400 59650 35410 59670
rect 35580 59650 35590 59670
rect 35760 59650 35770 59670
rect 35940 59650 35950 59670
rect 36120 59650 36130 59670
rect 36300 59650 36310 59670
rect 36480 59650 36490 59670
rect 36660 59650 36670 59670
rect 36840 59650 36850 59670
rect 37020 59650 37030 59670
rect 19880 59580 19960 59590
rect 20060 59580 20140 59590
rect 20240 59580 20320 59590
rect 20420 59580 20500 59590
rect 20600 59580 20680 59590
rect 20780 59580 20860 59590
rect 20960 59580 21040 59590
rect 21140 59580 21220 59590
rect 21320 59580 21400 59590
rect 21500 59580 21580 59590
rect 21680 59580 21760 59590
rect 21860 59580 21940 59590
rect 22040 59580 22120 59590
rect 22220 59580 22300 59590
rect 22400 59580 22480 59590
rect 22580 59580 22660 59590
rect 22760 59580 22840 59590
rect 22940 59580 23020 59590
rect 23120 59580 23200 59590
rect 23300 59580 23380 59590
rect 23480 59580 23560 59590
rect 23660 59580 23740 59590
rect 23840 59580 23920 59590
rect 24020 59580 24100 59590
rect 24200 59580 24280 59590
rect 24380 59580 24460 59590
rect 24560 59580 24640 59590
rect 24740 59580 24820 59590
rect 24920 59580 25000 59590
rect 25100 59580 25180 59590
rect 25280 59580 25360 59590
rect 25460 59580 25540 59590
rect 25640 59580 25720 59590
rect 31180 59580 31260 59590
rect 31360 59580 31440 59590
rect 31540 59580 31620 59590
rect 31720 59580 31800 59590
rect 31900 59580 31980 59590
rect 32080 59580 32160 59590
rect 32260 59580 32340 59590
rect 32440 59580 32520 59590
rect 32620 59580 32700 59590
rect 32800 59580 32880 59590
rect 32980 59580 33060 59590
rect 33160 59580 33240 59590
rect 33340 59580 33420 59590
rect 33520 59580 33600 59590
rect 33700 59580 33780 59590
rect 33880 59580 33960 59590
rect 34060 59580 34140 59590
rect 34240 59580 34320 59590
rect 34420 59580 34500 59590
rect 34600 59580 34680 59590
rect 34780 59580 34860 59590
rect 34960 59580 35040 59590
rect 35140 59580 35220 59590
rect 35320 59580 35400 59590
rect 35500 59580 35580 59590
rect 35680 59580 35760 59590
rect 35860 59580 35940 59590
rect 36040 59580 36120 59590
rect 36220 59580 36300 59590
rect 36400 59580 36480 59590
rect 36580 59580 36660 59590
rect 36760 59580 36840 59590
rect 36940 59580 37020 59590
rect 19130 59550 19160 59580
rect 19250 59550 19280 59580
rect 19010 59520 19070 59550
rect 19130 59520 19190 59550
rect 19250 59520 19310 59550
rect 19960 59500 19970 59580
rect 20140 59500 20150 59580
rect 20320 59500 20330 59580
rect 20500 59500 20510 59580
rect 20680 59500 20690 59580
rect 20860 59500 20870 59580
rect 21040 59500 21050 59580
rect 21220 59500 21230 59580
rect 21400 59500 21410 59580
rect 21580 59500 21590 59580
rect 21760 59500 21770 59580
rect 21940 59500 21950 59580
rect 22120 59500 22130 59580
rect 22300 59500 22310 59580
rect 22480 59500 22490 59580
rect 22660 59500 22670 59580
rect 22840 59500 22850 59580
rect 23020 59500 23030 59580
rect 23200 59500 23210 59580
rect 23380 59500 23390 59580
rect 23560 59500 23570 59580
rect 23740 59500 23750 59580
rect 23920 59500 23930 59580
rect 24100 59500 24110 59580
rect 24280 59500 24290 59580
rect 24460 59500 24470 59580
rect 24640 59500 24650 59580
rect 24820 59500 24830 59580
rect 25000 59500 25010 59580
rect 25180 59500 25190 59580
rect 25360 59500 25370 59580
rect 25540 59500 25550 59580
rect 25720 59500 25730 59580
rect 26420 59550 26450 59580
rect 26540 59550 26570 59580
rect 30420 59550 30450 59580
rect 30540 59550 30570 59580
rect 26300 59520 26360 59550
rect 26420 59520 26480 59550
rect 26540 59520 26600 59550
rect 30300 59520 30360 59550
rect 30420 59520 30480 59550
rect 30540 59520 30600 59550
rect 31260 59500 31270 59580
rect 31440 59500 31450 59580
rect 31620 59500 31630 59580
rect 31800 59500 31810 59580
rect 31980 59500 31990 59580
rect 32160 59500 32170 59580
rect 32340 59500 32350 59580
rect 32520 59500 32530 59580
rect 32700 59500 32710 59580
rect 32880 59500 32890 59580
rect 33060 59500 33070 59580
rect 33240 59500 33250 59580
rect 33420 59500 33430 59580
rect 33600 59500 33610 59580
rect 33780 59500 33790 59580
rect 33960 59500 33970 59580
rect 34140 59500 34150 59580
rect 34320 59500 34330 59580
rect 34500 59500 34510 59580
rect 34680 59500 34690 59580
rect 34860 59500 34870 59580
rect 35040 59500 35050 59580
rect 35220 59500 35230 59580
rect 35400 59500 35410 59580
rect 35580 59500 35590 59580
rect 35760 59500 35770 59580
rect 35940 59500 35950 59580
rect 36120 59500 36130 59580
rect 36300 59500 36310 59580
rect 36480 59500 36490 59580
rect 36660 59500 36670 59580
rect 36840 59500 36850 59580
rect 37020 59500 37030 59580
rect 19130 59430 19160 59460
rect 19250 59430 19280 59460
rect 19880 59430 19960 59440
rect 20060 59430 20140 59440
rect 20240 59430 20320 59440
rect 20420 59430 20500 59440
rect 20600 59430 20680 59440
rect 20780 59430 20860 59440
rect 20960 59430 21040 59440
rect 21140 59430 21220 59440
rect 21320 59430 21400 59440
rect 21500 59430 21580 59440
rect 21680 59430 21760 59440
rect 21860 59430 21940 59440
rect 22040 59430 22120 59440
rect 22220 59430 22300 59440
rect 22400 59430 22480 59440
rect 22580 59430 22660 59440
rect 22760 59430 22840 59440
rect 22940 59430 23020 59440
rect 23120 59430 23200 59440
rect 23300 59430 23380 59440
rect 23480 59430 23560 59440
rect 23660 59430 23740 59440
rect 23840 59430 23920 59440
rect 24020 59430 24100 59440
rect 24200 59430 24280 59440
rect 24380 59430 24460 59440
rect 24560 59430 24640 59440
rect 24740 59430 24820 59440
rect 24920 59430 25000 59440
rect 25100 59430 25180 59440
rect 25280 59430 25360 59440
rect 25460 59430 25540 59440
rect 25640 59430 25720 59440
rect 26420 59430 26450 59460
rect 26540 59430 26570 59460
rect 30420 59430 30450 59460
rect 30540 59430 30570 59460
rect 37100 59440 37190 59670
rect 37600 59640 37660 59670
rect 37720 59640 37780 59670
rect 37840 59640 37900 59670
rect 40060 59590 40120 59620
rect 41540 59590 41600 59620
rect 42360 59590 42420 59620
rect 43840 59590 43900 59620
rect 37720 59550 37750 59580
rect 37840 59550 37870 59580
rect 146100 59550 146160 59580
rect 37600 59520 37660 59550
rect 37720 59520 37780 59550
rect 37840 59520 37900 59550
rect 40060 59470 40120 59500
rect 41540 59470 41600 59500
rect 42360 59470 42420 59500
rect 43840 59470 43900 59500
rect 19010 59400 19070 59430
rect 19130 59400 19190 59430
rect 19250 59400 19310 59430
rect 19960 59350 19970 59430
rect 20140 59350 20150 59430
rect 20320 59350 20330 59430
rect 20500 59350 20510 59430
rect 20680 59350 20690 59430
rect 20860 59350 20870 59430
rect 21040 59350 21050 59430
rect 21220 59350 21230 59430
rect 21400 59350 21410 59430
rect 21580 59350 21590 59430
rect 21760 59350 21770 59430
rect 21940 59350 21950 59430
rect 22120 59350 22130 59430
rect 22300 59350 22310 59430
rect 22480 59350 22490 59430
rect 22660 59350 22670 59430
rect 22840 59350 22850 59430
rect 23020 59350 23030 59430
rect 23200 59350 23210 59430
rect 23380 59350 23390 59430
rect 23560 59350 23570 59430
rect 23740 59350 23750 59430
rect 23920 59350 23930 59430
rect 24100 59350 24110 59430
rect 24280 59350 24290 59430
rect 24460 59350 24470 59430
rect 24640 59350 24650 59430
rect 24820 59350 24830 59430
rect 25000 59350 25010 59430
rect 25180 59350 25190 59430
rect 25360 59350 25370 59430
rect 25540 59350 25550 59430
rect 25720 59350 25730 59430
rect 26300 59400 26360 59430
rect 26420 59400 26480 59430
rect 26540 59400 26600 59430
rect 30300 59400 30360 59430
rect 30420 59400 30480 59430
rect 30540 59400 30600 59430
rect 31100 59410 37190 59440
rect 37720 59430 37750 59460
rect 37840 59430 37870 59460
rect 146100 59430 146160 59460
rect 31260 59350 31270 59410
rect 31440 59350 31450 59410
rect 31620 59350 31630 59410
rect 31800 59350 31810 59410
rect 31980 59350 31990 59410
rect 32160 59350 32170 59410
rect 32340 59350 32350 59410
rect 32520 59350 32530 59410
rect 32700 59350 32710 59410
rect 32880 59350 32890 59410
rect 33060 59350 33070 59410
rect 33240 59350 33250 59410
rect 33420 59350 33430 59410
rect 33600 59350 33610 59410
rect 33780 59350 33790 59410
rect 33960 59350 33970 59410
rect 34140 59350 34150 59410
rect 34320 59350 34330 59410
rect 34500 59350 34510 59410
rect 34680 59350 34690 59410
rect 34860 59350 34870 59410
rect 35040 59350 35050 59410
rect 35220 59350 35230 59410
rect 35400 59350 35410 59410
rect 35580 59350 35590 59410
rect 35760 59350 35770 59410
rect 35940 59350 35950 59410
rect 36120 59350 36130 59410
rect 36300 59350 36310 59410
rect 36480 59350 36490 59410
rect 36660 59350 36670 59410
rect 36840 59350 36850 59410
rect 37020 59350 37030 59410
rect 37100 59340 37190 59410
rect 37600 59400 37660 59430
rect 37720 59400 37780 59430
rect 37840 59400 37900 59430
rect 40060 59350 40120 59380
rect 41540 59350 41600 59380
rect 42360 59350 42420 59380
rect 43840 59350 43900 59380
rect 19130 59310 19160 59340
rect 19250 59310 19280 59340
rect 26420 59310 26450 59340
rect 26540 59310 26570 59340
rect 30420 59310 30450 59340
rect 30540 59310 30570 59340
rect 31100 59310 37190 59340
rect 37720 59310 37750 59340
rect 37840 59310 37870 59340
rect 146100 59310 146160 59340
rect 19010 59280 19070 59310
rect 19130 59280 19190 59310
rect 19250 59280 19310 59310
rect 19800 59290 25800 59300
rect 26300 59280 26360 59310
rect 26420 59280 26480 59310
rect 26540 59280 26600 59310
rect 30300 59280 30360 59310
rect 30420 59280 30480 59310
rect 30540 59280 30600 59310
rect 37100 59300 37190 59310
rect 31100 59290 37190 59300
rect 19130 59190 19160 59220
rect 19250 59190 19280 59220
rect 26420 59190 26450 59220
rect 26540 59190 26570 59220
rect 30420 59190 30450 59220
rect 30540 59190 30570 59220
rect 19010 59160 19070 59190
rect 19130 59160 19190 59190
rect 19250 59160 19310 59190
rect 26300 59160 26360 59190
rect 26420 59160 26480 59190
rect 26540 59160 26600 59190
rect 30300 59160 30360 59190
rect 30420 59160 30480 59190
rect 30540 59160 30600 59190
rect 31180 59110 31260 59120
rect 31360 59110 31440 59120
rect 31540 59110 31620 59120
rect 31720 59110 31800 59120
rect 31900 59110 31980 59120
rect 32080 59110 32160 59120
rect 32260 59110 32340 59120
rect 32440 59110 32520 59120
rect 32620 59110 32700 59120
rect 32800 59110 32880 59120
rect 32980 59110 33060 59120
rect 33160 59110 33240 59120
rect 33340 59110 33420 59120
rect 33520 59110 33600 59120
rect 33700 59110 33780 59120
rect 33880 59110 33960 59120
rect 34060 59110 34140 59120
rect 34240 59110 34320 59120
rect 34420 59110 34500 59120
rect 34600 59110 34680 59120
rect 34780 59110 34860 59120
rect 34960 59110 35040 59120
rect 35140 59110 35220 59120
rect 35320 59110 35400 59120
rect 35500 59110 35580 59120
rect 35680 59110 35760 59120
rect 35860 59110 35940 59120
rect 36040 59110 36120 59120
rect 36220 59110 36300 59120
rect 36400 59110 36480 59120
rect 36580 59110 36660 59120
rect 36760 59110 36840 59120
rect 36940 59110 37020 59120
rect 19130 59070 19160 59100
rect 19250 59070 19280 59100
rect 19880 59090 19960 59100
rect 20060 59090 20140 59100
rect 20240 59090 20320 59100
rect 20420 59090 20500 59100
rect 20600 59090 20680 59100
rect 20780 59090 20860 59100
rect 20960 59090 21040 59100
rect 21140 59090 21220 59100
rect 21320 59090 21400 59100
rect 21500 59090 21580 59100
rect 21680 59090 21760 59100
rect 21860 59090 21940 59100
rect 22040 59090 22120 59100
rect 22220 59090 22300 59100
rect 22400 59090 22480 59100
rect 22580 59090 22660 59100
rect 22760 59090 22840 59100
rect 22940 59090 23020 59100
rect 23120 59090 23200 59100
rect 23300 59090 23380 59100
rect 23480 59090 23560 59100
rect 23660 59090 23740 59100
rect 23840 59090 23920 59100
rect 24020 59090 24100 59100
rect 24200 59090 24280 59100
rect 24380 59090 24460 59100
rect 24560 59090 24640 59100
rect 24740 59090 24820 59100
rect 24920 59090 25000 59100
rect 25100 59090 25180 59100
rect 25280 59090 25360 59100
rect 25460 59090 25540 59100
rect 25640 59090 25720 59100
rect 19010 59040 19070 59070
rect 19130 59040 19190 59070
rect 19250 59040 19310 59070
rect 19960 59010 19970 59090
rect 20140 59010 20150 59090
rect 20320 59010 20330 59090
rect 20500 59010 20510 59090
rect 20680 59010 20690 59090
rect 20860 59010 20870 59090
rect 21040 59010 21050 59090
rect 21220 59010 21230 59090
rect 21400 59010 21410 59090
rect 21580 59010 21590 59090
rect 21760 59010 21770 59090
rect 21940 59010 21950 59090
rect 22120 59010 22130 59090
rect 22300 59010 22310 59090
rect 22480 59010 22490 59090
rect 22660 59010 22670 59090
rect 22840 59010 22850 59090
rect 23020 59010 23030 59090
rect 23200 59010 23210 59090
rect 23380 59010 23390 59090
rect 23560 59010 23570 59090
rect 23740 59010 23750 59090
rect 23920 59010 23930 59090
rect 24100 59010 24110 59090
rect 24280 59010 24290 59090
rect 24460 59010 24470 59090
rect 24640 59010 24650 59090
rect 24820 59010 24830 59090
rect 25000 59010 25010 59090
rect 25180 59010 25190 59090
rect 25360 59010 25370 59090
rect 25540 59010 25550 59090
rect 25720 59010 25730 59090
rect 26420 59070 26450 59100
rect 26540 59070 26570 59100
rect 30420 59070 30450 59100
rect 30540 59070 30570 59100
rect 26300 59040 26360 59070
rect 26420 59040 26480 59070
rect 26540 59040 26600 59070
rect 30300 59040 30360 59070
rect 30420 59040 30480 59070
rect 30540 59040 30600 59070
rect 31260 59030 31270 59110
rect 31440 59030 31450 59110
rect 31620 59030 31630 59110
rect 31800 59030 31810 59110
rect 31980 59030 31990 59110
rect 32160 59030 32170 59110
rect 32340 59030 32350 59110
rect 32520 59030 32530 59110
rect 32700 59030 32710 59110
rect 32880 59030 32890 59110
rect 33060 59030 33070 59110
rect 33240 59030 33250 59110
rect 33420 59030 33430 59110
rect 33600 59030 33610 59110
rect 33780 59030 33790 59110
rect 33960 59030 33970 59110
rect 34140 59030 34150 59110
rect 34320 59030 34330 59110
rect 34500 59030 34510 59110
rect 34680 59030 34690 59110
rect 34860 59030 34870 59110
rect 35040 59030 35050 59110
rect 35220 59030 35230 59110
rect 35400 59030 35410 59110
rect 35580 59030 35590 59110
rect 35760 59030 35770 59110
rect 35940 59030 35950 59110
rect 36120 59030 36130 59110
rect 36300 59030 36310 59110
rect 36480 59030 36490 59110
rect 36660 59030 36670 59110
rect 36840 59030 36850 59110
rect 37020 59030 37030 59110
rect 19130 58950 19160 58980
rect 19250 58950 19280 58980
rect 26420 58950 26450 58980
rect 26540 58950 26570 58980
rect 30420 58950 30450 58980
rect 30540 58950 30570 58980
rect 19010 58920 19070 58950
rect 19130 58920 19190 58950
rect 19250 58920 19310 58950
rect 26300 58920 26360 58950
rect 26420 58920 26480 58950
rect 26540 58920 26600 58950
rect 30300 58920 30360 58950
rect 30420 58920 30480 58950
rect 30540 58920 30600 58950
rect 19130 58830 19160 58860
rect 19250 58830 19280 58860
rect 26420 58830 26450 58860
rect 26540 58830 26570 58860
rect 30420 58830 30450 58860
rect 30540 58830 30570 58860
rect 19010 58800 19070 58830
rect 19130 58800 19190 58830
rect 19250 58800 19310 58830
rect 26300 58800 26360 58830
rect 26420 58800 26480 58830
rect 26540 58800 26600 58830
rect 30300 58800 30360 58830
rect 30420 58800 30480 58830
rect 30540 58800 30600 58830
rect 19880 58790 19960 58800
rect 20060 58790 20140 58800
rect 20240 58790 20320 58800
rect 20420 58790 20500 58800
rect 20600 58790 20680 58800
rect 20780 58790 20860 58800
rect 20960 58790 21040 58800
rect 21140 58790 21220 58800
rect 21320 58790 21400 58800
rect 21500 58790 21580 58800
rect 21680 58790 21760 58800
rect 21860 58790 21940 58800
rect 22040 58790 22120 58800
rect 22220 58790 22300 58800
rect 22400 58790 22480 58800
rect 22580 58790 22660 58800
rect 22760 58790 22840 58800
rect 22940 58790 23020 58800
rect 23120 58790 23200 58800
rect 23300 58790 23380 58800
rect 23480 58790 23560 58800
rect 23660 58790 23740 58800
rect 23840 58790 23920 58800
rect 24020 58790 24100 58800
rect 24200 58790 24280 58800
rect 24380 58790 24460 58800
rect 24560 58790 24640 58800
rect 24740 58790 24820 58800
rect 24920 58790 25000 58800
rect 25100 58790 25180 58800
rect 25280 58790 25360 58800
rect 25460 58790 25540 58800
rect 25640 58790 25720 58800
rect 31180 58790 31260 58800
rect 31360 58790 31440 58800
rect 31540 58790 31620 58800
rect 31720 58790 31800 58800
rect 31900 58790 31980 58800
rect 32080 58790 32160 58800
rect 32260 58790 32340 58800
rect 32440 58790 32520 58800
rect 32620 58790 32700 58800
rect 32800 58790 32880 58800
rect 32980 58790 33060 58800
rect 33160 58790 33240 58800
rect 33340 58790 33420 58800
rect 33520 58790 33600 58800
rect 33700 58790 33780 58800
rect 33880 58790 33960 58800
rect 34060 58790 34140 58800
rect 34240 58790 34320 58800
rect 34420 58790 34500 58800
rect 34600 58790 34680 58800
rect 34780 58790 34860 58800
rect 34960 58790 35040 58800
rect 35140 58790 35220 58800
rect 35320 58790 35400 58800
rect 35500 58790 35580 58800
rect 35680 58790 35760 58800
rect 35860 58790 35940 58800
rect 36040 58790 36120 58800
rect 36220 58790 36300 58800
rect 36400 58790 36480 58800
rect 36580 58790 36660 58800
rect 36760 58790 36840 58800
rect 36940 58790 37020 58800
rect 19130 58710 19160 58740
rect 19250 58710 19280 58740
rect 19960 58710 19970 58790
rect 20140 58710 20150 58790
rect 20320 58710 20330 58790
rect 20500 58710 20510 58790
rect 20680 58710 20690 58790
rect 20860 58710 20870 58790
rect 21040 58710 21050 58790
rect 21220 58710 21230 58790
rect 21400 58710 21410 58790
rect 21580 58710 21590 58790
rect 21760 58710 21770 58790
rect 21940 58710 21950 58790
rect 22120 58710 22130 58790
rect 22300 58710 22310 58790
rect 22480 58710 22490 58790
rect 22660 58710 22670 58790
rect 22840 58710 22850 58790
rect 23020 58710 23030 58790
rect 23200 58710 23210 58790
rect 23380 58710 23390 58790
rect 23560 58710 23570 58790
rect 23740 58710 23750 58790
rect 23920 58710 23930 58790
rect 24100 58710 24110 58790
rect 24280 58710 24290 58790
rect 24460 58710 24470 58790
rect 24640 58710 24650 58790
rect 24820 58710 24830 58790
rect 25000 58710 25010 58790
rect 25180 58710 25190 58790
rect 25360 58710 25370 58790
rect 25540 58710 25550 58790
rect 25720 58710 25730 58790
rect 26420 58710 26450 58740
rect 26540 58710 26570 58740
rect 30420 58710 30450 58740
rect 30540 58710 30570 58740
rect 31260 58710 31270 58790
rect 31440 58710 31450 58790
rect 31620 58710 31630 58790
rect 31800 58710 31810 58790
rect 31980 58710 31990 58790
rect 32160 58710 32170 58790
rect 32340 58710 32350 58790
rect 32520 58710 32530 58790
rect 32700 58710 32710 58790
rect 32880 58710 32890 58790
rect 33060 58710 33070 58790
rect 33240 58710 33250 58790
rect 33420 58710 33430 58790
rect 33600 58710 33610 58790
rect 33780 58710 33790 58790
rect 33960 58710 33970 58790
rect 34140 58710 34150 58790
rect 34320 58710 34330 58790
rect 34500 58710 34510 58790
rect 34680 58710 34690 58790
rect 34860 58710 34870 58790
rect 35040 58710 35050 58790
rect 35220 58710 35230 58790
rect 35400 58710 35410 58790
rect 35580 58710 35590 58790
rect 35760 58710 35770 58790
rect 35940 58710 35950 58790
rect 36120 58710 36130 58790
rect 36300 58710 36310 58790
rect 36480 58710 36490 58790
rect 36660 58710 36670 58790
rect 36840 58710 36850 58790
rect 37020 58710 37030 58790
rect 19010 58680 19070 58710
rect 19130 58680 19190 58710
rect 19250 58680 19310 58710
rect 26300 58680 26360 58710
rect 26420 58680 26480 58710
rect 26540 58680 26600 58710
rect 30300 58680 30360 58710
rect 30420 58680 30480 58710
rect 30540 58680 30600 58710
rect 37100 58620 37190 59290
rect 37600 59280 37660 59310
rect 37720 59280 37780 59310
rect 37840 59280 37900 59310
rect 40060 59230 40120 59260
rect 41540 59230 41600 59260
rect 42360 59230 42420 59260
rect 43840 59230 43900 59260
rect 37720 59190 37750 59220
rect 37840 59190 37870 59220
rect 146100 59190 146160 59220
rect 37600 59160 37660 59190
rect 37720 59160 37780 59190
rect 37840 59160 37900 59190
rect 40060 59110 40120 59140
rect 41540 59110 41600 59140
rect 42360 59110 42420 59140
rect 43840 59110 43900 59140
rect 37720 59070 37750 59100
rect 37840 59070 37870 59100
rect 146100 59070 146160 59100
rect 37600 59040 37660 59070
rect 37720 59040 37780 59070
rect 37840 59040 37900 59070
rect 40060 58990 40120 59020
rect 41540 58990 41600 59020
rect 42360 58990 42420 59020
rect 43840 58990 43900 59020
rect 37720 58950 37750 58980
rect 37840 58950 37870 58980
rect 146100 58950 146160 58980
rect 37600 58920 37660 58950
rect 37720 58920 37780 58950
rect 37840 58920 37900 58950
rect 40060 58870 40120 58900
rect 41540 58870 41600 58900
rect 42360 58870 42420 58900
rect 43840 58870 43900 58900
rect 37720 58830 37750 58860
rect 37840 58830 37870 58860
rect 146100 58830 146160 58860
rect 37600 58800 37660 58830
rect 37720 58800 37780 58830
rect 37840 58800 37900 58830
rect 40060 58750 40120 58780
rect 41540 58750 41600 58780
rect 42360 58750 42420 58780
rect 43840 58750 43900 58780
rect 37720 58710 37750 58740
rect 37840 58710 37870 58740
rect 146100 58710 146160 58740
rect 37600 58680 37660 58710
rect 37720 58680 37780 58710
rect 37840 58680 37900 58710
rect 40060 58630 40120 58660
rect 41540 58630 41600 58660
rect 42360 58630 42420 58660
rect 43840 58630 43900 58660
rect 146300 58650 146310 60040
rect 146690 60000 146810 60060
rect 146970 60000 147090 60060
rect 147580 60030 147640 60060
rect 148400 60030 148460 60060
rect 148820 60050 149620 60140
rect 148950 60020 149070 60050
rect 149230 60020 149350 60050
rect 149070 60010 149130 60020
rect 149350 60010 149410 60020
rect 149070 60000 149190 60010
rect 149350 60000 149470 60010
rect 146810 59990 146870 60000
rect 146570 59980 146650 59990
rect 146810 59980 146930 59990
rect 146650 59900 146660 59980
rect 146810 59880 146870 59980
rect 146930 59900 146940 59980
rect 147090 59880 147150 60000
rect 146410 59830 147140 59840
rect 146410 59750 146420 59830
rect 147220 59825 147230 59880
rect 147270 59850 147390 59910
rect 146460 59815 147250 59825
rect 146450 59765 146460 59815
rect 146500 59560 146510 59750
rect 146690 59700 146810 59760
rect 146970 59700 147090 59760
rect 146810 59690 146870 59700
rect 146570 59680 146650 59690
rect 146710 59680 146790 59690
rect 146810 59680 146930 59690
rect 146990 59680 147070 59690
rect 146650 59600 146660 59680
rect 146790 59600 146800 59680
rect 146810 59580 146870 59680
rect 146930 59600 146940 59680
rect 147070 59600 147080 59680
rect 147090 59580 147150 59700
rect 146500 59550 147130 59560
rect 146500 59540 146510 59550
rect 146690 59410 146810 59470
rect 146970 59410 147090 59470
rect 146690 59320 146700 59410
rect 146800 59380 146870 59410
rect 146810 59290 146870 59380
rect 146970 59320 146980 59410
rect 147090 59290 147150 59410
rect 146410 59240 147140 59250
rect 146410 59160 146420 59240
rect 147220 59235 147230 59815
rect 147390 59730 147450 59850
rect 147300 59620 147380 59630
rect 147380 59540 147390 59620
rect 147300 59440 147380 59450
rect 147380 59360 147390 59440
rect 147270 59260 147390 59320
rect 146460 59225 147250 59235
rect 146450 59175 146460 59225
rect 146500 58970 146510 59160
rect 146690 59110 146810 59170
rect 146970 59110 147090 59170
rect 146810 59100 146870 59110
rect 146570 59090 146650 59100
rect 146710 59090 146790 59100
rect 146810 59090 146930 59100
rect 146990 59090 147070 59100
rect 146650 59010 146660 59090
rect 146790 59010 146800 59090
rect 146810 58990 146870 59090
rect 146930 59010 146940 59090
rect 147070 59010 147080 59090
rect 147090 58990 147150 59110
rect 146500 58960 147130 58970
rect 146500 58950 146510 58960
rect 146690 58820 146810 58880
rect 146970 58820 147090 58880
rect 146690 58730 146700 58820
rect 146800 58790 146870 58820
rect 146810 58700 146870 58790
rect 146970 58730 146980 58820
rect 147090 58700 147150 58820
rect 146410 58650 147140 58660
rect 147220 58645 147230 59225
rect 147390 59140 147450 59260
rect 147300 59020 147380 59030
rect 147380 58940 147390 59020
rect 147300 58840 147380 58850
rect 147380 58760 147390 58840
rect 147270 58670 147390 58730
rect 146460 58635 147250 58645
rect 19130 58590 19160 58620
rect 19250 58590 19280 58620
rect 19800 58610 25800 58620
rect 26420 58590 26450 58620
rect 26540 58590 26570 58620
rect 30420 58590 30450 58620
rect 30540 58590 30570 58620
rect 31100 58610 37190 58620
rect 19010 58560 19070 58590
rect 19130 58560 19190 58590
rect 19250 58560 19310 58590
rect 26300 58560 26360 58590
rect 26420 58560 26480 58590
rect 26540 58560 26600 58590
rect 30300 58560 30360 58590
rect 30420 58560 30480 58590
rect 30540 58560 30600 58590
rect 37100 58510 37190 58610
rect 37720 58590 37750 58620
rect 37840 58590 37870 58620
rect 146100 58590 146160 58620
rect 37600 58560 37660 58590
rect 37720 58560 37780 58590
rect 37840 58560 37900 58590
rect 146450 58585 146460 58635
rect 40060 58510 40120 58540
rect 41540 58510 41600 58540
rect 42360 58510 42420 58540
rect 43840 58510 43900 58540
rect 19130 58470 19160 58500
rect 19250 58470 19280 58500
rect 19880 58470 19960 58480
rect 20060 58470 20140 58480
rect 20240 58470 20320 58480
rect 20420 58470 20500 58480
rect 20600 58470 20680 58480
rect 20780 58470 20860 58480
rect 20960 58470 21040 58480
rect 21140 58470 21220 58480
rect 21320 58470 21400 58480
rect 21500 58470 21580 58480
rect 21680 58470 21760 58480
rect 21860 58470 21940 58480
rect 22040 58470 22120 58480
rect 22220 58470 22300 58480
rect 22400 58470 22480 58480
rect 22580 58470 22660 58480
rect 22760 58470 22840 58480
rect 22940 58470 23020 58480
rect 23120 58470 23200 58480
rect 23300 58470 23380 58480
rect 23480 58470 23560 58480
rect 23660 58470 23740 58480
rect 23840 58470 23920 58480
rect 24020 58470 24100 58480
rect 24200 58470 24280 58480
rect 24380 58470 24460 58480
rect 24560 58470 24640 58480
rect 24740 58470 24820 58480
rect 24920 58470 25000 58480
rect 25100 58470 25180 58480
rect 25280 58470 25360 58480
rect 25460 58470 25540 58480
rect 25640 58470 25720 58480
rect 26420 58470 26450 58500
rect 26540 58470 26570 58500
rect 30420 58470 30450 58500
rect 30540 58470 30570 58500
rect 31100 58480 37190 58510
rect 31180 58470 31260 58480
rect 31360 58470 31440 58480
rect 31540 58470 31620 58480
rect 31720 58470 31800 58480
rect 31900 58470 31980 58480
rect 32080 58470 32160 58480
rect 32260 58470 32340 58480
rect 32440 58470 32520 58480
rect 32620 58470 32700 58480
rect 32800 58470 32880 58480
rect 32980 58470 33060 58480
rect 33160 58470 33240 58480
rect 33340 58470 33420 58480
rect 33520 58470 33600 58480
rect 33700 58470 33780 58480
rect 33880 58470 33960 58480
rect 34060 58470 34140 58480
rect 34240 58470 34320 58480
rect 34420 58470 34500 58480
rect 34600 58470 34680 58480
rect 34780 58470 34860 58480
rect 34960 58470 35040 58480
rect 35140 58470 35220 58480
rect 35320 58470 35400 58480
rect 35500 58470 35580 58480
rect 35680 58470 35760 58480
rect 35860 58470 35940 58480
rect 36040 58470 36120 58480
rect 36220 58470 36300 58480
rect 36400 58470 36480 58480
rect 36580 58470 36660 58480
rect 36760 58470 36840 58480
rect 36940 58470 37020 58480
rect 19010 58440 19070 58470
rect 19130 58440 19190 58470
rect 19250 58440 19310 58470
rect 19960 58390 19970 58470
rect 20140 58390 20150 58470
rect 20320 58390 20330 58470
rect 20500 58390 20510 58470
rect 20680 58390 20690 58470
rect 20860 58390 20870 58470
rect 21040 58390 21050 58470
rect 21220 58390 21230 58470
rect 21400 58390 21410 58470
rect 21580 58390 21590 58470
rect 21760 58390 21770 58470
rect 21940 58390 21950 58470
rect 22120 58390 22130 58470
rect 22300 58390 22310 58470
rect 22480 58390 22490 58470
rect 22660 58390 22670 58470
rect 22840 58390 22850 58470
rect 23020 58390 23030 58470
rect 23200 58390 23210 58470
rect 23380 58390 23390 58470
rect 23560 58390 23570 58470
rect 23740 58390 23750 58470
rect 23920 58390 23930 58470
rect 24100 58390 24110 58470
rect 24280 58390 24290 58470
rect 24460 58390 24470 58470
rect 24640 58390 24650 58470
rect 24820 58390 24830 58470
rect 25000 58390 25010 58470
rect 25180 58390 25190 58470
rect 25360 58390 25370 58470
rect 25540 58390 25550 58470
rect 25720 58390 25730 58470
rect 26300 58440 26360 58470
rect 26420 58440 26480 58470
rect 26540 58440 26600 58470
rect 30300 58440 30360 58470
rect 30420 58440 30480 58470
rect 30540 58440 30600 58470
rect 31260 58410 31270 58470
rect 31440 58410 31450 58470
rect 31620 58410 31630 58470
rect 31800 58410 31810 58470
rect 31980 58410 31990 58470
rect 32160 58410 32170 58470
rect 32340 58410 32350 58470
rect 32520 58410 32530 58470
rect 32700 58410 32710 58470
rect 32880 58410 32890 58470
rect 33060 58410 33070 58470
rect 33240 58410 33250 58470
rect 33420 58410 33430 58470
rect 33600 58410 33610 58470
rect 33780 58410 33790 58470
rect 33960 58410 33970 58470
rect 34140 58410 34150 58470
rect 34320 58410 34330 58470
rect 34500 58410 34510 58470
rect 34680 58410 34690 58470
rect 34860 58410 34870 58470
rect 35040 58410 35050 58470
rect 35220 58410 35230 58470
rect 35400 58410 35410 58470
rect 35580 58410 35590 58470
rect 35760 58410 35770 58470
rect 35940 58410 35950 58470
rect 36120 58410 36130 58470
rect 36300 58410 36310 58470
rect 36480 58410 36490 58470
rect 36660 58410 36670 58470
rect 36840 58410 36850 58470
rect 37020 58410 37030 58470
rect 37100 58410 37190 58480
rect 37720 58470 37750 58500
rect 37840 58470 37870 58500
rect 37600 58440 37660 58470
rect 37720 58440 37780 58470
rect 37840 58440 37900 58470
rect 31100 58380 37190 58410
rect 40060 58390 40120 58420
rect 41540 58390 41600 58420
rect 42360 58390 42420 58420
rect 43840 58390 43900 58420
rect 19130 58350 19160 58380
rect 19250 58350 19280 58380
rect 26420 58350 26450 58380
rect 26540 58350 26570 58380
rect 30420 58350 30450 58380
rect 30540 58350 30570 58380
rect 19010 58320 19070 58350
rect 19130 58320 19190 58350
rect 19250 58320 19310 58350
rect 19880 58320 19960 58330
rect 20060 58320 20140 58330
rect 20240 58320 20320 58330
rect 20420 58320 20500 58330
rect 20600 58320 20680 58330
rect 20780 58320 20860 58330
rect 20960 58320 21040 58330
rect 21140 58320 21220 58330
rect 21320 58320 21400 58330
rect 21500 58320 21580 58330
rect 21680 58320 21760 58330
rect 21860 58320 21940 58330
rect 22040 58320 22120 58330
rect 22220 58320 22300 58330
rect 22400 58320 22480 58330
rect 22580 58320 22660 58330
rect 22760 58320 22840 58330
rect 22940 58320 23020 58330
rect 23120 58320 23200 58330
rect 23300 58320 23380 58330
rect 23480 58320 23560 58330
rect 23660 58320 23740 58330
rect 23840 58320 23920 58330
rect 24020 58320 24100 58330
rect 24200 58320 24280 58330
rect 24380 58320 24460 58330
rect 24560 58320 24640 58330
rect 24740 58320 24820 58330
rect 24920 58320 25000 58330
rect 25100 58320 25180 58330
rect 25280 58320 25360 58330
rect 25460 58320 25540 58330
rect 25640 58320 25720 58330
rect 26300 58320 26360 58350
rect 26420 58320 26480 58350
rect 26540 58320 26600 58350
rect 30300 58320 30360 58350
rect 30420 58320 30480 58350
rect 30540 58320 30600 58350
rect 31180 58320 31260 58330
rect 31360 58320 31440 58330
rect 31540 58320 31620 58330
rect 31720 58320 31800 58330
rect 31900 58320 31980 58330
rect 32080 58320 32160 58330
rect 32260 58320 32340 58330
rect 32440 58320 32520 58330
rect 32620 58320 32700 58330
rect 32800 58320 32880 58330
rect 32980 58320 33060 58330
rect 33160 58320 33240 58330
rect 33340 58320 33420 58330
rect 33520 58320 33600 58330
rect 33700 58320 33780 58330
rect 33880 58320 33960 58330
rect 34060 58320 34140 58330
rect 34240 58320 34320 58330
rect 34420 58320 34500 58330
rect 34600 58320 34680 58330
rect 34780 58320 34860 58330
rect 34960 58320 35040 58330
rect 35140 58320 35220 58330
rect 35320 58320 35400 58330
rect 35500 58320 35580 58330
rect 35680 58320 35760 58330
rect 35860 58320 35940 58330
rect 36040 58320 36120 58330
rect 36220 58320 36300 58330
rect 36400 58320 36480 58330
rect 36580 58320 36660 58330
rect 36760 58320 36840 58330
rect 36940 58320 37020 58330
rect 19130 58230 19160 58260
rect 19250 58230 19280 58260
rect 19960 58240 19970 58320
rect 20140 58240 20150 58320
rect 20320 58240 20330 58320
rect 20500 58240 20510 58320
rect 20680 58240 20690 58320
rect 20860 58240 20870 58320
rect 21040 58240 21050 58320
rect 21220 58240 21230 58320
rect 21400 58240 21410 58320
rect 21580 58240 21590 58320
rect 21760 58240 21770 58320
rect 21940 58240 21950 58320
rect 22120 58240 22130 58320
rect 22300 58240 22310 58320
rect 22480 58240 22490 58320
rect 22660 58240 22670 58320
rect 22840 58240 22850 58320
rect 23020 58240 23030 58320
rect 23200 58240 23210 58320
rect 23380 58240 23390 58320
rect 23560 58240 23570 58320
rect 23740 58240 23750 58320
rect 23920 58240 23930 58320
rect 24100 58240 24110 58320
rect 24280 58240 24290 58320
rect 24460 58240 24470 58320
rect 24640 58240 24650 58320
rect 24820 58240 24830 58320
rect 25000 58240 25010 58320
rect 25180 58240 25190 58320
rect 25360 58240 25370 58320
rect 25540 58240 25550 58320
rect 25720 58240 25730 58320
rect 26420 58230 26450 58260
rect 26540 58230 26570 58260
rect 30420 58230 30450 58260
rect 30540 58230 30570 58260
rect 31260 58240 31270 58320
rect 31440 58240 31450 58320
rect 31620 58240 31630 58320
rect 31800 58240 31810 58320
rect 31980 58240 31990 58320
rect 32160 58240 32170 58320
rect 32340 58240 32350 58320
rect 32520 58240 32530 58320
rect 32700 58240 32710 58320
rect 32880 58240 32890 58320
rect 33060 58240 33070 58320
rect 33240 58240 33250 58320
rect 33420 58240 33430 58320
rect 33600 58240 33610 58320
rect 33780 58240 33790 58320
rect 33960 58240 33970 58320
rect 34140 58240 34150 58320
rect 34320 58240 34330 58320
rect 34500 58240 34510 58320
rect 34680 58240 34690 58320
rect 34860 58240 34870 58320
rect 35040 58240 35050 58320
rect 35220 58240 35230 58320
rect 35400 58240 35410 58320
rect 35580 58240 35590 58320
rect 35760 58240 35770 58320
rect 35940 58240 35950 58320
rect 36120 58240 36130 58320
rect 36300 58240 36310 58320
rect 36480 58240 36490 58320
rect 36660 58240 36670 58320
rect 36840 58240 36850 58320
rect 37020 58240 37030 58320
rect 19010 58200 19070 58230
rect 19130 58200 19190 58230
rect 19250 58200 19310 58230
rect 26300 58200 26360 58230
rect 26420 58200 26480 58230
rect 26540 58200 26600 58230
rect 30300 58200 30360 58230
rect 30420 58200 30480 58230
rect 30540 58200 30600 58230
rect 37100 58180 37190 58380
rect 37720 58350 37750 58380
rect 37840 58350 37870 58380
rect 146690 58520 146810 58580
rect 146970 58520 147090 58580
rect 147220 58520 147230 58635
rect 147390 58550 147450 58670
rect 147520 58520 147530 59970
rect 147580 59910 147640 59940
rect 148400 59910 148460 59940
rect 148510 59900 148520 59990
rect 147580 59790 147640 59820
rect 148400 59790 148460 59820
rect 147580 59670 147640 59700
rect 148400 59670 148460 59700
rect 147580 59550 147640 59580
rect 148400 59550 148460 59580
rect 147580 59430 147640 59460
rect 148400 59430 148460 59460
rect 147580 59310 147640 59340
rect 148400 59310 148460 59340
rect 147580 59190 147640 59220
rect 148400 59190 148460 59220
rect 147580 59070 147640 59100
rect 148400 59070 148460 59100
rect 147580 58950 147640 58980
rect 148400 58950 148460 58980
rect 147580 58830 147640 58860
rect 148400 58830 148460 58860
rect 147580 58710 147640 58740
rect 148400 58710 148460 58740
rect 147580 58590 147640 58620
rect 148400 58590 148460 58620
rect 146810 58510 146870 58520
rect 146570 58500 146650 58510
rect 146710 58500 146790 58510
rect 146810 58500 146930 58510
rect 146990 58500 147070 58510
rect 146100 58470 146160 58500
rect 146650 58420 146660 58500
rect 146790 58420 146800 58500
rect 146810 58400 146870 58500
rect 146930 58420 146940 58500
rect 147070 58420 147080 58500
rect 147090 58400 147150 58520
rect 147580 58470 147640 58500
rect 148400 58470 148460 58500
rect 146100 58350 146160 58380
rect 147580 58350 147640 58380
rect 148400 58350 148460 58380
rect 37600 58320 37660 58350
rect 37720 58320 37780 58350
rect 37840 58320 37900 58350
rect 40060 58270 40120 58300
rect 41540 58270 41600 58300
rect 42360 58270 42420 58300
rect 43840 58270 43900 58300
rect 37720 58230 37750 58260
rect 37840 58230 37870 58260
rect 146100 58230 146160 58260
rect 147580 58230 147640 58260
rect 148400 58230 148460 58260
rect 37600 58200 37660 58230
rect 37720 58200 37780 58230
rect 37840 58200 37900 58230
rect 148600 58220 148610 59900
rect 148650 59870 148770 59930
rect 149070 59900 149130 60000
rect 149190 59920 149200 60000
rect 149350 59900 149410 60000
rect 149470 59920 149480 60000
rect 148770 59845 148830 59870
rect 149530 59865 149620 60050
rect 148910 59860 149620 59865
rect 148900 59850 149630 59860
rect 148910 59845 149630 59850
rect 148770 59835 149630 59845
rect 148770 59750 148830 59835
rect 149530 59785 149630 59835
rect 148910 59755 149630 59785
rect 148950 59720 149070 59755
rect 149230 59720 149350 59755
rect 148660 59710 148740 59720
rect 149070 59710 149130 59720
rect 149350 59710 149410 59720
rect 148740 59630 148750 59710
rect 148970 59700 149050 59710
rect 149070 59700 149190 59710
rect 149250 59700 149330 59710
rect 149350 59700 149470 59710
rect 148650 59570 148770 59630
rect 149050 59620 149060 59700
rect 149070 59600 149130 59700
rect 149190 59620 149200 59700
rect 149330 59620 149340 59700
rect 149350 59600 149410 59700
rect 149470 59620 149480 59700
rect 148770 59545 148830 59570
rect 149530 59565 149630 59755
rect 148910 59550 149630 59565
rect 148910 59545 149620 59550
rect 148770 59535 149620 59545
rect 148770 59450 148830 59535
rect 149530 59485 149620 59535
rect 148910 59455 149620 59485
rect 148950 59420 149070 59455
rect 149230 59420 149350 59455
rect 148660 59400 148740 59410
rect 148740 59330 148750 59400
rect 149060 59390 149130 59420
rect 148650 59270 148770 59330
rect 149070 59300 149130 59390
rect 149230 59330 149240 59420
rect 149340 59390 149410 59420
rect 149350 59300 149410 59390
rect 148770 59245 148830 59270
rect 149530 59265 149620 59455
rect 148910 59260 149620 59265
rect 148900 59250 149630 59260
rect 148910 59245 149630 59250
rect 148770 59235 149630 59245
rect 148770 59150 148830 59235
rect 149530 59185 149630 59235
rect 148910 59155 149630 59185
rect 148950 59120 149070 59155
rect 149230 59120 149350 59155
rect 149070 59110 149130 59120
rect 149350 59110 149410 59120
rect 148660 59100 148740 59110
rect 148970 59100 149050 59110
rect 149070 59100 149190 59110
rect 149250 59100 149330 59110
rect 149350 59100 149470 59110
rect 148740 59030 148750 59100
rect 148650 58970 148770 59030
rect 149050 59020 149060 59100
rect 149070 59000 149130 59100
rect 149190 59020 149200 59100
rect 149330 59020 149340 59100
rect 149350 59000 149410 59100
rect 149470 59020 149480 59100
rect 148770 58945 148830 58970
rect 149530 58965 149630 59155
rect 148910 58950 149630 58965
rect 148910 58945 149620 58950
rect 148770 58935 149620 58945
rect 148770 58850 148830 58935
rect 149530 58885 149620 58935
rect 148910 58855 149620 58885
rect 148950 58820 149070 58855
rect 149230 58820 149350 58855
rect 148660 58800 148740 58810
rect 148740 58730 148750 58800
rect 149060 58790 149130 58820
rect 148650 58670 148770 58730
rect 149070 58700 149130 58790
rect 149230 58730 149240 58820
rect 149340 58790 149410 58820
rect 149350 58700 149410 58790
rect 148770 58645 148830 58670
rect 149530 58665 149620 58855
rect 148910 58660 149620 58665
rect 148900 58650 149630 58660
rect 148910 58645 149630 58650
rect 148770 58635 149630 58645
rect 148770 58550 148830 58635
rect 149530 58585 149630 58635
rect 148910 58555 149630 58585
rect 148950 58520 149070 58555
rect 149230 58520 149350 58555
rect 149070 58510 149130 58520
rect 149350 58510 149410 58520
rect 148660 58500 148740 58510
rect 148970 58500 149050 58510
rect 149070 58500 149190 58510
rect 149250 58500 149330 58510
rect 149350 58500 149470 58510
rect 148740 58430 148750 58500
rect 148650 58370 148770 58430
rect 149050 58420 149060 58500
rect 149070 58400 149130 58500
rect 149190 58420 149200 58500
rect 149330 58420 149340 58500
rect 149350 58400 149410 58500
rect 149470 58420 149480 58500
rect 148770 58345 148830 58370
rect 149530 58365 149630 58555
rect 148910 58360 149630 58365
rect 148900 58350 149630 58360
rect 148910 58345 149620 58350
rect 148770 58335 149620 58345
rect 148770 58250 148830 58335
rect 149530 58285 149620 58335
rect 148910 58255 149620 58285
rect 148950 58220 149070 58255
rect 149230 58220 149350 58255
rect 149060 58190 149130 58220
rect 19880 58170 19960 58180
rect 20060 58170 20140 58180
rect 20240 58170 20320 58180
rect 20420 58170 20500 58180
rect 20600 58170 20680 58180
rect 20780 58170 20860 58180
rect 20960 58170 21040 58180
rect 21140 58170 21220 58180
rect 21320 58170 21400 58180
rect 21500 58170 21580 58180
rect 21680 58170 21760 58180
rect 21860 58170 21940 58180
rect 22040 58170 22120 58180
rect 22220 58170 22300 58180
rect 22400 58170 22480 58180
rect 22580 58170 22660 58180
rect 22760 58170 22840 58180
rect 22940 58170 23020 58180
rect 23120 58170 23200 58180
rect 23300 58170 23380 58180
rect 23480 58170 23560 58180
rect 23660 58170 23740 58180
rect 23840 58170 23920 58180
rect 24020 58170 24100 58180
rect 24200 58170 24280 58180
rect 24380 58170 24460 58180
rect 24560 58170 24640 58180
rect 24740 58170 24820 58180
rect 24920 58170 25000 58180
rect 25100 58170 25180 58180
rect 25280 58170 25360 58180
rect 25460 58170 25540 58180
rect 25640 58170 25720 58180
rect 19130 58110 19160 58140
rect 19250 58110 19280 58140
rect 19010 58080 19070 58110
rect 19130 58080 19190 58110
rect 19250 58080 19310 58110
rect 19960 58090 19970 58170
rect 20140 58090 20150 58170
rect 20320 58090 20330 58170
rect 20500 58090 20510 58170
rect 20680 58090 20690 58170
rect 20860 58090 20870 58170
rect 21040 58090 21050 58170
rect 21220 58090 21230 58170
rect 21400 58090 21410 58170
rect 21580 58090 21590 58170
rect 21760 58090 21770 58170
rect 21940 58090 21950 58170
rect 22120 58090 22130 58170
rect 22300 58090 22310 58170
rect 22480 58090 22490 58170
rect 22660 58090 22670 58170
rect 22840 58090 22850 58170
rect 23020 58090 23030 58170
rect 23200 58090 23210 58170
rect 23380 58090 23390 58170
rect 23560 58090 23570 58170
rect 23740 58090 23750 58170
rect 23920 58090 23930 58170
rect 24100 58090 24110 58170
rect 24280 58090 24290 58170
rect 24460 58090 24470 58170
rect 24640 58090 24650 58170
rect 24820 58090 24830 58170
rect 25000 58090 25010 58170
rect 25180 58090 25190 58170
rect 25360 58090 25370 58170
rect 25540 58090 25550 58170
rect 25720 58090 25730 58170
rect 31100 58150 37190 58180
rect 40060 58150 40120 58180
rect 41540 58150 41600 58180
rect 42360 58150 42420 58180
rect 43840 58150 43900 58180
rect 26420 58110 26450 58140
rect 26540 58110 26570 58140
rect 30420 58110 30450 58140
rect 30540 58110 30570 58140
rect 26300 58080 26360 58110
rect 26420 58080 26480 58110
rect 26540 58080 26600 58110
rect 30300 58080 30360 58110
rect 30420 58080 30480 58110
rect 30540 58080 30600 58110
rect 31260 58090 31270 58150
rect 31440 58090 31450 58150
rect 31620 58090 31630 58150
rect 31800 58090 31810 58150
rect 31980 58090 31990 58150
rect 32160 58090 32170 58150
rect 32340 58090 32350 58150
rect 32520 58090 32530 58150
rect 32700 58090 32710 58150
rect 32880 58090 32890 58150
rect 33060 58090 33070 58150
rect 33240 58090 33250 58150
rect 33420 58090 33430 58150
rect 33600 58090 33610 58150
rect 33780 58090 33790 58150
rect 33960 58090 33970 58150
rect 34140 58090 34150 58150
rect 34320 58090 34330 58150
rect 34500 58090 34510 58150
rect 34680 58090 34690 58150
rect 34860 58090 34870 58150
rect 35040 58090 35050 58150
rect 35220 58090 35230 58150
rect 35400 58090 35410 58150
rect 35580 58090 35590 58150
rect 35760 58090 35770 58150
rect 35940 58090 35950 58150
rect 36120 58090 36130 58150
rect 36300 58090 36310 58150
rect 36480 58090 36490 58150
rect 36660 58090 36670 58150
rect 36840 58090 36850 58150
rect 37020 58090 37030 58150
rect 37100 58080 37190 58150
rect 37720 58110 37750 58140
rect 37840 58110 37870 58140
rect 146100 58110 146160 58140
rect 147580 58110 147640 58140
rect 148400 58110 148460 58140
rect 37600 58080 37660 58110
rect 37720 58080 37780 58110
rect 37840 58080 37900 58110
rect 149070 58100 149130 58190
rect 149230 58130 149240 58220
rect 149340 58190 149410 58220
rect 149350 58100 149410 58190
rect 149530 58090 149620 58255
rect 31100 58050 37190 58080
rect 148910 58070 149620 58090
rect 148900 58060 149740 58070
rect 37100 58040 37190 58050
rect 19800 58030 25800 58040
rect 31100 58030 37190 58040
rect 40060 58030 40120 58060
rect 41540 58030 41600 58060
rect 42360 58030 42420 58060
rect 43840 58030 43900 58060
rect 19130 57990 19160 58020
rect 19250 57990 19280 58020
rect 26420 57990 26450 58020
rect 26540 57990 26570 58020
rect 30420 57990 30450 58020
rect 30540 57990 30570 58020
rect 19010 57960 19070 57990
rect 19130 57960 19190 57990
rect 19250 57960 19310 57990
rect 26300 57960 26360 57990
rect 26420 57960 26480 57990
rect 26540 57960 26600 57990
rect 30300 57960 30360 57990
rect 30420 57960 30480 57990
rect 30540 57960 30600 57990
rect 19130 57870 19160 57900
rect 19250 57870 19280 57900
rect 26420 57870 26450 57900
rect 26540 57870 26570 57900
rect 30420 57870 30450 57900
rect 30540 57870 30570 57900
rect 19010 57840 19070 57870
rect 19130 57840 19190 57870
rect 19250 57840 19310 57870
rect 26300 57840 26360 57870
rect 26420 57840 26480 57870
rect 26540 57840 26600 57870
rect 30300 57840 30360 57870
rect 30420 57840 30480 57870
rect 30540 57840 30600 57870
rect 31180 57850 31260 57860
rect 31360 57850 31440 57860
rect 31540 57850 31620 57860
rect 31720 57850 31800 57860
rect 31900 57850 31980 57860
rect 32080 57850 32160 57860
rect 32260 57850 32340 57860
rect 32440 57850 32520 57860
rect 32620 57850 32700 57860
rect 32800 57850 32880 57860
rect 32980 57850 33060 57860
rect 33160 57850 33240 57860
rect 33340 57850 33420 57860
rect 33520 57850 33600 57860
rect 33700 57850 33780 57860
rect 33880 57850 33960 57860
rect 34060 57850 34140 57860
rect 34240 57850 34320 57860
rect 34420 57850 34500 57860
rect 34600 57850 34680 57860
rect 34780 57850 34860 57860
rect 34960 57850 35040 57860
rect 35140 57850 35220 57860
rect 35320 57850 35400 57860
rect 35500 57850 35580 57860
rect 35680 57850 35760 57860
rect 35860 57850 35940 57860
rect 36040 57850 36120 57860
rect 36220 57850 36300 57860
rect 36400 57850 36480 57860
rect 36580 57850 36660 57860
rect 36760 57850 36840 57860
rect 36940 57850 37020 57860
rect 19880 57830 19960 57840
rect 20060 57830 20140 57840
rect 20240 57830 20320 57840
rect 20420 57830 20500 57840
rect 20600 57830 20680 57840
rect 20780 57830 20860 57840
rect 20960 57830 21040 57840
rect 21140 57830 21220 57840
rect 21320 57830 21400 57840
rect 21500 57830 21580 57840
rect 21680 57830 21760 57840
rect 21860 57830 21940 57840
rect 22040 57830 22120 57840
rect 22220 57830 22300 57840
rect 22400 57830 22480 57840
rect 22580 57830 22660 57840
rect 22760 57830 22840 57840
rect 22940 57830 23020 57840
rect 23120 57830 23200 57840
rect 23300 57830 23380 57840
rect 23480 57830 23560 57840
rect 23660 57830 23740 57840
rect 23840 57830 23920 57840
rect 24020 57830 24100 57840
rect 24200 57830 24280 57840
rect 24380 57830 24460 57840
rect 24560 57830 24640 57840
rect 24740 57830 24820 57840
rect 24920 57830 25000 57840
rect 25100 57830 25180 57840
rect 25280 57830 25360 57840
rect 25460 57830 25540 57840
rect 25640 57830 25720 57840
rect 19130 57750 19160 57780
rect 19250 57750 19280 57780
rect 19960 57750 19970 57830
rect 20140 57750 20150 57830
rect 20320 57750 20330 57830
rect 20500 57750 20510 57830
rect 20680 57750 20690 57830
rect 20860 57750 20870 57830
rect 21040 57750 21050 57830
rect 21220 57750 21230 57830
rect 21400 57750 21410 57830
rect 21580 57750 21590 57830
rect 21760 57750 21770 57830
rect 21940 57750 21950 57830
rect 22120 57750 22130 57830
rect 22300 57750 22310 57830
rect 22480 57750 22490 57830
rect 22660 57750 22670 57830
rect 22840 57750 22850 57830
rect 23020 57750 23030 57830
rect 23200 57750 23210 57830
rect 23380 57750 23390 57830
rect 23560 57750 23570 57830
rect 23740 57750 23750 57830
rect 23920 57750 23930 57830
rect 24100 57750 24110 57830
rect 24280 57750 24290 57830
rect 24460 57750 24470 57830
rect 24640 57750 24650 57830
rect 24820 57750 24830 57830
rect 25000 57750 25010 57830
rect 25180 57750 25190 57830
rect 25360 57750 25370 57830
rect 25540 57750 25550 57830
rect 25720 57750 25730 57830
rect 26420 57750 26450 57780
rect 26540 57750 26570 57780
rect 30420 57750 30450 57780
rect 30540 57750 30570 57780
rect 31260 57770 31270 57850
rect 31440 57770 31450 57850
rect 31620 57770 31630 57850
rect 31800 57770 31810 57850
rect 31980 57770 31990 57850
rect 32160 57770 32170 57850
rect 32340 57770 32350 57850
rect 32520 57770 32530 57850
rect 32700 57770 32710 57850
rect 32880 57770 32890 57850
rect 33060 57770 33070 57850
rect 33240 57770 33250 57850
rect 33420 57770 33430 57850
rect 33600 57770 33610 57850
rect 33780 57770 33790 57850
rect 33960 57770 33970 57850
rect 34140 57770 34150 57850
rect 34320 57770 34330 57850
rect 34500 57770 34510 57850
rect 34680 57770 34690 57850
rect 34860 57770 34870 57850
rect 35040 57770 35050 57850
rect 35220 57770 35230 57850
rect 35400 57770 35410 57850
rect 35580 57770 35590 57850
rect 35760 57770 35770 57850
rect 35940 57770 35950 57850
rect 36120 57770 36130 57850
rect 36300 57770 36310 57850
rect 36480 57770 36490 57850
rect 36660 57770 36670 57850
rect 36840 57770 36850 57850
rect 37020 57770 37030 57850
rect 19010 57720 19070 57750
rect 19130 57720 19190 57750
rect 19250 57720 19310 57750
rect 26300 57720 26360 57750
rect 26420 57720 26480 57750
rect 26540 57720 26600 57750
rect 30300 57720 30360 57750
rect 30420 57720 30480 57750
rect 30540 57720 30600 57750
rect 19130 57630 19160 57660
rect 19250 57630 19280 57660
rect 26420 57630 26450 57660
rect 26540 57630 26570 57660
rect 30420 57630 30450 57660
rect 30540 57630 30570 57660
rect 19010 57600 19070 57630
rect 19130 57600 19190 57630
rect 19250 57600 19310 57630
rect 26300 57600 26360 57630
rect 26420 57600 26480 57630
rect 26540 57600 26600 57630
rect 30300 57600 30360 57630
rect 30420 57600 30480 57630
rect 30540 57600 30600 57630
rect 19130 57510 19160 57540
rect 19250 57510 19280 57540
rect 19880 57530 19960 57540
rect 20060 57530 20140 57540
rect 20240 57530 20320 57540
rect 20420 57530 20500 57540
rect 20600 57530 20680 57540
rect 20780 57530 20860 57540
rect 20960 57530 21040 57540
rect 21140 57530 21220 57540
rect 21320 57530 21400 57540
rect 21500 57530 21580 57540
rect 21680 57530 21760 57540
rect 21860 57530 21940 57540
rect 22040 57530 22120 57540
rect 22220 57530 22300 57540
rect 22400 57530 22480 57540
rect 22580 57530 22660 57540
rect 22760 57530 22840 57540
rect 22940 57530 23020 57540
rect 23120 57530 23200 57540
rect 23300 57530 23380 57540
rect 23480 57530 23560 57540
rect 23660 57530 23740 57540
rect 23840 57530 23920 57540
rect 24020 57530 24100 57540
rect 24200 57530 24280 57540
rect 24380 57530 24460 57540
rect 24560 57530 24640 57540
rect 24740 57530 24820 57540
rect 24920 57530 25000 57540
rect 25100 57530 25180 57540
rect 25280 57530 25360 57540
rect 25460 57530 25540 57540
rect 25640 57530 25720 57540
rect 19010 57480 19070 57510
rect 19130 57480 19190 57510
rect 19250 57480 19310 57510
rect 19960 57450 19970 57530
rect 20140 57450 20150 57530
rect 20320 57450 20330 57530
rect 20500 57450 20510 57530
rect 20680 57450 20690 57530
rect 20860 57450 20870 57530
rect 21040 57450 21050 57530
rect 21220 57450 21230 57530
rect 21400 57450 21410 57530
rect 21580 57450 21590 57530
rect 21760 57450 21770 57530
rect 21940 57450 21950 57530
rect 22120 57450 22130 57530
rect 22300 57450 22310 57530
rect 22480 57450 22490 57530
rect 22660 57450 22670 57530
rect 22840 57450 22850 57530
rect 23020 57450 23030 57530
rect 23200 57450 23210 57530
rect 23380 57450 23390 57530
rect 23560 57450 23570 57530
rect 23740 57450 23750 57530
rect 23920 57450 23930 57530
rect 24100 57450 24110 57530
rect 24280 57450 24290 57530
rect 24460 57450 24470 57530
rect 24640 57450 24650 57530
rect 24820 57450 24830 57530
rect 25000 57450 25010 57530
rect 25180 57450 25190 57530
rect 25360 57450 25370 57530
rect 25540 57450 25550 57530
rect 25720 57450 25730 57530
rect 26420 57510 26450 57540
rect 26540 57510 26570 57540
rect 30420 57510 30450 57540
rect 30540 57510 30570 57540
rect 31180 57530 31260 57540
rect 31360 57530 31440 57540
rect 31540 57530 31620 57540
rect 31720 57530 31800 57540
rect 31900 57530 31980 57540
rect 32080 57530 32160 57540
rect 32260 57530 32340 57540
rect 32440 57530 32520 57540
rect 32620 57530 32700 57540
rect 32800 57530 32880 57540
rect 32980 57530 33060 57540
rect 33160 57530 33240 57540
rect 33340 57530 33420 57540
rect 33520 57530 33600 57540
rect 33700 57530 33780 57540
rect 33880 57530 33960 57540
rect 34060 57530 34140 57540
rect 34240 57530 34320 57540
rect 34420 57530 34500 57540
rect 34600 57530 34680 57540
rect 34780 57530 34860 57540
rect 34960 57530 35040 57540
rect 35140 57530 35220 57540
rect 35320 57530 35400 57540
rect 35500 57530 35580 57540
rect 35680 57530 35760 57540
rect 35860 57530 35940 57540
rect 36040 57530 36120 57540
rect 36220 57530 36300 57540
rect 36400 57530 36480 57540
rect 36580 57530 36660 57540
rect 36760 57530 36840 57540
rect 36940 57530 37020 57540
rect 26300 57480 26360 57510
rect 26420 57480 26480 57510
rect 26540 57480 26600 57510
rect 30300 57480 30360 57510
rect 30420 57480 30480 57510
rect 30540 57480 30600 57510
rect 31260 57450 31270 57530
rect 31440 57450 31450 57530
rect 31620 57450 31630 57530
rect 31800 57450 31810 57530
rect 31980 57450 31990 57530
rect 32160 57450 32170 57530
rect 32340 57450 32350 57530
rect 32520 57450 32530 57530
rect 32700 57450 32710 57530
rect 32880 57450 32890 57530
rect 33060 57450 33070 57530
rect 33240 57450 33250 57530
rect 33420 57450 33430 57530
rect 33600 57450 33610 57530
rect 33780 57450 33790 57530
rect 33960 57450 33970 57530
rect 34140 57450 34150 57530
rect 34320 57450 34330 57530
rect 34500 57450 34510 57530
rect 34680 57450 34690 57530
rect 34860 57450 34870 57530
rect 35040 57450 35050 57530
rect 35220 57450 35230 57530
rect 35400 57450 35410 57530
rect 35580 57450 35590 57530
rect 35760 57450 35770 57530
rect 35940 57450 35950 57530
rect 36120 57450 36130 57530
rect 36300 57450 36310 57530
rect 36480 57450 36490 57530
rect 36660 57450 36670 57530
rect 36840 57450 36850 57530
rect 37020 57450 37030 57530
rect 19130 57390 19160 57420
rect 19250 57390 19280 57420
rect 26420 57390 26450 57420
rect 26540 57390 26570 57420
rect 30420 57390 30450 57420
rect 30540 57390 30570 57420
rect 19010 57360 19070 57390
rect 19130 57360 19190 57390
rect 19250 57360 19310 57390
rect 26300 57360 26360 57390
rect 26420 57360 26480 57390
rect 26540 57360 26600 57390
rect 30300 57360 30360 57390
rect 30420 57360 30480 57390
rect 30540 57360 30600 57390
rect 37100 57360 37190 58030
rect 37720 57990 37750 58020
rect 37840 57990 37870 58020
rect 146100 57990 146160 58020
rect 37600 57960 37660 57990
rect 37720 57960 37780 57990
rect 37840 57960 37900 57990
rect 146690 57940 146810 58000
rect 146970 57940 147090 58000
rect 147580 57990 147640 58020
rect 148400 57990 148460 58020
rect 148820 57970 149620 58060
rect 148950 57940 149070 57970
rect 149230 57940 149350 57970
rect 40060 57910 40120 57940
rect 41540 57910 41600 57940
rect 42360 57910 42420 57940
rect 43840 57910 43900 57940
rect 146810 57930 146870 57940
rect 146570 57920 146650 57930
rect 146810 57920 146930 57930
rect 37720 57870 37750 57900
rect 37840 57870 37870 57900
rect 146100 57870 146160 57900
rect 37600 57840 37660 57870
rect 37720 57840 37780 57870
rect 37840 57840 37900 57870
rect 146650 57840 146660 57920
rect 146810 57820 146870 57920
rect 146930 57840 146940 57920
rect 147090 57820 147150 57940
rect 149070 57930 149130 57940
rect 149350 57930 149410 57940
rect 149070 57920 149190 57930
rect 149350 57920 149470 57930
rect 40060 57790 40120 57820
rect 41540 57790 41600 57820
rect 42360 57790 42420 57820
rect 43840 57790 43900 57820
rect 37720 57750 37750 57780
rect 37840 57750 37870 57780
rect 146100 57750 146160 57780
rect 146500 57770 147140 57780
rect 147220 57765 147230 57820
rect 147270 57790 147390 57850
rect 146460 57755 147250 57765
rect 37600 57720 37660 57750
rect 37720 57720 37780 57750
rect 37840 57720 37900 57750
rect 146450 57705 146460 57755
rect 40060 57670 40120 57700
rect 41540 57670 41600 57700
rect 42360 57670 42420 57700
rect 43840 57670 43900 57700
rect 37720 57630 37750 57660
rect 37840 57630 37870 57660
rect 146100 57630 146160 57660
rect 146690 57640 146810 57700
rect 146970 57640 147090 57700
rect 146810 57630 146870 57640
rect 37600 57600 37660 57630
rect 37720 57600 37780 57630
rect 37840 57600 37900 57630
rect 146570 57620 146650 57630
rect 146710 57620 146790 57630
rect 146810 57620 146930 57630
rect 146990 57620 147070 57630
rect 40060 57550 40120 57580
rect 41540 57550 41600 57580
rect 42360 57550 42420 57580
rect 43840 57550 43900 57580
rect 146650 57540 146660 57620
rect 146790 57540 146800 57620
rect 37720 57510 37750 57540
rect 37840 57510 37870 57540
rect 146100 57510 146160 57540
rect 146810 57520 146870 57620
rect 146930 57540 146940 57620
rect 147070 57540 147080 57620
rect 147090 57520 147150 57640
rect 37600 57480 37660 57510
rect 37720 57480 37780 57510
rect 37840 57480 37900 57510
rect 146510 57490 147130 57500
rect 147220 57480 147230 57755
rect 147390 57670 147450 57790
rect 147300 57640 147380 57650
rect 147380 57570 147390 57640
rect 147300 57560 147390 57570
rect 147300 57480 147380 57490
rect 40060 57430 40120 57460
rect 41540 57430 41600 57460
rect 42360 57430 42420 57460
rect 43840 57430 43900 57460
rect 37720 57390 37750 57420
rect 37840 57390 37870 57420
rect 146100 57390 146160 57420
rect 37600 57360 37660 57390
rect 37720 57360 37780 57390
rect 37840 57360 37900 57390
rect 146610 57360 146970 57420
rect 147380 57400 147390 57480
rect 19800 57350 25800 57360
rect 31100 57350 37190 57360
rect 19130 57270 19160 57300
rect 19250 57270 19280 57300
rect 26420 57270 26450 57300
rect 26540 57270 26570 57300
rect 30420 57270 30450 57300
rect 30540 57270 30570 57300
rect 19010 57240 19070 57270
rect 19130 57240 19190 57270
rect 19250 57240 19310 57270
rect 26300 57240 26360 57270
rect 26420 57240 26480 57270
rect 26540 57240 26600 57270
rect 30300 57240 30360 57270
rect 30420 57240 30480 57270
rect 30540 57240 30600 57270
rect 37100 57250 37190 57350
rect 147520 57340 147530 57910
rect 147580 57870 147640 57900
rect 148400 57870 148460 57900
rect 148510 57820 148520 57910
rect 147580 57750 147640 57780
rect 148400 57750 148460 57780
rect 147580 57630 147640 57660
rect 148400 57630 148460 57660
rect 147580 57510 147640 57540
rect 148400 57510 148460 57540
rect 147580 57390 147640 57420
rect 148400 57390 148460 57420
rect 40060 57310 40120 57340
rect 41540 57310 41600 57340
rect 42360 57310 42420 57340
rect 43840 57310 43900 57340
rect 37720 57270 37750 57300
rect 37840 57270 37870 57300
rect 146100 57270 146160 57300
rect 31100 57220 37190 57250
rect 37600 57240 37660 57270
rect 37720 57240 37780 57270
rect 37840 57240 37900 57270
rect 146300 57230 146420 57290
rect 147580 57270 147640 57300
rect 148400 57270 148460 57300
rect 146420 57220 146480 57230
rect 19880 57210 19960 57220
rect 20060 57210 20140 57220
rect 20240 57210 20320 57220
rect 20420 57210 20500 57220
rect 20600 57210 20680 57220
rect 20780 57210 20860 57220
rect 20960 57210 21040 57220
rect 21140 57210 21220 57220
rect 21320 57210 21400 57220
rect 21500 57210 21580 57220
rect 21680 57210 21760 57220
rect 21860 57210 21940 57220
rect 22040 57210 22120 57220
rect 22220 57210 22300 57220
rect 22400 57210 22480 57220
rect 22580 57210 22660 57220
rect 22760 57210 22840 57220
rect 22940 57210 23020 57220
rect 23120 57210 23200 57220
rect 23300 57210 23380 57220
rect 23480 57210 23560 57220
rect 23660 57210 23740 57220
rect 23840 57210 23920 57220
rect 24020 57210 24100 57220
rect 24200 57210 24280 57220
rect 24380 57210 24460 57220
rect 24560 57210 24640 57220
rect 24740 57210 24820 57220
rect 24920 57210 25000 57220
rect 25100 57210 25180 57220
rect 25280 57210 25360 57220
rect 25460 57210 25540 57220
rect 25640 57210 25720 57220
rect 31180 57210 31260 57220
rect 31360 57210 31440 57220
rect 31540 57210 31620 57220
rect 31720 57210 31800 57220
rect 31900 57210 31980 57220
rect 32080 57210 32160 57220
rect 32260 57210 32340 57220
rect 32440 57210 32520 57220
rect 32620 57210 32700 57220
rect 32800 57210 32880 57220
rect 32980 57210 33060 57220
rect 33160 57210 33240 57220
rect 33340 57210 33420 57220
rect 33520 57210 33600 57220
rect 33700 57210 33780 57220
rect 33880 57210 33960 57220
rect 34060 57210 34140 57220
rect 34240 57210 34320 57220
rect 34420 57210 34500 57220
rect 34600 57210 34680 57220
rect 34780 57210 34860 57220
rect 34960 57210 35040 57220
rect 35140 57210 35220 57220
rect 35320 57210 35400 57220
rect 35500 57210 35580 57220
rect 35680 57210 35760 57220
rect 35860 57210 35940 57220
rect 36040 57210 36120 57220
rect 36220 57210 36300 57220
rect 36400 57210 36480 57220
rect 36580 57210 36660 57220
rect 36760 57210 36840 57220
rect 36940 57210 37020 57220
rect 19130 57150 19160 57180
rect 19250 57150 19280 57180
rect 19010 57120 19070 57150
rect 19130 57120 19190 57150
rect 19250 57120 19310 57150
rect 19960 57130 19970 57210
rect 20140 57130 20150 57210
rect 20320 57130 20330 57210
rect 20500 57130 20510 57210
rect 20680 57130 20690 57210
rect 20860 57130 20870 57210
rect 21040 57130 21050 57210
rect 21220 57130 21230 57210
rect 21400 57130 21410 57210
rect 21580 57130 21590 57210
rect 21760 57130 21770 57210
rect 21940 57130 21950 57210
rect 22120 57130 22130 57210
rect 22300 57130 22310 57210
rect 22480 57130 22490 57210
rect 22660 57130 22670 57210
rect 22840 57130 22850 57210
rect 23020 57130 23030 57210
rect 23200 57130 23210 57210
rect 23380 57130 23390 57210
rect 23560 57130 23570 57210
rect 23740 57130 23750 57210
rect 23920 57130 23930 57210
rect 24100 57130 24110 57210
rect 24280 57130 24290 57210
rect 24460 57130 24470 57210
rect 24640 57130 24650 57210
rect 24820 57130 24830 57210
rect 25000 57130 25010 57210
rect 25180 57130 25190 57210
rect 25360 57130 25370 57210
rect 25540 57130 25550 57210
rect 25720 57130 25730 57210
rect 26420 57150 26450 57180
rect 26540 57150 26570 57180
rect 30420 57150 30450 57180
rect 30540 57150 30570 57180
rect 31260 57150 31270 57210
rect 31440 57150 31450 57210
rect 31620 57150 31630 57210
rect 31800 57150 31810 57210
rect 31980 57150 31990 57210
rect 32160 57150 32170 57210
rect 32340 57150 32350 57210
rect 32520 57150 32530 57210
rect 32700 57150 32710 57210
rect 32880 57150 32890 57210
rect 33060 57150 33070 57210
rect 33240 57150 33250 57210
rect 33420 57150 33430 57210
rect 33600 57150 33610 57210
rect 33780 57150 33790 57210
rect 33960 57150 33970 57210
rect 34140 57150 34150 57210
rect 34320 57150 34330 57210
rect 34500 57150 34510 57210
rect 34680 57150 34690 57210
rect 34860 57150 34870 57210
rect 35040 57150 35050 57210
rect 35220 57150 35230 57210
rect 35400 57150 35410 57210
rect 35580 57150 35590 57210
rect 35760 57150 35770 57210
rect 35940 57150 35950 57210
rect 36120 57150 36130 57210
rect 36300 57150 36310 57210
rect 36480 57150 36490 57210
rect 36660 57150 36670 57210
rect 36840 57150 36850 57210
rect 37020 57150 37030 57210
rect 37100 57150 37190 57220
rect 40060 57190 40120 57220
rect 41540 57190 41600 57220
rect 42360 57190 42420 57220
rect 43840 57190 43900 57220
rect 146420 57210 147050 57220
rect 146420 57205 146480 57210
rect 146420 57195 147090 57205
rect 148600 57200 148610 57820
rect 148650 57790 148770 57850
rect 149070 57820 149130 57920
rect 149190 57840 149200 57920
rect 149350 57820 149410 57920
rect 149470 57840 149480 57920
rect 148770 57765 148830 57790
rect 149530 57785 149620 57970
rect 148910 57780 149620 57785
rect 148900 57770 149630 57780
rect 148910 57765 149630 57770
rect 148770 57755 149630 57765
rect 148770 57670 148830 57755
rect 149530 57705 149630 57755
rect 148910 57675 149630 57705
rect 148950 57640 149070 57675
rect 149230 57640 149350 57675
rect 149070 57630 149130 57640
rect 149350 57630 149410 57640
rect 148660 57620 148740 57630
rect 148970 57620 149050 57630
rect 149070 57620 149190 57630
rect 149250 57620 149330 57630
rect 149350 57620 149470 57630
rect 148740 57550 148750 57620
rect 148650 57490 148770 57550
rect 149050 57540 149060 57620
rect 149070 57520 149130 57620
rect 149190 57540 149200 57620
rect 149330 57540 149340 57620
rect 149350 57520 149410 57620
rect 149470 57540 149480 57620
rect 148770 57465 148830 57490
rect 149530 57485 149630 57675
rect 148910 57480 149630 57485
rect 148900 57470 149630 57480
rect 148910 57465 149620 57470
rect 148770 57455 149620 57465
rect 148770 57370 148830 57455
rect 149530 57405 149620 57455
rect 148910 57375 149620 57405
rect 148660 57340 148740 57350
rect 148950 57340 149070 57375
rect 149230 57340 149350 57375
rect 148740 57260 148750 57340
rect 149060 57310 149130 57340
rect 149070 57220 149130 57310
rect 149230 57250 149240 57340
rect 149340 57310 149410 57340
rect 149350 57220 149410 57310
rect 37720 57150 37750 57180
rect 37840 57150 37870 57180
rect 146100 57150 146160 57180
rect 26300 57120 26360 57150
rect 26420 57120 26480 57150
rect 26540 57120 26600 57150
rect 30300 57120 30360 57150
rect 30420 57120 30480 57150
rect 30540 57120 30600 57150
rect 31100 57120 37190 57150
rect 37600 57120 37660 57150
rect 37720 57120 37780 57150
rect 37840 57120 37900 57150
rect 19880 57060 19960 57070
rect 20060 57060 20140 57070
rect 20240 57060 20320 57070
rect 20420 57060 20500 57070
rect 20600 57060 20680 57070
rect 20780 57060 20860 57070
rect 20960 57060 21040 57070
rect 21140 57060 21220 57070
rect 21320 57060 21400 57070
rect 21500 57060 21580 57070
rect 21680 57060 21760 57070
rect 21860 57060 21940 57070
rect 22040 57060 22120 57070
rect 22220 57060 22300 57070
rect 22400 57060 22480 57070
rect 22580 57060 22660 57070
rect 22760 57060 22840 57070
rect 22940 57060 23020 57070
rect 23120 57060 23200 57070
rect 23300 57060 23380 57070
rect 23480 57060 23560 57070
rect 23660 57060 23740 57070
rect 23840 57060 23920 57070
rect 24020 57060 24100 57070
rect 24200 57060 24280 57070
rect 24380 57060 24460 57070
rect 24560 57060 24640 57070
rect 24740 57060 24820 57070
rect 24920 57060 25000 57070
rect 25100 57060 25180 57070
rect 25280 57060 25360 57070
rect 25460 57060 25540 57070
rect 25640 57060 25720 57070
rect 31180 57060 31260 57070
rect 31360 57060 31440 57070
rect 31540 57060 31620 57070
rect 31720 57060 31800 57070
rect 31900 57060 31980 57070
rect 32080 57060 32160 57070
rect 32260 57060 32340 57070
rect 32440 57060 32520 57070
rect 32620 57060 32700 57070
rect 32800 57060 32880 57070
rect 32980 57060 33060 57070
rect 33160 57060 33240 57070
rect 33340 57060 33420 57070
rect 33520 57060 33600 57070
rect 33700 57060 33780 57070
rect 33880 57060 33960 57070
rect 34060 57060 34140 57070
rect 34240 57060 34320 57070
rect 34420 57060 34500 57070
rect 34600 57060 34680 57070
rect 34780 57060 34860 57070
rect 34960 57060 35040 57070
rect 35140 57060 35220 57070
rect 35320 57060 35400 57070
rect 35500 57060 35580 57070
rect 35680 57060 35760 57070
rect 35860 57060 35940 57070
rect 36040 57060 36120 57070
rect 36220 57060 36300 57070
rect 36400 57060 36480 57070
rect 36580 57060 36660 57070
rect 36760 57060 36840 57070
rect 36940 57060 37020 57070
rect 19130 57030 19160 57060
rect 19250 57030 19280 57060
rect 19010 57000 19070 57030
rect 19130 57000 19190 57030
rect 19250 57000 19310 57030
rect 19960 56980 19970 57060
rect 20140 56980 20150 57060
rect 20320 56980 20330 57060
rect 20500 56980 20510 57060
rect 20680 56980 20690 57060
rect 20860 56980 20870 57060
rect 21040 56980 21050 57060
rect 21220 56980 21230 57060
rect 21400 56980 21410 57060
rect 21580 56980 21590 57060
rect 21760 56980 21770 57060
rect 21940 56980 21950 57060
rect 22120 56980 22130 57060
rect 22300 56980 22310 57060
rect 22480 56980 22490 57060
rect 22660 56980 22670 57060
rect 22840 56980 22850 57060
rect 23020 56980 23030 57060
rect 23200 56980 23210 57060
rect 23380 56980 23390 57060
rect 23560 56980 23570 57060
rect 23740 56980 23750 57060
rect 23920 56980 23930 57060
rect 24100 56980 24110 57060
rect 24280 56980 24290 57060
rect 24460 56980 24470 57060
rect 24640 56980 24650 57060
rect 24820 56980 24830 57060
rect 25000 56980 25010 57060
rect 25180 56980 25190 57060
rect 25360 56980 25370 57060
rect 25540 56980 25550 57060
rect 25720 56980 25730 57060
rect 26420 57030 26450 57060
rect 26540 57030 26570 57060
rect 30420 57030 30450 57060
rect 30540 57030 30570 57060
rect 26300 57000 26360 57030
rect 26420 57000 26480 57030
rect 26540 57000 26600 57030
rect 30300 57000 30360 57030
rect 30420 57000 30480 57030
rect 30540 57000 30600 57030
rect 31260 56980 31270 57060
rect 31440 56980 31450 57060
rect 31620 56980 31630 57060
rect 31800 56980 31810 57060
rect 31980 56980 31990 57060
rect 32160 56980 32170 57060
rect 32340 56980 32350 57060
rect 32520 56980 32530 57060
rect 32700 56980 32710 57060
rect 32880 56980 32890 57060
rect 33060 56980 33070 57060
rect 33240 56980 33250 57060
rect 33420 56980 33430 57060
rect 33600 56980 33610 57060
rect 33780 56980 33790 57060
rect 33960 56980 33970 57060
rect 34140 56980 34150 57060
rect 34320 56980 34330 57060
rect 34500 56980 34510 57060
rect 34680 56980 34690 57060
rect 34860 56980 34870 57060
rect 35040 56980 35050 57060
rect 35220 56980 35230 57060
rect 35400 56980 35410 57060
rect 35580 56980 35590 57060
rect 35760 56980 35770 57060
rect 35940 56980 35950 57060
rect 36120 56980 36130 57060
rect 36300 56980 36310 57060
rect 36480 56980 36490 57060
rect 36660 56980 36670 57060
rect 36840 56980 36850 57060
rect 37020 56980 37030 57060
rect 19130 56910 19160 56940
rect 19250 56910 19280 56940
rect 19880 56910 19960 56920
rect 20060 56910 20140 56920
rect 20240 56910 20320 56920
rect 20420 56910 20500 56920
rect 20600 56910 20680 56920
rect 20780 56910 20860 56920
rect 20960 56910 21040 56920
rect 21140 56910 21220 56920
rect 21320 56910 21400 56920
rect 21500 56910 21580 56920
rect 21680 56910 21760 56920
rect 21860 56910 21940 56920
rect 22040 56910 22120 56920
rect 22220 56910 22300 56920
rect 22400 56910 22480 56920
rect 22580 56910 22660 56920
rect 22760 56910 22840 56920
rect 22940 56910 23020 56920
rect 23120 56910 23200 56920
rect 23300 56910 23380 56920
rect 23480 56910 23560 56920
rect 23660 56910 23740 56920
rect 23840 56910 23920 56920
rect 24020 56910 24100 56920
rect 24200 56910 24280 56920
rect 24380 56910 24460 56920
rect 24560 56910 24640 56920
rect 24740 56910 24820 56920
rect 24920 56910 25000 56920
rect 25100 56910 25180 56920
rect 25280 56910 25360 56920
rect 25460 56910 25540 56920
rect 25640 56910 25720 56920
rect 26420 56910 26450 56940
rect 26540 56910 26570 56940
rect 30420 56910 30450 56940
rect 30540 56910 30570 56940
rect 37100 56920 37190 57120
rect 146420 57110 146480 57195
rect 40060 57070 40120 57100
rect 41540 57070 41600 57100
rect 42360 57070 42420 57100
rect 43840 57070 43900 57100
rect 37720 57030 37750 57060
rect 37840 57030 37870 57060
rect 146100 57030 146160 57060
rect 37600 57000 37660 57030
rect 37720 57000 37780 57030
rect 37840 57000 37900 57030
rect 40060 56950 40120 56980
rect 41540 56950 41600 56980
rect 42360 56950 42420 56980
rect 43840 56950 43900 56980
rect 146300 56970 146420 57030
rect 146420 56945 146480 56970
rect 146530 56960 146540 57130
rect 146610 57100 146970 57160
rect 147090 57145 147100 57195
rect 149530 57190 149620 57375
rect 149820 57180 149830 60150
rect 152080 60140 152160 60150
rect 152260 60140 152340 60150
rect 152440 60140 152520 60150
rect 152620 60140 152700 60150
rect 152800 60140 152880 60150
rect 152980 60140 153060 60150
rect 153160 60140 153240 60150
rect 153340 60140 153420 60150
rect 153520 60140 153600 60150
rect 153700 60140 153780 60150
rect 153880 60140 153960 60150
rect 154060 60140 154140 60150
rect 154240 60140 154320 60150
rect 154420 60140 154500 60150
rect 154600 60140 154680 60150
rect 154780 60140 154860 60150
rect 154960 60140 155040 60150
rect 155140 60140 155220 60150
rect 155320 60140 155400 60150
rect 155500 60140 155580 60150
rect 155680 60140 155760 60150
rect 155860 60140 155940 60150
rect 156040 60140 156120 60150
rect 156220 60140 156300 60150
rect 156400 60140 156480 60150
rect 156580 60140 156660 60150
rect 156760 60140 156840 60150
rect 156940 60140 157020 60150
rect 157120 60140 157200 60150
rect 157300 60140 157380 60150
rect 157480 60140 157560 60150
rect 157660 60140 157740 60150
rect 157840 60140 157920 60150
rect 158020 60140 158100 60150
rect 158200 60140 158280 60150
rect 158380 60140 158460 60150
rect 158560 60140 158640 60150
rect 158740 60140 158820 60150
rect 158920 60140 159000 60150
rect 159100 60140 159180 60150
rect 159280 60140 159360 60150
rect 159460 60140 159540 60150
rect 159640 60140 159720 60150
rect 152160 60060 152170 60140
rect 152340 60060 152350 60140
rect 152520 60060 152530 60140
rect 152700 60060 152710 60140
rect 152880 60060 152890 60140
rect 153060 60060 153070 60140
rect 153240 60060 153250 60140
rect 153420 60060 153430 60140
rect 153600 60060 153610 60140
rect 153780 60060 153790 60140
rect 153960 60060 153970 60140
rect 154140 60060 154150 60140
rect 154320 60060 154330 60140
rect 154500 60060 154510 60140
rect 154680 60060 154690 60140
rect 154860 60060 154870 60140
rect 155040 60060 155050 60140
rect 155220 60060 155230 60140
rect 155400 60060 155410 60140
rect 155580 60060 155590 60140
rect 155760 60060 155770 60140
rect 155940 60060 155950 60140
rect 156120 60060 156130 60140
rect 156300 60060 156310 60140
rect 156480 60060 156490 60140
rect 156660 60060 156670 60140
rect 156840 60060 156850 60140
rect 157020 60060 157030 60140
rect 157200 60060 157210 60140
rect 157380 60060 157390 60140
rect 157560 60060 157570 60140
rect 157740 60060 157750 60140
rect 157920 60060 157930 60140
rect 158100 60060 158110 60140
rect 158280 60060 158290 60140
rect 158460 60060 158470 60140
rect 158640 60060 158650 60140
rect 158820 60060 158830 60140
rect 159000 60060 159010 60140
rect 159180 60060 159190 60140
rect 159360 60060 159370 60140
rect 159540 60060 159550 60140
rect 159720 60060 159730 60140
rect 161965 60085 161975 60165
rect 162145 60085 162155 60165
rect 162325 60085 162335 60165
rect 162505 60085 162515 60165
rect 162685 60085 162695 60165
rect 163380 60140 163460 60150
rect 163560 60140 163640 60150
rect 163740 60140 163820 60150
rect 163920 60140 164000 60150
rect 164100 60140 164180 60150
rect 164280 60140 164360 60150
rect 164460 60140 164540 60150
rect 164640 60140 164720 60150
rect 164820 60140 164900 60150
rect 165000 60140 165080 60150
rect 165180 60140 165260 60150
rect 165360 60140 165440 60150
rect 165540 60140 165620 60150
rect 165720 60140 165800 60150
rect 165900 60140 165980 60150
rect 166080 60140 166160 60150
rect 166260 60140 166340 60150
rect 166440 60140 166520 60150
rect 166620 60140 166700 60150
rect 166800 60140 166880 60150
rect 166980 60140 167060 60150
rect 167160 60140 167240 60150
rect 167340 60140 167420 60150
rect 167520 60140 167600 60150
rect 167700 60140 167780 60150
rect 167880 60140 167960 60150
rect 168060 60140 168140 60150
rect 168240 60140 168320 60150
rect 168420 60140 168500 60150
rect 168600 60140 168680 60150
rect 168780 60140 168860 60150
rect 168960 60140 169040 60150
rect 169140 60140 169220 60150
rect 169320 60140 169400 60150
rect 169500 60140 169580 60150
rect 169680 60140 169760 60150
rect 169860 60140 169940 60150
rect 170040 60140 170120 60150
rect 170220 60140 170300 60150
rect 170400 60140 170480 60150
rect 170580 60140 170660 60150
rect 170760 60140 170840 60150
rect 170940 60140 171020 60150
rect 163460 60060 163470 60140
rect 163640 60060 163650 60140
rect 163820 60060 163830 60140
rect 164000 60060 164010 60140
rect 164180 60060 164190 60140
rect 164360 60060 164370 60140
rect 164540 60060 164550 60140
rect 164720 60060 164730 60140
rect 164900 60060 164910 60140
rect 165080 60060 165090 60140
rect 165260 60060 165270 60140
rect 165440 60060 165450 60140
rect 165620 60060 165630 60140
rect 165800 60060 165810 60140
rect 165980 60060 165990 60140
rect 166160 60060 166170 60140
rect 166340 60060 166350 60140
rect 166520 60060 166530 60140
rect 166700 60060 166710 60140
rect 166880 60060 166890 60140
rect 167060 60060 167070 60140
rect 167240 60060 167250 60140
rect 167420 60060 167430 60140
rect 167600 60060 167610 60140
rect 167780 60060 167790 60140
rect 167960 60060 167970 60140
rect 168140 60060 168150 60140
rect 168320 60060 168330 60140
rect 168500 60060 168510 60140
rect 168680 60060 168690 60140
rect 168860 60060 168870 60140
rect 169040 60060 169050 60140
rect 169220 60060 169230 60140
rect 169400 60060 169410 60140
rect 169580 60060 169590 60140
rect 169760 60060 169770 60140
rect 169940 60060 169950 60140
rect 170120 60060 170130 60140
rect 170300 60060 170310 60140
rect 170480 60060 170490 60140
rect 170660 60060 170670 60140
rect 170840 60060 170850 60140
rect 171020 60060 171030 60140
rect 149880 60030 149940 60060
rect 149880 59910 149940 59940
rect 152220 59890 152250 59920
rect 152340 59890 152370 59920
rect 159520 59890 159550 59920
rect 159640 59890 159670 59920
rect 152100 59860 152160 59890
rect 152220 59860 152280 59890
rect 152340 59860 152400 59890
rect 159400 59860 159460 59890
rect 159520 59860 159580 59890
rect 159640 59860 159700 59890
rect 149880 59790 149940 59820
rect 152220 59770 152250 59800
rect 152340 59770 152370 59800
rect 159520 59770 159550 59800
rect 159640 59770 159670 59800
rect 163520 59770 163550 59800
rect 163640 59770 163670 59800
rect 170810 59770 170840 59800
rect 170930 59770 170960 59800
rect 152100 59740 152160 59770
rect 152220 59740 152280 59770
rect 152340 59740 152400 59770
rect 149880 59670 149940 59700
rect 152220 59650 152250 59680
rect 152340 59650 152370 59680
rect 152810 59670 158990 59760
rect 159400 59740 159460 59770
rect 159520 59740 159580 59770
rect 159640 59740 159700 59770
rect 163400 59740 163460 59770
rect 163520 59740 163580 59770
rect 163640 59740 163700 59770
rect 170690 59740 170750 59770
rect 170810 59740 170870 59770
rect 170930 59740 170990 59770
rect 164280 59730 164360 59740
rect 164460 59730 164540 59740
rect 164640 59730 164720 59740
rect 164820 59730 164900 59740
rect 165000 59730 165080 59740
rect 165180 59730 165260 59740
rect 165360 59730 165440 59740
rect 165540 59730 165620 59740
rect 165720 59730 165800 59740
rect 165900 59730 165980 59740
rect 166080 59730 166160 59740
rect 166260 59730 166340 59740
rect 166440 59730 166520 59740
rect 166620 59730 166700 59740
rect 166800 59730 166880 59740
rect 166980 59730 167060 59740
rect 167160 59730 167240 59740
rect 167340 59730 167420 59740
rect 167520 59730 167600 59740
rect 167700 59730 167780 59740
rect 167880 59730 167960 59740
rect 168060 59730 168140 59740
rect 168240 59730 168320 59740
rect 168420 59730 168500 59740
rect 168600 59730 168680 59740
rect 168780 59730 168860 59740
rect 168960 59730 169040 59740
rect 169140 59730 169220 59740
rect 169320 59730 169400 59740
rect 169500 59730 169580 59740
rect 169680 59730 169760 59740
rect 169860 59730 169940 59740
rect 170040 59730 170120 59740
rect 153060 59650 153070 59670
rect 153240 59650 153250 59670
rect 153420 59650 153430 59670
rect 153600 59650 153610 59670
rect 153780 59650 153790 59670
rect 153960 59650 153970 59670
rect 154140 59650 154150 59670
rect 154320 59650 154330 59670
rect 154500 59650 154510 59670
rect 154680 59650 154690 59670
rect 154860 59650 154870 59670
rect 155040 59650 155050 59670
rect 155220 59650 155230 59670
rect 155400 59650 155410 59670
rect 155580 59650 155590 59670
rect 155760 59650 155770 59670
rect 155940 59650 155950 59670
rect 156120 59650 156130 59670
rect 156300 59650 156310 59670
rect 156480 59650 156490 59670
rect 156660 59650 156670 59670
rect 156840 59650 156850 59670
rect 157020 59650 157030 59670
rect 157200 59650 157210 59670
rect 157380 59650 157390 59670
rect 157560 59650 157570 59670
rect 157740 59650 157750 59670
rect 157920 59650 157930 59670
rect 158100 59650 158110 59670
rect 158280 59650 158290 59670
rect 158460 59650 158470 59670
rect 158640 59650 158650 59670
rect 158820 59650 158830 59670
rect 152100 59620 152160 59650
rect 152220 59620 152280 59650
rect 152340 59620 152400 59650
rect 152980 59580 153060 59590
rect 153160 59580 153240 59590
rect 153340 59580 153420 59590
rect 153520 59580 153600 59590
rect 153700 59580 153780 59590
rect 153880 59580 153960 59590
rect 154060 59580 154140 59590
rect 154240 59580 154320 59590
rect 154420 59580 154500 59590
rect 154600 59580 154680 59590
rect 154780 59580 154860 59590
rect 154960 59580 155040 59590
rect 155140 59580 155220 59590
rect 155320 59580 155400 59590
rect 155500 59580 155580 59590
rect 155680 59580 155760 59590
rect 155860 59580 155940 59590
rect 156040 59580 156120 59590
rect 156220 59580 156300 59590
rect 156400 59580 156480 59590
rect 156580 59580 156660 59590
rect 156760 59580 156840 59590
rect 156940 59580 157020 59590
rect 157120 59580 157200 59590
rect 157300 59580 157380 59590
rect 157480 59580 157560 59590
rect 157660 59580 157740 59590
rect 157840 59580 157920 59590
rect 158020 59580 158100 59590
rect 158200 59580 158280 59590
rect 158380 59580 158460 59590
rect 158560 59580 158640 59590
rect 158740 59580 158820 59590
rect 149880 59550 149940 59580
rect 152220 59530 152250 59560
rect 152340 59530 152370 59560
rect 152100 59500 152160 59530
rect 152220 59500 152280 59530
rect 152340 59500 152400 59530
rect 153060 59500 153070 59580
rect 153240 59500 153250 59580
rect 153420 59500 153430 59580
rect 153600 59500 153610 59580
rect 153780 59500 153790 59580
rect 153960 59500 153970 59580
rect 154140 59500 154150 59580
rect 154320 59500 154330 59580
rect 154500 59500 154510 59580
rect 154680 59500 154690 59580
rect 154860 59500 154870 59580
rect 155040 59500 155050 59580
rect 155220 59500 155230 59580
rect 155400 59500 155410 59580
rect 155580 59500 155590 59580
rect 155760 59500 155770 59580
rect 155940 59500 155950 59580
rect 156120 59500 156130 59580
rect 156300 59500 156310 59580
rect 156480 59500 156490 59580
rect 156660 59500 156670 59580
rect 156840 59500 156850 59580
rect 157020 59500 157030 59580
rect 157200 59500 157210 59580
rect 157380 59500 157390 59580
rect 157560 59500 157570 59580
rect 157740 59500 157750 59580
rect 157920 59500 157930 59580
rect 158100 59500 158110 59580
rect 158280 59500 158290 59580
rect 158460 59500 158470 59580
rect 158640 59500 158650 59580
rect 158820 59500 158830 59580
rect 149880 59430 149940 59460
rect 158900 59440 158990 59670
rect 159520 59650 159550 59680
rect 159640 59650 159670 59680
rect 163520 59650 163550 59680
rect 163640 59650 163670 59680
rect 164360 59650 164370 59730
rect 164540 59650 164550 59730
rect 164720 59650 164730 59730
rect 164900 59650 164910 59730
rect 165080 59650 165090 59730
rect 165260 59650 165270 59730
rect 165440 59650 165450 59730
rect 165620 59650 165630 59730
rect 165800 59650 165810 59730
rect 165980 59650 165990 59730
rect 166160 59650 166170 59730
rect 166340 59650 166350 59730
rect 166520 59650 166530 59730
rect 166700 59650 166710 59730
rect 166880 59650 166890 59730
rect 167060 59650 167070 59730
rect 167240 59650 167250 59730
rect 167420 59650 167430 59730
rect 167600 59650 167610 59730
rect 167780 59650 167790 59730
rect 167960 59650 167970 59730
rect 168140 59650 168150 59730
rect 168320 59650 168330 59730
rect 168500 59650 168510 59730
rect 168680 59650 168690 59730
rect 168860 59650 168870 59730
rect 169040 59650 169050 59730
rect 169220 59650 169230 59730
rect 169400 59650 169410 59730
rect 169580 59650 169590 59730
rect 169760 59650 169770 59730
rect 169940 59650 169950 59730
rect 170120 59650 170130 59730
rect 170810 59650 170840 59680
rect 170930 59650 170960 59680
rect 159400 59620 159460 59650
rect 159520 59620 159580 59650
rect 159640 59620 159700 59650
rect 163400 59620 163460 59650
rect 163520 59620 163580 59650
rect 163640 59620 163700 59650
rect 170690 59620 170750 59650
rect 170810 59620 170870 59650
rect 170930 59620 170990 59650
rect 164280 59580 164360 59590
rect 164460 59580 164540 59590
rect 164640 59580 164720 59590
rect 164820 59580 164900 59590
rect 165000 59580 165080 59590
rect 165180 59580 165260 59590
rect 165360 59580 165440 59590
rect 165540 59580 165620 59590
rect 165720 59580 165800 59590
rect 165900 59580 165980 59590
rect 166080 59580 166160 59590
rect 166260 59580 166340 59590
rect 166440 59580 166520 59590
rect 166620 59580 166700 59590
rect 166800 59580 166880 59590
rect 166980 59580 167060 59590
rect 167160 59580 167240 59590
rect 167340 59580 167420 59590
rect 167520 59580 167600 59590
rect 167700 59580 167780 59590
rect 167880 59580 167960 59590
rect 168060 59580 168140 59590
rect 168240 59580 168320 59590
rect 168420 59580 168500 59590
rect 168600 59580 168680 59590
rect 168780 59580 168860 59590
rect 168960 59580 169040 59590
rect 169140 59580 169220 59590
rect 169320 59580 169400 59590
rect 169500 59580 169580 59590
rect 169680 59580 169760 59590
rect 169860 59580 169940 59590
rect 170040 59580 170120 59590
rect 159520 59530 159550 59560
rect 159640 59530 159670 59560
rect 163520 59530 163550 59560
rect 163640 59530 163670 59560
rect 159400 59500 159460 59530
rect 159520 59500 159580 59530
rect 159640 59500 159700 59530
rect 163400 59500 163460 59530
rect 163520 59500 163580 59530
rect 163640 59500 163700 59530
rect 164360 59500 164370 59580
rect 164540 59500 164550 59580
rect 164720 59500 164730 59580
rect 164900 59500 164910 59580
rect 165080 59500 165090 59580
rect 165260 59500 165270 59580
rect 165440 59500 165450 59580
rect 165620 59500 165630 59580
rect 165800 59500 165810 59580
rect 165980 59500 165990 59580
rect 166160 59500 166170 59580
rect 166340 59500 166350 59580
rect 166520 59500 166530 59580
rect 166700 59500 166710 59580
rect 166880 59500 166890 59580
rect 167060 59500 167070 59580
rect 167240 59500 167250 59580
rect 167420 59500 167430 59580
rect 167600 59500 167610 59580
rect 167780 59500 167790 59580
rect 167960 59500 167970 59580
rect 168140 59500 168150 59580
rect 168320 59500 168330 59580
rect 168500 59500 168510 59580
rect 168680 59500 168690 59580
rect 168860 59500 168870 59580
rect 169040 59500 169050 59580
rect 169220 59500 169230 59580
rect 169400 59500 169410 59580
rect 169580 59500 169590 59580
rect 169760 59500 169770 59580
rect 169940 59500 169950 59580
rect 170120 59500 170130 59580
rect 170810 59530 170840 59560
rect 170930 59530 170960 59560
rect 170690 59500 170750 59530
rect 170810 59500 170870 59530
rect 170930 59500 170990 59530
rect 152220 59410 152250 59440
rect 152340 59410 152370 59440
rect 152900 59410 158990 59440
rect 159520 59410 159550 59440
rect 159640 59410 159670 59440
rect 163520 59410 163550 59440
rect 163640 59410 163670 59440
rect 164280 59430 164360 59440
rect 164460 59430 164540 59440
rect 164640 59430 164720 59440
rect 164820 59430 164900 59440
rect 165000 59430 165080 59440
rect 165180 59430 165260 59440
rect 165360 59430 165440 59440
rect 165540 59430 165620 59440
rect 165720 59430 165800 59440
rect 165900 59430 165980 59440
rect 166080 59430 166160 59440
rect 166260 59430 166340 59440
rect 166440 59430 166520 59440
rect 166620 59430 166700 59440
rect 166800 59430 166880 59440
rect 166980 59430 167060 59440
rect 167160 59430 167240 59440
rect 167340 59430 167420 59440
rect 167520 59430 167600 59440
rect 167700 59430 167780 59440
rect 167880 59430 167960 59440
rect 168060 59430 168140 59440
rect 168240 59430 168320 59440
rect 168420 59430 168500 59440
rect 168600 59430 168680 59440
rect 168780 59430 168860 59440
rect 168960 59430 169040 59440
rect 169140 59430 169220 59440
rect 169320 59430 169400 59440
rect 169500 59430 169580 59440
rect 169680 59430 169760 59440
rect 169860 59430 169940 59440
rect 170040 59430 170120 59440
rect 152100 59380 152160 59410
rect 152220 59380 152280 59410
rect 152340 59380 152400 59410
rect 153060 59350 153070 59410
rect 153240 59350 153250 59410
rect 153420 59350 153430 59410
rect 153600 59350 153610 59410
rect 153780 59350 153790 59410
rect 153960 59350 153970 59410
rect 154140 59350 154150 59410
rect 154320 59350 154330 59410
rect 154500 59350 154510 59410
rect 154680 59350 154690 59410
rect 154860 59350 154870 59410
rect 155040 59350 155050 59410
rect 155220 59350 155230 59410
rect 155400 59350 155410 59410
rect 155580 59350 155590 59410
rect 155760 59350 155770 59410
rect 155940 59350 155950 59410
rect 156120 59350 156130 59410
rect 156300 59350 156310 59410
rect 156480 59350 156490 59410
rect 156660 59350 156670 59410
rect 156840 59350 156850 59410
rect 157020 59350 157030 59410
rect 157200 59350 157210 59410
rect 157380 59350 157390 59410
rect 157560 59350 157570 59410
rect 157740 59350 157750 59410
rect 157920 59350 157930 59410
rect 158100 59350 158110 59410
rect 158280 59350 158290 59410
rect 158460 59350 158470 59410
rect 158640 59350 158650 59410
rect 158820 59350 158830 59410
rect 158900 59340 158990 59410
rect 159400 59380 159460 59410
rect 159520 59380 159580 59410
rect 159640 59380 159700 59410
rect 163400 59380 163460 59410
rect 163520 59380 163580 59410
rect 163640 59380 163700 59410
rect 164360 59350 164370 59430
rect 164540 59350 164550 59430
rect 164720 59350 164730 59430
rect 164900 59350 164910 59430
rect 165080 59350 165090 59430
rect 165260 59350 165270 59430
rect 165440 59350 165450 59430
rect 165620 59350 165630 59430
rect 165800 59350 165810 59430
rect 165980 59350 165990 59430
rect 166160 59350 166170 59430
rect 166340 59350 166350 59430
rect 166520 59350 166530 59430
rect 166700 59350 166710 59430
rect 166880 59350 166890 59430
rect 167060 59350 167070 59430
rect 167240 59350 167250 59430
rect 167420 59350 167430 59430
rect 167600 59350 167610 59430
rect 167780 59350 167790 59430
rect 167960 59350 167970 59430
rect 168140 59350 168150 59430
rect 168320 59350 168330 59430
rect 168500 59350 168510 59430
rect 168680 59350 168690 59430
rect 168860 59350 168870 59430
rect 169040 59350 169050 59430
rect 169220 59350 169230 59430
rect 169400 59350 169410 59430
rect 169580 59350 169590 59430
rect 169760 59350 169770 59430
rect 169940 59350 169950 59430
rect 170120 59350 170130 59430
rect 170810 59410 170840 59440
rect 170930 59410 170960 59440
rect 170690 59380 170750 59410
rect 170810 59380 170870 59410
rect 170930 59380 170990 59410
rect 149880 59310 149940 59340
rect 152220 59290 152250 59320
rect 152340 59290 152370 59320
rect 152900 59310 158990 59340
rect 158900 59300 158990 59310
rect 152900 59290 158990 59300
rect 159520 59290 159550 59320
rect 159640 59290 159670 59320
rect 163520 59290 163550 59320
rect 163640 59290 163670 59320
rect 164200 59290 170200 59300
rect 170810 59290 170840 59320
rect 170930 59290 170960 59320
rect 152100 59260 152160 59290
rect 152220 59260 152280 59290
rect 152340 59260 152400 59290
rect 149880 59190 149940 59220
rect 152220 59170 152250 59200
rect 152340 59170 152370 59200
rect 152100 59140 152160 59170
rect 152220 59140 152280 59170
rect 152340 59140 152400 59170
rect 152980 59110 153060 59120
rect 153160 59110 153240 59120
rect 153340 59110 153420 59120
rect 153520 59110 153600 59120
rect 153700 59110 153780 59120
rect 153880 59110 153960 59120
rect 154060 59110 154140 59120
rect 154240 59110 154320 59120
rect 154420 59110 154500 59120
rect 154600 59110 154680 59120
rect 154780 59110 154860 59120
rect 154960 59110 155040 59120
rect 155140 59110 155220 59120
rect 155320 59110 155400 59120
rect 155500 59110 155580 59120
rect 155680 59110 155760 59120
rect 155860 59110 155940 59120
rect 156040 59110 156120 59120
rect 156220 59110 156300 59120
rect 156400 59110 156480 59120
rect 156580 59110 156660 59120
rect 156760 59110 156840 59120
rect 156940 59110 157020 59120
rect 157120 59110 157200 59120
rect 157300 59110 157380 59120
rect 157480 59110 157560 59120
rect 157660 59110 157740 59120
rect 157840 59110 157920 59120
rect 158020 59110 158100 59120
rect 158200 59110 158280 59120
rect 158380 59110 158460 59120
rect 158560 59110 158640 59120
rect 158740 59110 158820 59120
rect 149880 59070 149940 59100
rect 152220 59050 152250 59080
rect 152340 59050 152370 59080
rect 152100 59020 152160 59050
rect 152220 59020 152280 59050
rect 152340 59020 152400 59050
rect 153060 59030 153070 59110
rect 153240 59030 153250 59110
rect 153420 59030 153430 59110
rect 153600 59030 153610 59110
rect 153780 59030 153790 59110
rect 153960 59030 153970 59110
rect 154140 59030 154150 59110
rect 154320 59030 154330 59110
rect 154500 59030 154510 59110
rect 154680 59030 154690 59110
rect 154860 59030 154870 59110
rect 155040 59030 155050 59110
rect 155220 59030 155230 59110
rect 155400 59030 155410 59110
rect 155580 59030 155590 59110
rect 155760 59030 155770 59110
rect 155940 59030 155950 59110
rect 156120 59030 156130 59110
rect 156300 59030 156310 59110
rect 156480 59030 156490 59110
rect 156660 59030 156670 59110
rect 156840 59030 156850 59110
rect 157020 59030 157030 59110
rect 157200 59030 157210 59110
rect 157380 59030 157390 59110
rect 157560 59030 157570 59110
rect 157740 59030 157750 59110
rect 157920 59030 157930 59110
rect 158100 59030 158110 59110
rect 158280 59030 158290 59110
rect 158460 59030 158470 59110
rect 158640 59030 158650 59110
rect 158820 59030 158830 59110
rect 149880 58950 149940 58980
rect 152220 58930 152250 58960
rect 152340 58930 152370 58960
rect 152100 58900 152160 58930
rect 152220 58900 152280 58930
rect 152340 58900 152400 58930
rect 149880 58830 149940 58860
rect 152220 58810 152250 58840
rect 152340 58810 152370 58840
rect 152100 58780 152160 58810
rect 152220 58780 152280 58810
rect 152340 58780 152400 58810
rect 152980 58790 153060 58800
rect 153160 58790 153240 58800
rect 153340 58790 153420 58800
rect 153520 58790 153600 58800
rect 153700 58790 153780 58800
rect 153880 58790 153960 58800
rect 154060 58790 154140 58800
rect 154240 58790 154320 58800
rect 154420 58790 154500 58800
rect 154600 58790 154680 58800
rect 154780 58790 154860 58800
rect 154960 58790 155040 58800
rect 155140 58790 155220 58800
rect 155320 58790 155400 58800
rect 155500 58790 155580 58800
rect 155680 58790 155760 58800
rect 155860 58790 155940 58800
rect 156040 58790 156120 58800
rect 156220 58790 156300 58800
rect 156400 58790 156480 58800
rect 156580 58790 156660 58800
rect 156760 58790 156840 58800
rect 156940 58790 157020 58800
rect 157120 58790 157200 58800
rect 157300 58790 157380 58800
rect 157480 58790 157560 58800
rect 157660 58790 157740 58800
rect 157840 58790 157920 58800
rect 158020 58790 158100 58800
rect 158200 58790 158280 58800
rect 158380 58790 158460 58800
rect 158560 58790 158640 58800
rect 158740 58790 158820 58800
rect 149880 58710 149940 58740
rect 152220 58690 152250 58720
rect 152340 58690 152370 58720
rect 153060 58710 153070 58790
rect 153240 58710 153250 58790
rect 153420 58710 153430 58790
rect 153600 58710 153610 58790
rect 153780 58710 153790 58790
rect 153960 58710 153970 58790
rect 154140 58710 154150 58790
rect 154320 58710 154330 58790
rect 154500 58710 154510 58790
rect 154680 58710 154690 58790
rect 154860 58710 154870 58790
rect 155040 58710 155050 58790
rect 155220 58710 155230 58790
rect 155400 58710 155410 58790
rect 155580 58710 155590 58790
rect 155760 58710 155770 58790
rect 155940 58710 155950 58790
rect 156120 58710 156130 58790
rect 156300 58710 156310 58790
rect 156480 58710 156490 58790
rect 156660 58710 156670 58790
rect 156840 58710 156850 58790
rect 157020 58710 157030 58790
rect 157200 58710 157210 58790
rect 157380 58710 157390 58790
rect 157560 58710 157570 58790
rect 157740 58710 157750 58790
rect 157920 58710 157930 58790
rect 158100 58710 158110 58790
rect 158280 58710 158290 58790
rect 158460 58710 158470 58790
rect 158640 58710 158650 58790
rect 158820 58710 158830 58790
rect 152100 58660 152160 58690
rect 152220 58660 152280 58690
rect 152340 58660 152400 58690
rect 158900 58620 158990 59290
rect 159400 59260 159460 59290
rect 159520 59260 159580 59290
rect 159640 59260 159700 59290
rect 163400 59260 163460 59290
rect 163520 59260 163580 59290
rect 163640 59260 163700 59290
rect 170690 59260 170750 59290
rect 170810 59260 170870 59290
rect 170930 59260 170990 59290
rect 159520 59170 159550 59200
rect 159640 59170 159670 59200
rect 163520 59170 163550 59200
rect 163640 59170 163670 59200
rect 170810 59170 170840 59200
rect 170930 59170 170960 59200
rect 159400 59140 159460 59170
rect 159520 59140 159580 59170
rect 159640 59140 159700 59170
rect 163400 59140 163460 59170
rect 163520 59140 163580 59170
rect 163640 59140 163700 59170
rect 170690 59140 170750 59170
rect 170810 59140 170870 59170
rect 170930 59140 170990 59170
rect 164280 59110 164360 59120
rect 164460 59110 164540 59120
rect 164640 59110 164720 59120
rect 164820 59110 164900 59120
rect 165000 59110 165080 59120
rect 165180 59110 165260 59120
rect 165360 59110 165440 59120
rect 165540 59110 165620 59120
rect 165720 59110 165800 59120
rect 165900 59110 165980 59120
rect 166080 59110 166160 59120
rect 166260 59110 166340 59120
rect 166440 59110 166520 59120
rect 166620 59110 166700 59120
rect 166800 59110 166880 59120
rect 166980 59110 167060 59120
rect 167160 59110 167240 59120
rect 167340 59110 167420 59120
rect 167520 59110 167600 59120
rect 167700 59110 167780 59120
rect 167880 59110 167960 59120
rect 168060 59110 168140 59120
rect 168240 59110 168320 59120
rect 168420 59110 168500 59120
rect 168600 59110 168680 59120
rect 168780 59110 168860 59120
rect 168960 59110 169040 59120
rect 169140 59110 169220 59120
rect 169320 59110 169400 59120
rect 169500 59110 169580 59120
rect 169680 59110 169760 59120
rect 169860 59110 169940 59120
rect 170040 59110 170120 59120
rect 159520 59050 159550 59080
rect 159640 59050 159670 59080
rect 163520 59050 163550 59080
rect 163640 59050 163670 59080
rect 159400 59020 159460 59050
rect 159520 59020 159580 59050
rect 159640 59020 159700 59050
rect 163400 59020 163460 59050
rect 163520 59020 163580 59050
rect 163640 59020 163700 59050
rect 164360 59030 164370 59110
rect 164540 59030 164550 59110
rect 164720 59030 164730 59110
rect 164900 59030 164910 59110
rect 165080 59030 165090 59110
rect 165260 59030 165270 59110
rect 165440 59030 165450 59110
rect 165620 59030 165630 59110
rect 165800 59030 165810 59110
rect 165980 59030 165990 59110
rect 166160 59030 166170 59110
rect 166340 59030 166350 59110
rect 166520 59030 166530 59110
rect 166700 59030 166710 59110
rect 166880 59030 166890 59110
rect 167060 59030 167070 59110
rect 167240 59030 167250 59110
rect 167420 59030 167430 59110
rect 167600 59030 167610 59110
rect 167780 59030 167790 59110
rect 167960 59030 167970 59110
rect 168140 59030 168150 59110
rect 168320 59030 168330 59110
rect 168500 59030 168510 59110
rect 168680 59030 168690 59110
rect 168860 59030 168870 59110
rect 169040 59030 169050 59110
rect 169220 59030 169230 59110
rect 169400 59030 169410 59110
rect 169580 59030 169590 59110
rect 169760 59030 169770 59110
rect 169940 59030 169950 59110
rect 170120 59030 170130 59110
rect 170810 59050 170840 59080
rect 170930 59050 170960 59080
rect 170690 59020 170750 59050
rect 170810 59020 170870 59050
rect 170930 59020 170990 59050
rect 159520 58930 159550 58960
rect 159640 58930 159670 58960
rect 163520 58930 163550 58960
rect 163640 58930 163670 58960
rect 170810 58930 170840 58960
rect 170930 58930 170960 58960
rect 159400 58900 159460 58930
rect 159520 58900 159580 58930
rect 159640 58900 159700 58930
rect 163400 58900 163460 58930
rect 163520 58900 163580 58930
rect 163640 58900 163700 58930
rect 170690 58900 170750 58930
rect 170810 58900 170870 58930
rect 170930 58900 170990 58930
rect 159520 58810 159550 58840
rect 159640 58810 159670 58840
rect 163520 58810 163550 58840
rect 163640 58810 163670 58840
rect 164280 58810 164360 58820
rect 164460 58810 164540 58820
rect 164640 58810 164720 58820
rect 164820 58810 164900 58820
rect 165000 58810 165080 58820
rect 165180 58810 165260 58820
rect 165360 58810 165440 58820
rect 165540 58810 165620 58820
rect 165720 58810 165800 58820
rect 165900 58810 165980 58820
rect 166080 58810 166160 58820
rect 166260 58810 166340 58820
rect 166440 58810 166520 58820
rect 166620 58810 166700 58820
rect 166800 58810 166880 58820
rect 166980 58810 167060 58820
rect 167160 58810 167240 58820
rect 167340 58810 167420 58820
rect 167520 58810 167600 58820
rect 167700 58810 167780 58820
rect 167880 58810 167960 58820
rect 168060 58810 168140 58820
rect 168240 58810 168320 58820
rect 168420 58810 168500 58820
rect 168600 58810 168680 58820
rect 168780 58810 168860 58820
rect 168960 58810 169040 58820
rect 169140 58810 169220 58820
rect 169320 58810 169400 58820
rect 169500 58810 169580 58820
rect 169680 58810 169760 58820
rect 169860 58810 169940 58820
rect 170040 58810 170120 58820
rect 170810 58810 170840 58840
rect 170930 58810 170960 58840
rect 159400 58780 159460 58810
rect 159520 58780 159580 58810
rect 159640 58780 159700 58810
rect 163400 58780 163460 58810
rect 163520 58780 163580 58810
rect 163640 58780 163700 58810
rect 164360 58730 164370 58810
rect 164540 58730 164550 58810
rect 164720 58730 164730 58810
rect 164900 58730 164910 58810
rect 165080 58730 165090 58810
rect 165260 58730 165270 58810
rect 165440 58730 165450 58810
rect 165620 58730 165630 58810
rect 165800 58730 165810 58810
rect 165980 58730 165990 58810
rect 166160 58730 166170 58810
rect 166340 58730 166350 58810
rect 166520 58730 166530 58810
rect 166700 58730 166710 58810
rect 166880 58730 166890 58810
rect 167060 58730 167070 58810
rect 167240 58730 167250 58810
rect 167420 58730 167430 58810
rect 167600 58730 167610 58810
rect 167780 58730 167790 58810
rect 167960 58730 167970 58810
rect 168140 58730 168150 58810
rect 168320 58730 168330 58810
rect 168500 58730 168510 58810
rect 168680 58730 168690 58810
rect 168860 58730 168870 58810
rect 169040 58730 169050 58810
rect 169220 58730 169230 58810
rect 169400 58730 169410 58810
rect 169580 58730 169590 58810
rect 169760 58730 169770 58810
rect 169940 58730 169950 58810
rect 170120 58730 170130 58810
rect 170690 58780 170750 58810
rect 170810 58780 170870 58810
rect 170930 58780 170990 58810
rect 159520 58690 159550 58720
rect 159640 58690 159670 58720
rect 163520 58690 163550 58720
rect 163640 58690 163670 58720
rect 170810 58690 170840 58720
rect 170930 58690 170960 58720
rect 159400 58660 159460 58690
rect 159520 58660 159580 58690
rect 159640 58660 159700 58690
rect 163400 58660 163460 58690
rect 163520 58660 163580 58690
rect 163640 58660 163700 58690
rect 170690 58660 170750 58690
rect 170810 58660 170870 58690
rect 170930 58660 170990 58690
rect 149880 58590 149940 58620
rect 152900 58610 158990 58620
rect 164200 58610 170200 58620
rect 152220 58570 152250 58600
rect 152340 58570 152370 58600
rect 152100 58540 152160 58570
rect 152220 58540 152280 58570
rect 152340 58540 152400 58570
rect 158900 58510 158990 58610
rect 159520 58570 159550 58600
rect 159640 58570 159670 58600
rect 163520 58570 163550 58600
rect 163640 58570 163670 58600
rect 170810 58570 170840 58600
rect 170930 58570 170960 58600
rect 159400 58540 159460 58570
rect 159520 58540 159580 58570
rect 159640 58540 159700 58570
rect 163400 58540 163460 58570
rect 163520 58540 163580 58570
rect 163640 58540 163700 58570
rect 170690 58540 170750 58570
rect 170810 58540 170870 58570
rect 170930 58540 170990 58570
rect 149880 58470 149940 58500
rect 152900 58480 158990 58510
rect 152220 58450 152250 58480
rect 152340 58450 152370 58480
rect 152980 58470 153060 58480
rect 153160 58470 153240 58480
rect 153340 58470 153420 58480
rect 153520 58470 153600 58480
rect 153700 58470 153780 58480
rect 153880 58470 153960 58480
rect 154060 58470 154140 58480
rect 154240 58470 154320 58480
rect 154420 58470 154500 58480
rect 154600 58470 154680 58480
rect 154780 58470 154860 58480
rect 154960 58470 155040 58480
rect 155140 58470 155220 58480
rect 155320 58470 155400 58480
rect 155500 58470 155580 58480
rect 155680 58470 155760 58480
rect 155860 58470 155940 58480
rect 156040 58470 156120 58480
rect 156220 58470 156300 58480
rect 156400 58470 156480 58480
rect 156580 58470 156660 58480
rect 156760 58470 156840 58480
rect 156940 58470 157020 58480
rect 157120 58470 157200 58480
rect 157300 58470 157380 58480
rect 157480 58470 157560 58480
rect 157660 58470 157740 58480
rect 157840 58470 157920 58480
rect 158020 58470 158100 58480
rect 158200 58470 158280 58480
rect 158380 58470 158460 58480
rect 158560 58470 158640 58480
rect 158740 58470 158820 58480
rect 152100 58420 152160 58450
rect 152220 58420 152280 58450
rect 152340 58420 152400 58450
rect 153060 58410 153070 58470
rect 153240 58410 153250 58470
rect 153420 58410 153430 58470
rect 153600 58410 153610 58470
rect 153780 58410 153790 58470
rect 153960 58410 153970 58470
rect 154140 58410 154150 58470
rect 154320 58410 154330 58470
rect 154500 58410 154510 58470
rect 154680 58410 154690 58470
rect 154860 58410 154870 58470
rect 155040 58410 155050 58470
rect 155220 58410 155230 58470
rect 155400 58410 155410 58470
rect 155580 58410 155590 58470
rect 155760 58410 155770 58470
rect 155940 58410 155950 58470
rect 156120 58410 156130 58470
rect 156300 58410 156310 58470
rect 156480 58410 156490 58470
rect 156660 58410 156670 58470
rect 156840 58410 156850 58470
rect 157020 58410 157030 58470
rect 157200 58410 157210 58470
rect 157380 58410 157390 58470
rect 157560 58410 157570 58470
rect 157740 58410 157750 58470
rect 157920 58410 157930 58470
rect 158100 58410 158110 58470
rect 158280 58410 158290 58470
rect 158460 58410 158470 58470
rect 158640 58410 158650 58470
rect 158820 58410 158830 58470
rect 158900 58410 158990 58480
rect 159520 58450 159550 58480
rect 159640 58450 159670 58480
rect 163520 58450 163550 58480
rect 163640 58450 163670 58480
rect 164280 58470 164360 58480
rect 164460 58470 164540 58480
rect 164640 58470 164720 58480
rect 164820 58470 164900 58480
rect 165000 58470 165080 58480
rect 165180 58470 165260 58480
rect 165360 58470 165440 58480
rect 165540 58470 165620 58480
rect 165720 58470 165800 58480
rect 165900 58470 165980 58480
rect 166080 58470 166160 58480
rect 166260 58470 166340 58480
rect 166440 58470 166520 58480
rect 166620 58470 166700 58480
rect 166800 58470 166880 58480
rect 166980 58470 167060 58480
rect 167160 58470 167240 58480
rect 167340 58470 167420 58480
rect 167520 58470 167600 58480
rect 167700 58470 167780 58480
rect 167880 58470 167960 58480
rect 168060 58470 168140 58480
rect 168240 58470 168320 58480
rect 168420 58470 168500 58480
rect 168600 58470 168680 58480
rect 168780 58470 168860 58480
rect 168960 58470 169040 58480
rect 169140 58470 169220 58480
rect 169320 58470 169400 58480
rect 169500 58470 169580 58480
rect 169680 58470 169760 58480
rect 169860 58470 169940 58480
rect 170040 58470 170120 58480
rect 159400 58420 159460 58450
rect 159520 58420 159580 58450
rect 159640 58420 159700 58450
rect 163400 58420 163460 58450
rect 163520 58420 163580 58450
rect 163640 58420 163700 58450
rect 152900 58380 158990 58410
rect 164360 58390 164370 58470
rect 164540 58390 164550 58470
rect 164720 58390 164730 58470
rect 164900 58390 164910 58470
rect 165080 58390 165090 58470
rect 165260 58390 165270 58470
rect 165440 58390 165450 58470
rect 165620 58390 165630 58470
rect 165800 58390 165810 58470
rect 165980 58390 165990 58470
rect 166160 58390 166170 58470
rect 166340 58390 166350 58470
rect 166520 58390 166530 58470
rect 166700 58390 166710 58470
rect 166880 58390 166890 58470
rect 167060 58390 167070 58470
rect 167240 58390 167250 58470
rect 167420 58390 167430 58470
rect 167600 58390 167610 58470
rect 167780 58390 167790 58470
rect 167960 58390 167970 58470
rect 168140 58390 168150 58470
rect 168320 58390 168330 58470
rect 168500 58390 168510 58470
rect 168680 58390 168690 58470
rect 168860 58390 168870 58470
rect 169040 58390 169050 58470
rect 169220 58390 169230 58470
rect 169400 58390 169410 58470
rect 169580 58390 169590 58470
rect 169760 58390 169770 58470
rect 169940 58390 169950 58470
rect 170120 58390 170130 58470
rect 170810 58450 170840 58480
rect 170930 58450 170960 58480
rect 170690 58420 170750 58450
rect 170810 58420 170870 58450
rect 170930 58420 170990 58450
rect 149880 58350 149940 58380
rect 152220 58330 152250 58360
rect 152340 58330 152370 58360
rect 152100 58300 152160 58330
rect 152220 58300 152280 58330
rect 152340 58300 152400 58330
rect 152980 58320 153060 58330
rect 153160 58320 153240 58330
rect 153340 58320 153420 58330
rect 153520 58320 153600 58330
rect 153700 58320 153780 58330
rect 153880 58320 153960 58330
rect 154060 58320 154140 58330
rect 154240 58320 154320 58330
rect 154420 58320 154500 58330
rect 154600 58320 154680 58330
rect 154780 58320 154860 58330
rect 154960 58320 155040 58330
rect 155140 58320 155220 58330
rect 155320 58320 155400 58330
rect 155500 58320 155580 58330
rect 155680 58320 155760 58330
rect 155860 58320 155940 58330
rect 156040 58320 156120 58330
rect 156220 58320 156300 58330
rect 156400 58320 156480 58330
rect 156580 58320 156660 58330
rect 156760 58320 156840 58330
rect 156940 58320 157020 58330
rect 157120 58320 157200 58330
rect 157300 58320 157380 58330
rect 157480 58320 157560 58330
rect 157660 58320 157740 58330
rect 157840 58320 157920 58330
rect 158020 58320 158100 58330
rect 158200 58320 158280 58330
rect 158380 58320 158460 58330
rect 158560 58320 158640 58330
rect 158740 58320 158820 58330
rect 149880 58230 149940 58260
rect 153060 58240 153070 58320
rect 153240 58240 153250 58320
rect 153420 58240 153430 58320
rect 153600 58240 153610 58320
rect 153780 58240 153790 58320
rect 153960 58240 153970 58320
rect 154140 58240 154150 58320
rect 154320 58240 154330 58320
rect 154500 58240 154510 58320
rect 154680 58240 154690 58320
rect 154860 58240 154870 58320
rect 155040 58240 155050 58320
rect 155220 58240 155230 58320
rect 155400 58240 155410 58320
rect 155580 58240 155590 58320
rect 155760 58240 155770 58320
rect 155940 58240 155950 58320
rect 156120 58240 156130 58320
rect 156300 58240 156310 58320
rect 156480 58240 156490 58320
rect 156660 58240 156670 58320
rect 156840 58240 156850 58320
rect 157020 58240 157030 58320
rect 157200 58240 157210 58320
rect 157380 58240 157390 58320
rect 157560 58240 157570 58320
rect 157740 58240 157750 58320
rect 157920 58240 157930 58320
rect 158100 58240 158110 58320
rect 158280 58240 158290 58320
rect 158460 58240 158470 58320
rect 158640 58240 158650 58320
rect 158820 58240 158830 58320
rect 152220 58210 152250 58240
rect 152340 58210 152370 58240
rect 152100 58180 152160 58210
rect 152220 58180 152280 58210
rect 152340 58180 152400 58210
rect 158900 58180 158990 58380
rect 159520 58330 159550 58360
rect 159640 58330 159670 58360
rect 163520 58330 163550 58360
rect 163640 58330 163670 58360
rect 170810 58330 170840 58360
rect 170930 58330 170960 58360
rect 159400 58300 159460 58330
rect 159520 58300 159580 58330
rect 159640 58300 159700 58330
rect 163400 58300 163460 58330
rect 163520 58300 163580 58330
rect 163640 58300 163700 58330
rect 164280 58320 164360 58330
rect 164460 58320 164540 58330
rect 164640 58320 164720 58330
rect 164820 58320 164900 58330
rect 165000 58320 165080 58330
rect 165180 58320 165260 58330
rect 165360 58320 165440 58330
rect 165540 58320 165620 58330
rect 165720 58320 165800 58330
rect 165900 58320 165980 58330
rect 166080 58320 166160 58330
rect 166260 58320 166340 58330
rect 166440 58320 166520 58330
rect 166620 58320 166700 58330
rect 166800 58320 166880 58330
rect 166980 58320 167060 58330
rect 167160 58320 167240 58330
rect 167340 58320 167420 58330
rect 167520 58320 167600 58330
rect 167700 58320 167780 58330
rect 167880 58320 167960 58330
rect 168060 58320 168140 58330
rect 168240 58320 168320 58330
rect 168420 58320 168500 58330
rect 168600 58320 168680 58330
rect 168780 58320 168860 58330
rect 168960 58320 169040 58330
rect 169140 58320 169220 58330
rect 169320 58320 169400 58330
rect 169500 58320 169580 58330
rect 169680 58320 169760 58330
rect 169860 58320 169940 58330
rect 170040 58320 170120 58330
rect 164360 58240 164370 58320
rect 164540 58240 164550 58320
rect 164720 58240 164730 58320
rect 164900 58240 164910 58320
rect 165080 58240 165090 58320
rect 165260 58240 165270 58320
rect 165440 58240 165450 58320
rect 165620 58240 165630 58320
rect 165800 58240 165810 58320
rect 165980 58240 165990 58320
rect 166160 58240 166170 58320
rect 166340 58240 166350 58320
rect 166520 58240 166530 58320
rect 166700 58240 166710 58320
rect 166880 58240 166890 58320
rect 167060 58240 167070 58320
rect 167240 58240 167250 58320
rect 167420 58240 167430 58320
rect 167600 58240 167610 58320
rect 167780 58240 167790 58320
rect 167960 58240 167970 58320
rect 168140 58240 168150 58320
rect 168320 58240 168330 58320
rect 168500 58240 168510 58320
rect 168680 58240 168690 58320
rect 168860 58240 168870 58320
rect 169040 58240 169050 58320
rect 169220 58240 169230 58320
rect 169400 58240 169410 58320
rect 169580 58240 169590 58320
rect 169760 58240 169770 58320
rect 169940 58240 169950 58320
rect 170120 58240 170130 58320
rect 170690 58300 170750 58330
rect 170810 58300 170870 58330
rect 170930 58300 170990 58330
rect 159520 58210 159550 58240
rect 159640 58210 159670 58240
rect 163520 58210 163550 58240
rect 163640 58210 163670 58240
rect 170810 58210 170840 58240
rect 170930 58210 170960 58240
rect 159400 58180 159460 58210
rect 159520 58180 159580 58210
rect 159640 58180 159700 58210
rect 163400 58180 163460 58210
rect 163520 58180 163580 58210
rect 163640 58180 163700 58210
rect 170690 58180 170750 58210
rect 170810 58180 170870 58210
rect 170930 58180 170990 58210
rect 152900 58150 158990 58180
rect 164280 58170 164360 58180
rect 164460 58170 164540 58180
rect 164640 58170 164720 58180
rect 164820 58170 164900 58180
rect 165000 58170 165080 58180
rect 165180 58170 165260 58180
rect 165360 58170 165440 58180
rect 165540 58170 165620 58180
rect 165720 58170 165800 58180
rect 165900 58170 165980 58180
rect 166080 58170 166160 58180
rect 166260 58170 166340 58180
rect 166440 58170 166520 58180
rect 166620 58170 166700 58180
rect 166800 58170 166880 58180
rect 166980 58170 167060 58180
rect 167160 58170 167240 58180
rect 167340 58170 167420 58180
rect 167520 58170 167600 58180
rect 167700 58170 167780 58180
rect 167880 58170 167960 58180
rect 168060 58170 168140 58180
rect 168240 58170 168320 58180
rect 168420 58170 168500 58180
rect 168600 58170 168680 58180
rect 168780 58170 168860 58180
rect 168960 58170 169040 58180
rect 169140 58170 169220 58180
rect 169320 58170 169400 58180
rect 169500 58170 169580 58180
rect 169680 58170 169760 58180
rect 169860 58170 169940 58180
rect 170040 58170 170120 58180
rect 149880 58110 149940 58140
rect 152220 58090 152250 58120
rect 152340 58090 152370 58120
rect 153060 58090 153070 58150
rect 153240 58090 153250 58150
rect 153420 58090 153430 58150
rect 153600 58090 153610 58150
rect 153780 58090 153790 58150
rect 153960 58090 153970 58150
rect 154140 58090 154150 58150
rect 154320 58090 154330 58150
rect 154500 58090 154510 58150
rect 154680 58090 154690 58150
rect 154860 58090 154870 58150
rect 155040 58090 155050 58150
rect 155220 58090 155230 58150
rect 155400 58090 155410 58150
rect 155580 58090 155590 58150
rect 155760 58090 155770 58150
rect 155940 58090 155950 58150
rect 156120 58090 156130 58150
rect 156300 58090 156310 58150
rect 156480 58090 156490 58150
rect 156660 58090 156670 58150
rect 156840 58090 156850 58150
rect 157020 58090 157030 58150
rect 157200 58090 157210 58150
rect 157380 58090 157390 58150
rect 157560 58090 157570 58150
rect 157740 58090 157750 58150
rect 157920 58090 157930 58150
rect 158100 58090 158110 58150
rect 158280 58090 158290 58150
rect 158460 58090 158470 58150
rect 158640 58090 158650 58150
rect 158820 58090 158830 58150
rect 152100 58060 152160 58090
rect 152220 58060 152280 58090
rect 152340 58060 152400 58090
rect 158900 58080 158990 58150
rect 159520 58090 159550 58120
rect 159640 58090 159670 58120
rect 163520 58090 163550 58120
rect 163640 58090 163670 58120
rect 164360 58090 164370 58170
rect 164540 58090 164550 58170
rect 164720 58090 164730 58170
rect 164900 58090 164910 58170
rect 165080 58090 165090 58170
rect 165260 58090 165270 58170
rect 165440 58090 165450 58170
rect 165620 58090 165630 58170
rect 165800 58090 165810 58170
rect 165980 58090 165990 58170
rect 166160 58090 166170 58170
rect 166340 58090 166350 58170
rect 166520 58090 166530 58170
rect 166700 58090 166710 58170
rect 166880 58090 166890 58170
rect 167060 58090 167070 58170
rect 167240 58090 167250 58170
rect 167420 58090 167430 58170
rect 167600 58090 167610 58170
rect 167780 58090 167790 58170
rect 167960 58090 167970 58170
rect 168140 58090 168150 58170
rect 168320 58090 168330 58170
rect 168500 58090 168510 58170
rect 168680 58090 168690 58170
rect 168860 58090 168870 58170
rect 169040 58090 169050 58170
rect 169220 58090 169230 58170
rect 169400 58090 169410 58170
rect 169580 58090 169590 58170
rect 169760 58090 169770 58170
rect 169940 58090 169950 58170
rect 170120 58090 170130 58170
rect 170810 58090 170840 58120
rect 170930 58090 170960 58120
rect 152900 58050 158990 58080
rect 159400 58060 159460 58090
rect 159520 58060 159580 58090
rect 159640 58060 159700 58090
rect 163400 58060 163460 58090
rect 163520 58060 163580 58090
rect 163640 58060 163700 58090
rect 170690 58060 170750 58090
rect 170810 58060 170870 58090
rect 170930 58060 170990 58090
rect 158900 58040 158990 58050
rect 152900 58030 158990 58040
rect 164200 58030 170200 58040
rect 149880 57990 149940 58020
rect 152220 57970 152250 58000
rect 152340 57970 152370 58000
rect 152100 57940 152160 57970
rect 152220 57940 152280 57970
rect 152340 57940 152400 57970
rect 149880 57870 149940 57900
rect 152220 57850 152250 57880
rect 152340 57850 152370 57880
rect 152980 57850 153060 57860
rect 153160 57850 153240 57860
rect 153340 57850 153420 57860
rect 153520 57850 153600 57860
rect 153700 57850 153780 57860
rect 153880 57850 153960 57860
rect 154060 57850 154140 57860
rect 154240 57850 154320 57860
rect 154420 57850 154500 57860
rect 154600 57850 154680 57860
rect 154780 57850 154860 57860
rect 154960 57850 155040 57860
rect 155140 57850 155220 57860
rect 155320 57850 155400 57860
rect 155500 57850 155580 57860
rect 155680 57850 155760 57860
rect 155860 57850 155940 57860
rect 156040 57850 156120 57860
rect 156220 57850 156300 57860
rect 156400 57850 156480 57860
rect 156580 57850 156660 57860
rect 156760 57850 156840 57860
rect 156940 57850 157020 57860
rect 157120 57850 157200 57860
rect 157300 57850 157380 57860
rect 157480 57850 157560 57860
rect 157660 57850 157740 57860
rect 157840 57850 157920 57860
rect 158020 57850 158100 57860
rect 158200 57850 158280 57860
rect 158380 57850 158460 57860
rect 158560 57850 158640 57860
rect 158740 57850 158820 57860
rect 152100 57820 152160 57850
rect 152220 57820 152280 57850
rect 152340 57820 152400 57850
rect 149880 57750 149940 57780
rect 153060 57770 153070 57850
rect 153240 57770 153250 57850
rect 153420 57770 153430 57850
rect 153600 57770 153610 57850
rect 153780 57770 153790 57850
rect 153960 57770 153970 57850
rect 154140 57770 154150 57850
rect 154320 57770 154330 57850
rect 154500 57770 154510 57850
rect 154680 57770 154690 57850
rect 154860 57770 154870 57850
rect 155040 57770 155050 57850
rect 155220 57770 155230 57850
rect 155400 57770 155410 57850
rect 155580 57770 155590 57850
rect 155760 57770 155770 57850
rect 155940 57770 155950 57850
rect 156120 57770 156130 57850
rect 156300 57770 156310 57850
rect 156480 57770 156490 57850
rect 156660 57770 156670 57850
rect 156840 57770 156850 57850
rect 157020 57770 157030 57850
rect 157200 57770 157210 57850
rect 157380 57770 157390 57850
rect 157560 57770 157570 57850
rect 157740 57770 157750 57850
rect 157920 57770 157930 57850
rect 158100 57770 158110 57850
rect 158280 57770 158290 57850
rect 158460 57770 158470 57850
rect 158640 57770 158650 57850
rect 158820 57770 158830 57850
rect 152220 57730 152250 57760
rect 152340 57730 152370 57760
rect 152100 57700 152160 57730
rect 152220 57700 152280 57730
rect 152340 57700 152400 57730
rect 149880 57630 149940 57660
rect 152220 57610 152250 57640
rect 152340 57610 152370 57640
rect 152100 57580 152160 57610
rect 152220 57580 152280 57610
rect 152340 57580 152400 57610
rect 149880 57510 149940 57540
rect 152980 57530 153060 57540
rect 153160 57530 153240 57540
rect 153340 57530 153420 57540
rect 153520 57530 153600 57540
rect 153700 57530 153780 57540
rect 153880 57530 153960 57540
rect 154060 57530 154140 57540
rect 154240 57530 154320 57540
rect 154420 57530 154500 57540
rect 154600 57530 154680 57540
rect 154780 57530 154860 57540
rect 154960 57530 155040 57540
rect 155140 57530 155220 57540
rect 155320 57530 155400 57540
rect 155500 57530 155580 57540
rect 155680 57530 155760 57540
rect 155860 57530 155940 57540
rect 156040 57530 156120 57540
rect 156220 57530 156300 57540
rect 156400 57530 156480 57540
rect 156580 57530 156660 57540
rect 156760 57530 156840 57540
rect 156940 57530 157020 57540
rect 157120 57530 157200 57540
rect 157300 57530 157380 57540
rect 157480 57530 157560 57540
rect 157660 57530 157740 57540
rect 157840 57530 157920 57540
rect 158020 57530 158100 57540
rect 158200 57530 158280 57540
rect 158380 57530 158460 57540
rect 158560 57530 158640 57540
rect 158740 57530 158820 57540
rect 152220 57490 152250 57520
rect 152340 57490 152370 57520
rect 152100 57460 152160 57490
rect 152220 57460 152280 57490
rect 152340 57460 152400 57490
rect 153060 57450 153070 57530
rect 153240 57450 153250 57530
rect 153420 57450 153430 57530
rect 153600 57450 153610 57530
rect 153780 57450 153790 57530
rect 153960 57450 153970 57530
rect 154140 57450 154150 57530
rect 154320 57450 154330 57530
rect 154500 57450 154510 57530
rect 154680 57450 154690 57530
rect 154860 57450 154870 57530
rect 155040 57450 155050 57530
rect 155220 57450 155230 57530
rect 155400 57450 155410 57530
rect 155580 57450 155590 57530
rect 155760 57450 155770 57530
rect 155940 57450 155950 57530
rect 156120 57450 156130 57530
rect 156300 57450 156310 57530
rect 156480 57450 156490 57530
rect 156660 57450 156670 57530
rect 156840 57450 156850 57530
rect 157020 57450 157030 57530
rect 157200 57450 157210 57530
rect 157380 57450 157390 57530
rect 157560 57450 157570 57530
rect 157740 57450 157750 57530
rect 157920 57450 157930 57530
rect 158100 57450 158110 57530
rect 158280 57450 158290 57530
rect 158460 57450 158470 57530
rect 158640 57450 158650 57530
rect 158820 57450 158830 57530
rect 149880 57390 149940 57420
rect 152220 57370 152250 57400
rect 152340 57370 152370 57400
rect 152100 57340 152160 57370
rect 152220 57340 152280 57370
rect 152340 57340 152400 57370
rect 158900 57360 158990 58030
rect 159520 57970 159550 58000
rect 159640 57970 159670 58000
rect 163520 57970 163550 58000
rect 163640 57970 163670 58000
rect 170810 57970 170840 58000
rect 170930 57970 170960 58000
rect 159400 57940 159460 57970
rect 159520 57940 159580 57970
rect 159640 57940 159700 57970
rect 163400 57940 163460 57970
rect 163520 57940 163580 57970
rect 163640 57940 163700 57970
rect 170690 57940 170750 57970
rect 170810 57940 170870 57970
rect 170930 57940 170990 57970
rect 159520 57850 159550 57880
rect 159640 57850 159670 57880
rect 163520 57850 163550 57880
rect 163640 57850 163670 57880
rect 164280 57850 164360 57860
rect 164460 57850 164540 57860
rect 164640 57850 164720 57860
rect 164820 57850 164900 57860
rect 165000 57850 165080 57860
rect 165180 57850 165260 57860
rect 165360 57850 165440 57860
rect 165540 57850 165620 57860
rect 165720 57850 165800 57860
rect 165900 57850 165980 57860
rect 166080 57850 166160 57860
rect 166260 57850 166340 57860
rect 166440 57850 166520 57860
rect 166620 57850 166700 57860
rect 166800 57850 166880 57860
rect 166980 57850 167060 57860
rect 167160 57850 167240 57860
rect 167340 57850 167420 57860
rect 167520 57850 167600 57860
rect 167700 57850 167780 57860
rect 167880 57850 167960 57860
rect 168060 57850 168140 57860
rect 168240 57850 168320 57860
rect 168420 57850 168500 57860
rect 168600 57850 168680 57860
rect 168780 57850 168860 57860
rect 168960 57850 169040 57860
rect 169140 57850 169220 57860
rect 169320 57850 169400 57860
rect 169500 57850 169580 57860
rect 169680 57850 169760 57860
rect 169860 57850 169940 57860
rect 170040 57850 170120 57860
rect 170810 57850 170840 57880
rect 170930 57850 170960 57880
rect 159400 57820 159460 57850
rect 159520 57820 159580 57850
rect 159640 57820 159700 57850
rect 163400 57820 163460 57850
rect 163520 57820 163580 57850
rect 163640 57820 163700 57850
rect 164360 57770 164370 57850
rect 164540 57770 164550 57850
rect 164720 57770 164730 57850
rect 164900 57770 164910 57850
rect 165080 57770 165090 57850
rect 165260 57770 165270 57850
rect 165440 57770 165450 57850
rect 165620 57770 165630 57850
rect 165800 57770 165810 57850
rect 165980 57770 165990 57850
rect 166160 57770 166170 57850
rect 166340 57770 166350 57850
rect 166520 57770 166530 57850
rect 166700 57770 166710 57850
rect 166880 57770 166890 57850
rect 167060 57770 167070 57850
rect 167240 57770 167250 57850
rect 167420 57770 167430 57850
rect 167600 57770 167610 57850
rect 167780 57770 167790 57850
rect 167960 57770 167970 57850
rect 168140 57770 168150 57850
rect 168320 57770 168330 57850
rect 168500 57770 168510 57850
rect 168680 57770 168690 57850
rect 168860 57770 168870 57850
rect 169040 57770 169050 57850
rect 169220 57770 169230 57850
rect 169400 57770 169410 57850
rect 169580 57770 169590 57850
rect 169760 57770 169770 57850
rect 169940 57770 169950 57850
rect 170120 57770 170130 57850
rect 170690 57820 170750 57850
rect 170810 57820 170870 57850
rect 170930 57820 170990 57850
rect 159520 57730 159550 57760
rect 159640 57730 159670 57760
rect 163520 57730 163550 57760
rect 163640 57730 163670 57760
rect 170810 57730 170840 57760
rect 170930 57730 170960 57760
rect 159400 57700 159460 57730
rect 159520 57700 159580 57730
rect 159640 57700 159700 57730
rect 163400 57700 163460 57730
rect 163520 57700 163580 57730
rect 163640 57700 163700 57730
rect 170690 57700 170750 57730
rect 170810 57700 170870 57730
rect 170930 57700 170990 57730
rect 159520 57610 159550 57640
rect 159640 57610 159670 57640
rect 163520 57610 163550 57640
rect 163640 57610 163670 57640
rect 170810 57610 170840 57640
rect 170930 57610 170960 57640
rect 159400 57580 159460 57610
rect 159520 57580 159580 57610
rect 159640 57580 159700 57610
rect 163400 57580 163460 57610
rect 163520 57580 163580 57610
rect 163640 57580 163700 57610
rect 170690 57580 170750 57610
rect 170810 57580 170870 57610
rect 170930 57580 170990 57610
rect 164280 57550 164360 57560
rect 164460 57550 164540 57560
rect 164640 57550 164720 57560
rect 164820 57550 164900 57560
rect 165000 57550 165080 57560
rect 165180 57550 165260 57560
rect 165360 57550 165440 57560
rect 165540 57550 165620 57560
rect 165720 57550 165800 57560
rect 165900 57550 165980 57560
rect 166080 57550 166160 57560
rect 166260 57550 166340 57560
rect 166440 57550 166520 57560
rect 166620 57550 166700 57560
rect 166800 57550 166880 57560
rect 166980 57550 167060 57560
rect 167160 57550 167240 57560
rect 167340 57550 167420 57560
rect 167520 57550 167600 57560
rect 167700 57550 167780 57560
rect 167880 57550 167960 57560
rect 168060 57550 168140 57560
rect 168240 57550 168320 57560
rect 168420 57550 168500 57560
rect 168600 57550 168680 57560
rect 168780 57550 168860 57560
rect 168960 57550 169040 57560
rect 169140 57550 169220 57560
rect 169320 57550 169400 57560
rect 169500 57550 169580 57560
rect 169680 57550 169760 57560
rect 169860 57550 169940 57560
rect 170040 57550 170120 57560
rect 159520 57490 159550 57520
rect 159640 57490 159670 57520
rect 163520 57490 163550 57520
rect 163640 57490 163670 57520
rect 159400 57460 159460 57490
rect 159520 57460 159580 57490
rect 159640 57460 159700 57490
rect 163400 57460 163460 57490
rect 163520 57460 163580 57490
rect 163640 57460 163700 57490
rect 164360 57470 164370 57550
rect 164540 57470 164550 57550
rect 164720 57470 164730 57550
rect 164900 57470 164910 57550
rect 165080 57470 165090 57550
rect 165260 57470 165270 57550
rect 165440 57470 165450 57550
rect 165620 57470 165630 57550
rect 165800 57470 165810 57550
rect 165980 57470 165990 57550
rect 166160 57470 166170 57550
rect 166340 57470 166350 57550
rect 166520 57470 166530 57550
rect 166700 57470 166710 57550
rect 166880 57470 166890 57550
rect 167060 57470 167070 57550
rect 167240 57470 167250 57550
rect 167420 57470 167430 57550
rect 167600 57470 167610 57550
rect 167780 57470 167790 57550
rect 167960 57470 167970 57550
rect 168140 57470 168150 57550
rect 168320 57470 168330 57550
rect 168500 57470 168510 57550
rect 168680 57470 168690 57550
rect 168860 57470 168870 57550
rect 169040 57470 169050 57550
rect 169220 57470 169230 57550
rect 169400 57470 169410 57550
rect 169580 57470 169590 57550
rect 169760 57470 169770 57550
rect 169940 57470 169950 57550
rect 170120 57470 170130 57550
rect 170810 57490 170840 57520
rect 170930 57490 170960 57520
rect 170690 57460 170750 57490
rect 170810 57460 170870 57490
rect 170930 57460 170990 57490
rect 159520 57370 159550 57400
rect 159640 57370 159670 57400
rect 163520 57370 163550 57400
rect 163640 57370 163670 57400
rect 170810 57370 170840 57400
rect 170930 57370 170960 57400
rect 152900 57350 158990 57360
rect 149880 57270 149940 57300
rect 152220 57250 152250 57280
rect 152340 57250 152370 57280
rect 158900 57250 158990 57350
rect 159400 57340 159460 57370
rect 159520 57340 159580 57370
rect 159640 57340 159700 57370
rect 163400 57340 163460 57370
rect 163520 57340 163580 57370
rect 163640 57340 163700 57370
rect 164200 57350 170200 57360
rect 170690 57340 170750 57370
rect 170810 57340 170870 57370
rect 170930 57340 170990 57370
rect 159520 57250 159550 57280
rect 159640 57250 159670 57280
rect 163520 57250 163550 57280
rect 163640 57250 163670 57280
rect 170810 57250 170840 57280
rect 170930 57250 170960 57280
rect 152100 57220 152160 57250
rect 152220 57220 152280 57250
rect 152340 57220 152400 57250
rect 152900 57220 158990 57250
rect 159400 57220 159460 57250
rect 159520 57220 159580 57250
rect 159640 57220 159700 57250
rect 163400 57220 163460 57250
rect 163520 57220 163580 57250
rect 163640 57220 163700 57250
rect 170690 57220 170750 57250
rect 170810 57220 170870 57250
rect 170930 57220 170990 57250
rect 152980 57210 153060 57220
rect 153160 57210 153240 57220
rect 153340 57210 153420 57220
rect 153520 57210 153600 57220
rect 153700 57210 153780 57220
rect 153880 57210 153960 57220
rect 154060 57210 154140 57220
rect 154240 57210 154320 57220
rect 154420 57210 154500 57220
rect 154600 57210 154680 57220
rect 154780 57210 154860 57220
rect 154960 57210 155040 57220
rect 155140 57210 155220 57220
rect 155320 57210 155400 57220
rect 155500 57210 155580 57220
rect 155680 57210 155760 57220
rect 155860 57210 155940 57220
rect 156040 57210 156120 57220
rect 156220 57210 156300 57220
rect 156400 57210 156480 57220
rect 156580 57210 156660 57220
rect 156760 57210 156840 57220
rect 156940 57210 157020 57220
rect 157120 57210 157200 57220
rect 157300 57210 157380 57220
rect 157480 57210 157560 57220
rect 157660 57210 157740 57220
rect 157840 57210 157920 57220
rect 158020 57210 158100 57220
rect 158200 57210 158280 57220
rect 158380 57210 158460 57220
rect 158560 57210 158640 57220
rect 158740 57210 158820 57220
rect 147580 57150 147640 57180
rect 148400 57150 148460 57180
rect 149880 57150 149940 57180
rect 147178 57080 147318 57150
rect 152220 57130 152250 57160
rect 152340 57130 152370 57160
rect 153060 57150 153070 57210
rect 153240 57150 153250 57210
rect 153420 57150 153430 57210
rect 153600 57150 153610 57210
rect 153780 57150 153790 57210
rect 153960 57150 153970 57210
rect 154140 57150 154150 57210
rect 154320 57150 154330 57210
rect 154500 57150 154510 57210
rect 154680 57150 154690 57210
rect 154860 57150 154870 57210
rect 155040 57150 155050 57210
rect 155220 57150 155230 57210
rect 155400 57150 155410 57210
rect 155580 57150 155590 57210
rect 155760 57150 155770 57210
rect 155940 57150 155950 57210
rect 156120 57150 156130 57210
rect 156300 57150 156310 57210
rect 156480 57150 156490 57210
rect 156660 57150 156670 57210
rect 156840 57150 156850 57210
rect 157020 57150 157030 57210
rect 157200 57150 157210 57210
rect 157380 57150 157390 57210
rect 157560 57150 157570 57210
rect 157740 57150 157750 57210
rect 157920 57150 157930 57210
rect 158100 57150 158110 57210
rect 158280 57150 158290 57210
rect 158460 57150 158470 57210
rect 158640 57150 158650 57210
rect 158820 57150 158830 57210
rect 158900 57150 158990 57220
rect 164280 57210 164360 57220
rect 164460 57210 164540 57220
rect 164640 57210 164720 57220
rect 164820 57210 164900 57220
rect 165000 57210 165080 57220
rect 165180 57210 165260 57220
rect 165360 57210 165440 57220
rect 165540 57210 165620 57220
rect 165720 57210 165800 57220
rect 165900 57210 165980 57220
rect 166080 57210 166160 57220
rect 166260 57210 166340 57220
rect 166440 57210 166520 57220
rect 166620 57210 166700 57220
rect 166800 57210 166880 57220
rect 166980 57210 167060 57220
rect 167160 57210 167240 57220
rect 167340 57210 167420 57220
rect 167520 57210 167600 57220
rect 167700 57210 167780 57220
rect 167880 57210 167960 57220
rect 168060 57210 168140 57220
rect 168240 57210 168320 57220
rect 168420 57210 168500 57220
rect 168600 57210 168680 57220
rect 168780 57210 168860 57220
rect 168960 57210 169040 57220
rect 169140 57210 169220 57220
rect 169320 57210 169400 57220
rect 169500 57210 169580 57220
rect 169680 57210 169760 57220
rect 169860 57210 169940 57220
rect 170040 57210 170120 57220
rect 152100 57100 152160 57130
rect 152220 57100 152280 57130
rect 152340 57100 152400 57130
rect 152900 57120 158990 57150
rect 159520 57130 159550 57160
rect 159640 57130 159670 57160
rect 163520 57130 163550 57160
rect 163640 57130 163670 57160
rect 164360 57130 164370 57210
rect 164540 57130 164550 57210
rect 164720 57130 164730 57210
rect 164900 57130 164910 57210
rect 165080 57130 165090 57210
rect 165260 57130 165270 57210
rect 165440 57130 165450 57210
rect 165620 57130 165630 57210
rect 165800 57130 165810 57210
rect 165980 57130 165990 57210
rect 166160 57130 166170 57210
rect 166340 57130 166350 57210
rect 166520 57130 166530 57210
rect 166700 57130 166710 57210
rect 166880 57130 166890 57210
rect 167060 57130 167070 57210
rect 167240 57130 167250 57210
rect 167420 57130 167430 57210
rect 167600 57130 167610 57210
rect 167780 57130 167790 57210
rect 167960 57130 167970 57210
rect 168140 57130 168150 57210
rect 168320 57130 168330 57210
rect 168500 57130 168510 57210
rect 168680 57130 168690 57210
rect 168860 57130 168870 57210
rect 169040 57130 169050 57210
rect 169220 57130 169230 57210
rect 169400 57130 169410 57210
rect 169580 57130 169590 57210
rect 169760 57130 169770 57210
rect 169940 57130 169950 57210
rect 170120 57130 170130 57210
rect 170810 57130 170840 57160
rect 170930 57130 170960 57160
rect 150605 57085 150685 57095
rect 150785 57085 150865 57095
rect 150965 57085 151045 57095
rect 151145 57085 151225 57095
rect 151325 57085 151405 57095
rect 146530 56950 147140 56960
rect 19010 56880 19070 56910
rect 19130 56880 19190 56910
rect 19250 56880 19310 56910
rect 19960 56830 19970 56910
rect 20140 56830 20150 56910
rect 20320 56830 20330 56910
rect 20500 56830 20510 56910
rect 20680 56830 20690 56910
rect 20860 56830 20870 56910
rect 21040 56830 21050 56910
rect 21220 56830 21230 56910
rect 21400 56830 21410 56910
rect 21580 56830 21590 56910
rect 21760 56830 21770 56910
rect 21940 56830 21950 56910
rect 22120 56830 22130 56910
rect 22300 56830 22310 56910
rect 22480 56830 22490 56910
rect 22660 56830 22670 56910
rect 22840 56830 22850 56910
rect 23020 56830 23030 56910
rect 23200 56830 23210 56910
rect 23380 56830 23390 56910
rect 23560 56830 23570 56910
rect 23740 56830 23750 56910
rect 23920 56830 23930 56910
rect 24100 56830 24110 56910
rect 24280 56830 24290 56910
rect 24460 56830 24470 56910
rect 24640 56830 24650 56910
rect 24820 56830 24830 56910
rect 25000 56830 25010 56910
rect 25180 56830 25190 56910
rect 25360 56830 25370 56910
rect 25540 56830 25550 56910
rect 25720 56830 25730 56910
rect 26300 56880 26360 56910
rect 26420 56880 26480 56910
rect 26540 56880 26600 56910
rect 30300 56880 30360 56910
rect 30420 56880 30480 56910
rect 30540 56880 30600 56910
rect 31100 56890 37190 56920
rect 37720 56910 37750 56940
rect 37840 56910 37870 56940
rect 146100 56910 146160 56940
rect 146420 56935 147090 56945
rect 147318 56940 147388 57080
rect 147580 57030 147640 57060
rect 148400 57030 148460 57060
rect 149880 57030 149940 57060
rect 150685 57005 150695 57085
rect 150865 57005 150875 57085
rect 151045 57005 151055 57085
rect 151225 57005 151235 57085
rect 151405 57005 151415 57085
rect 152980 57060 153060 57070
rect 153160 57060 153240 57070
rect 153340 57060 153420 57070
rect 153520 57060 153600 57070
rect 153700 57060 153780 57070
rect 153880 57060 153960 57070
rect 154060 57060 154140 57070
rect 154240 57060 154320 57070
rect 154420 57060 154500 57070
rect 154600 57060 154680 57070
rect 154780 57060 154860 57070
rect 154960 57060 155040 57070
rect 155140 57060 155220 57070
rect 155320 57060 155400 57070
rect 155500 57060 155580 57070
rect 155680 57060 155760 57070
rect 155860 57060 155940 57070
rect 156040 57060 156120 57070
rect 156220 57060 156300 57070
rect 156400 57060 156480 57070
rect 156580 57060 156660 57070
rect 156760 57060 156840 57070
rect 156940 57060 157020 57070
rect 157120 57060 157200 57070
rect 157300 57060 157380 57070
rect 157480 57060 157560 57070
rect 157660 57060 157740 57070
rect 157840 57060 157920 57070
rect 158020 57060 158100 57070
rect 158200 57060 158280 57070
rect 158380 57060 158460 57070
rect 158560 57060 158640 57070
rect 158740 57060 158820 57070
rect 152220 57010 152250 57040
rect 152340 57010 152370 57040
rect 152100 56980 152160 57010
rect 152220 56980 152280 57010
rect 152340 56980 152400 57010
rect 153060 56980 153070 57060
rect 153240 56980 153250 57060
rect 153420 56980 153430 57060
rect 153600 56980 153610 57060
rect 153780 56980 153790 57060
rect 153960 56980 153970 57060
rect 154140 56980 154150 57060
rect 154320 56980 154330 57060
rect 154500 56980 154510 57060
rect 154680 56980 154690 57060
rect 154860 56980 154870 57060
rect 155040 56980 155050 57060
rect 155220 56980 155230 57060
rect 155400 56980 155410 57060
rect 155580 56980 155590 57060
rect 155760 56980 155770 57060
rect 155940 56980 155950 57060
rect 156120 56980 156130 57060
rect 156300 56980 156310 57060
rect 156480 56980 156490 57060
rect 156660 56980 156670 57060
rect 156840 56980 156850 57060
rect 157020 56980 157030 57060
rect 157200 56980 157210 57060
rect 157380 56980 157390 57060
rect 157560 56980 157570 57060
rect 157740 56980 157750 57060
rect 157920 56980 157930 57060
rect 158100 56980 158110 57060
rect 158280 56980 158290 57060
rect 158460 56980 158470 57060
rect 158640 56980 158650 57060
rect 158820 56980 158830 57060
rect 149082 56951 149162 56961
rect 149242 56951 149322 56961
rect 31260 56830 31270 56890
rect 31440 56830 31450 56890
rect 31620 56830 31630 56890
rect 31800 56830 31810 56890
rect 31980 56830 31990 56890
rect 32160 56830 32170 56890
rect 32340 56830 32350 56890
rect 32520 56830 32530 56890
rect 32700 56830 32710 56890
rect 32880 56830 32890 56890
rect 33060 56830 33070 56890
rect 33240 56830 33250 56890
rect 33420 56830 33430 56890
rect 33600 56830 33610 56890
rect 33780 56830 33790 56890
rect 33960 56830 33970 56890
rect 34140 56830 34150 56890
rect 34320 56830 34330 56890
rect 34500 56830 34510 56890
rect 34680 56830 34690 56890
rect 34860 56830 34870 56890
rect 35040 56830 35050 56890
rect 35220 56830 35230 56890
rect 35400 56830 35410 56890
rect 35580 56830 35590 56890
rect 35760 56830 35770 56890
rect 35940 56830 35950 56890
rect 36120 56830 36130 56890
rect 36300 56830 36310 56890
rect 36480 56830 36490 56890
rect 36660 56830 36670 56890
rect 36840 56830 36850 56890
rect 37020 56830 37030 56890
rect 37100 56820 37190 56890
rect 37600 56880 37660 56910
rect 37720 56880 37780 56910
rect 37840 56880 37900 56910
rect 40060 56830 40120 56860
rect 41540 56830 41600 56860
rect 42360 56830 42420 56860
rect 43840 56830 43900 56860
rect 146420 56850 146480 56935
rect 146610 56840 146970 56900
rect 147090 56885 147100 56935
rect 147178 56880 147318 56940
rect 147580 56910 147640 56940
rect 148400 56910 148460 56940
rect 19130 56790 19160 56820
rect 19250 56790 19280 56820
rect 26420 56790 26450 56820
rect 26540 56790 26570 56820
rect 30420 56790 30450 56820
rect 30540 56790 30570 56820
rect 31100 56790 37190 56820
rect 37720 56790 37750 56820
rect 37840 56790 37870 56820
rect 146100 56790 146160 56820
rect 19010 56760 19070 56790
rect 19130 56760 19190 56790
rect 19250 56760 19310 56790
rect 19800 56770 25800 56780
rect 26300 56760 26360 56790
rect 26420 56760 26480 56790
rect 26540 56760 26600 56790
rect 30300 56760 30360 56790
rect 30420 56760 30480 56790
rect 30540 56760 30600 56790
rect 37100 56780 37190 56790
rect 31100 56770 37190 56780
rect 19130 56670 19160 56700
rect 19250 56670 19280 56700
rect 26420 56670 26450 56700
rect 26540 56670 26570 56700
rect 30420 56670 30450 56700
rect 30540 56670 30570 56700
rect 19010 56640 19070 56670
rect 19130 56640 19190 56670
rect 19250 56640 19310 56670
rect 26300 56640 26360 56670
rect 26420 56640 26480 56670
rect 26540 56640 26600 56670
rect 30300 56640 30360 56670
rect 30420 56640 30480 56670
rect 30540 56640 30600 56670
rect 31180 56590 31260 56600
rect 31360 56590 31440 56600
rect 31540 56590 31620 56600
rect 31720 56590 31800 56600
rect 31900 56590 31980 56600
rect 32080 56590 32160 56600
rect 32260 56590 32340 56600
rect 32440 56590 32520 56600
rect 32620 56590 32700 56600
rect 32800 56590 32880 56600
rect 32980 56590 33060 56600
rect 33160 56590 33240 56600
rect 33340 56590 33420 56600
rect 33520 56590 33600 56600
rect 33700 56590 33780 56600
rect 33880 56590 33960 56600
rect 34060 56590 34140 56600
rect 34240 56590 34320 56600
rect 34420 56590 34500 56600
rect 34600 56590 34680 56600
rect 34780 56590 34860 56600
rect 34960 56590 35040 56600
rect 35140 56590 35220 56600
rect 35320 56590 35400 56600
rect 35500 56590 35580 56600
rect 35680 56590 35760 56600
rect 35860 56590 35940 56600
rect 36040 56590 36120 56600
rect 36220 56590 36300 56600
rect 36400 56590 36480 56600
rect 36580 56590 36660 56600
rect 36760 56590 36840 56600
rect 36940 56590 37020 56600
rect 19130 56550 19160 56580
rect 19250 56550 19280 56580
rect 19880 56570 19960 56580
rect 20060 56570 20140 56580
rect 20240 56570 20320 56580
rect 20420 56570 20500 56580
rect 20600 56570 20680 56580
rect 20780 56570 20860 56580
rect 20960 56570 21040 56580
rect 21140 56570 21220 56580
rect 21320 56570 21400 56580
rect 21500 56570 21580 56580
rect 21680 56570 21760 56580
rect 21860 56570 21940 56580
rect 22040 56570 22120 56580
rect 22220 56570 22300 56580
rect 22400 56570 22480 56580
rect 22580 56570 22660 56580
rect 22760 56570 22840 56580
rect 22940 56570 23020 56580
rect 23120 56570 23200 56580
rect 23300 56570 23380 56580
rect 23480 56570 23560 56580
rect 23660 56570 23740 56580
rect 23840 56570 23920 56580
rect 24020 56570 24100 56580
rect 24200 56570 24280 56580
rect 24380 56570 24460 56580
rect 24560 56570 24640 56580
rect 24740 56570 24820 56580
rect 24920 56570 25000 56580
rect 25100 56570 25180 56580
rect 25280 56570 25360 56580
rect 25460 56570 25540 56580
rect 25640 56570 25720 56580
rect 19010 56520 19070 56550
rect 19130 56520 19190 56550
rect 19250 56520 19310 56550
rect 19960 56490 19970 56570
rect 20140 56490 20150 56570
rect 20320 56490 20330 56570
rect 20500 56490 20510 56570
rect 20680 56490 20690 56570
rect 20860 56490 20870 56570
rect 21040 56490 21050 56570
rect 21220 56490 21230 56570
rect 21400 56490 21410 56570
rect 21580 56490 21590 56570
rect 21760 56490 21770 56570
rect 21940 56490 21950 56570
rect 22120 56490 22130 56570
rect 22300 56490 22310 56570
rect 22480 56490 22490 56570
rect 22660 56490 22670 56570
rect 22840 56490 22850 56570
rect 23020 56490 23030 56570
rect 23200 56490 23210 56570
rect 23380 56490 23390 56570
rect 23560 56490 23570 56570
rect 23740 56490 23750 56570
rect 23920 56490 23930 56570
rect 24100 56490 24110 56570
rect 24280 56490 24290 56570
rect 24460 56490 24470 56570
rect 24640 56490 24650 56570
rect 24820 56490 24830 56570
rect 25000 56490 25010 56570
rect 25180 56490 25190 56570
rect 25360 56490 25370 56570
rect 25540 56490 25550 56570
rect 25720 56490 25730 56570
rect 26420 56550 26450 56580
rect 26540 56550 26570 56580
rect 30420 56550 30450 56580
rect 30540 56550 30570 56580
rect 26300 56520 26360 56550
rect 26420 56520 26480 56550
rect 26540 56520 26600 56550
rect 30300 56520 30360 56550
rect 30420 56520 30480 56550
rect 30540 56520 30600 56550
rect 31260 56510 31270 56590
rect 31440 56510 31450 56590
rect 31620 56510 31630 56590
rect 31800 56510 31810 56590
rect 31980 56510 31990 56590
rect 32160 56510 32170 56590
rect 32340 56510 32350 56590
rect 32520 56510 32530 56590
rect 32700 56510 32710 56590
rect 32880 56510 32890 56590
rect 33060 56510 33070 56590
rect 33240 56510 33250 56590
rect 33420 56510 33430 56590
rect 33600 56510 33610 56590
rect 33780 56510 33790 56590
rect 33960 56510 33970 56590
rect 34140 56510 34150 56590
rect 34320 56510 34330 56590
rect 34500 56510 34510 56590
rect 34680 56510 34690 56590
rect 34860 56510 34870 56590
rect 35040 56510 35050 56590
rect 35220 56510 35230 56590
rect 35400 56510 35410 56590
rect 35580 56510 35590 56590
rect 35760 56510 35770 56590
rect 35940 56510 35950 56590
rect 36120 56510 36130 56590
rect 36300 56510 36310 56590
rect 36480 56510 36490 56590
rect 36660 56510 36670 56590
rect 36840 56510 36850 56590
rect 37020 56510 37030 56590
rect 19130 56430 19160 56460
rect 19250 56430 19280 56460
rect 26420 56430 26450 56460
rect 26540 56430 26570 56460
rect 30420 56430 30450 56460
rect 30540 56430 30570 56460
rect 19010 56400 19070 56430
rect 19130 56400 19190 56430
rect 19250 56400 19310 56430
rect 26300 56400 26360 56430
rect 26420 56400 26480 56430
rect 26540 56400 26600 56430
rect 30300 56400 30360 56430
rect 30420 56400 30480 56430
rect 30540 56400 30600 56430
rect 19130 56310 19160 56340
rect 19250 56310 19280 56340
rect 26420 56310 26450 56340
rect 26540 56310 26570 56340
rect 30420 56310 30450 56340
rect 30540 56310 30570 56340
rect 19010 56280 19070 56310
rect 19130 56280 19190 56310
rect 19250 56280 19310 56310
rect 26300 56280 26360 56310
rect 26420 56280 26480 56310
rect 26540 56280 26600 56310
rect 30300 56280 30360 56310
rect 30420 56280 30480 56310
rect 30540 56280 30600 56310
rect 19880 56270 19960 56280
rect 20060 56270 20140 56280
rect 20240 56270 20320 56280
rect 20420 56270 20500 56280
rect 20600 56270 20680 56280
rect 20780 56270 20860 56280
rect 20960 56270 21040 56280
rect 21140 56270 21220 56280
rect 21320 56270 21400 56280
rect 21500 56270 21580 56280
rect 21680 56270 21760 56280
rect 21860 56270 21940 56280
rect 22040 56270 22120 56280
rect 22220 56270 22300 56280
rect 22400 56270 22480 56280
rect 22580 56270 22660 56280
rect 22760 56270 22840 56280
rect 22940 56270 23020 56280
rect 23120 56270 23200 56280
rect 23300 56270 23380 56280
rect 23480 56270 23560 56280
rect 23660 56270 23740 56280
rect 23840 56270 23920 56280
rect 24020 56270 24100 56280
rect 24200 56270 24280 56280
rect 24380 56270 24460 56280
rect 24560 56270 24640 56280
rect 24740 56270 24820 56280
rect 24920 56270 25000 56280
rect 25100 56270 25180 56280
rect 25280 56270 25360 56280
rect 25460 56270 25540 56280
rect 25640 56270 25720 56280
rect 31180 56270 31260 56280
rect 31360 56270 31440 56280
rect 31540 56270 31620 56280
rect 31720 56270 31800 56280
rect 31900 56270 31980 56280
rect 32080 56270 32160 56280
rect 32260 56270 32340 56280
rect 32440 56270 32520 56280
rect 32620 56270 32700 56280
rect 32800 56270 32880 56280
rect 32980 56270 33060 56280
rect 33160 56270 33240 56280
rect 33340 56270 33420 56280
rect 33520 56270 33600 56280
rect 33700 56270 33780 56280
rect 33880 56270 33960 56280
rect 34060 56270 34140 56280
rect 34240 56270 34320 56280
rect 34420 56270 34500 56280
rect 34600 56270 34680 56280
rect 34780 56270 34860 56280
rect 34960 56270 35040 56280
rect 35140 56270 35220 56280
rect 35320 56270 35400 56280
rect 35500 56270 35580 56280
rect 35680 56270 35760 56280
rect 35860 56270 35940 56280
rect 36040 56270 36120 56280
rect 36220 56270 36300 56280
rect 36400 56270 36480 56280
rect 36580 56270 36660 56280
rect 36760 56270 36840 56280
rect 36940 56270 37020 56280
rect 19130 56190 19160 56220
rect 19250 56190 19280 56220
rect 19960 56190 19970 56270
rect 20140 56190 20150 56270
rect 20320 56190 20330 56270
rect 20500 56190 20510 56270
rect 20680 56190 20690 56270
rect 20860 56190 20870 56270
rect 21040 56190 21050 56270
rect 21220 56190 21230 56270
rect 21400 56190 21410 56270
rect 21580 56190 21590 56270
rect 21760 56190 21770 56270
rect 21940 56190 21950 56270
rect 22120 56190 22130 56270
rect 22300 56190 22310 56270
rect 22480 56190 22490 56270
rect 22660 56190 22670 56270
rect 22840 56190 22850 56270
rect 23020 56190 23030 56270
rect 23200 56190 23210 56270
rect 23380 56190 23390 56270
rect 23560 56190 23570 56270
rect 23740 56190 23750 56270
rect 23920 56190 23930 56270
rect 24100 56190 24110 56270
rect 24280 56190 24290 56270
rect 24460 56190 24470 56270
rect 24640 56190 24650 56270
rect 24820 56190 24830 56270
rect 25000 56190 25010 56270
rect 25180 56190 25190 56270
rect 25360 56190 25370 56270
rect 25540 56190 25550 56270
rect 25720 56190 25730 56270
rect 26420 56190 26450 56220
rect 26540 56190 26570 56220
rect 30420 56190 30450 56220
rect 30540 56190 30570 56220
rect 31260 56190 31270 56270
rect 31440 56190 31450 56270
rect 31620 56190 31630 56270
rect 31800 56190 31810 56270
rect 31980 56190 31990 56270
rect 32160 56190 32170 56270
rect 32340 56190 32350 56270
rect 32520 56190 32530 56270
rect 32700 56190 32710 56270
rect 32880 56190 32890 56270
rect 33060 56190 33070 56270
rect 33240 56190 33250 56270
rect 33420 56190 33430 56270
rect 33600 56190 33610 56270
rect 33780 56190 33790 56270
rect 33960 56190 33970 56270
rect 34140 56190 34150 56270
rect 34320 56190 34330 56270
rect 34500 56190 34510 56270
rect 34680 56190 34690 56270
rect 34860 56190 34870 56270
rect 35040 56190 35050 56270
rect 35220 56190 35230 56270
rect 35400 56190 35410 56270
rect 35580 56190 35590 56270
rect 35760 56190 35770 56270
rect 35940 56190 35950 56270
rect 36120 56190 36130 56270
rect 36300 56190 36310 56270
rect 36480 56190 36490 56270
rect 36660 56190 36670 56270
rect 36840 56190 36850 56270
rect 37020 56190 37030 56270
rect 19010 56160 19070 56190
rect 19130 56160 19190 56190
rect 19250 56160 19310 56190
rect 26300 56160 26360 56190
rect 26420 56160 26480 56190
rect 26540 56160 26600 56190
rect 30300 56160 30360 56190
rect 30420 56160 30480 56190
rect 30540 56160 30600 56190
rect 37100 56100 37190 56770
rect 37600 56760 37660 56790
rect 37720 56760 37780 56790
rect 37840 56760 37900 56790
rect 40060 56710 40120 56740
rect 41540 56710 41600 56740
rect 42360 56710 42420 56740
rect 43840 56710 43900 56740
rect 146300 56710 146420 56770
rect 147318 56740 147388 56880
rect 149162 56871 149172 56951
rect 149242 56871 149252 56951
rect 149322 56871 149332 56951
rect 149880 56910 149940 56940
rect 158900 56920 158990 57120
rect 159400 57100 159460 57130
rect 159520 57100 159580 57130
rect 159640 57100 159700 57130
rect 163400 57100 163460 57130
rect 163520 57100 163580 57130
rect 163640 57100 163700 57130
rect 170690 57100 170750 57130
rect 170810 57100 170870 57130
rect 170930 57100 170990 57130
rect 164280 57060 164360 57070
rect 164460 57060 164540 57070
rect 164640 57060 164720 57070
rect 164820 57060 164900 57070
rect 165000 57060 165080 57070
rect 165180 57060 165260 57070
rect 165360 57060 165440 57070
rect 165540 57060 165620 57070
rect 165720 57060 165800 57070
rect 165900 57060 165980 57070
rect 166080 57060 166160 57070
rect 166260 57060 166340 57070
rect 166440 57060 166520 57070
rect 166620 57060 166700 57070
rect 166800 57060 166880 57070
rect 166980 57060 167060 57070
rect 167160 57060 167240 57070
rect 167340 57060 167420 57070
rect 167520 57060 167600 57070
rect 167700 57060 167780 57070
rect 167880 57060 167960 57070
rect 168060 57060 168140 57070
rect 168240 57060 168320 57070
rect 168420 57060 168500 57070
rect 168600 57060 168680 57070
rect 168780 57060 168860 57070
rect 168960 57060 169040 57070
rect 169140 57060 169220 57070
rect 169320 57060 169400 57070
rect 169500 57060 169580 57070
rect 169680 57060 169760 57070
rect 169860 57060 169940 57070
rect 170040 57060 170120 57070
rect 159520 57010 159550 57040
rect 159640 57010 159670 57040
rect 163520 57010 163550 57040
rect 163640 57010 163670 57040
rect 159400 56980 159460 57010
rect 159520 56980 159580 57010
rect 159640 56980 159700 57010
rect 163400 56980 163460 57010
rect 163520 56980 163580 57010
rect 163640 56980 163700 57010
rect 164360 56980 164370 57060
rect 164540 56980 164550 57060
rect 164720 56980 164730 57060
rect 164900 56980 164910 57060
rect 165080 56980 165090 57060
rect 165260 56980 165270 57060
rect 165440 56980 165450 57060
rect 165620 56980 165630 57060
rect 165800 56980 165810 57060
rect 165980 56980 165990 57060
rect 166160 56980 166170 57060
rect 166340 56980 166350 57060
rect 166520 56980 166530 57060
rect 166700 56980 166710 57060
rect 166880 56980 166890 57060
rect 167060 56980 167070 57060
rect 167240 56980 167250 57060
rect 167420 56980 167430 57060
rect 167600 56980 167610 57060
rect 167780 56980 167790 57060
rect 167960 56980 167970 57060
rect 168140 56980 168150 57060
rect 168320 56980 168330 57060
rect 168500 56980 168510 57060
rect 168680 56980 168690 57060
rect 168860 56980 168870 57060
rect 169040 56980 169050 57060
rect 169220 56980 169230 57060
rect 169400 56980 169410 57060
rect 169580 56980 169590 57060
rect 169760 56980 169770 57060
rect 169940 56980 169950 57060
rect 170120 56980 170130 57060
rect 170810 57010 170840 57040
rect 170930 57010 170960 57040
rect 170690 56980 170750 57010
rect 170810 56980 170870 57010
rect 170930 56980 170990 57010
rect 150605 56905 150685 56915
rect 150785 56905 150865 56915
rect 150965 56905 151045 56915
rect 151145 56905 151225 56915
rect 151325 56905 151405 56915
rect 147580 56790 147640 56820
rect 148400 56790 148460 56820
rect 149075 56810 149315 56840
rect 150685 56825 150695 56905
rect 150865 56825 150875 56905
rect 151045 56825 151055 56905
rect 151225 56825 151235 56905
rect 151405 56825 151415 56905
rect 152220 56890 152250 56920
rect 152340 56890 152370 56920
rect 152900 56890 158990 56920
rect 159520 56890 159550 56920
rect 159640 56890 159670 56920
rect 163520 56890 163550 56920
rect 163640 56890 163670 56920
rect 164280 56910 164360 56920
rect 164460 56910 164540 56920
rect 164640 56910 164720 56920
rect 164820 56910 164900 56920
rect 165000 56910 165080 56920
rect 165180 56910 165260 56920
rect 165360 56910 165440 56920
rect 165540 56910 165620 56920
rect 165720 56910 165800 56920
rect 165900 56910 165980 56920
rect 166080 56910 166160 56920
rect 166260 56910 166340 56920
rect 166440 56910 166520 56920
rect 166620 56910 166700 56920
rect 166800 56910 166880 56920
rect 166980 56910 167060 56920
rect 167160 56910 167240 56920
rect 167340 56910 167420 56920
rect 167520 56910 167600 56920
rect 167700 56910 167780 56920
rect 167880 56910 167960 56920
rect 168060 56910 168140 56920
rect 168240 56910 168320 56920
rect 168420 56910 168500 56920
rect 168600 56910 168680 56920
rect 168780 56910 168860 56920
rect 168960 56910 169040 56920
rect 169140 56910 169220 56920
rect 169320 56910 169400 56920
rect 169500 56910 169580 56920
rect 169680 56910 169760 56920
rect 169860 56910 169940 56920
rect 170040 56910 170120 56920
rect 152100 56860 152160 56890
rect 152220 56860 152280 56890
rect 152340 56860 152400 56890
rect 153060 56830 153070 56890
rect 153240 56830 153250 56890
rect 153420 56830 153430 56890
rect 153600 56830 153610 56890
rect 153780 56830 153790 56890
rect 153960 56830 153970 56890
rect 154140 56830 154150 56890
rect 154320 56830 154330 56890
rect 154500 56830 154510 56890
rect 154680 56830 154690 56890
rect 154860 56830 154870 56890
rect 155040 56830 155050 56890
rect 155220 56830 155230 56890
rect 155400 56830 155410 56890
rect 155580 56830 155590 56890
rect 155760 56830 155770 56890
rect 155940 56830 155950 56890
rect 156120 56830 156130 56890
rect 156300 56830 156310 56890
rect 156480 56830 156490 56890
rect 156660 56830 156670 56890
rect 156840 56830 156850 56890
rect 157020 56830 157030 56890
rect 157200 56830 157210 56890
rect 157380 56830 157390 56890
rect 157560 56830 157570 56890
rect 157740 56830 157750 56890
rect 157920 56830 157930 56890
rect 158100 56830 158110 56890
rect 158280 56830 158290 56890
rect 158460 56830 158470 56890
rect 158640 56830 158650 56890
rect 158820 56830 158830 56890
rect 158900 56820 158990 56890
rect 159400 56860 159460 56890
rect 159520 56860 159580 56890
rect 159640 56860 159700 56890
rect 163400 56860 163460 56890
rect 163520 56860 163580 56890
rect 163640 56860 163700 56890
rect 164360 56830 164370 56910
rect 164540 56830 164550 56910
rect 164720 56830 164730 56910
rect 164900 56830 164910 56910
rect 165080 56830 165090 56910
rect 165260 56830 165270 56910
rect 165440 56830 165450 56910
rect 165620 56830 165630 56910
rect 165800 56830 165810 56910
rect 165980 56830 165990 56910
rect 166160 56830 166170 56910
rect 166340 56830 166350 56910
rect 166520 56830 166530 56910
rect 166700 56830 166710 56910
rect 166880 56830 166890 56910
rect 167060 56830 167070 56910
rect 167240 56830 167250 56910
rect 167420 56830 167430 56910
rect 167600 56830 167610 56910
rect 167780 56830 167790 56910
rect 167960 56830 167970 56910
rect 168140 56830 168150 56910
rect 168320 56830 168330 56910
rect 168500 56830 168510 56910
rect 168680 56830 168690 56910
rect 168860 56830 168870 56910
rect 169040 56830 169050 56910
rect 169220 56830 169230 56910
rect 169400 56830 169410 56910
rect 169580 56830 169590 56910
rect 169760 56830 169770 56910
rect 169940 56830 169950 56910
rect 170120 56830 170130 56910
rect 170810 56890 170840 56920
rect 170930 56890 170960 56920
rect 170690 56860 170750 56890
rect 170810 56860 170870 56890
rect 170930 56860 170990 56890
rect 149075 56750 149105 56810
rect 149165 56750 149255 56810
rect 149285 56750 149315 56810
rect 149880 56790 149940 56820
rect 152220 56770 152250 56800
rect 152340 56770 152370 56800
rect 152900 56790 158990 56820
rect 158900 56780 158990 56790
rect 152900 56770 158990 56780
rect 159520 56770 159550 56800
rect 159640 56770 159670 56800
rect 163520 56770 163550 56800
rect 163640 56770 163670 56800
rect 164200 56770 170200 56780
rect 170810 56770 170840 56800
rect 170930 56770 170960 56800
rect 146420 56700 146480 56710
rect 37720 56670 37750 56700
rect 37840 56670 37870 56700
rect 146100 56670 146160 56700
rect 146420 56690 147050 56700
rect 146420 56685 146480 56690
rect 146420 56675 147090 56685
rect 147178 56680 147318 56740
rect 149075 56720 149315 56750
rect 152100 56740 152160 56770
rect 152220 56740 152280 56770
rect 152340 56740 152400 56770
rect 150605 56725 150685 56735
rect 150785 56725 150865 56735
rect 150965 56725 151045 56735
rect 151145 56725 151225 56735
rect 151325 56725 151405 56735
rect 37600 56640 37660 56670
rect 37720 56640 37780 56670
rect 37840 56640 37900 56670
rect 40060 56590 40120 56620
rect 41540 56590 41600 56620
rect 42360 56590 42420 56620
rect 43840 56590 43900 56620
rect 146420 56590 146480 56675
rect 37720 56550 37750 56580
rect 37840 56550 37870 56580
rect 146100 56550 146160 56580
rect 37600 56520 37660 56550
rect 37720 56520 37780 56550
rect 37840 56520 37900 56550
rect 40060 56470 40120 56500
rect 41540 56470 41600 56500
rect 42360 56470 42420 56500
rect 43840 56470 43900 56500
rect 37720 56430 37750 56460
rect 37840 56430 37870 56460
rect 146100 56430 146160 56460
rect 146300 56450 146420 56510
rect 37600 56400 37660 56430
rect 37720 56400 37780 56430
rect 37840 56400 37900 56430
rect 146420 56425 146480 56450
rect 146530 56440 146540 56610
rect 146610 56580 146970 56640
rect 147090 56625 147100 56675
rect 147318 56540 147388 56680
rect 147580 56670 147640 56700
rect 148400 56670 148460 56700
rect 149082 56681 149162 56691
rect 149242 56681 149322 56691
rect 149162 56601 149172 56681
rect 149242 56601 149252 56681
rect 149322 56601 149332 56681
rect 149880 56670 149940 56700
rect 150685 56645 150695 56725
rect 150865 56645 150875 56725
rect 151045 56645 151055 56725
rect 151225 56645 151235 56725
rect 151405 56645 151415 56725
rect 152220 56650 152250 56680
rect 152340 56650 152370 56680
rect 152100 56620 152160 56650
rect 152220 56620 152280 56650
rect 152340 56620 152400 56650
rect 152980 56590 153060 56600
rect 153160 56590 153240 56600
rect 153340 56590 153420 56600
rect 153520 56590 153600 56600
rect 153700 56590 153780 56600
rect 153880 56590 153960 56600
rect 154060 56590 154140 56600
rect 154240 56590 154320 56600
rect 154420 56590 154500 56600
rect 154600 56590 154680 56600
rect 154780 56590 154860 56600
rect 154960 56590 155040 56600
rect 155140 56590 155220 56600
rect 155320 56590 155400 56600
rect 155500 56590 155580 56600
rect 155680 56590 155760 56600
rect 155860 56590 155940 56600
rect 156040 56590 156120 56600
rect 156220 56590 156300 56600
rect 156400 56590 156480 56600
rect 156580 56590 156660 56600
rect 156760 56590 156840 56600
rect 156940 56590 157020 56600
rect 157120 56590 157200 56600
rect 157300 56590 157380 56600
rect 157480 56590 157560 56600
rect 157660 56590 157740 56600
rect 157840 56590 157920 56600
rect 158020 56590 158100 56600
rect 158200 56590 158280 56600
rect 158380 56590 158460 56600
rect 158560 56590 158640 56600
rect 158740 56590 158820 56600
rect 147580 56550 147640 56580
rect 148400 56550 148460 56580
rect 149880 56550 149940 56580
rect 150605 56545 150685 56555
rect 150785 56545 150865 56555
rect 150965 56545 151045 56555
rect 151145 56545 151225 56555
rect 151325 56545 151405 56555
rect 150685 56465 150695 56545
rect 150865 56465 150875 56545
rect 151045 56465 151055 56545
rect 151225 56465 151235 56545
rect 151405 56465 151415 56545
rect 152220 56530 152250 56560
rect 152340 56530 152370 56560
rect 152100 56500 152160 56530
rect 152220 56500 152280 56530
rect 152340 56500 152400 56530
rect 153060 56510 153070 56590
rect 153240 56510 153250 56590
rect 153420 56510 153430 56590
rect 153600 56510 153610 56590
rect 153780 56510 153790 56590
rect 153960 56510 153970 56590
rect 154140 56510 154150 56590
rect 154320 56510 154330 56590
rect 154500 56510 154510 56590
rect 154680 56510 154690 56590
rect 154860 56510 154870 56590
rect 155040 56510 155050 56590
rect 155220 56510 155230 56590
rect 155400 56510 155410 56590
rect 155580 56510 155590 56590
rect 155760 56510 155770 56590
rect 155940 56510 155950 56590
rect 156120 56510 156130 56590
rect 156300 56510 156310 56590
rect 156480 56510 156490 56590
rect 156660 56510 156670 56590
rect 156840 56510 156850 56590
rect 157020 56510 157030 56590
rect 157200 56510 157210 56590
rect 157380 56510 157390 56590
rect 157560 56510 157570 56590
rect 157740 56510 157750 56590
rect 157920 56510 157930 56590
rect 158100 56510 158110 56590
rect 158280 56510 158290 56590
rect 158460 56510 158470 56590
rect 158640 56510 158650 56590
rect 158820 56510 158830 56590
rect 146530 56430 147140 56440
rect 147580 56430 147640 56460
rect 148400 56430 148460 56460
rect 149880 56430 149940 56460
rect 146420 56415 147090 56425
rect 40060 56350 40120 56380
rect 41540 56350 41600 56380
rect 42360 56350 42420 56380
rect 43840 56350 43900 56380
rect 37720 56310 37750 56340
rect 37840 56310 37870 56340
rect 146100 56310 146160 56340
rect 146420 56330 146480 56415
rect 146610 56320 146970 56380
rect 147090 56365 147100 56415
rect 152220 56410 152250 56440
rect 152340 56410 152370 56440
rect 152100 56380 152160 56410
rect 152220 56380 152280 56410
rect 152340 56380 152400 56410
rect 150605 56365 150685 56375
rect 150785 56365 150865 56375
rect 150965 56365 151045 56375
rect 151145 56365 151225 56375
rect 151325 56365 151405 56375
rect 147580 56310 147640 56340
rect 148400 56310 148460 56340
rect 149880 56310 149940 56340
rect 37600 56280 37660 56310
rect 37720 56280 37780 56310
rect 37840 56280 37900 56310
rect 150685 56285 150695 56365
rect 150865 56285 150875 56365
rect 151045 56285 151055 56365
rect 151225 56285 151235 56365
rect 151405 56285 151415 56365
rect 152220 56290 152250 56320
rect 152340 56290 152370 56320
rect 147325 56265 147405 56275
rect 40060 56230 40120 56260
rect 41540 56230 41600 56260
rect 42360 56230 42420 56260
rect 43840 56230 43900 56260
rect 37720 56190 37750 56220
rect 37840 56190 37870 56220
rect 146100 56190 146160 56220
rect 147405 56195 147415 56265
rect 152100 56260 152160 56290
rect 152220 56260 152280 56290
rect 152340 56260 152400 56290
rect 152980 56270 153060 56280
rect 153160 56270 153240 56280
rect 153340 56270 153420 56280
rect 153520 56270 153600 56280
rect 153700 56270 153780 56280
rect 153880 56270 153960 56280
rect 154060 56270 154140 56280
rect 154240 56270 154320 56280
rect 154420 56270 154500 56280
rect 154600 56270 154680 56280
rect 154780 56270 154860 56280
rect 154960 56270 155040 56280
rect 155140 56270 155220 56280
rect 155320 56270 155400 56280
rect 155500 56270 155580 56280
rect 155680 56270 155760 56280
rect 155860 56270 155940 56280
rect 156040 56270 156120 56280
rect 156220 56270 156300 56280
rect 156400 56270 156480 56280
rect 156580 56270 156660 56280
rect 156760 56270 156840 56280
rect 156940 56270 157020 56280
rect 157120 56270 157200 56280
rect 157300 56270 157380 56280
rect 157480 56270 157560 56280
rect 157660 56270 157740 56280
rect 157840 56270 157920 56280
rect 158020 56270 158100 56280
rect 158200 56270 158280 56280
rect 158380 56270 158460 56280
rect 158560 56270 158640 56280
rect 158740 56270 158820 56280
rect 37600 56160 37660 56190
rect 37720 56160 37780 56190
rect 37840 56160 37900 56190
rect 147325 56185 147415 56195
rect 147580 56190 147640 56220
rect 148400 56190 148460 56220
rect 149880 56190 149940 56220
rect 152220 56170 152250 56200
rect 152340 56170 152370 56200
rect 153060 56190 153070 56270
rect 153240 56190 153250 56270
rect 153420 56190 153430 56270
rect 153600 56190 153610 56270
rect 153780 56190 153790 56270
rect 153960 56190 153970 56270
rect 154140 56190 154150 56270
rect 154320 56190 154330 56270
rect 154500 56190 154510 56270
rect 154680 56190 154690 56270
rect 154860 56190 154870 56270
rect 155040 56190 155050 56270
rect 155220 56190 155230 56270
rect 155400 56190 155410 56270
rect 155580 56190 155590 56270
rect 155760 56190 155770 56270
rect 155940 56190 155950 56270
rect 156120 56190 156130 56270
rect 156300 56190 156310 56270
rect 156480 56190 156490 56270
rect 156660 56190 156670 56270
rect 156840 56190 156850 56270
rect 157020 56190 157030 56270
rect 157200 56190 157210 56270
rect 157380 56190 157390 56270
rect 157560 56190 157570 56270
rect 157740 56190 157750 56270
rect 157920 56190 157930 56270
rect 158100 56190 158110 56270
rect 158280 56190 158290 56270
rect 158460 56190 158470 56270
rect 158640 56190 158650 56270
rect 158820 56190 158830 56270
rect 152100 56140 152160 56170
rect 152220 56140 152280 56170
rect 152340 56140 152400 56170
rect 40060 56110 40120 56140
rect 41540 56110 41600 56140
rect 42360 56110 42420 56140
rect 43840 56110 43900 56140
rect 147325 56105 147405 56115
rect 19130 56070 19160 56100
rect 19250 56070 19280 56100
rect 19800 56090 25800 56100
rect 26420 56070 26450 56100
rect 26540 56070 26570 56100
rect 30420 56070 30450 56100
rect 30540 56070 30570 56100
rect 31100 56090 37190 56100
rect 19010 56040 19070 56070
rect 19130 56040 19190 56070
rect 19250 56040 19310 56070
rect 26300 56040 26360 56070
rect 26420 56040 26480 56070
rect 26540 56040 26600 56070
rect 30300 56040 30360 56070
rect 30420 56040 30480 56070
rect 30540 56040 30600 56070
rect 37100 55990 37190 56090
rect 37720 56070 37750 56100
rect 37840 56070 37870 56100
rect 146100 56070 146160 56100
rect 37600 56040 37660 56070
rect 37720 56040 37780 56070
rect 37840 56040 37900 56070
rect 147405 56025 147415 56105
rect 158900 56100 158990 56770
rect 159400 56740 159460 56770
rect 159520 56740 159580 56770
rect 159640 56740 159700 56770
rect 163400 56740 163460 56770
rect 163520 56740 163580 56770
rect 163640 56740 163700 56770
rect 170690 56740 170750 56770
rect 170810 56740 170870 56770
rect 170930 56740 170990 56770
rect 159520 56650 159550 56680
rect 159640 56650 159670 56680
rect 163520 56650 163550 56680
rect 163640 56650 163670 56680
rect 170810 56650 170840 56680
rect 170930 56650 170960 56680
rect 159400 56620 159460 56650
rect 159520 56620 159580 56650
rect 159640 56620 159700 56650
rect 163400 56620 163460 56650
rect 163520 56620 163580 56650
rect 163640 56620 163700 56650
rect 170690 56620 170750 56650
rect 170810 56620 170870 56650
rect 170930 56620 170990 56650
rect 164280 56590 164360 56600
rect 164460 56590 164540 56600
rect 164640 56590 164720 56600
rect 164820 56590 164900 56600
rect 165000 56590 165080 56600
rect 165180 56590 165260 56600
rect 165360 56590 165440 56600
rect 165540 56590 165620 56600
rect 165720 56590 165800 56600
rect 165900 56590 165980 56600
rect 166080 56590 166160 56600
rect 166260 56590 166340 56600
rect 166440 56590 166520 56600
rect 166620 56590 166700 56600
rect 166800 56590 166880 56600
rect 166980 56590 167060 56600
rect 167160 56590 167240 56600
rect 167340 56590 167420 56600
rect 167520 56590 167600 56600
rect 167700 56590 167780 56600
rect 167880 56590 167960 56600
rect 168060 56590 168140 56600
rect 168240 56590 168320 56600
rect 168420 56590 168500 56600
rect 168600 56590 168680 56600
rect 168780 56590 168860 56600
rect 168960 56590 169040 56600
rect 169140 56590 169220 56600
rect 169320 56590 169400 56600
rect 169500 56590 169580 56600
rect 169680 56590 169760 56600
rect 169860 56590 169940 56600
rect 170040 56590 170120 56600
rect 159520 56530 159550 56560
rect 159640 56530 159670 56560
rect 163520 56530 163550 56560
rect 163640 56530 163670 56560
rect 159400 56500 159460 56530
rect 159520 56500 159580 56530
rect 159640 56500 159700 56530
rect 163400 56500 163460 56530
rect 163520 56500 163580 56530
rect 163640 56500 163700 56530
rect 164360 56510 164370 56590
rect 164540 56510 164550 56590
rect 164720 56510 164730 56590
rect 164900 56510 164910 56590
rect 165080 56510 165090 56590
rect 165260 56510 165270 56590
rect 165440 56510 165450 56590
rect 165620 56510 165630 56590
rect 165800 56510 165810 56590
rect 165980 56510 165990 56590
rect 166160 56510 166170 56590
rect 166340 56510 166350 56590
rect 166520 56510 166530 56590
rect 166700 56510 166710 56590
rect 166880 56510 166890 56590
rect 167060 56510 167070 56590
rect 167240 56510 167250 56590
rect 167420 56510 167430 56590
rect 167600 56510 167610 56590
rect 167780 56510 167790 56590
rect 167960 56510 167970 56590
rect 168140 56510 168150 56590
rect 168320 56510 168330 56590
rect 168500 56510 168510 56590
rect 168680 56510 168690 56590
rect 168860 56510 168870 56590
rect 169040 56510 169050 56590
rect 169220 56510 169230 56590
rect 169400 56510 169410 56590
rect 169580 56510 169590 56590
rect 169760 56510 169770 56590
rect 169940 56510 169950 56590
rect 170120 56510 170130 56590
rect 170810 56530 170840 56560
rect 170930 56530 170960 56560
rect 170690 56500 170750 56530
rect 170810 56500 170870 56530
rect 170930 56500 170990 56530
rect 159520 56410 159550 56440
rect 159640 56410 159670 56440
rect 163520 56410 163550 56440
rect 163640 56410 163670 56440
rect 170810 56410 170840 56440
rect 170930 56410 170960 56440
rect 159400 56380 159460 56410
rect 159520 56380 159580 56410
rect 159640 56380 159700 56410
rect 163400 56380 163460 56410
rect 163520 56380 163580 56410
rect 163640 56380 163700 56410
rect 170690 56380 170750 56410
rect 170810 56380 170870 56410
rect 170930 56380 170990 56410
rect 159520 56290 159550 56320
rect 159640 56290 159670 56320
rect 163520 56290 163550 56320
rect 163640 56290 163670 56320
rect 164280 56290 164360 56300
rect 164460 56290 164540 56300
rect 164640 56290 164720 56300
rect 164820 56290 164900 56300
rect 165000 56290 165080 56300
rect 165180 56290 165260 56300
rect 165360 56290 165440 56300
rect 165540 56290 165620 56300
rect 165720 56290 165800 56300
rect 165900 56290 165980 56300
rect 166080 56290 166160 56300
rect 166260 56290 166340 56300
rect 166440 56290 166520 56300
rect 166620 56290 166700 56300
rect 166800 56290 166880 56300
rect 166980 56290 167060 56300
rect 167160 56290 167240 56300
rect 167340 56290 167420 56300
rect 167520 56290 167600 56300
rect 167700 56290 167780 56300
rect 167880 56290 167960 56300
rect 168060 56290 168140 56300
rect 168240 56290 168320 56300
rect 168420 56290 168500 56300
rect 168600 56290 168680 56300
rect 168780 56290 168860 56300
rect 168960 56290 169040 56300
rect 169140 56290 169220 56300
rect 169320 56290 169400 56300
rect 169500 56290 169580 56300
rect 169680 56290 169760 56300
rect 169860 56290 169940 56300
rect 170040 56290 170120 56300
rect 170810 56290 170840 56320
rect 170930 56290 170960 56320
rect 159400 56260 159460 56290
rect 159520 56260 159580 56290
rect 159640 56260 159700 56290
rect 163400 56260 163460 56290
rect 163520 56260 163580 56290
rect 163640 56260 163700 56290
rect 164360 56210 164370 56290
rect 164540 56210 164550 56290
rect 164720 56210 164730 56290
rect 164900 56210 164910 56290
rect 165080 56210 165090 56290
rect 165260 56210 165270 56290
rect 165440 56210 165450 56290
rect 165620 56210 165630 56290
rect 165800 56210 165810 56290
rect 165980 56210 165990 56290
rect 166160 56210 166170 56290
rect 166340 56210 166350 56290
rect 166520 56210 166530 56290
rect 166700 56210 166710 56290
rect 166880 56210 166890 56290
rect 167060 56210 167070 56290
rect 167240 56210 167250 56290
rect 167420 56210 167430 56290
rect 167600 56210 167610 56290
rect 167780 56210 167790 56290
rect 167960 56210 167970 56290
rect 168140 56210 168150 56290
rect 168320 56210 168330 56290
rect 168500 56210 168510 56290
rect 168680 56210 168690 56290
rect 168860 56210 168870 56290
rect 169040 56210 169050 56290
rect 169220 56210 169230 56290
rect 169400 56210 169410 56290
rect 169580 56210 169590 56290
rect 169760 56210 169770 56290
rect 169940 56210 169950 56290
rect 170120 56210 170130 56290
rect 170690 56260 170750 56290
rect 170810 56260 170870 56290
rect 170930 56260 170990 56290
rect 159520 56170 159550 56200
rect 159640 56170 159670 56200
rect 163520 56170 163550 56200
rect 163640 56170 163670 56200
rect 170810 56170 170840 56200
rect 170930 56170 170960 56200
rect 159400 56140 159460 56170
rect 159520 56140 159580 56170
rect 159640 56140 159700 56170
rect 163400 56140 163460 56170
rect 163520 56140 163580 56170
rect 163640 56140 163700 56170
rect 170690 56140 170750 56170
rect 170810 56140 170870 56170
rect 170930 56140 170990 56170
rect 147580 56070 147640 56100
rect 148400 56070 148460 56100
rect 149880 56070 149940 56100
rect 152900 56090 158990 56100
rect 164200 56090 170200 56100
rect 152220 56050 152250 56080
rect 152340 56050 152370 56080
rect 152100 56020 152160 56050
rect 152220 56020 152280 56050
rect 152340 56020 152400 56050
rect 40060 55990 40120 56020
rect 41540 55990 41600 56020
rect 42360 55990 42420 56020
rect 43840 55990 43900 56020
rect 158900 55990 158990 56090
rect 159520 56050 159550 56080
rect 159640 56050 159670 56080
rect 163520 56050 163550 56080
rect 163640 56050 163670 56080
rect 170810 56050 170840 56080
rect 170930 56050 170960 56080
rect 159400 56020 159460 56050
rect 159520 56020 159580 56050
rect 159640 56020 159700 56050
rect 163400 56020 163460 56050
rect 163520 56020 163580 56050
rect 163640 56020 163700 56050
rect 170690 56020 170750 56050
rect 170810 56020 170870 56050
rect 170930 56020 170990 56050
rect 19130 55950 19160 55980
rect 19250 55950 19280 55980
rect 19880 55950 19960 55960
rect 20060 55950 20140 55960
rect 20240 55950 20320 55960
rect 20420 55950 20500 55960
rect 20600 55950 20680 55960
rect 20780 55950 20860 55960
rect 20960 55950 21040 55960
rect 21140 55950 21220 55960
rect 21320 55950 21400 55960
rect 21500 55950 21580 55960
rect 21680 55950 21760 55960
rect 21860 55950 21940 55960
rect 22040 55950 22120 55960
rect 22220 55950 22300 55960
rect 22400 55950 22480 55960
rect 22580 55950 22660 55960
rect 22760 55950 22840 55960
rect 22940 55950 23020 55960
rect 23120 55950 23200 55960
rect 23300 55950 23380 55960
rect 23480 55950 23560 55960
rect 23660 55950 23740 55960
rect 23840 55950 23920 55960
rect 24020 55950 24100 55960
rect 24200 55950 24280 55960
rect 24380 55950 24460 55960
rect 24560 55950 24640 55960
rect 24740 55950 24820 55960
rect 24920 55950 25000 55960
rect 25100 55950 25180 55960
rect 25280 55950 25360 55960
rect 25460 55950 25540 55960
rect 25640 55950 25720 55960
rect 26420 55950 26450 55980
rect 26540 55950 26570 55980
rect 30420 55950 30450 55980
rect 30540 55950 30570 55980
rect 31100 55960 37190 55990
rect 31180 55950 31260 55960
rect 31360 55950 31440 55960
rect 31540 55950 31620 55960
rect 31720 55950 31800 55960
rect 31900 55950 31980 55960
rect 32080 55950 32160 55960
rect 32260 55950 32340 55960
rect 32440 55950 32520 55960
rect 32620 55950 32700 55960
rect 32800 55950 32880 55960
rect 32980 55950 33060 55960
rect 33160 55950 33240 55960
rect 33340 55950 33420 55960
rect 33520 55950 33600 55960
rect 33700 55950 33780 55960
rect 33880 55950 33960 55960
rect 34060 55950 34140 55960
rect 34240 55950 34320 55960
rect 34420 55950 34500 55960
rect 34600 55950 34680 55960
rect 34780 55950 34860 55960
rect 34960 55950 35040 55960
rect 35140 55950 35220 55960
rect 35320 55950 35400 55960
rect 35500 55950 35580 55960
rect 35680 55950 35760 55960
rect 35860 55950 35940 55960
rect 36040 55950 36120 55960
rect 36220 55950 36300 55960
rect 36400 55950 36480 55960
rect 36580 55950 36660 55960
rect 36760 55950 36840 55960
rect 36940 55950 37020 55960
rect 19010 55920 19070 55950
rect 19130 55920 19190 55950
rect 19250 55920 19310 55950
rect 19960 55870 19970 55950
rect 20140 55870 20150 55950
rect 20320 55870 20330 55950
rect 20500 55870 20510 55950
rect 20680 55870 20690 55950
rect 20860 55870 20870 55950
rect 21040 55870 21050 55950
rect 21220 55870 21230 55950
rect 21400 55870 21410 55950
rect 21580 55870 21590 55950
rect 21760 55870 21770 55950
rect 21940 55870 21950 55950
rect 22120 55870 22130 55950
rect 22300 55870 22310 55950
rect 22480 55870 22490 55950
rect 22660 55870 22670 55950
rect 22840 55870 22850 55950
rect 23020 55870 23030 55950
rect 23200 55870 23210 55950
rect 23380 55870 23390 55950
rect 23560 55870 23570 55950
rect 23740 55870 23750 55950
rect 23920 55870 23930 55950
rect 24100 55870 24110 55950
rect 24280 55870 24290 55950
rect 24460 55870 24470 55950
rect 24640 55870 24650 55950
rect 24820 55870 24830 55950
rect 25000 55870 25010 55950
rect 25180 55870 25190 55950
rect 25360 55870 25370 55950
rect 25540 55870 25550 55950
rect 25720 55870 25730 55950
rect 26300 55920 26360 55950
rect 26420 55920 26480 55950
rect 26540 55920 26600 55950
rect 30300 55920 30360 55950
rect 30420 55920 30480 55950
rect 30540 55920 30600 55950
rect 31260 55890 31270 55950
rect 31440 55890 31450 55950
rect 31620 55890 31630 55950
rect 31800 55890 31810 55950
rect 31980 55890 31990 55950
rect 32160 55890 32170 55950
rect 32340 55890 32350 55950
rect 32520 55890 32530 55950
rect 32700 55890 32710 55950
rect 32880 55890 32890 55950
rect 33060 55890 33070 55950
rect 33240 55890 33250 55950
rect 33420 55890 33430 55950
rect 33600 55890 33610 55950
rect 33780 55890 33790 55950
rect 33960 55890 33970 55950
rect 34140 55890 34150 55950
rect 34320 55890 34330 55950
rect 34500 55890 34510 55950
rect 34680 55890 34690 55950
rect 34860 55890 34870 55950
rect 35040 55890 35050 55950
rect 35220 55890 35230 55950
rect 35400 55890 35410 55950
rect 35580 55890 35590 55950
rect 35760 55890 35770 55950
rect 35940 55890 35950 55950
rect 36120 55890 36130 55950
rect 36300 55890 36310 55950
rect 36480 55890 36490 55950
rect 36660 55890 36670 55950
rect 36840 55890 36850 55950
rect 37020 55890 37030 55950
rect 37100 55890 37190 55960
rect 37720 55950 37750 55980
rect 37840 55950 37870 55980
rect 146100 55950 146160 55980
rect 147580 55950 147640 55980
rect 148400 55950 148460 55980
rect 149880 55950 149940 55980
rect 152900 55960 158990 55990
rect 37600 55920 37660 55950
rect 37720 55920 37780 55950
rect 37840 55920 37900 55950
rect 152220 55930 152250 55960
rect 152340 55930 152370 55960
rect 152980 55950 153060 55960
rect 153160 55950 153240 55960
rect 153340 55950 153420 55960
rect 153520 55950 153600 55960
rect 153700 55950 153780 55960
rect 153880 55950 153960 55960
rect 154060 55950 154140 55960
rect 154240 55950 154320 55960
rect 154420 55950 154500 55960
rect 154600 55950 154680 55960
rect 154780 55950 154860 55960
rect 154960 55950 155040 55960
rect 155140 55950 155220 55960
rect 155320 55950 155400 55960
rect 155500 55950 155580 55960
rect 155680 55950 155760 55960
rect 155860 55950 155940 55960
rect 156040 55950 156120 55960
rect 156220 55950 156300 55960
rect 156400 55950 156480 55960
rect 156580 55950 156660 55960
rect 156760 55950 156840 55960
rect 156940 55950 157020 55960
rect 157120 55950 157200 55960
rect 157300 55950 157380 55960
rect 157480 55950 157560 55960
rect 157660 55950 157740 55960
rect 157840 55950 157920 55960
rect 158020 55950 158100 55960
rect 158200 55950 158280 55960
rect 158380 55950 158460 55960
rect 158560 55950 158640 55960
rect 158740 55950 158820 55960
rect 152100 55900 152160 55930
rect 152220 55900 152280 55930
rect 152340 55900 152400 55930
rect 31100 55860 37190 55890
rect 40060 55870 40120 55900
rect 41540 55870 41600 55900
rect 42360 55870 42420 55900
rect 43840 55870 43900 55900
rect 153060 55890 153070 55950
rect 153240 55890 153250 55950
rect 153420 55890 153430 55950
rect 153600 55890 153610 55950
rect 153780 55890 153790 55950
rect 153960 55890 153970 55950
rect 154140 55890 154150 55950
rect 154320 55890 154330 55950
rect 154500 55890 154510 55950
rect 154680 55890 154690 55950
rect 154860 55890 154870 55950
rect 155040 55890 155050 55950
rect 155220 55890 155230 55950
rect 155400 55890 155410 55950
rect 155580 55890 155590 55950
rect 155760 55890 155770 55950
rect 155940 55890 155950 55950
rect 156120 55890 156130 55950
rect 156300 55890 156310 55950
rect 156480 55890 156490 55950
rect 156660 55890 156670 55950
rect 156840 55890 156850 55950
rect 157020 55890 157030 55950
rect 157200 55890 157210 55950
rect 157380 55890 157390 55950
rect 157560 55890 157570 55950
rect 157740 55890 157750 55950
rect 157920 55890 157930 55950
rect 158100 55890 158110 55950
rect 158280 55890 158290 55950
rect 158460 55890 158470 55950
rect 158640 55890 158650 55950
rect 158820 55890 158830 55950
rect 158900 55890 158990 55960
rect 159520 55930 159550 55960
rect 159640 55930 159670 55960
rect 163520 55930 163550 55960
rect 163640 55930 163670 55960
rect 164280 55950 164360 55960
rect 164460 55950 164540 55960
rect 164640 55950 164720 55960
rect 164820 55950 164900 55960
rect 165000 55950 165080 55960
rect 165180 55950 165260 55960
rect 165360 55950 165440 55960
rect 165540 55950 165620 55960
rect 165720 55950 165800 55960
rect 165900 55950 165980 55960
rect 166080 55950 166160 55960
rect 166260 55950 166340 55960
rect 166440 55950 166520 55960
rect 166620 55950 166700 55960
rect 166800 55950 166880 55960
rect 166980 55950 167060 55960
rect 167160 55950 167240 55960
rect 167340 55950 167420 55960
rect 167520 55950 167600 55960
rect 167700 55950 167780 55960
rect 167880 55950 167960 55960
rect 168060 55950 168140 55960
rect 168240 55950 168320 55960
rect 168420 55950 168500 55960
rect 168600 55950 168680 55960
rect 168780 55950 168860 55960
rect 168960 55950 169040 55960
rect 169140 55950 169220 55960
rect 169320 55950 169400 55960
rect 169500 55950 169580 55960
rect 169680 55950 169760 55960
rect 169860 55950 169940 55960
rect 170040 55950 170120 55960
rect 159400 55900 159460 55930
rect 159520 55900 159580 55930
rect 159640 55900 159700 55930
rect 163400 55900 163460 55930
rect 163520 55900 163580 55930
rect 163640 55900 163700 55930
rect 152900 55860 158990 55890
rect 164360 55870 164370 55950
rect 164540 55870 164550 55950
rect 164720 55870 164730 55950
rect 164900 55870 164910 55950
rect 165080 55870 165090 55950
rect 165260 55870 165270 55950
rect 165440 55870 165450 55950
rect 165620 55870 165630 55950
rect 165800 55870 165810 55950
rect 165980 55870 165990 55950
rect 166160 55870 166170 55950
rect 166340 55870 166350 55950
rect 166520 55870 166530 55950
rect 166700 55870 166710 55950
rect 166880 55870 166890 55950
rect 167060 55870 167070 55950
rect 167240 55870 167250 55950
rect 167420 55870 167430 55950
rect 167600 55870 167610 55950
rect 167780 55870 167790 55950
rect 167960 55870 167970 55950
rect 168140 55870 168150 55950
rect 168320 55870 168330 55950
rect 168500 55870 168510 55950
rect 168680 55870 168690 55950
rect 168860 55870 168870 55950
rect 169040 55870 169050 55950
rect 169220 55870 169230 55950
rect 169400 55870 169410 55950
rect 169580 55870 169590 55950
rect 169760 55870 169770 55950
rect 169940 55870 169950 55950
rect 170120 55870 170130 55950
rect 170810 55930 170840 55960
rect 170930 55930 170960 55960
rect 170690 55900 170750 55930
rect 170810 55900 170870 55930
rect 170930 55900 170990 55930
rect 19130 55830 19160 55860
rect 19250 55830 19280 55860
rect 26420 55830 26450 55860
rect 26540 55830 26570 55860
rect 30420 55830 30450 55860
rect 30540 55830 30570 55860
rect 19010 55800 19070 55830
rect 19130 55800 19190 55830
rect 19250 55800 19310 55830
rect 19880 55800 19960 55810
rect 20060 55800 20140 55810
rect 20240 55800 20320 55810
rect 20420 55800 20500 55810
rect 20600 55800 20680 55810
rect 20780 55800 20860 55810
rect 20960 55800 21040 55810
rect 21140 55800 21220 55810
rect 21320 55800 21400 55810
rect 21500 55800 21580 55810
rect 21680 55800 21760 55810
rect 21860 55800 21940 55810
rect 22040 55800 22120 55810
rect 22220 55800 22300 55810
rect 22400 55800 22480 55810
rect 22580 55800 22660 55810
rect 22760 55800 22840 55810
rect 22940 55800 23020 55810
rect 23120 55800 23200 55810
rect 23300 55800 23380 55810
rect 23480 55800 23560 55810
rect 23660 55800 23740 55810
rect 23840 55800 23920 55810
rect 24020 55800 24100 55810
rect 24200 55800 24280 55810
rect 24380 55800 24460 55810
rect 24560 55800 24640 55810
rect 24740 55800 24820 55810
rect 24920 55800 25000 55810
rect 25100 55800 25180 55810
rect 25280 55800 25360 55810
rect 25460 55800 25540 55810
rect 25640 55800 25720 55810
rect 26300 55800 26360 55830
rect 26420 55800 26480 55830
rect 26540 55800 26600 55830
rect 30300 55800 30360 55830
rect 30420 55800 30480 55830
rect 30540 55800 30600 55830
rect 31180 55800 31260 55810
rect 31360 55800 31440 55810
rect 31540 55800 31620 55810
rect 31720 55800 31800 55810
rect 31900 55800 31980 55810
rect 32080 55800 32160 55810
rect 32260 55800 32340 55810
rect 32440 55800 32520 55810
rect 32620 55800 32700 55810
rect 32800 55800 32880 55810
rect 32980 55800 33060 55810
rect 33160 55800 33240 55810
rect 33340 55800 33420 55810
rect 33520 55800 33600 55810
rect 33700 55800 33780 55810
rect 33880 55800 33960 55810
rect 34060 55800 34140 55810
rect 34240 55800 34320 55810
rect 34420 55800 34500 55810
rect 34600 55800 34680 55810
rect 34780 55800 34860 55810
rect 34960 55800 35040 55810
rect 35140 55800 35220 55810
rect 35320 55800 35400 55810
rect 35500 55800 35580 55810
rect 35680 55800 35760 55810
rect 35860 55800 35940 55810
rect 36040 55800 36120 55810
rect 36220 55800 36300 55810
rect 36400 55800 36480 55810
rect 36580 55800 36660 55810
rect 36760 55800 36840 55810
rect 36940 55800 37020 55810
rect 19130 55710 19160 55740
rect 19250 55710 19280 55740
rect 19960 55720 19970 55800
rect 20140 55720 20150 55800
rect 20320 55720 20330 55800
rect 20500 55720 20510 55800
rect 20680 55720 20690 55800
rect 20860 55720 20870 55800
rect 21040 55720 21050 55800
rect 21220 55720 21230 55800
rect 21400 55720 21410 55800
rect 21580 55720 21590 55800
rect 21760 55720 21770 55800
rect 21940 55720 21950 55800
rect 22120 55720 22130 55800
rect 22300 55720 22310 55800
rect 22480 55720 22490 55800
rect 22660 55720 22670 55800
rect 22840 55720 22850 55800
rect 23020 55720 23030 55800
rect 23200 55720 23210 55800
rect 23380 55720 23390 55800
rect 23560 55720 23570 55800
rect 23740 55720 23750 55800
rect 23920 55720 23930 55800
rect 24100 55720 24110 55800
rect 24280 55720 24290 55800
rect 24460 55720 24470 55800
rect 24640 55720 24650 55800
rect 24820 55720 24830 55800
rect 25000 55720 25010 55800
rect 25180 55720 25190 55800
rect 25360 55720 25370 55800
rect 25540 55720 25550 55800
rect 25720 55720 25730 55800
rect 26420 55710 26450 55740
rect 26540 55710 26570 55740
rect 30420 55710 30450 55740
rect 30540 55710 30570 55740
rect 31260 55720 31270 55800
rect 31440 55720 31450 55800
rect 31620 55720 31630 55800
rect 31800 55720 31810 55800
rect 31980 55720 31990 55800
rect 32160 55720 32170 55800
rect 32340 55720 32350 55800
rect 32520 55720 32530 55800
rect 32700 55720 32710 55800
rect 32880 55720 32890 55800
rect 33060 55720 33070 55800
rect 33240 55720 33250 55800
rect 33420 55720 33430 55800
rect 33600 55720 33610 55800
rect 33780 55720 33790 55800
rect 33960 55720 33970 55800
rect 34140 55720 34150 55800
rect 34320 55720 34330 55800
rect 34500 55720 34510 55800
rect 34680 55720 34690 55800
rect 34860 55720 34870 55800
rect 35040 55720 35050 55800
rect 35220 55720 35230 55800
rect 35400 55720 35410 55800
rect 35580 55720 35590 55800
rect 35760 55720 35770 55800
rect 35940 55720 35950 55800
rect 36120 55720 36130 55800
rect 36300 55720 36310 55800
rect 36480 55720 36490 55800
rect 36660 55720 36670 55800
rect 36840 55720 36850 55800
rect 37020 55720 37030 55800
rect 19010 55680 19070 55710
rect 19130 55680 19190 55710
rect 19250 55680 19310 55710
rect 26300 55680 26360 55710
rect 26420 55680 26480 55710
rect 26540 55680 26600 55710
rect 30300 55680 30360 55710
rect 30420 55680 30480 55710
rect 30540 55680 30600 55710
rect 37100 55660 37190 55860
rect 37720 55830 37750 55860
rect 37840 55830 37870 55860
rect 146100 55830 146160 55860
rect 147580 55830 147640 55860
rect 148400 55830 148460 55860
rect 149880 55830 149940 55860
rect 37600 55800 37660 55830
rect 37720 55800 37780 55830
rect 37840 55800 37900 55830
rect 152220 55810 152250 55840
rect 152340 55810 152370 55840
rect 152100 55780 152160 55810
rect 152220 55780 152280 55810
rect 152340 55780 152400 55810
rect 152980 55800 153060 55810
rect 153160 55800 153240 55810
rect 153340 55800 153420 55810
rect 153520 55800 153600 55810
rect 153700 55800 153780 55810
rect 153880 55800 153960 55810
rect 154060 55800 154140 55810
rect 154240 55800 154320 55810
rect 154420 55800 154500 55810
rect 154600 55800 154680 55810
rect 154780 55800 154860 55810
rect 154960 55800 155040 55810
rect 155140 55800 155220 55810
rect 155320 55800 155400 55810
rect 155500 55800 155580 55810
rect 155680 55800 155760 55810
rect 155860 55800 155940 55810
rect 156040 55800 156120 55810
rect 156220 55800 156300 55810
rect 156400 55800 156480 55810
rect 156580 55800 156660 55810
rect 156760 55800 156840 55810
rect 156940 55800 157020 55810
rect 157120 55800 157200 55810
rect 157300 55800 157380 55810
rect 157480 55800 157560 55810
rect 157660 55800 157740 55810
rect 157840 55800 157920 55810
rect 158020 55800 158100 55810
rect 158200 55800 158280 55810
rect 158380 55800 158460 55810
rect 158560 55800 158640 55810
rect 158740 55800 158820 55810
rect 40060 55750 40120 55780
rect 41540 55750 41600 55780
rect 42360 55750 42420 55780
rect 43840 55750 43900 55780
rect 37720 55710 37750 55740
rect 37840 55710 37870 55740
rect 146100 55710 146160 55740
rect 147580 55710 147640 55740
rect 148400 55710 148460 55740
rect 149880 55710 149940 55740
rect 153060 55720 153070 55800
rect 153240 55720 153250 55800
rect 153420 55720 153430 55800
rect 153600 55720 153610 55800
rect 153780 55720 153790 55800
rect 153960 55720 153970 55800
rect 154140 55720 154150 55800
rect 154320 55720 154330 55800
rect 154500 55720 154510 55800
rect 154680 55720 154690 55800
rect 154860 55720 154870 55800
rect 155040 55720 155050 55800
rect 155220 55720 155230 55800
rect 155400 55720 155410 55800
rect 155580 55720 155590 55800
rect 155760 55720 155770 55800
rect 155940 55720 155950 55800
rect 156120 55720 156130 55800
rect 156300 55720 156310 55800
rect 156480 55720 156490 55800
rect 156660 55720 156670 55800
rect 156840 55720 156850 55800
rect 157020 55720 157030 55800
rect 157200 55720 157210 55800
rect 157380 55720 157390 55800
rect 157560 55720 157570 55800
rect 157740 55720 157750 55800
rect 157920 55720 157930 55800
rect 158100 55720 158110 55800
rect 158280 55720 158290 55800
rect 158460 55720 158470 55800
rect 158640 55720 158650 55800
rect 158820 55720 158830 55800
rect 37600 55680 37660 55710
rect 37720 55680 37780 55710
rect 37840 55680 37900 55710
rect 152220 55690 152250 55720
rect 152340 55690 152370 55720
rect 152100 55660 152160 55690
rect 152220 55660 152280 55690
rect 152340 55660 152400 55690
rect 158900 55660 158990 55860
rect 159520 55810 159550 55840
rect 159640 55810 159670 55840
rect 163520 55810 163550 55840
rect 163640 55810 163670 55840
rect 170810 55810 170840 55840
rect 170930 55810 170960 55840
rect 159400 55780 159460 55810
rect 159520 55780 159580 55810
rect 159640 55780 159700 55810
rect 163400 55780 163460 55810
rect 163520 55780 163580 55810
rect 163640 55780 163700 55810
rect 164280 55800 164360 55810
rect 164460 55800 164540 55810
rect 164640 55800 164720 55810
rect 164820 55800 164900 55810
rect 165000 55800 165080 55810
rect 165180 55800 165260 55810
rect 165360 55800 165440 55810
rect 165540 55800 165620 55810
rect 165720 55800 165800 55810
rect 165900 55800 165980 55810
rect 166080 55800 166160 55810
rect 166260 55800 166340 55810
rect 166440 55800 166520 55810
rect 166620 55800 166700 55810
rect 166800 55800 166880 55810
rect 166980 55800 167060 55810
rect 167160 55800 167240 55810
rect 167340 55800 167420 55810
rect 167520 55800 167600 55810
rect 167700 55800 167780 55810
rect 167880 55800 167960 55810
rect 168060 55800 168140 55810
rect 168240 55800 168320 55810
rect 168420 55800 168500 55810
rect 168600 55800 168680 55810
rect 168780 55800 168860 55810
rect 168960 55800 169040 55810
rect 169140 55800 169220 55810
rect 169320 55800 169400 55810
rect 169500 55800 169580 55810
rect 169680 55800 169760 55810
rect 169860 55800 169940 55810
rect 170040 55800 170120 55810
rect 164360 55720 164370 55800
rect 164540 55720 164550 55800
rect 164720 55720 164730 55800
rect 164900 55720 164910 55800
rect 165080 55720 165090 55800
rect 165260 55720 165270 55800
rect 165440 55720 165450 55800
rect 165620 55720 165630 55800
rect 165800 55720 165810 55800
rect 165980 55720 165990 55800
rect 166160 55720 166170 55800
rect 166340 55720 166350 55800
rect 166520 55720 166530 55800
rect 166700 55720 166710 55800
rect 166880 55720 166890 55800
rect 167060 55720 167070 55800
rect 167240 55720 167250 55800
rect 167420 55720 167430 55800
rect 167600 55720 167610 55800
rect 167780 55720 167790 55800
rect 167960 55720 167970 55800
rect 168140 55720 168150 55800
rect 168320 55720 168330 55800
rect 168500 55720 168510 55800
rect 168680 55720 168690 55800
rect 168860 55720 168870 55800
rect 169040 55720 169050 55800
rect 169220 55720 169230 55800
rect 169400 55720 169410 55800
rect 169580 55720 169590 55800
rect 169760 55720 169770 55800
rect 169940 55720 169950 55800
rect 170120 55720 170130 55800
rect 170690 55780 170750 55810
rect 170810 55780 170870 55810
rect 170930 55780 170990 55810
rect 159520 55690 159550 55720
rect 159640 55690 159670 55720
rect 163520 55690 163550 55720
rect 163640 55690 163670 55720
rect 170810 55690 170840 55720
rect 170930 55690 170960 55720
rect 159400 55660 159460 55690
rect 159520 55660 159580 55690
rect 159640 55660 159700 55690
rect 163400 55660 163460 55690
rect 163520 55660 163580 55690
rect 163640 55660 163700 55690
rect 170690 55660 170750 55690
rect 170810 55660 170870 55690
rect 170930 55660 170990 55690
rect 19880 55650 19960 55660
rect 20060 55650 20140 55660
rect 20240 55650 20320 55660
rect 20420 55650 20500 55660
rect 20600 55650 20680 55660
rect 20780 55650 20860 55660
rect 20960 55650 21040 55660
rect 21140 55650 21220 55660
rect 21320 55650 21400 55660
rect 21500 55650 21580 55660
rect 21680 55650 21760 55660
rect 21860 55650 21940 55660
rect 22040 55650 22120 55660
rect 22220 55650 22300 55660
rect 22400 55650 22480 55660
rect 22580 55650 22660 55660
rect 22760 55650 22840 55660
rect 22940 55650 23020 55660
rect 23120 55650 23200 55660
rect 23300 55650 23380 55660
rect 23480 55650 23560 55660
rect 23660 55650 23740 55660
rect 23840 55650 23920 55660
rect 24020 55650 24100 55660
rect 24200 55650 24280 55660
rect 24380 55650 24460 55660
rect 24560 55650 24640 55660
rect 24740 55650 24820 55660
rect 24920 55650 25000 55660
rect 25100 55650 25180 55660
rect 25280 55650 25360 55660
rect 25460 55650 25540 55660
rect 25640 55650 25720 55660
rect 19130 55590 19160 55620
rect 19250 55590 19280 55620
rect 19010 55560 19070 55590
rect 19130 55560 19190 55590
rect 19250 55560 19310 55590
rect 19960 55570 19970 55650
rect 20140 55570 20150 55650
rect 20320 55570 20330 55650
rect 20500 55570 20510 55650
rect 20680 55570 20690 55650
rect 20860 55570 20870 55650
rect 21040 55570 21050 55650
rect 21220 55570 21230 55650
rect 21400 55570 21410 55650
rect 21580 55570 21590 55650
rect 21760 55570 21770 55650
rect 21940 55570 21950 55650
rect 22120 55570 22130 55650
rect 22300 55570 22310 55650
rect 22480 55570 22490 55650
rect 22660 55570 22670 55650
rect 22840 55570 22850 55650
rect 23020 55570 23030 55650
rect 23200 55570 23210 55650
rect 23380 55570 23390 55650
rect 23560 55570 23570 55650
rect 23740 55570 23750 55650
rect 23920 55570 23930 55650
rect 24100 55570 24110 55650
rect 24280 55570 24290 55650
rect 24460 55570 24470 55650
rect 24640 55570 24650 55650
rect 24820 55570 24830 55650
rect 25000 55570 25010 55650
rect 25180 55570 25190 55650
rect 25360 55570 25370 55650
rect 25540 55570 25550 55650
rect 25720 55570 25730 55650
rect 31100 55630 37190 55660
rect 40060 55630 40120 55660
rect 41540 55630 41600 55660
rect 42360 55630 42420 55660
rect 43840 55630 43900 55660
rect 152900 55630 158990 55660
rect 164280 55650 164360 55660
rect 164460 55650 164540 55660
rect 164640 55650 164720 55660
rect 164820 55650 164900 55660
rect 165000 55650 165080 55660
rect 165180 55650 165260 55660
rect 165360 55650 165440 55660
rect 165540 55650 165620 55660
rect 165720 55650 165800 55660
rect 165900 55650 165980 55660
rect 166080 55650 166160 55660
rect 166260 55650 166340 55660
rect 166440 55650 166520 55660
rect 166620 55650 166700 55660
rect 166800 55650 166880 55660
rect 166980 55650 167060 55660
rect 167160 55650 167240 55660
rect 167340 55650 167420 55660
rect 167520 55650 167600 55660
rect 167700 55650 167780 55660
rect 167880 55650 167960 55660
rect 168060 55650 168140 55660
rect 168240 55650 168320 55660
rect 168420 55650 168500 55660
rect 168600 55650 168680 55660
rect 168780 55650 168860 55660
rect 168960 55650 169040 55660
rect 169140 55650 169220 55660
rect 169320 55650 169400 55660
rect 169500 55650 169580 55660
rect 169680 55650 169760 55660
rect 169860 55650 169940 55660
rect 170040 55650 170120 55660
rect 26420 55590 26450 55620
rect 26540 55590 26570 55620
rect 30420 55590 30450 55620
rect 30540 55590 30570 55620
rect 26300 55560 26360 55590
rect 26420 55560 26480 55590
rect 26540 55560 26600 55590
rect 30300 55560 30360 55590
rect 30420 55560 30480 55590
rect 30540 55560 30600 55590
rect 31260 55570 31270 55630
rect 31440 55570 31450 55630
rect 31620 55570 31630 55630
rect 31800 55570 31810 55630
rect 31980 55570 31990 55630
rect 32160 55570 32170 55630
rect 32340 55570 32350 55630
rect 32520 55570 32530 55630
rect 32700 55570 32710 55630
rect 32880 55570 32890 55630
rect 33060 55570 33070 55630
rect 33240 55570 33250 55630
rect 33420 55570 33430 55630
rect 33600 55570 33610 55630
rect 33780 55570 33790 55630
rect 33960 55570 33970 55630
rect 34140 55570 34150 55630
rect 34320 55570 34330 55630
rect 34500 55570 34510 55630
rect 34680 55570 34690 55630
rect 34860 55570 34870 55630
rect 35040 55570 35050 55630
rect 35220 55570 35230 55630
rect 35400 55570 35410 55630
rect 35580 55570 35590 55630
rect 35760 55570 35770 55630
rect 35940 55570 35950 55630
rect 36120 55570 36130 55630
rect 36300 55570 36310 55630
rect 36480 55570 36490 55630
rect 36660 55570 36670 55630
rect 36840 55570 36850 55630
rect 37020 55570 37030 55630
rect 37100 55560 37190 55630
rect 37720 55590 37750 55620
rect 37840 55590 37870 55620
rect 146100 55590 146160 55620
rect 147580 55590 147640 55620
rect 148400 55590 148460 55620
rect 149880 55590 149940 55620
rect 37600 55560 37660 55590
rect 37720 55560 37780 55590
rect 37840 55560 37900 55590
rect 152220 55570 152250 55600
rect 152340 55570 152370 55600
rect 153060 55570 153070 55630
rect 153240 55570 153250 55630
rect 153420 55570 153430 55630
rect 153600 55570 153610 55630
rect 153780 55570 153790 55630
rect 153960 55570 153970 55630
rect 154140 55570 154150 55630
rect 154320 55570 154330 55630
rect 154500 55570 154510 55630
rect 154680 55570 154690 55630
rect 154860 55570 154870 55630
rect 155040 55570 155050 55630
rect 155220 55570 155230 55630
rect 155400 55570 155410 55630
rect 155580 55570 155590 55630
rect 155760 55570 155770 55630
rect 155940 55570 155950 55630
rect 156120 55570 156130 55630
rect 156300 55570 156310 55630
rect 156480 55570 156490 55630
rect 156660 55570 156670 55630
rect 156840 55570 156850 55630
rect 157020 55570 157030 55630
rect 157200 55570 157210 55630
rect 157380 55570 157390 55630
rect 157560 55570 157570 55630
rect 157740 55570 157750 55630
rect 157920 55570 157930 55630
rect 158100 55570 158110 55630
rect 158280 55570 158290 55630
rect 158460 55570 158470 55630
rect 158640 55570 158650 55630
rect 158820 55570 158830 55630
rect 31100 55530 37190 55560
rect 152100 55540 152160 55570
rect 152220 55540 152280 55570
rect 152340 55540 152400 55570
rect 158900 55560 158990 55630
rect 159520 55570 159550 55600
rect 159640 55570 159670 55600
rect 163520 55570 163550 55600
rect 163640 55570 163670 55600
rect 164360 55570 164370 55650
rect 164540 55570 164550 55650
rect 164720 55570 164730 55650
rect 164900 55570 164910 55650
rect 165080 55570 165090 55650
rect 165260 55570 165270 55650
rect 165440 55570 165450 55650
rect 165620 55570 165630 55650
rect 165800 55570 165810 55650
rect 165980 55570 165990 55650
rect 166160 55570 166170 55650
rect 166340 55570 166350 55650
rect 166520 55570 166530 55650
rect 166700 55570 166710 55650
rect 166880 55570 166890 55650
rect 167060 55570 167070 55650
rect 167240 55570 167250 55650
rect 167420 55570 167430 55650
rect 167600 55570 167610 55650
rect 167780 55570 167790 55650
rect 167960 55570 167970 55650
rect 168140 55570 168150 55650
rect 168320 55570 168330 55650
rect 168500 55570 168510 55650
rect 168680 55570 168690 55650
rect 168860 55570 168870 55650
rect 169040 55570 169050 55650
rect 169220 55570 169230 55650
rect 169400 55570 169410 55650
rect 169580 55570 169590 55650
rect 169760 55570 169770 55650
rect 169940 55570 169950 55650
rect 170120 55570 170130 55650
rect 170810 55570 170840 55600
rect 170930 55570 170960 55600
rect 37100 55520 37190 55530
rect 19800 55510 25800 55520
rect 31100 55510 37190 55520
rect 40060 55510 40120 55540
rect 41540 55510 41600 55540
rect 42360 55510 42420 55540
rect 43840 55510 43900 55540
rect 152900 55530 158990 55560
rect 159400 55540 159460 55570
rect 159520 55540 159580 55570
rect 159640 55540 159700 55570
rect 163400 55540 163460 55570
rect 163520 55540 163580 55570
rect 163640 55540 163700 55570
rect 170690 55540 170750 55570
rect 170810 55540 170870 55570
rect 170930 55540 170990 55570
rect 158900 55520 158990 55530
rect 152900 55510 158990 55520
rect 164200 55510 170200 55520
rect 19130 55470 19160 55500
rect 19250 55470 19280 55500
rect 26420 55470 26450 55500
rect 26540 55470 26570 55500
rect 30420 55470 30450 55500
rect 30540 55470 30570 55500
rect 19010 55440 19070 55470
rect 19130 55440 19190 55470
rect 19250 55440 19310 55470
rect 26300 55440 26360 55470
rect 26420 55440 26480 55470
rect 26540 55440 26600 55470
rect 30300 55440 30360 55470
rect 30420 55440 30480 55470
rect 30540 55440 30600 55470
rect 19130 55350 19160 55380
rect 19250 55350 19280 55380
rect 26420 55350 26450 55380
rect 26540 55350 26570 55380
rect 30420 55350 30450 55380
rect 30540 55350 30570 55380
rect 19010 55320 19070 55350
rect 19130 55320 19190 55350
rect 19250 55320 19310 55350
rect 26300 55320 26360 55350
rect 26420 55320 26480 55350
rect 26540 55320 26600 55350
rect 30300 55320 30360 55350
rect 30420 55320 30480 55350
rect 30540 55320 30600 55350
rect 31180 55330 31260 55340
rect 31360 55330 31440 55340
rect 31540 55330 31620 55340
rect 31720 55330 31800 55340
rect 31900 55330 31980 55340
rect 32080 55330 32160 55340
rect 32260 55330 32340 55340
rect 32440 55330 32520 55340
rect 32620 55330 32700 55340
rect 32800 55330 32880 55340
rect 32980 55330 33060 55340
rect 33160 55330 33240 55340
rect 33340 55330 33420 55340
rect 33520 55330 33600 55340
rect 33700 55330 33780 55340
rect 33880 55330 33960 55340
rect 34060 55330 34140 55340
rect 34240 55330 34320 55340
rect 34420 55330 34500 55340
rect 34600 55330 34680 55340
rect 34780 55330 34860 55340
rect 34960 55330 35040 55340
rect 35140 55330 35220 55340
rect 35320 55330 35400 55340
rect 35500 55330 35580 55340
rect 35680 55330 35760 55340
rect 35860 55330 35940 55340
rect 36040 55330 36120 55340
rect 36220 55330 36300 55340
rect 36400 55330 36480 55340
rect 36580 55330 36660 55340
rect 36760 55330 36840 55340
rect 36940 55330 37020 55340
rect 19880 55310 19960 55320
rect 20060 55310 20140 55320
rect 20240 55310 20320 55320
rect 20420 55310 20500 55320
rect 20600 55310 20680 55320
rect 20780 55310 20860 55320
rect 20960 55310 21040 55320
rect 21140 55310 21220 55320
rect 21320 55310 21400 55320
rect 21500 55310 21580 55320
rect 21680 55310 21760 55320
rect 21860 55310 21940 55320
rect 22040 55310 22120 55320
rect 22220 55310 22300 55320
rect 22400 55310 22480 55320
rect 22580 55310 22660 55320
rect 22760 55310 22840 55320
rect 22940 55310 23020 55320
rect 23120 55310 23200 55320
rect 23300 55310 23380 55320
rect 23480 55310 23560 55320
rect 23660 55310 23740 55320
rect 23840 55310 23920 55320
rect 24020 55310 24100 55320
rect 24200 55310 24280 55320
rect 24380 55310 24460 55320
rect 24560 55310 24640 55320
rect 24740 55310 24820 55320
rect 24920 55310 25000 55320
rect 25100 55310 25180 55320
rect 25280 55310 25360 55320
rect 25460 55310 25540 55320
rect 25640 55310 25720 55320
rect 19130 55230 19160 55260
rect 19250 55230 19280 55260
rect 19960 55230 19970 55310
rect 20140 55230 20150 55310
rect 20320 55230 20330 55310
rect 20500 55230 20510 55310
rect 20680 55230 20690 55310
rect 20860 55230 20870 55310
rect 21040 55230 21050 55310
rect 21220 55230 21230 55310
rect 21400 55230 21410 55310
rect 21580 55230 21590 55310
rect 21760 55230 21770 55310
rect 21940 55230 21950 55310
rect 22120 55230 22130 55310
rect 22300 55230 22310 55310
rect 22480 55230 22490 55310
rect 22660 55230 22670 55310
rect 22840 55230 22850 55310
rect 23020 55230 23030 55310
rect 23200 55230 23210 55310
rect 23380 55230 23390 55310
rect 23560 55230 23570 55310
rect 23740 55230 23750 55310
rect 23920 55230 23930 55310
rect 24100 55230 24110 55310
rect 24280 55230 24290 55310
rect 24460 55230 24470 55310
rect 24640 55230 24650 55310
rect 24820 55230 24830 55310
rect 25000 55230 25010 55310
rect 25180 55230 25190 55310
rect 25360 55230 25370 55310
rect 25540 55230 25550 55310
rect 25720 55230 25730 55310
rect 26420 55230 26450 55260
rect 26540 55230 26570 55260
rect 30420 55230 30450 55260
rect 30540 55230 30570 55260
rect 31260 55250 31270 55330
rect 31440 55250 31450 55330
rect 31620 55250 31630 55330
rect 31800 55250 31810 55330
rect 31980 55250 31990 55330
rect 32160 55250 32170 55330
rect 32340 55250 32350 55330
rect 32520 55250 32530 55330
rect 32700 55250 32710 55330
rect 32880 55250 32890 55330
rect 33060 55250 33070 55330
rect 33240 55250 33250 55330
rect 33420 55250 33430 55330
rect 33600 55250 33610 55330
rect 33780 55250 33790 55330
rect 33960 55250 33970 55330
rect 34140 55250 34150 55330
rect 34320 55250 34330 55330
rect 34500 55250 34510 55330
rect 34680 55250 34690 55330
rect 34860 55250 34870 55330
rect 35040 55250 35050 55330
rect 35220 55250 35230 55330
rect 35400 55250 35410 55330
rect 35580 55250 35590 55330
rect 35760 55250 35770 55330
rect 35940 55250 35950 55330
rect 36120 55250 36130 55330
rect 36300 55250 36310 55330
rect 36480 55250 36490 55330
rect 36660 55250 36670 55330
rect 36840 55250 36850 55330
rect 37020 55250 37030 55330
rect 19010 55200 19070 55230
rect 19130 55200 19190 55230
rect 19250 55200 19310 55230
rect 26300 55200 26360 55230
rect 26420 55200 26480 55230
rect 26540 55200 26600 55230
rect 30300 55200 30360 55230
rect 30420 55200 30480 55230
rect 30540 55200 30600 55230
rect 19130 55110 19160 55140
rect 19250 55110 19280 55140
rect 26420 55110 26450 55140
rect 26540 55110 26570 55140
rect 30420 55110 30450 55140
rect 30540 55110 30570 55140
rect 19010 55080 19070 55110
rect 19130 55080 19190 55110
rect 19250 55080 19310 55110
rect 26300 55080 26360 55110
rect 26420 55080 26480 55110
rect 26540 55080 26600 55110
rect 30300 55080 30360 55110
rect 30420 55080 30480 55110
rect 30540 55080 30600 55110
rect 19130 54990 19160 55020
rect 19250 54990 19280 55020
rect 19880 55010 19960 55020
rect 20060 55010 20140 55020
rect 20240 55010 20320 55020
rect 20420 55010 20500 55020
rect 20600 55010 20680 55020
rect 20780 55010 20860 55020
rect 20960 55010 21040 55020
rect 21140 55010 21220 55020
rect 21320 55010 21400 55020
rect 21500 55010 21580 55020
rect 21680 55010 21760 55020
rect 21860 55010 21940 55020
rect 22040 55010 22120 55020
rect 22220 55010 22300 55020
rect 22400 55010 22480 55020
rect 22580 55010 22660 55020
rect 22760 55010 22840 55020
rect 22940 55010 23020 55020
rect 23120 55010 23200 55020
rect 23300 55010 23380 55020
rect 23480 55010 23560 55020
rect 23660 55010 23740 55020
rect 23840 55010 23920 55020
rect 24020 55010 24100 55020
rect 24200 55010 24280 55020
rect 24380 55010 24460 55020
rect 24560 55010 24640 55020
rect 24740 55010 24820 55020
rect 24920 55010 25000 55020
rect 25100 55010 25180 55020
rect 25280 55010 25360 55020
rect 25460 55010 25540 55020
rect 25640 55010 25720 55020
rect 19010 54960 19070 54990
rect 19130 54960 19190 54990
rect 19250 54960 19310 54990
rect 19960 54930 19970 55010
rect 20140 54930 20150 55010
rect 20320 54930 20330 55010
rect 20500 54930 20510 55010
rect 20680 54930 20690 55010
rect 20860 54930 20870 55010
rect 21040 54930 21050 55010
rect 21220 54930 21230 55010
rect 21400 54930 21410 55010
rect 21580 54930 21590 55010
rect 21760 54930 21770 55010
rect 21940 54930 21950 55010
rect 22120 54930 22130 55010
rect 22300 54930 22310 55010
rect 22480 54930 22490 55010
rect 22660 54930 22670 55010
rect 22840 54930 22850 55010
rect 23020 54930 23030 55010
rect 23200 54930 23210 55010
rect 23380 54930 23390 55010
rect 23560 54930 23570 55010
rect 23740 54930 23750 55010
rect 23920 54930 23930 55010
rect 24100 54930 24110 55010
rect 24280 54930 24290 55010
rect 24460 54930 24470 55010
rect 24640 54930 24650 55010
rect 24820 54930 24830 55010
rect 25000 54930 25010 55010
rect 25180 54930 25190 55010
rect 25360 54930 25370 55010
rect 25540 54930 25550 55010
rect 25720 54930 25730 55010
rect 26420 54990 26450 55020
rect 26540 54990 26570 55020
rect 30420 54990 30450 55020
rect 30540 54990 30570 55020
rect 31180 55010 31260 55020
rect 31360 55010 31440 55020
rect 31540 55010 31620 55020
rect 31720 55010 31800 55020
rect 31900 55010 31980 55020
rect 32080 55010 32160 55020
rect 32260 55010 32340 55020
rect 32440 55010 32520 55020
rect 32620 55010 32700 55020
rect 32800 55010 32880 55020
rect 32980 55010 33060 55020
rect 33160 55010 33240 55020
rect 33340 55010 33420 55020
rect 33520 55010 33600 55020
rect 33700 55010 33780 55020
rect 33880 55010 33960 55020
rect 34060 55010 34140 55020
rect 34240 55010 34320 55020
rect 34420 55010 34500 55020
rect 34600 55010 34680 55020
rect 34780 55010 34860 55020
rect 34960 55010 35040 55020
rect 35140 55010 35220 55020
rect 35320 55010 35400 55020
rect 35500 55010 35580 55020
rect 35680 55010 35760 55020
rect 35860 55010 35940 55020
rect 36040 55010 36120 55020
rect 36220 55010 36300 55020
rect 36400 55010 36480 55020
rect 36580 55010 36660 55020
rect 36760 55010 36840 55020
rect 36940 55010 37020 55020
rect 26300 54960 26360 54990
rect 26420 54960 26480 54990
rect 26540 54960 26600 54990
rect 30300 54960 30360 54990
rect 30420 54960 30480 54990
rect 30540 54960 30600 54990
rect 31260 54930 31270 55010
rect 31440 54930 31450 55010
rect 31620 54930 31630 55010
rect 31800 54930 31810 55010
rect 31980 54930 31990 55010
rect 32160 54930 32170 55010
rect 32340 54930 32350 55010
rect 32520 54930 32530 55010
rect 32700 54930 32710 55010
rect 32880 54930 32890 55010
rect 33060 54930 33070 55010
rect 33240 54930 33250 55010
rect 33420 54930 33430 55010
rect 33600 54930 33610 55010
rect 33780 54930 33790 55010
rect 33960 54930 33970 55010
rect 34140 54930 34150 55010
rect 34320 54930 34330 55010
rect 34500 54930 34510 55010
rect 34680 54930 34690 55010
rect 34860 54930 34870 55010
rect 35040 54930 35050 55010
rect 35220 54930 35230 55010
rect 35400 54930 35410 55010
rect 35580 54930 35590 55010
rect 35760 54930 35770 55010
rect 35940 54930 35950 55010
rect 36120 54930 36130 55010
rect 36300 54930 36310 55010
rect 36480 54930 36490 55010
rect 36660 54930 36670 55010
rect 36840 54930 36850 55010
rect 37020 54930 37030 55010
rect 19130 54870 19160 54900
rect 19250 54870 19280 54900
rect 26420 54870 26450 54900
rect 26540 54870 26570 54900
rect 30420 54870 30450 54900
rect 30540 54870 30570 54900
rect 19010 54840 19070 54870
rect 19130 54840 19190 54870
rect 19250 54840 19310 54870
rect 26300 54840 26360 54870
rect 26420 54840 26480 54870
rect 26540 54840 26600 54870
rect 30300 54840 30360 54870
rect 30420 54840 30480 54870
rect 30540 54840 30600 54870
rect 37100 54840 37190 55510
rect 37720 55470 37750 55500
rect 37840 55470 37870 55500
rect 146100 55470 146160 55500
rect 147580 55470 147640 55500
rect 148400 55470 148460 55500
rect 149880 55470 149940 55500
rect 37600 55440 37660 55470
rect 37720 55440 37780 55470
rect 37840 55440 37900 55470
rect 152220 55450 152250 55480
rect 152340 55450 152370 55480
rect 152100 55420 152160 55450
rect 152220 55420 152280 55450
rect 152340 55420 152400 55450
rect 40060 55390 40120 55420
rect 41540 55390 41600 55420
rect 42360 55390 42420 55420
rect 43840 55390 43900 55420
rect 37720 55350 37750 55380
rect 37840 55350 37870 55380
rect 146100 55350 146160 55380
rect 147580 55350 147640 55380
rect 148400 55350 148460 55380
rect 149880 55350 149940 55380
rect 37600 55320 37660 55350
rect 37720 55320 37780 55350
rect 37840 55320 37900 55350
rect 152220 55330 152250 55360
rect 152340 55330 152370 55360
rect 152980 55330 153060 55340
rect 153160 55330 153240 55340
rect 153340 55330 153420 55340
rect 153520 55330 153600 55340
rect 153700 55330 153780 55340
rect 153880 55330 153960 55340
rect 154060 55330 154140 55340
rect 154240 55330 154320 55340
rect 154420 55330 154500 55340
rect 154600 55330 154680 55340
rect 154780 55330 154860 55340
rect 154960 55330 155040 55340
rect 155140 55330 155220 55340
rect 155320 55330 155400 55340
rect 155500 55330 155580 55340
rect 155680 55330 155760 55340
rect 155860 55330 155940 55340
rect 156040 55330 156120 55340
rect 156220 55330 156300 55340
rect 156400 55330 156480 55340
rect 156580 55330 156660 55340
rect 156760 55330 156840 55340
rect 156940 55330 157020 55340
rect 157120 55330 157200 55340
rect 157300 55330 157380 55340
rect 157480 55330 157560 55340
rect 157660 55330 157740 55340
rect 157840 55330 157920 55340
rect 158020 55330 158100 55340
rect 158200 55330 158280 55340
rect 158380 55330 158460 55340
rect 158560 55330 158640 55340
rect 158740 55330 158820 55340
rect 152100 55300 152160 55330
rect 152220 55300 152280 55330
rect 152340 55300 152400 55330
rect 40060 55270 40120 55300
rect 41540 55270 41600 55300
rect 42360 55270 42420 55300
rect 43840 55270 43900 55300
rect 37720 55230 37750 55260
rect 37840 55230 37870 55260
rect 146100 55230 146160 55260
rect 147580 55230 147640 55260
rect 148400 55230 148460 55260
rect 149082 55236 149162 55246
rect 149242 55236 149322 55246
rect 37600 55200 37660 55230
rect 37720 55200 37780 55230
rect 37840 55200 37900 55230
rect 40060 55150 40120 55180
rect 41540 55150 41600 55180
rect 42360 55150 42420 55180
rect 43840 55150 43900 55180
rect 149162 55166 149172 55236
rect 149082 55156 149172 55166
rect 149242 55166 149252 55236
rect 149322 55166 149332 55236
rect 149880 55230 149940 55260
rect 153060 55250 153070 55330
rect 153240 55250 153250 55330
rect 153420 55250 153430 55330
rect 153600 55250 153610 55330
rect 153780 55250 153790 55330
rect 153960 55250 153970 55330
rect 154140 55250 154150 55330
rect 154320 55250 154330 55330
rect 154500 55250 154510 55330
rect 154680 55250 154690 55330
rect 154860 55250 154870 55330
rect 155040 55250 155050 55330
rect 155220 55250 155230 55330
rect 155400 55250 155410 55330
rect 155580 55250 155590 55330
rect 155760 55250 155770 55330
rect 155940 55250 155950 55330
rect 156120 55250 156130 55330
rect 156300 55250 156310 55330
rect 156480 55250 156490 55330
rect 156660 55250 156670 55330
rect 156840 55250 156850 55330
rect 157020 55250 157030 55330
rect 157200 55250 157210 55330
rect 157380 55250 157390 55330
rect 157560 55250 157570 55330
rect 157740 55250 157750 55330
rect 157920 55250 157930 55330
rect 158100 55250 158110 55330
rect 158280 55250 158290 55330
rect 158460 55250 158470 55330
rect 158640 55250 158650 55330
rect 158820 55250 158830 55330
rect 152220 55210 152250 55240
rect 152340 55210 152370 55240
rect 152100 55180 152160 55210
rect 152220 55180 152280 55210
rect 152340 55180 152400 55210
rect 149242 55156 149332 55166
rect 37720 55110 37750 55140
rect 37840 55110 37870 55140
rect 146100 55110 146160 55140
rect 147580 55110 147640 55140
rect 148400 55110 148460 55140
rect 149880 55110 149940 55140
rect 37600 55080 37660 55110
rect 37720 55080 37780 55110
rect 37840 55080 37900 55110
rect 152220 55090 152250 55120
rect 152340 55090 152370 55120
rect 149082 55076 149162 55086
rect 149242 55076 149322 55086
rect 40060 55030 40120 55060
rect 41540 55030 41600 55060
rect 42360 55030 42420 55060
rect 43840 55030 43900 55060
rect 37720 54990 37750 55020
rect 37840 54990 37870 55020
rect 146100 54990 146160 55020
rect 147580 54990 147640 55020
rect 148400 54990 148460 55020
rect 149162 54996 149172 55076
rect 149242 54996 149252 55076
rect 149322 54996 149332 55076
rect 152100 55060 152160 55090
rect 152220 55060 152280 55090
rect 152340 55060 152400 55090
rect 149880 54990 149940 55020
rect 152980 55010 153060 55020
rect 153160 55010 153240 55020
rect 153340 55010 153420 55020
rect 153520 55010 153600 55020
rect 153700 55010 153780 55020
rect 153880 55010 153960 55020
rect 154060 55010 154140 55020
rect 154240 55010 154320 55020
rect 154420 55010 154500 55020
rect 154600 55010 154680 55020
rect 154780 55010 154860 55020
rect 154960 55010 155040 55020
rect 155140 55010 155220 55020
rect 155320 55010 155400 55020
rect 155500 55010 155580 55020
rect 155680 55010 155760 55020
rect 155860 55010 155940 55020
rect 156040 55010 156120 55020
rect 156220 55010 156300 55020
rect 156400 55010 156480 55020
rect 156580 55010 156660 55020
rect 156760 55010 156840 55020
rect 156940 55010 157020 55020
rect 157120 55010 157200 55020
rect 157300 55010 157380 55020
rect 157480 55010 157560 55020
rect 157660 55010 157740 55020
rect 157840 55010 157920 55020
rect 158020 55010 158100 55020
rect 158200 55010 158280 55020
rect 158380 55010 158460 55020
rect 158560 55010 158640 55020
rect 158740 55010 158820 55020
rect 37600 54960 37660 54990
rect 37720 54960 37780 54990
rect 37840 54960 37900 54990
rect 152220 54970 152250 55000
rect 152340 54970 152370 55000
rect 152100 54940 152160 54970
rect 152220 54940 152280 54970
rect 152340 54940 152400 54970
rect 40060 54910 40120 54940
rect 41540 54910 41600 54940
rect 42360 54910 42420 54940
rect 43840 54910 43900 54940
rect 153060 54930 153070 55010
rect 153240 54930 153250 55010
rect 153420 54930 153430 55010
rect 153600 54930 153610 55010
rect 153780 54930 153790 55010
rect 153960 54930 153970 55010
rect 154140 54930 154150 55010
rect 154320 54930 154330 55010
rect 154500 54930 154510 55010
rect 154680 54930 154690 55010
rect 154860 54930 154870 55010
rect 155040 54930 155050 55010
rect 155220 54930 155230 55010
rect 155400 54930 155410 55010
rect 155580 54930 155590 55010
rect 155760 54930 155770 55010
rect 155940 54930 155950 55010
rect 156120 54930 156130 55010
rect 156300 54930 156310 55010
rect 156480 54930 156490 55010
rect 156660 54930 156670 55010
rect 156840 54930 156850 55010
rect 157020 54930 157030 55010
rect 157200 54930 157210 55010
rect 157380 54930 157390 55010
rect 157560 54930 157570 55010
rect 157740 54930 157750 55010
rect 157920 54930 157930 55010
rect 158100 54930 158110 55010
rect 158280 54930 158290 55010
rect 158460 54930 158470 55010
rect 158640 54930 158650 55010
rect 158820 54930 158830 55010
rect 37720 54870 37750 54900
rect 37840 54870 37870 54900
rect 146100 54870 146160 54900
rect 147580 54870 147640 54900
rect 148400 54870 148460 54900
rect 149880 54870 149940 54900
rect 37600 54840 37660 54870
rect 37720 54840 37780 54870
rect 37840 54840 37900 54870
rect 152220 54850 152250 54880
rect 152340 54850 152370 54880
rect 19800 54830 25800 54840
rect 31100 54830 37190 54840
rect 19130 54750 19160 54780
rect 19250 54750 19280 54780
rect 26420 54750 26450 54780
rect 26540 54750 26570 54780
rect 30420 54750 30450 54780
rect 30540 54750 30570 54780
rect 19010 54720 19070 54750
rect 19130 54720 19190 54750
rect 19250 54720 19310 54750
rect 26300 54720 26360 54750
rect 26420 54720 26480 54750
rect 26540 54720 26600 54750
rect 30300 54720 30360 54750
rect 30420 54720 30480 54750
rect 30540 54720 30600 54750
rect 37100 54730 37190 54830
rect 152100 54820 152160 54850
rect 152220 54820 152280 54850
rect 152340 54820 152400 54850
rect 158900 54840 158990 55510
rect 159520 55450 159550 55480
rect 159640 55450 159670 55480
rect 163520 55450 163550 55480
rect 163640 55450 163670 55480
rect 170810 55450 170840 55480
rect 170930 55450 170960 55480
rect 159400 55420 159460 55450
rect 159520 55420 159580 55450
rect 159640 55420 159700 55450
rect 163400 55420 163460 55450
rect 163520 55420 163580 55450
rect 163640 55420 163700 55450
rect 170690 55420 170750 55450
rect 170810 55420 170870 55450
rect 170930 55420 170990 55450
rect 159520 55330 159550 55360
rect 159640 55330 159670 55360
rect 163520 55330 163550 55360
rect 163640 55330 163670 55360
rect 164280 55330 164360 55340
rect 164460 55330 164540 55340
rect 164640 55330 164720 55340
rect 164820 55330 164900 55340
rect 165000 55330 165080 55340
rect 165180 55330 165260 55340
rect 165360 55330 165440 55340
rect 165540 55330 165620 55340
rect 165720 55330 165800 55340
rect 165900 55330 165980 55340
rect 166080 55330 166160 55340
rect 166260 55330 166340 55340
rect 166440 55330 166520 55340
rect 166620 55330 166700 55340
rect 166800 55330 166880 55340
rect 166980 55330 167060 55340
rect 167160 55330 167240 55340
rect 167340 55330 167420 55340
rect 167520 55330 167600 55340
rect 167700 55330 167780 55340
rect 167880 55330 167960 55340
rect 168060 55330 168140 55340
rect 168240 55330 168320 55340
rect 168420 55330 168500 55340
rect 168600 55330 168680 55340
rect 168780 55330 168860 55340
rect 168960 55330 169040 55340
rect 169140 55330 169220 55340
rect 169320 55330 169400 55340
rect 169500 55330 169580 55340
rect 169680 55330 169760 55340
rect 169860 55330 169940 55340
rect 170040 55330 170120 55340
rect 170810 55330 170840 55360
rect 170930 55330 170960 55360
rect 159400 55300 159460 55330
rect 159520 55300 159580 55330
rect 159640 55300 159700 55330
rect 163400 55300 163460 55330
rect 163520 55300 163580 55330
rect 163640 55300 163700 55330
rect 164360 55250 164370 55330
rect 164540 55250 164550 55330
rect 164720 55250 164730 55330
rect 164900 55250 164910 55330
rect 165080 55250 165090 55330
rect 165260 55250 165270 55330
rect 165440 55250 165450 55330
rect 165620 55250 165630 55330
rect 165800 55250 165810 55330
rect 165980 55250 165990 55330
rect 166160 55250 166170 55330
rect 166340 55250 166350 55330
rect 166520 55250 166530 55330
rect 166700 55250 166710 55330
rect 166880 55250 166890 55330
rect 167060 55250 167070 55330
rect 167240 55250 167250 55330
rect 167420 55250 167430 55330
rect 167600 55250 167610 55330
rect 167780 55250 167790 55330
rect 167960 55250 167970 55330
rect 168140 55250 168150 55330
rect 168320 55250 168330 55330
rect 168500 55250 168510 55330
rect 168680 55250 168690 55330
rect 168860 55250 168870 55330
rect 169040 55250 169050 55330
rect 169220 55250 169230 55330
rect 169400 55250 169410 55330
rect 169580 55250 169590 55330
rect 169760 55250 169770 55330
rect 169940 55250 169950 55330
rect 170120 55250 170130 55330
rect 170690 55300 170750 55330
rect 170810 55300 170870 55330
rect 170930 55300 170990 55330
rect 159520 55210 159550 55240
rect 159640 55210 159670 55240
rect 163520 55210 163550 55240
rect 163640 55210 163670 55240
rect 170810 55210 170840 55240
rect 170930 55210 170960 55240
rect 159400 55180 159460 55210
rect 159520 55180 159580 55210
rect 159640 55180 159700 55210
rect 163400 55180 163460 55210
rect 163520 55180 163580 55210
rect 163640 55180 163700 55210
rect 170690 55180 170750 55210
rect 170810 55180 170870 55210
rect 170930 55180 170990 55210
rect 159520 55090 159550 55120
rect 159640 55090 159670 55120
rect 163520 55090 163550 55120
rect 163640 55090 163670 55120
rect 170810 55090 170840 55120
rect 170930 55090 170960 55120
rect 159400 55060 159460 55090
rect 159520 55060 159580 55090
rect 159640 55060 159700 55090
rect 163400 55060 163460 55090
rect 163520 55060 163580 55090
rect 163640 55060 163700 55090
rect 170690 55060 170750 55090
rect 170810 55060 170870 55090
rect 170930 55060 170990 55090
rect 164280 55030 164360 55040
rect 164460 55030 164540 55040
rect 164640 55030 164720 55040
rect 164820 55030 164900 55040
rect 165000 55030 165080 55040
rect 165180 55030 165260 55040
rect 165360 55030 165440 55040
rect 165540 55030 165620 55040
rect 165720 55030 165800 55040
rect 165900 55030 165980 55040
rect 166080 55030 166160 55040
rect 166260 55030 166340 55040
rect 166440 55030 166520 55040
rect 166620 55030 166700 55040
rect 166800 55030 166880 55040
rect 166980 55030 167060 55040
rect 167160 55030 167240 55040
rect 167340 55030 167420 55040
rect 167520 55030 167600 55040
rect 167700 55030 167780 55040
rect 167880 55030 167960 55040
rect 168060 55030 168140 55040
rect 168240 55030 168320 55040
rect 168420 55030 168500 55040
rect 168600 55030 168680 55040
rect 168780 55030 168860 55040
rect 168960 55030 169040 55040
rect 169140 55030 169220 55040
rect 169320 55030 169400 55040
rect 169500 55030 169580 55040
rect 169680 55030 169760 55040
rect 169860 55030 169940 55040
rect 170040 55030 170120 55040
rect 159520 54970 159550 55000
rect 159640 54970 159670 55000
rect 163520 54970 163550 55000
rect 163640 54970 163670 55000
rect 159400 54940 159460 54970
rect 159520 54940 159580 54970
rect 159640 54940 159700 54970
rect 163400 54940 163460 54970
rect 163520 54940 163580 54970
rect 163640 54940 163700 54970
rect 164360 54950 164370 55030
rect 164540 54950 164550 55030
rect 164720 54950 164730 55030
rect 164900 54950 164910 55030
rect 165080 54950 165090 55030
rect 165260 54950 165270 55030
rect 165440 54950 165450 55030
rect 165620 54950 165630 55030
rect 165800 54950 165810 55030
rect 165980 54950 165990 55030
rect 166160 54950 166170 55030
rect 166340 54950 166350 55030
rect 166520 54950 166530 55030
rect 166700 54950 166710 55030
rect 166880 54950 166890 55030
rect 167060 54950 167070 55030
rect 167240 54950 167250 55030
rect 167420 54950 167430 55030
rect 167600 54950 167610 55030
rect 167780 54950 167790 55030
rect 167960 54950 167970 55030
rect 168140 54950 168150 55030
rect 168320 54950 168330 55030
rect 168500 54950 168510 55030
rect 168680 54950 168690 55030
rect 168860 54950 168870 55030
rect 169040 54950 169050 55030
rect 169220 54950 169230 55030
rect 169400 54950 169410 55030
rect 169580 54950 169590 55030
rect 169760 54950 169770 55030
rect 169940 54950 169950 55030
rect 170120 54950 170130 55030
rect 170810 54970 170840 55000
rect 170930 54970 170960 55000
rect 170690 54940 170750 54970
rect 170810 54940 170870 54970
rect 170930 54940 170990 54970
rect 159520 54850 159550 54880
rect 159640 54850 159670 54880
rect 163520 54850 163550 54880
rect 163640 54850 163670 54880
rect 170810 54850 170840 54880
rect 170930 54850 170960 54880
rect 152900 54830 158990 54840
rect 40060 54790 40120 54820
rect 41540 54790 41600 54820
rect 42360 54790 42420 54820
rect 43840 54790 43900 54820
rect 37720 54750 37750 54780
rect 37840 54750 37870 54780
rect 146100 54750 146160 54780
rect 147580 54750 147640 54780
rect 148400 54750 148460 54780
rect 149880 54750 149940 54780
rect 31100 54700 37190 54730
rect 37600 54720 37660 54750
rect 37720 54720 37780 54750
rect 37840 54720 37900 54750
rect 40685 54710 40925 54740
rect 152220 54730 152250 54760
rect 152340 54730 152370 54760
rect 158900 54730 158990 54830
rect 159400 54820 159460 54850
rect 159520 54820 159580 54850
rect 159640 54820 159700 54850
rect 163400 54820 163460 54850
rect 163520 54820 163580 54850
rect 163640 54820 163700 54850
rect 164200 54830 170200 54840
rect 170690 54820 170750 54850
rect 170810 54820 170870 54850
rect 170930 54820 170990 54850
rect 159520 54730 159550 54760
rect 159640 54730 159670 54760
rect 163520 54730 163550 54760
rect 163640 54730 163670 54760
rect 170810 54730 170840 54760
rect 170930 54730 170960 54760
rect 19880 54690 19960 54700
rect 20060 54690 20140 54700
rect 20240 54690 20320 54700
rect 20420 54690 20500 54700
rect 20600 54690 20680 54700
rect 20780 54690 20860 54700
rect 20960 54690 21040 54700
rect 21140 54690 21220 54700
rect 21320 54690 21400 54700
rect 21500 54690 21580 54700
rect 21680 54690 21760 54700
rect 21860 54690 21940 54700
rect 22040 54690 22120 54700
rect 22220 54690 22300 54700
rect 22400 54690 22480 54700
rect 22580 54690 22660 54700
rect 22760 54690 22840 54700
rect 22940 54690 23020 54700
rect 23120 54690 23200 54700
rect 23300 54690 23380 54700
rect 23480 54690 23560 54700
rect 23660 54690 23740 54700
rect 23840 54690 23920 54700
rect 24020 54690 24100 54700
rect 24200 54690 24280 54700
rect 24380 54690 24460 54700
rect 24560 54690 24640 54700
rect 24740 54690 24820 54700
rect 24920 54690 25000 54700
rect 25100 54690 25180 54700
rect 25280 54690 25360 54700
rect 25460 54690 25540 54700
rect 25640 54690 25720 54700
rect 31180 54690 31260 54700
rect 31360 54690 31440 54700
rect 31540 54690 31620 54700
rect 31720 54690 31800 54700
rect 31900 54690 31980 54700
rect 32080 54690 32160 54700
rect 32260 54690 32340 54700
rect 32440 54690 32520 54700
rect 32620 54690 32700 54700
rect 32800 54690 32880 54700
rect 32980 54690 33060 54700
rect 33160 54690 33240 54700
rect 33340 54690 33420 54700
rect 33520 54690 33600 54700
rect 33700 54690 33780 54700
rect 33880 54690 33960 54700
rect 34060 54690 34140 54700
rect 34240 54690 34320 54700
rect 34420 54690 34500 54700
rect 34600 54690 34680 54700
rect 34780 54690 34860 54700
rect 34960 54690 35040 54700
rect 35140 54690 35220 54700
rect 35320 54690 35400 54700
rect 35500 54690 35580 54700
rect 35680 54690 35760 54700
rect 35860 54690 35940 54700
rect 36040 54690 36120 54700
rect 36220 54690 36300 54700
rect 36400 54690 36480 54700
rect 36580 54690 36660 54700
rect 36760 54690 36840 54700
rect 36940 54690 37020 54700
rect 19130 54630 19160 54660
rect 19250 54630 19280 54660
rect 19010 54600 19070 54630
rect 19130 54600 19190 54630
rect 19250 54600 19310 54630
rect 19960 54610 19970 54690
rect 20140 54610 20150 54690
rect 20320 54610 20330 54690
rect 20500 54610 20510 54690
rect 20680 54610 20690 54690
rect 20860 54610 20870 54690
rect 21040 54610 21050 54690
rect 21220 54610 21230 54690
rect 21400 54610 21410 54690
rect 21580 54610 21590 54690
rect 21760 54610 21770 54690
rect 21940 54610 21950 54690
rect 22120 54610 22130 54690
rect 22300 54610 22310 54690
rect 22480 54610 22490 54690
rect 22660 54610 22670 54690
rect 22840 54610 22850 54690
rect 23020 54610 23030 54690
rect 23200 54610 23210 54690
rect 23380 54610 23390 54690
rect 23560 54610 23570 54690
rect 23740 54610 23750 54690
rect 23920 54610 23930 54690
rect 24100 54610 24110 54690
rect 24280 54610 24290 54690
rect 24460 54610 24470 54690
rect 24640 54610 24650 54690
rect 24820 54610 24830 54690
rect 25000 54610 25010 54690
rect 25180 54610 25190 54690
rect 25360 54610 25370 54690
rect 25540 54610 25550 54690
rect 25720 54610 25730 54690
rect 26420 54630 26450 54660
rect 26540 54630 26570 54660
rect 30420 54630 30450 54660
rect 30540 54630 30570 54660
rect 31260 54630 31270 54690
rect 31440 54630 31450 54690
rect 31620 54630 31630 54690
rect 31800 54630 31810 54690
rect 31980 54630 31990 54690
rect 32160 54630 32170 54690
rect 32340 54630 32350 54690
rect 32520 54630 32530 54690
rect 32700 54630 32710 54690
rect 32880 54630 32890 54690
rect 33060 54630 33070 54690
rect 33240 54630 33250 54690
rect 33420 54630 33430 54690
rect 33600 54630 33610 54690
rect 33780 54630 33790 54690
rect 33960 54630 33970 54690
rect 34140 54630 34150 54690
rect 34320 54630 34330 54690
rect 34500 54630 34510 54690
rect 34680 54630 34690 54690
rect 34860 54630 34870 54690
rect 35040 54630 35050 54690
rect 35220 54630 35230 54690
rect 35400 54630 35410 54690
rect 35580 54630 35590 54690
rect 35760 54630 35770 54690
rect 35940 54630 35950 54690
rect 36120 54630 36130 54690
rect 36300 54630 36310 54690
rect 36480 54630 36490 54690
rect 36660 54630 36670 54690
rect 36840 54630 36850 54690
rect 37020 54630 37030 54690
rect 37100 54630 37190 54700
rect 40060 54670 40120 54700
rect 37720 54630 37750 54660
rect 37840 54630 37870 54660
rect 40685 54650 40715 54710
rect 40775 54650 40865 54710
rect 40895 54650 40925 54710
rect 152100 54700 152160 54730
rect 152220 54700 152280 54730
rect 152340 54700 152400 54730
rect 152900 54700 158990 54730
rect 159400 54700 159460 54730
rect 159520 54700 159580 54730
rect 159640 54700 159700 54730
rect 163400 54700 163460 54730
rect 163520 54700 163580 54730
rect 163640 54700 163700 54730
rect 170690 54700 170750 54730
rect 170810 54700 170870 54730
rect 170930 54700 170990 54730
rect 41540 54670 41600 54700
rect 42360 54670 42420 54700
rect 43840 54670 43900 54700
rect 152980 54690 153060 54700
rect 153160 54690 153240 54700
rect 153340 54690 153420 54700
rect 153520 54690 153600 54700
rect 153700 54690 153780 54700
rect 153880 54690 153960 54700
rect 154060 54690 154140 54700
rect 154240 54690 154320 54700
rect 154420 54690 154500 54700
rect 154600 54690 154680 54700
rect 154780 54690 154860 54700
rect 154960 54690 155040 54700
rect 155140 54690 155220 54700
rect 155320 54690 155400 54700
rect 155500 54690 155580 54700
rect 155680 54690 155760 54700
rect 155860 54690 155940 54700
rect 156040 54690 156120 54700
rect 156220 54690 156300 54700
rect 156400 54690 156480 54700
rect 156580 54690 156660 54700
rect 156760 54690 156840 54700
rect 156940 54690 157020 54700
rect 157120 54690 157200 54700
rect 157300 54690 157380 54700
rect 157480 54690 157560 54700
rect 157660 54690 157740 54700
rect 157840 54690 157920 54700
rect 158020 54690 158100 54700
rect 158200 54690 158280 54700
rect 158380 54690 158460 54700
rect 158560 54690 158640 54700
rect 158740 54690 158820 54700
rect 26300 54600 26360 54630
rect 26420 54600 26480 54630
rect 26540 54600 26600 54630
rect 30300 54600 30360 54630
rect 30420 54600 30480 54630
rect 30540 54600 30600 54630
rect 31100 54600 37190 54630
rect 37600 54600 37660 54630
rect 37720 54600 37780 54630
rect 37840 54600 37900 54630
rect 40685 54620 40925 54650
rect 19880 54540 19960 54550
rect 20060 54540 20140 54550
rect 20240 54540 20320 54550
rect 20420 54540 20500 54550
rect 20600 54540 20680 54550
rect 20780 54540 20860 54550
rect 20960 54540 21040 54550
rect 21140 54540 21220 54550
rect 21320 54540 21400 54550
rect 21500 54540 21580 54550
rect 21680 54540 21760 54550
rect 21860 54540 21940 54550
rect 22040 54540 22120 54550
rect 22220 54540 22300 54550
rect 22400 54540 22480 54550
rect 22580 54540 22660 54550
rect 22760 54540 22840 54550
rect 22940 54540 23020 54550
rect 23120 54540 23200 54550
rect 23300 54540 23380 54550
rect 23480 54540 23560 54550
rect 23660 54540 23740 54550
rect 23840 54540 23920 54550
rect 24020 54540 24100 54550
rect 24200 54540 24280 54550
rect 24380 54540 24460 54550
rect 24560 54540 24640 54550
rect 24740 54540 24820 54550
rect 24920 54540 25000 54550
rect 25100 54540 25180 54550
rect 25280 54540 25360 54550
rect 25460 54540 25540 54550
rect 25640 54540 25720 54550
rect 31180 54540 31260 54550
rect 31360 54540 31440 54550
rect 31540 54540 31620 54550
rect 31720 54540 31800 54550
rect 31900 54540 31980 54550
rect 32080 54540 32160 54550
rect 32260 54540 32340 54550
rect 32440 54540 32520 54550
rect 32620 54540 32700 54550
rect 32800 54540 32880 54550
rect 32980 54540 33060 54550
rect 33160 54540 33240 54550
rect 33340 54540 33420 54550
rect 33520 54540 33600 54550
rect 33700 54540 33780 54550
rect 33880 54540 33960 54550
rect 34060 54540 34140 54550
rect 34240 54540 34320 54550
rect 34420 54540 34500 54550
rect 34600 54540 34680 54550
rect 34780 54540 34860 54550
rect 34960 54540 35040 54550
rect 35140 54540 35220 54550
rect 35320 54540 35400 54550
rect 35500 54540 35580 54550
rect 35680 54540 35760 54550
rect 35860 54540 35940 54550
rect 36040 54540 36120 54550
rect 36220 54540 36300 54550
rect 36400 54540 36480 54550
rect 36580 54540 36660 54550
rect 36760 54540 36840 54550
rect 36940 54540 37020 54550
rect 19130 54510 19160 54540
rect 19250 54510 19280 54540
rect 19010 54480 19070 54510
rect 19130 54480 19190 54510
rect 19250 54480 19310 54510
rect 19960 54460 19970 54540
rect 20140 54460 20150 54540
rect 20320 54460 20330 54540
rect 20500 54460 20510 54540
rect 20680 54460 20690 54540
rect 20860 54460 20870 54540
rect 21040 54460 21050 54540
rect 21220 54460 21230 54540
rect 21400 54460 21410 54540
rect 21580 54460 21590 54540
rect 21760 54460 21770 54540
rect 21940 54460 21950 54540
rect 22120 54460 22130 54540
rect 22300 54460 22310 54540
rect 22480 54460 22490 54540
rect 22660 54460 22670 54540
rect 22840 54460 22850 54540
rect 23020 54460 23030 54540
rect 23200 54460 23210 54540
rect 23380 54460 23390 54540
rect 23560 54460 23570 54540
rect 23740 54460 23750 54540
rect 23920 54460 23930 54540
rect 24100 54460 24110 54540
rect 24280 54460 24290 54540
rect 24460 54460 24470 54540
rect 24640 54460 24650 54540
rect 24820 54460 24830 54540
rect 25000 54460 25010 54540
rect 25180 54460 25190 54540
rect 25360 54460 25370 54540
rect 25540 54460 25550 54540
rect 25720 54460 25730 54540
rect 26420 54510 26450 54540
rect 26540 54510 26570 54540
rect 30420 54510 30450 54540
rect 30540 54510 30570 54540
rect 26300 54480 26360 54510
rect 26420 54480 26480 54510
rect 26540 54480 26600 54510
rect 30300 54480 30360 54510
rect 30420 54480 30480 54510
rect 30540 54480 30600 54510
rect 31260 54460 31270 54540
rect 31440 54460 31450 54540
rect 31620 54460 31630 54540
rect 31800 54460 31810 54540
rect 31980 54460 31990 54540
rect 32160 54460 32170 54540
rect 32340 54460 32350 54540
rect 32520 54460 32530 54540
rect 32700 54460 32710 54540
rect 32880 54460 32890 54540
rect 33060 54460 33070 54540
rect 33240 54460 33250 54540
rect 33420 54460 33430 54540
rect 33600 54460 33610 54540
rect 33780 54460 33790 54540
rect 33960 54460 33970 54540
rect 34140 54460 34150 54540
rect 34320 54460 34330 54540
rect 34500 54460 34510 54540
rect 34680 54460 34690 54540
rect 34860 54460 34870 54540
rect 35040 54460 35050 54540
rect 35220 54460 35230 54540
rect 35400 54460 35410 54540
rect 35580 54460 35590 54540
rect 35760 54460 35770 54540
rect 35940 54460 35950 54540
rect 36120 54460 36130 54540
rect 36300 54460 36310 54540
rect 36480 54460 36490 54540
rect 36660 54460 36670 54540
rect 36840 54460 36850 54540
rect 37020 54460 37030 54540
rect 19130 54390 19160 54420
rect 19250 54390 19280 54420
rect 19880 54390 19960 54400
rect 20060 54390 20140 54400
rect 20240 54390 20320 54400
rect 20420 54390 20500 54400
rect 20600 54390 20680 54400
rect 20780 54390 20860 54400
rect 20960 54390 21040 54400
rect 21140 54390 21220 54400
rect 21320 54390 21400 54400
rect 21500 54390 21580 54400
rect 21680 54390 21760 54400
rect 21860 54390 21940 54400
rect 22040 54390 22120 54400
rect 22220 54390 22300 54400
rect 22400 54390 22480 54400
rect 22580 54390 22660 54400
rect 22760 54390 22840 54400
rect 22940 54390 23020 54400
rect 23120 54390 23200 54400
rect 23300 54390 23380 54400
rect 23480 54390 23560 54400
rect 23660 54390 23740 54400
rect 23840 54390 23920 54400
rect 24020 54390 24100 54400
rect 24200 54390 24280 54400
rect 24380 54390 24460 54400
rect 24560 54390 24640 54400
rect 24740 54390 24820 54400
rect 24920 54390 25000 54400
rect 25100 54390 25180 54400
rect 25280 54390 25360 54400
rect 25460 54390 25540 54400
rect 25640 54390 25720 54400
rect 26420 54390 26450 54420
rect 26540 54390 26570 54420
rect 30420 54390 30450 54420
rect 30540 54390 30570 54420
rect 37100 54400 37190 54600
rect 40060 54550 40120 54580
rect 41540 54550 41600 54580
rect 42360 54550 42420 54580
rect 43840 54550 43900 54580
rect 37720 54510 37750 54540
rect 37840 54510 37870 54540
rect 37600 54480 37660 54510
rect 37720 54480 37780 54510
rect 37840 54480 37900 54510
rect 146100 54630 146160 54660
rect 147580 54630 147640 54660
rect 148400 54630 148460 54660
rect 149880 54630 149940 54660
rect 152220 54610 152250 54640
rect 152340 54610 152370 54640
rect 153060 54630 153070 54690
rect 153240 54630 153250 54690
rect 153420 54630 153430 54690
rect 153600 54630 153610 54690
rect 153780 54630 153790 54690
rect 153960 54630 153970 54690
rect 154140 54630 154150 54690
rect 154320 54630 154330 54690
rect 154500 54630 154510 54690
rect 154680 54630 154690 54690
rect 154860 54630 154870 54690
rect 155040 54630 155050 54690
rect 155220 54630 155230 54690
rect 155400 54630 155410 54690
rect 155580 54630 155590 54690
rect 155760 54630 155770 54690
rect 155940 54630 155950 54690
rect 156120 54630 156130 54690
rect 156300 54630 156310 54690
rect 156480 54630 156490 54690
rect 156660 54630 156670 54690
rect 156840 54630 156850 54690
rect 157020 54630 157030 54690
rect 157200 54630 157210 54690
rect 157380 54630 157390 54690
rect 157560 54630 157570 54690
rect 157740 54630 157750 54690
rect 157920 54630 157930 54690
rect 158100 54630 158110 54690
rect 158280 54630 158290 54690
rect 158460 54630 158470 54690
rect 158640 54630 158650 54690
rect 158820 54630 158830 54690
rect 158900 54630 158990 54700
rect 164280 54690 164360 54700
rect 164460 54690 164540 54700
rect 164640 54690 164720 54700
rect 164820 54690 164900 54700
rect 165000 54690 165080 54700
rect 165180 54690 165260 54700
rect 165360 54690 165440 54700
rect 165540 54690 165620 54700
rect 165720 54690 165800 54700
rect 165900 54690 165980 54700
rect 166080 54690 166160 54700
rect 166260 54690 166340 54700
rect 166440 54690 166520 54700
rect 166620 54690 166700 54700
rect 166800 54690 166880 54700
rect 166980 54690 167060 54700
rect 167160 54690 167240 54700
rect 167340 54690 167420 54700
rect 167520 54690 167600 54700
rect 167700 54690 167780 54700
rect 167880 54690 167960 54700
rect 168060 54690 168140 54700
rect 168240 54690 168320 54700
rect 168420 54690 168500 54700
rect 168600 54690 168680 54700
rect 168780 54690 168860 54700
rect 168960 54690 169040 54700
rect 169140 54690 169220 54700
rect 169320 54690 169400 54700
rect 169500 54690 169580 54700
rect 169680 54690 169760 54700
rect 169860 54690 169940 54700
rect 170040 54690 170120 54700
rect 152100 54580 152160 54610
rect 152220 54580 152280 54610
rect 152340 54580 152400 54610
rect 152900 54600 158990 54630
rect 159520 54610 159550 54640
rect 159640 54610 159670 54640
rect 163520 54610 163550 54640
rect 163640 54610 163670 54640
rect 164360 54610 164370 54690
rect 164540 54610 164550 54690
rect 164720 54610 164730 54690
rect 164900 54610 164910 54690
rect 165080 54610 165090 54690
rect 165260 54610 165270 54690
rect 165440 54610 165450 54690
rect 165620 54610 165630 54690
rect 165800 54610 165810 54690
rect 165980 54610 165990 54690
rect 166160 54610 166170 54690
rect 166340 54610 166350 54690
rect 166520 54610 166530 54690
rect 166700 54610 166710 54690
rect 166880 54610 166890 54690
rect 167060 54610 167070 54690
rect 167240 54610 167250 54690
rect 167420 54610 167430 54690
rect 167600 54610 167610 54690
rect 167780 54610 167790 54690
rect 167960 54610 167970 54690
rect 168140 54610 168150 54690
rect 168320 54610 168330 54690
rect 168500 54610 168510 54690
rect 168680 54610 168690 54690
rect 168860 54610 168870 54690
rect 169040 54610 169050 54690
rect 169220 54610 169230 54690
rect 169400 54610 169410 54690
rect 169580 54610 169590 54690
rect 169760 54610 169770 54690
rect 169940 54610 169950 54690
rect 170120 54610 170130 54690
rect 170810 54610 170840 54640
rect 170930 54610 170960 54640
rect 152980 54540 153060 54550
rect 153160 54540 153240 54550
rect 153340 54540 153420 54550
rect 153520 54540 153600 54550
rect 153700 54540 153780 54550
rect 153880 54540 153960 54550
rect 154060 54540 154140 54550
rect 154240 54540 154320 54550
rect 154420 54540 154500 54550
rect 154600 54540 154680 54550
rect 154780 54540 154860 54550
rect 154960 54540 155040 54550
rect 155140 54540 155220 54550
rect 155320 54540 155400 54550
rect 155500 54540 155580 54550
rect 155680 54540 155760 54550
rect 155860 54540 155940 54550
rect 156040 54540 156120 54550
rect 156220 54540 156300 54550
rect 156400 54540 156480 54550
rect 156580 54540 156660 54550
rect 156760 54540 156840 54550
rect 156940 54540 157020 54550
rect 157120 54540 157200 54550
rect 157300 54540 157380 54550
rect 157480 54540 157560 54550
rect 157660 54540 157740 54550
rect 157840 54540 157920 54550
rect 158020 54540 158100 54550
rect 158200 54540 158280 54550
rect 158380 54540 158460 54550
rect 158560 54540 158640 54550
rect 158740 54540 158820 54550
rect 146100 54510 146160 54540
rect 147580 54510 147640 54540
rect 148400 54510 148460 54540
rect 149880 54510 149940 54540
rect 152220 54490 152250 54520
rect 152340 54490 152370 54520
rect 152100 54460 152160 54490
rect 152220 54460 152280 54490
rect 152340 54460 152400 54490
rect 153060 54460 153070 54540
rect 153240 54460 153250 54540
rect 153420 54460 153430 54540
rect 153600 54460 153610 54540
rect 153780 54460 153790 54540
rect 153960 54460 153970 54540
rect 154140 54460 154150 54540
rect 154320 54460 154330 54540
rect 154500 54460 154510 54540
rect 154680 54460 154690 54540
rect 154860 54460 154870 54540
rect 155040 54460 155050 54540
rect 155220 54460 155230 54540
rect 155400 54460 155410 54540
rect 155580 54460 155590 54540
rect 155760 54460 155770 54540
rect 155940 54460 155950 54540
rect 156120 54460 156130 54540
rect 156300 54460 156310 54540
rect 156480 54460 156490 54540
rect 156660 54460 156670 54540
rect 156840 54460 156850 54540
rect 157020 54460 157030 54540
rect 157200 54460 157210 54540
rect 157380 54460 157390 54540
rect 157560 54460 157570 54540
rect 157740 54460 157750 54540
rect 157920 54460 157930 54540
rect 158100 54460 158110 54540
rect 158280 54460 158290 54540
rect 158460 54460 158470 54540
rect 158640 54460 158650 54540
rect 158820 54460 158830 54540
rect 40060 54430 40120 54460
rect 41540 54430 41600 54460
rect 42360 54430 42420 54460
rect 43840 54430 43900 54460
rect 19010 54360 19070 54390
rect 19130 54360 19190 54390
rect 19250 54360 19310 54390
rect 19960 54310 19970 54390
rect 20140 54310 20150 54390
rect 20320 54310 20330 54390
rect 20500 54310 20510 54390
rect 20680 54310 20690 54390
rect 20860 54310 20870 54390
rect 21040 54310 21050 54390
rect 21220 54310 21230 54390
rect 21400 54310 21410 54390
rect 21580 54310 21590 54390
rect 21760 54310 21770 54390
rect 21940 54310 21950 54390
rect 22120 54310 22130 54390
rect 22300 54310 22310 54390
rect 22480 54310 22490 54390
rect 22660 54310 22670 54390
rect 22840 54310 22850 54390
rect 23020 54310 23030 54390
rect 23200 54310 23210 54390
rect 23380 54310 23390 54390
rect 23560 54310 23570 54390
rect 23740 54310 23750 54390
rect 23920 54310 23930 54390
rect 24100 54310 24110 54390
rect 24280 54310 24290 54390
rect 24460 54310 24470 54390
rect 24640 54310 24650 54390
rect 24820 54310 24830 54390
rect 25000 54310 25010 54390
rect 25180 54310 25190 54390
rect 25360 54310 25370 54390
rect 25540 54310 25550 54390
rect 25720 54310 25730 54390
rect 26300 54360 26360 54390
rect 26420 54360 26480 54390
rect 26540 54360 26600 54390
rect 30300 54360 30360 54390
rect 30420 54360 30480 54390
rect 30540 54360 30600 54390
rect 31100 54370 37190 54400
rect 37720 54390 37750 54420
rect 37840 54390 37870 54420
rect 146100 54390 146160 54420
rect 147580 54390 147640 54420
rect 148400 54390 148460 54420
rect 149880 54390 149940 54420
rect 158900 54400 158990 54600
rect 159400 54580 159460 54610
rect 159520 54580 159580 54610
rect 159640 54580 159700 54610
rect 163400 54580 163460 54610
rect 163520 54580 163580 54610
rect 163640 54580 163700 54610
rect 170690 54580 170750 54610
rect 170810 54580 170870 54610
rect 170930 54580 170990 54610
rect 164280 54540 164360 54550
rect 164460 54540 164540 54550
rect 164640 54540 164720 54550
rect 164820 54540 164900 54550
rect 165000 54540 165080 54550
rect 165180 54540 165260 54550
rect 165360 54540 165440 54550
rect 165540 54540 165620 54550
rect 165720 54540 165800 54550
rect 165900 54540 165980 54550
rect 166080 54540 166160 54550
rect 166260 54540 166340 54550
rect 166440 54540 166520 54550
rect 166620 54540 166700 54550
rect 166800 54540 166880 54550
rect 166980 54540 167060 54550
rect 167160 54540 167240 54550
rect 167340 54540 167420 54550
rect 167520 54540 167600 54550
rect 167700 54540 167780 54550
rect 167880 54540 167960 54550
rect 168060 54540 168140 54550
rect 168240 54540 168320 54550
rect 168420 54540 168500 54550
rect 168600 54540 168680 54550
rect 168780 54540 168860 54550
rect 168960 54540 169040 54550
rect 169140 54540 169220 54550
rect 169320 54540 169400 54550
rect 169500 54540 169580 54550
rect 169680 54540 169760 54550
rect 169860 54540 169940 54550
rect 170040 54540 170120 54550
rect 159520 54490 159550 54520
rect 159640 54490 159670 54520
rect 163520 54490 163550 54520
rect 163640 54490 163670 54520
rect 159400 54460 159460 54490
rect 159520 54460 159580 54490
rect 159640 54460 159700 54490
rect 163400 54460 163460 54490
rect 163520 54460 163580 54490
rect 163640 54460 163700 54490
rect 164360 54460 164370 54540
rect 164540 54460 164550 54540
rect 164720 54460 164730 54540
rect 164900 54460 164910 54540
rect 165080 54460 165090 54540
rect 165260 54460 165270 54540
rect 165440 54460 165450 54540
rect 165620 54460 165630 54540
rect 165800 54460 165810 54540
rect 165980 54460 165990 54540
rect 166160 54460 166170 54540
rect 166340 54460 166350 54540
rect 166520 54460 166530 54540
rect 166700 54460 166710 54540
rect 166880 54460 166890 54540
rect 167060 54460 167070 54540
rect 167240 54460 167250 54540
rect 167420 54460 167430 54540
rect 167600 54460 167610 54540
rect 167780 54460 167790 54540
rect 167960 54460 167970 54540
rect 168140 54460 168150 54540
rect 168320 54460 168330 54540
rect 168500 54460 168510 54540
rect 168680 54460 168690 54540
rect 168860 54460 168870 54540
rect 169040 54460 169050 54540
rect 169220 54460 169230 54540
rect 169400 54460 169410 54540
rect 169580 54460 169590 54540
rect 169760 54460 169770 54540
rect 169940 54460 169950 54540
rect 170120 54460 170130 54540
rect 170810 54490 170840 54520
rect 170930 54490 170960 54520
rect 170690 54460 170750 54490
rect 170810 54460 170870 54490
rect 170930 54460 170990 54490
rect 31260 54310 31270 54370
rect 31440 54310 31450 54370
rect 31620 54310 31630 54370
rect 31800 54310 31810 54370
rect 31980 54310 31990 54370
rect 32160 54310 32170 54370
rect 32340 54310 32350 54370
rect 32520 54310 32530 54370
rect 32700 54310 32710 54370
rect 32880 54310 32890 54370
rect 33060 54310 33070 54370
rect 33240 54310 33250 54370
rect 33420 54310 33430 54370
rect 33600 54310 33610 54370
rect 33780 54310 33790 54370
rect 33960 54310 33970 54370
rect 34140 54310 34150 54370
rect 34320 54310 34330 54370
rect 34500 54310 34510 54370
rect 34680 54310 34690 54370
rect 34860 54310 34870 54370
rect 35040 54310 35050 54370
rect 35220 54310 35230 54370
rect 35400 54310 35410 54370
rect 35580 54310 35590 54370
rect 35760 54310 35770 54370
rect 35940 54310 35950 54370
rect 36120 54310 36130 54370
rect 36300 54310 36310 54370
rect 36480 54310 36490 54370
rect 36660 54310 36670 54370
rect 36840 54310 36850 54370
rect 37020 54310 37030 54370
rect 37100 54300 37190 54370
rect 37600 54360 37660 54390
rect 37720 54360 37780 54390
rect 37840 54360 37900 54390
rect 149075 54350 149315 54380
rect 152220 54370 152250 54400
rect 152340 54370 152370 54400
rect 152900 54370 158990 54400
rect 159520 54370 159550 54400
rect 159640 54370 159670 54400
rect 163520 54370 163550 54400
rect 163640 54370 163670 54400
rect 164280 54390 164360 54400
rect 164460 54390 164540 54400
rect 164640 54390 164720 54400
rect 164820 54390 164900 54400
rect 165000 54390 165080 54400
rect 165180 54390 165260 54400
rect 165360 54390 165440 54400
rect 165540 54390 165620 54400
rect 165720 54390 165800 54400
rect 165900 54390 165980 54400
rect 166080 54390 166160 54400
rect 166260 54390 166340 54400
rect 166440 54390 166520 54400
rect 166620 54390 166700 54400
rect 166800 54390 166880 54400
rect 166980 54390 167060 54400
rect 167160 54390 167240 54400
rect 167340 54390 167420 54400
rect 167520 54390 167600 54400
rect 167700 54390 167780 54400
rect 167880 54390 167960 54400
rect 168060 54390 168140 54400
rect 168240 54390 168320 54400
rect 168420 54390 168500 54400
rect 168600 54390 168680 54400
rect 168780 54390 168860 54400
rect 168960 54390 169040 54400
rect 169140 54390 169220 54400
rect 169320 54390 169400 54400
rect 169500 54390 169580 54400
rect 169680 54390 169760 54400
rect 169860 54390 169940 54400
rect 170040 54390 170120 54400
rect 40060 54310 40120 54340
rect 41540 54310 41600 54340
rect 42360 54310 42420 54340
rect 43840 54310 43900 54340
rect 19130 54270 19160 54300
rect 19250 54270 19280 54300
rect 26420 54270 26450 54300
rect 26540 54270 26570 54300
rect 30420 54270 30450 54300
rect 30540 54270 30570 54300
rect 31100 54270 37190 54300
rect 37720 54270 37750 54300
rect 37840 54270 37870 54300
rect 146100 54270 146160 54300
rect 147580 54270 147640 54300
rect 148400 54270 148460 54300
rect 149075 54290 149105 54350
rect 149165 54290 149255 54350
rect 149285 54290 149315 54350
rect 152100 54340 152160 54370
rect 152220 54340 152280 54370
rect 152340 54340 152400 54370
rect 153060 54310 153070 54370
rect 153240 54310 153250 54370
rect 153420 54310 153430 54370
rect 153600 54310 153610 54370
rect 153780 54310 153790 54370
rect 153960 54310 153970 54370
rect 154140 54310 154150 54370
rect 154320 54310 154330 54370
rect 154500 54310 154510 54370
rect 154680 54310 154690 54370
rect 154860 54310 154870 54370
rect 155040 54310 155050 54370
rect 155220 54310 155230 54370
rect 155400 54310 155410 54370
rect 155580 54310 155590 54370
rect 155760 54310 155770 54370
rect 155940 54310 155950 54370
rect 156120 54310 156130 54370
rect 156300 54310 156310 54370
rect 156480 54310 156490 54370
rect 156660 54310 156670 54370
rect 156840 54310 156850 54370
rect 157020 54310 157030 54370
rect 157200 54310 157210 54370
rect 157380 54310 157390 54370
rect 157560 54310 157570 54370
rect 157740 54310 157750 54370
rect 157920 54310 157930 54370
rect 158100 54310 158110 54370
rect 158280 54310 158290 54370
rect 158460 54310 158470 54370
rect 158640 54310 158650 54370
rect 158820 54310 158830 54370
rect 158900 54300 158990 54370
rect 159400 54340 159460 54370
rect 159520 54340 159580 54370
rect 159640 54340 159700 54370
rect 163400 54340 163460 54370
rect 163520 54340 163580 54370
rect 163640 54340 163700 54370
rect 164360 54310 164370 54390
rect 164540 54310 164550 54390
rect 164720 54310 164730 54390
rect 164900 54310 164910 54390
rect 165080 54310 165090 54390
rect 165260 54310 165270 54390
rect 165440 54310 165450 54390
rect 165620 54310 165630 54390
rect 165800 54310 165810 54390
rect 165980 54310 165990 54390
rect 166160 54310 166170 54390
rect 166340 54310 166350 54390
rect 166520 54310 166530 54390
rect 166700 54310 166710 54390
rect 166880 54310 166890 54390
rect 167060 54310 167070 54390
rect 167240 54310 167250 54390
rect 167420 54310 167430 54390
rect 167600 54310 167610 54390
rect 167780 54310 167790 54390
rect 167960 54310 167970 54390
rect 168140 54310 168150 54390
rect 168320 54310 168330 54390
rect 168500 54310 168510 54390
rect 168680 54310 168690 54390
rect 168860 54310 168870 54390
rect 169040 54310 169050 54390
rect 169220 54310 169230 54390
rect 169400 54310 169410 54390
rect 169580 54310 169590 54390
rect 169760 54310 169770 54390
rect 169940 54310 169950 54390
rect 170120 54310 170130 54390
rect 170810 54370 170840 54400
rect 170930 54370 170960 54400
rect 170690 54340 170750 54370
rect 170810 54340 170870 54370
rect 170930 54340 170990 54370
rect 19010 54240 19070 54270
rect 19130 54240 19190 54270
rect 19250 54240 19310 54270
rect 19800 54250 25800 54260
rect 26300 54240 26360 54270
rect 26420 54240 26480 54270
rect 26540 54240 26600 54270
rect 30300 54240 30360 54270
rect 30420 54240 30480 54270
rect 30540 54240 30600 54270
rect 37100 54260 37190 54270
rect 31100 54250 37190 54260
rect 19130 54150 19160 54180
rect 19250 54150 19280 54180
rect 26420 54150 26450 54180
rect 26540 54150 26570 54180
rect 30420 54150 30450 54180
rect 30540 54150 30570 54180
rect 19010 54120 19070 54150
rect 19130 54120 19190 54150
rect 19250 54120 19310 54150
rect 26300 54120 26360 54150
rect 26420 54120 26480 54150
rect 26540 54120 26600 54150
rect 30300 54120 30360 54150
rect 30420 54120 30480 54150
rect 30540 54120 30600 54150
rect 31180 54070 31260 54080
rect 31360 54070 31440 54080
rect 31540 54070 31620 54080
rect 31720 54070 31800 54080
rect 31900 54070 31980 54080
rect 32080 54070 32160 54080
rect 32260 54070 32340 54080
rect 32440 54070 32520 54080
rect 32620 54070 32700 54080
rect 32800 54070 32880 54080
rect 32980 54070 33060 54080
rect 33160 54070 33240 54080
rect 33340 54070 33420 54080
rect 33520 54070 33600 54080
rect 33700 54070 33780 54080
rect 33880 54070 33960 54080
rect 34060 54070 34140 54080
rect 34240 54070 34320 54080
rect 34420 54070 34500 54080
rect 34600 54070 34680 54080
rect 34780 54070 34860 54080
rect 34960 54070 35040 54080
rect 35140 54070 35220 54080
rect 35320 54070 35400 54080
rect 35500 54070 35580 54080
rect 35680 54070 35760 54080
rect 35860 54070 35940 54080
rect 36040 54070 36120 54080
rect 36220 54070 36300 54080
rect 36400 54070 36480 54080
rect 36580 54070 36660 54080
rect 36760 54070 36840 54080
rect 36940 54070 37020 54080
rect 19130 54030 19160 54060
rect 19250 54030 19280 54060
rect 19880 54050 19960 54060
rect 20060 54050 20140 54060
rect 20240 54050 20320 54060
rect 20420 54050 20500 54060
rect 20600 54050 20680 54060
rect 20780 54050 20860 54060
rect 20960 54050 21040 54060
rect 21140 54050 21220 54060
rect 21320 54050 21400 54060
rect 21500 54050 21580 54060
rect 21680 54050 21760 54060
rect 21860 54050 21940 54060
rect 22040 54050 22120 54060
rect 22220 54050 22300 54060
rect 22400 54050 22480 54060
rect 22580 54050 22660 54060
rect 22760 54050 22840 54060
rect 22940 54050 23020 54060
rect 23120 54050 23200 54060
rect 23300 54050 23380 54060
rect 23480 54050 23560 54060
rect 23660 54050 23740 54060
rect 23840 54050 23920 54060
rect 24020 54050 24100 54060
rect 24200 54050 24280 54060
rect 24380 54050 24460 54060
rect 24560 54050 24640 54060
rect 24740 54050 24820 54060
rect 24920 54050 25000 54060
rect 25100 54050 25180 54060
rect 25280 54050 25360 54060
rect 25460 54050 25540 54060
rect 25640 54050 25720 54060
rect 19010 54000 19070 54030
rect 19130 54000 19190 54030
rect 19250 54000 19310 54030
rect 19960 53970 19970 54050
rect 20140 53970 20150 54050
rect 20320 53970 20330 54050
rect 20500 53970 20510 54050
rect 20680 53970 20690 54050
rect 20860 53970 20870 54050
rect 21040 53970 21050 54050
rect 21220 53970 21230 54050
rect 21400 53970 21410 54050
rect 21580 53970 21590 54050
rect 21760 53970 21770 54050
rect 21940 53970 21950 54050
rect 22120 53970 22130 54050
rect 22300 53970 22310 54050
rect 22480 53970 22490 54050
rect 22660 53970 22670 54050
rect 22840 53970 22850 54050
rect 23020 53970 23030 54050
rect 23200 53970 23210 54050
rect 23380 53970 23390 54050
rect 23560 53970 23570 54050
rect 23740 53970 23750 54050
rect 23920 53970 23930 54050
rect 24100 53970 24110 54050
rect 24280 53970 24290 54050
rect 24460 53970 24470 54050
rect 24640 53970 24650 54050
rect 24820 53970 24830 54050
rect 25000 53970 25010 54050
rect 25180 53970 25190 54050
rect 25360 53970 25370 54050
rect 25540 53970 25550 54050
rect 25720 53970 25730 54050
rect 26420 54030 26450 54060
rect 26540 54030 26570 54060
rect 30420 54030 30450 54060
rect 30540 54030 30570 54060
rect 26300 54000 26360 54030
rect 26420 54000 26480 54030
rect 26540 54000 26600 54030
rect 30300 54000 30360 54030
rect 30420 54000 30480 54030
rect 30540 54000 30600 54030
rect 31260 53990 31270 54070
rect 31440 53990 31450 54070
rect 31620 53990 31630 54070
rect 31800 53990 31810 54070
rect 31980 53990 31990 54070
rect 32160 53990 32170 54070
rect 32340 53990 32350 54070
rect 32520 53990 32530 54070
rect 32700 53990 32710 54070
rect 32880 53990 32890 54070
rect 33060 53990 33070 54070
rect 33240 53990 33250 54070
rect 33420 53990 33430 54070
rect 33600 53990 33610 54070
rect 33780 53990 33790 54070
rect 33960 53990 33970 54070
rect 34140 53990 34150 54070
rect 34320 53990 34330 54070
rect 34500 53990 34510 54070
rect 34680 53990 34690 54070
rect 34860 53990 34870 54070
rect 35040 53990 35050 54070
rect 35220 53990 35230 54070
rect 35400 53990 35410 54070
rect 35580 53990 35590 54070
rect 35760 53990 35770 54070
rect 35940 53990 35950 54070
rect 36120 53990 36130 54070
rect 36300 53990 36310 54070
rect 36480 53990 36490 54070
rect 36660 53990 36670 54070
rect 36840 53990 36850 54070
rect 37020 53990 37030 54070
rect 19130 53910 19160 53940
rect 19250 53910 19280 53940
rect 26420 53910 26450 53940
rect 26540 53910 26570 53940
rect 30420 53910 30450 53940
rect 30540 53910 30570 53940
rect 19010 53880 19070 53910
rect 19130 53880 19190 53910
rect 19250 53880 19310 53910
rect 26300 53880 26360 53910
rect 26420 53880 26480 53910
rect 26540 53880 26600 53910
rect 30300 53880 30360 53910
rect 30420 53880 30480 53910
rect 30540 53880 30600 53910
rect 19130 53790 19160 53820
rect 19250 53790 19280 53820
rect 26420 53790 26450 53820
rect 26540 53790 26570 53820
rect 30420 53790 30450 53820
rect 30540 53790 30570 53820
rect 19010 53760 19070 53790
rect 19130 53760 19190 53790
rect 19250 53760 19310 53790
rect 26300 53760 26360 53790
rect 26420 53760 26480 53790
rect 26540 53760 26600 53790
rect 30300 53760 30360 53790
rect 30420 53760 30480 53790
rect 30540 53760 30600 53790
rect 19880 53750 19960 53760
rect 20060 53750 20140 53760
rect 20240 53750 20320 53760
rect 20420 53750 20500 53760
rect 20600 53750 20680 53760
rect 20780 53750 20860 53760
rect 20960 53750 21040 53760
rect 21140 53750 21220 53760
rect 21320 53750 21400 53760
rect 21500 53750 21580 53760
rect 21680 53750 21760 53760
rect 21860 53750 21940 53760
rect 22040 53750 22120 53760
rect 22220 53750 22300 53760
rect 22400 53750 22480 53760
rect 22580 53750 22660 53760
rect 22760 53750 22840 53760
rect 22940 53750 23020 53760
rect 23120 53750 23200 53760
rect 23300 53750 23380 53760
rect 23480 53750 23560 53760
rect 23660 53750 23740 53760
rect 23840 53750 23920 53760
rect 24020 53750 24100 53760
rect 24200 53750 24280 53760
rect 24380 53750 24460 53760
rect 24560 53750 24640 53760
rect 24740 53750 24820 53760
rect 24920 53750 25000 53760
rect 25100 53750 25180 53760
rect 25280 53750 25360 53760
rect 25460 53750 25540 53760
rect 25640 53750 25720 53760
rect 31180 53750 31260 53760
rect 31360 53750 31440 53760
rect 31540 53750 31620 53760
rect 31720 53750 31800 53760
rect 31900 53750 31980 53760
rect 32080 53750 32160 53760
rect 32260 53750 32340 53760
rect 32440 53750 32520 53760
rect 32620 53750 32700 53760
rect 32800 53750 32880 53760
rect 32980 53750 33060 53760
rect 33160 53750 33240 53760
rect 33340 53750 33420 53760
rect 33520 53750 33600 53760
rect 33700 53750 33780 53760
rect 33880 53750 33960 53760
rect 34060 53750 34140 53760
rect 34240 53750 34320 53760
rect 34420 53750 34500 53760
rect 34600 53750 34680 53760
rect 34780 53750 34860 53760
rect 34960 53750 35040 53760
rect 35140 53750 35220 53760
rect 35320 53750 35400 53760
rect 35500 53750 35580 53760
rect 35680 53750 35760 53760
rect 35860 53750 35940 53760
rect 36040 53750 36120 53760
rect 36220 53750 36300 53760
rect 36400 53750 36480 53760
rect 36580 53750 36660 53760
rect 36760 53750 36840 53760
rect 36940 53750 37020 53760
rect 19130 53670 19160 53700
rect 19250 53670 19280 53700
rect 19960 53670 19970 53750
rect 20140 53670 20150 53750
rect 20320 53670 20330 53750
rect 20500 53670 20510 53750
rect 20680 53670 20690 53750
rect 20860 53670 20870 53750
rect 21040 53670 21050 53750
rect 21220 53670 21230 53750
rect 21400 53670 21410 53750
rect 21580 53670 21590 53750
rect 21760 53670 21770 53750
rect 21940 53670 21950 53750
rect 22120 53670 22130 53750
rect 22300 53670 22310 53750
rect 22480 53670 22490 53750
rect 22660 53670 22670 53750
rect 22840 53670 22850 53750
rect 23020 53670 23030 53750
rect 23200 53670 23210 53750
rect 23380 53670 23390 53750
rect 23560 53670 23570 53750
rect 23740 53670 23750 53750
rect 23920 53670 23930 53750
rect 24100 53670 24110 53750
rect 24280 53670 24290 53750
rect 24460 53670 24470 53750
rect 24640 53670 24650 53750
rect 24820 53670 24830 53750
rect 25000 53670 25010 53750
rect 25180 53670 25190 53750
rect 25360 53670 25370 53750
rect 25540 53670 25550 53750
rect 25720 53670 25730 53750
rect 26420 53670 26450 53700
rect 26540 53670 26570 53700
rect 30420 53670 30450 53700
rect 30540 53670 30570 53700
rect 31260 53670 31270 53750
rect 31440 53670 31450 53750
rect 31620 53670 31630 53750
rect 31800 53670 31810 53750
rect 31980 53670 31990 53750
rect 32160 53670 32170 53750
rect 32340 53670 32350 53750
rect 32520 53670 32530 53750
rect 32700 53670 32710 53750
rect 32880 53670 32890 53750
rect 33060 53670 33070 53750
rect 33240 53670 33250 53750
rect 33420 53670 33430 53750
rect 33600 53670 33610 53750
rect 33780 53670 33790 53750
rect 33960 53670 33970 53750
rect 34140 53670 34150 53750
rect 34320 53670 34330 53750
rect 34500 53670 34510 53750
rect 34680 53670 34690 53750
rect 34860 53670 34870 53750
rect 35040 53670 35050 53750
rect 35220 53670 35230 53750
rect 35400 53670 35410 53750
rect 35580 53670 35590 53750
rect 35760 53670 35770 53750
rect 35940 53670 35950 53750
rect 36120 53670 36130 53750
rect 36300 53670 36310 53750
rect 36480 53670 36490 53750
rect 36660 53670 36670 53750
rect 36840 53670 36850 53750
rect 37020 53670 37030 53750
rect 19010 53640 19070 53670
rect 19130 53640 19190 53670
rect 19250 53640 19310 53670
rect 26300 53640 26360 53670
rect 26420 53640 26480 53670
rect 26540 53640 26600 53670
rect 30300 53640 30360 53670
rect 30420 53640 30480 53670
rect 30540 53640 30600 53670
rect 37100 53580 37190 54250
rect 37600 54240 37660 54270
rect 37720 54240 37780 54270
rect 37840 54240 37900 54270
rect 149075 54260 149315 54290
rect 149880 54270 149940 54300
rect 152220 54250 152250 54280
rect 152340 54250 152370 54280
rect 152900 54270 158990 54300
rect 158900 54260 158990 54270
rect 152900 54250 158990 54260
rect 159520 54250 159550 54280
rect 159640 54250 159670 54280
rect 163520 54250 163550 54280
rect 163640 54250 163670 54280
rect 164200 54250 170200 54260
rect 170810 54250 170840 54280
rect 170930 54250 170960 54280
rect 152100 54220 152160 54250
rect 152220 54220 152280 54250
rect 152340 54220 152400 54250
rect 40060 54190 40120 54220
rect 41540 54190 41600 54220
rect 42360 54190 42420 54220
rect 43840 54190 43900 54220
rect 37720 54150 37750 54180
rect 37840 54150 37870 54180
rect 146100 54150 146160 54180
rect 147580 54150 147640 54180
rect 148400 54150 148460 54180
rect 149880 54150 149940 54180
rect 37600 54120 37660 54150
rect 37720 54120 37780 54150
rect 37840 54120 37900 54150
rect 152220 54130 152250 54160
rect 152340 54130 152370 54160
rect 152100 54100 152160 54130
rect 152220 54100 152280 54130
rect 152340 54100 152400 54130
rect 40060 54070 40120 54100
rect 41540 54070 41600 54100
rect 42360 54070 42420 54100
rect 43840 54070 43900 54100
rect 152980 54070 153060 54080
rect 153160 54070 153240 54080
rect 153340 54070 153420 54080
rect 153520 54070 153600 54080
rect 153700 54070 153780 54080
rect 153880 54070 153960 54080
rect 154060 54070 154140 54080
rect 154240 54070 154320 54080
rect 154420 54070 154500 54080
rect 154600 54070 154680 54080
rect 154780 54070 154860 54080
rect 154960 54070 155040 54080
rect 155140 54070 155220 54080
rect 155320 54070 155400 54080
rect 155500 54070 155580 54080
rect 155680 54070 155760 54080
rect 155860 54070 155940 54080
rect 156040 54070 156120 54080
rect 156220 54070 156300 54080
rect 156400 54070 156480 54080
rect 156580 54070 156660 54080
rect 156760 54070 156840 54080
rect 156940 54070 157020 54080
rect 157120 54070 157200 54080
rect 157300 54070 157380 54080
rect 157480 54070 157560 54080
rect 157660 54070 157740 54080
rect 157840 54070 157920 54080
rect 158020 54070 158100 54080
rect 158200 54070 158280 54080
rect 158380 54070 158460 54080
rect 158560 54070 158640 54080
rect 158740 54070 158820 54080
rect 37720 54030 37750 54060
rect 37840 54030 37870 54060
rect 146100 54030 146160 54060
rect 147580 54030 147640 54060
rect 148400 54030 148460 54060
rect 149880 54030 149940 54060
rect 37600 54000 37660 54030
rect 37720 54000 37780 54030
rect 37840 54000 37900 54030
rect 40678 54004 40758 54014
rect 40838 54004 40918 54014
rect 152220 54010 152250 54040
rect 152340 54010 152370 54040
rect 40060 53950 40120 53980
rect 37720 53910 37750 53940
rect 37840 53910 37870 53940
rect 40758 53934 40768 54004
rect 40678 53924 40768 53934
rect 40838 53934 40848 54004
rect 40918 53934 40928 54004
rect 152100 53980 152160 54010
rect 152220 53980 152280 54010
rect 152340 53980 152400 54010
rect 153060 53990 153070 54070
rect 153240 53990 153250 54070
rect 153420 53990 153430 54070
rect 153600 53990 153610 54070
rect 153780 53990 153790 54070
rect 153960 53990 153970 54070
rect 154140 53990 154150 54070
rect 154320 53990 154330 54070
rect 154500 53990 154510 54070
rect 154680 53990 154690 54070
rect 154860 53990 154870 54070
rect 155040 53990 155050 54070
rect 155220 53990 155230 54070
rect 155400 53990 155410 54070
rect 155580 53990 155590 54070
rect 155760 53990 155770 54070
rect 155940 53990 155950 54070
rect 156120 53990 156130 54070
rect 156300 53990 156310 54070
rect 156480 53990 156490 54070
rect 156660 53990 156670 54070
rect 156840 53990 156850 54070
rect 157020 53990 157030 54070
rect 157200 53990 157210 54070
rect 157380 53990 157390 54070
rect 157560 53990 157570 54070
rect 157740 53990 157750 54070
rect 157920 53990 157930 54070
rect 158100 53990 158110 54070
rect 158280 53990 158290 54070
rect 158460 53990 158470 54070
rect 158640 53990 158650 54070
rect 158820 53990 158830 54070
rect 41540 53950 41600 53980
rect 42360 53950 42420 53980
rect 43840 53950 43900 53980
rect 40838 53924 40928 53934
rect 146100 53910 146160 53940
rect 147580 53910 147640 53940
rect 148400 53910 148460 53940
rect 149880 53910 149940 53940
rect 37600 53880 37660 53910
rect 37720 53880 37780 53910
rect 37840 53880 37900 53910
rect 152220 53890 152250 53920
rect 152340 53890 152370 53920
rect 152100 53860 152160 53890
rect 152220 53860 152280 53890
rect 152340 53860 152400 53890
rect 40060 53830 40120 53860
rect 40678 53844 40758 53854
rect 40838 53844 40918 53854
rect 37720 53790 37750 53820
rect 37840 53790 37870 53820
rect 37600 53760 37660 53790
rect 37720 53760 37780 53790
rect 37840 53760 37900 53790
rect 40758 53764 40768 53844
rect 40838 53764 40848 53844
rect 40918 53764 40928 53844
rect 41540 53830 41600 53860
rect 42360 53830 42420 53860
rect 43840 53830 43900 53860
rect 146100 53790 146160 53820
rect 147580 53790 147640 53820
rect 148400 53790 148460 53820
rect 149880 53790 149940 53820
rect 152220 53770 152250 53800
rect 152340 53770 152370 53800
rect 152100 53740 152160 53770
rect 152220 53740 152280 53770
rect 152340 53740 152400 53770
rect 152980 53750 153060 53760
rect 153160 53750 153240 53760
rect 153340 53750 153420 53760
rect 153520 53750 153600 53760
rect 153700 53750 153780 53760
rect 153880 53750 153960 53760
rect 154060 53750 154140 53760
rect 154240 53750 154320 53760
rect 154420 53750 154500 53760
rect 154600 53750 154680 53760
rect 154780 53750 154860 53760
rect 154960 53750 155040 53760
rect 155140 53750 155220 53760
rect 155320 53750 155400 53760
rect 155500 53750 155580 53760
rect 155680 53750 155760 53760
rect 155860 53750 155940 53760
rect 156040 53750 156120 53760
rect 156220 53750 156300 53760
rect 156400 53750 156480 53760
rect 156580 53750 156660 53760
rect 156760 53750 156840 53760
rect 156940 53750 157020 53760
rect 157120 53750 157200 53760
rect 157300 53750 157380 53760
rect 157480 53750 157560 53760
rect 157660 53750 157740 53760
rect 157840 53750 157920 53760
rect 158020 53750 158100 53760
rect 158200 53750 158280 53760
rect 158380 53750 158460 53760
rect 158560 53750 158640 53760
rect 158740 53750 158820 53760
rect 40060 53710 40120 53740
rect 41540 53710 41600 53740
rect 42360 53710 42420 53740
rect 43840 53710 43900 53740
rect 37720 53670 37750 53700
rect 37840 53670 37870 53700
rect 146100 53670 146160 53700
rect 147580 53670 147640 53700
rect 148400 53670 148460 53700
rect 149880 53670 149940 53700
rect 37600 53640 37660 53670
rect 37720 53640 37780 53670
rect 37840 53640 37900 53670
rect 152220 53650 152250 53680
rect 152340 53650 152370 53680
rect 153060 53670 153070 53750
rect 153240 53670 153250 53750
rect 153420 53670 153430 53750
rect 153600 53670 153610 53750
rect 153780 53670 153790 53750
rect 153960 53670 153970 53750
rect 154140 53670 154150 53750
rect 154320 53670 154330 53750
rect 154500 53670 154510 53750
rect 154680 53670 154690 53750
rect 154860 53670 154870 53750
rect 155040 53670 155050 53750
rect 155220 53670 155230 53750
rect 155400 53670 155410 53750
rect 155580 53670 155590 53750
rect 155760 53670 155770 53750
rect 155940 53670 155950 53750
rect 156120 53670 156130 53750
rect 156300 53670 156310 53750
rect 156480 53670 156490 53750
rect 156660 53670 156670 53750
rect 156840 53670 156850 53750
rect 157020 53670 157030 53750
rect 157200 53670 157210 53750
rect 157380 53670 157390 53750
rect 157560 53670 157570 53750
rect 157740 53670 157750 53750
rect 157920 53670 157930 53750
rect 158100 53670 158110 53750
rect 158280 53670 158290 53750
rect 158460 53670 158470 53750
rect 158640 53670 158650 53750
rect 158820 53670 158830 53750
rect 152100 53620 152160 53650
rect 152220 53620 152280 53650
rect 152340 53620 152400 53650
rect 40060 53590 40120 53620
rect 41540 53590 41600 53620
rect 42360 53590 42420 53620
rect 43840 53590 43900 53620
rect 158900 53580 158990 54250
rect 159400 54220 159460 54250
rect 159520 54220 159580 54250
rect 159640 54220 159700 54250
rect 163400 54220 163460 54250
rect 163520 54220 163580 54250
rect 163640 54220 163700 54250
rect 170690 54220 170750 54250
rect 170810 54220 170870 54250
rect 170930 54220 170990 54250
rect 159520 54130 159550 54160
rect 159640 54130 159670 54160
rect 163520 54130 163550 54160
rect 163640 54130 163670 54160
rect 170810 54130 170840 54160
rect 170930 54130 170960 54160
rect 159400 54100 159460 54130
rect 159520 54100 159580 54130
rect 159640 54100 159700 54130
rect 163400 54100 163460 54130
rect 163520 54100 163580 54130
rect 163640 54100 163700 54130
rect 170690 54100 170750 54130
rect 170810 54100 170870 54130
rect 170930 54100 170990 54130
rect 164280 54070 164360 54080
rect 164460 54070 164540 54080
rect 164640 54070 164720 54080
rect 164820 54070 164900 54080
rect 165000 54070 165080 54080
rect 165180 54070 165260 54080
rect 165360 54070 165440 54080
rect 165540 54070 165620 54080
rect 165720 54070 165800 54080
rect 165900 54070 165980 54080
rect 166080 54070 166160 54080
rect 166260 54070 166340 54080
rect 166440 54070 166520 54080
rect 166620 54070 166700 54080
rect 166800 54070 166880 54080
rect 166980 54070 167060 54080
rect 167160 54070 167240 54080
rect 167340 54070 167420 54080
rect 167520 54070 167600 54080
rect 167700 54070 167780 54080
rect 167880 54070 167960 54080
rect 168060 54070 168140 54080
rect 168240 54070 168320 54080
rect 168420 54070 168500 54080
rect 168600 54070 168680 54080
rect 168780 54070 168860 54080
rect 168960 54070 169040 54080
rect 169140 54070 169220 54080
rect 169320 54070 169400 54080
rect 169500 54070 169580 54080
rect 169680 54070 169760 54080
rect 169860 54070 169940 54080
rect 170040 54070 170120 54080
rect 159520 54010 159550 54040
rect 159640 54010 159670 54040
rect 163520 54010 163550 54040
rect 163640 54010 163670 54040
rect 159400 53980 159460 54010
rect 159520 53980 159580 54010
rect 159640 53980 159700 54010
rect 163400 53980 163460 54010
rect 163520 53980 163580 54010
rect 163640 53980 163700 54010
rect 164360 53990 164370 54070
rect 164540 53990 164550 54070
rect 164720 53990 164730 54070
rect 164900 53990 164910 54070
rect 165080 53990 165090 54070
rect 165260 53990 165270 54070
rect 165440 53990 165450 54070
rect 165620 53990 165630 54070
rect 165800 53990 165810 54070
rect 165980 53990 165990 54070
rect 166160 53990 166170 54070
rect 166340 53990 166350 54070
rect 166520 53990 166530 54070
rect 166700 53990 166710 54070
rect 166880 53990 166890 54070
rect 167060 53990 167070 54070
rect 167240 53990 167250 54070
rect 167420 53990 167430 54070
rect 167600 53990 167610 54070
rect 167780 53990 167790 54070
rect 167960 53990 167970 54070
rect 168140 53990 168150 54070
rect 168320 53990 168330 54070
rect 168500 53990 168510 54070
rect 168680 53990 168690 54070
rect 168860 53990 168870 54070
rect 169040 53990 169050 54070
rect 169220 53990 169230 54070
rect 169400 53990 169410 54070
rect 169580 53990 169590 54070
rect 169760 53990 169770 54070
rect 169940 53990 169950 54070
rect 170120 53990 170130 54070
rect 170810 54010 170840 54040
rect 170930 54010 170960 54040
rect 170690 53980 170750 54010
rect 170810 53980 170870 54010
rect 170930 53980 170990 54010
rect 159520 53890 159550 53920
rect 159640 53890 159670 53920
rect 163520 53890 163550 53920
rect 163640 53890 163670 53920
rect 170810 53890 170840 53920
rect 170930 53890 170960 53920
rect 159400 53860 159460 53890
rect 159520 53860 159580 53890
rect 159640 53860 159700 53890
rect 163400 53860 163460 53890
rect 163520 53860 163580 53890
rect 163640 53860 163700 53890
rect 170690 53860 170750 53890
rect 170810 53860 170870 53890
rect 170930 53860 170990 53890
rect 159520 53770 159550 53800
rect 159640 53770 159670 53800
rect 163520 53770 163550 53800
rect 163640 53770 163670 53800
rect 164280 53770 164360 53780
rect 164460 53770 164540 53780
rect 164640 53770 164720 53780
rect 164820 53770 164900 53780
rect 165000 53770 165080 53780
rect 165180 53770 165260 53780
rect 165360 53770 165440 53780
rect 165540 53770 165620 53780
rect 165720 53770 165800 53780
rect 165900 53770 165980 53780
rect 166080 53770 166160 53780
rect 166260 53770 166340 53780
rect 166440 53770 166520 53780
rect 166620 53770 166700 53780
rect 166800 53770 166880 53780
rect 166980 53770 167060 53780
rect 167160 53770 167240 53780
rect 167340 53770 167420 53780
rect 167520 53770 167600 53780
rect 167700 53770 167780 53780
rect 167880 53770 167960 53780
rect 168060 53770 168140 53780
rect 168240 53770 168320 53780
rect 168420 53770 168500 53780
rect 168600 53770 168680 53780
rect 168780 53770 168860 53780
rect 168960 53770 169040 53780
rect 169140 53770 169220 53780
rect 169320 53770 169400 53780
rect 169500 53770 169580 53780
rect 169680 53770 169760 53780
rect 169860 53770 169940 53780
rect 170040 53770 170120 53780
rect 170810 53770 170840 53800
rect 170930 53770 170960 53800
rect 159400 53740 159460 53770
rect 159520 53740 159580 53770
rect 159640 53740 159700 53770
rect 163400 53740 163460 53770
rect 163520 53740 163580 53770
rect 163640 53740 163700 53770
rect 164360 53690 164370 53770
rect 164540 53690 164550 53770
rect 164720 53690 164730 53770
rect 164900 53690 164910 53770
rect 165080 53690 165090 53770
rect 165260 53690 165270 53770
rect 165440 53690 165450 53770
rect 165620 53690 165630 53770
rect 165800 53690 165810 53770
rect 165980 53690 165990 53770
rect 166160 53690 166170 53770
rect 166340 53690 166350 53770
rect 166520 53690 166530 53770
rect 166700 53690 166710 53770
rect 166880 53690 166890 53770
rect 167060 53690 167070 53770
rect 167240 53690 167250 53770
rect 167420 53690 167430 53770
rect 167600 53690 167610 53770
rect 167780 53690 167790 53770
rect 167960 53690 167970 53770
rect 168140 53690 168150 53770
rect 168320 53690 168330 53770
rect 168500 53690 168510 53770
rect 168680 53690 168690 53770
rect 168860 53690 168870 53770
rect 169040 53690 169050 53770
rect 169220 53690 169230 53770
rect 169400 53690 169410 53770
rect 169580 53690 169590 53770
rect 169760 53690 169770 53770
rect 169940 53690 169950 53770
rect 170120 53690 170130 53770
rect 170690 53740 170750 53770
rect 170810 53740 170870 53770
rect 170930 53740 170990 53770
rect 159520 53650 159550 53680
rect 159640 53650 159670 53680
rect 163520 53650 163550 53680
rect 163640 53650 163670 53680
rect 170810 53650 170840 53680
rect 170930 53650 170960 53680
rect 159400 53620 159460 53650
rect 159520 53620 159580 53650
rect 159640 53620 159700 53650
rect 163400 53620 163460 53650
rect 163520 53620 163580 53650
rect 163640 53620 163700 53650
rect 170690 53620 170750 53650
rect 170810 53620 170870 53650
rect 170930 53620 170990 53650
rect 19130 53550 19160 53580
rect 19250 53550 19280 53580
rect 19800 53570 25800 53580
rect 26420 53550 26450 53580
rect 26540 53550 26570 53580
rect 30420 53550 30450 53580
rect 30540 53550 30570 53580
rect 31100 53570 37190 53580
rect 19010 53520 19070 53550
rect 19130 53520 19190 53550
rect 19250 53520 19310 53550
rect 26300 53520 26360 53550
rect 26420 53520 26480 53550
rect 26540 53520 26600 53550
rect 30300 53520 30360 53550
rect 30420 53520 30480 53550
rect 30540 53520 30600 53550
rect 37100 53470 37190 53570
rect 37720 53550 37750 53580
rect 37840 53550 37870 53580
rect 146100 53550 146160 53580
rect 147580 53550 147640 53580
rect 148400 53550 148460 53580
rect 149880 53550 149940 53580
rect 152900 53570 158990 53580
rect 164200 53570 170200 53580
rect 37600 53520 37660 53550
rect 37720 53520 37780 53550
rect 37840 53520 37900 53550
rect 152220 53530 152250 53560
rect 152340 53530 152370 53560
rect 152100 53500 152160 53530
rect 152220 53500 152280 53530
rect 152340 53500 152400 53530
rect 40060 53470 40120 53500
rect 41540 53470 41600 53500
rect 42360 53470 42420 53500
rect 43840 53470 43900 53500
rect 158900 53470 158990 53570
rect 159520 53530 159550 53560
rect 159640 53530 159670 53560
rect 163520 53530 163550 53560
rect 163640 53530 163670 53560
rect 170810 53530 170840 53560
rect 170930 53530 170960 53560
rect 159400 53500 159460 53530
rect 159520 53500 159580 53530
rect 159640 53500 159700 53530
rect 163400 53500 163460 53530
rect 163520 53500 163580 53530
rect 163640 53500 163700 53530
rect 170690 53500 170750 53530
rect 170810 53500 170870 53530
rect 170930 53500 170990 53530
rect 19130 53430 19160 53460
rect 19250 53430 19280 53460
rect 19880 53430 19960 53440
rect 20060 53430 20140 53440
rect 20240 53430 20320 53440
rect 20420 53430 20500 53440
rect 20600 53430 20680 53440
rect 20780 53430 20860 53440
rect 20960 53430 21040 53440
rect 21140 53430 21220 53440
rect 21320 53430 21400 53440
rect 21500 53430 21580 53440
rect 21680 53430 21760 53440
rect 21860 53430 21940 53440
rect 22040 53430 22120 53440
rect 22220 53430 22300 53440
rect 22400 53430 22480 53440
rect 22580 53430 22660 53440
rect 22760 53430 22840 53440
rect 22940 53430 23020 53440
rect 23120 53430 23200 53440
rect 23300 53430 23380 53440
rect 23480 53430 23560 53440
rect 23660 53430 23740 53440
rect 23840 53430 23920 53440
rect 24020 53430 24100 53440
rect 24200 53430 24280 53440
rect 24380 53430 24460 53440
rect 24560 53430 24640 53440
rect 24740 53430 24820 53440
rect 24920 53430 25000 53440
rect 25100 53430 25180 53440
rect 25280 53430 25360 53440
rect 25460 53430 25540 53440
rect 25640 53430 25720 53440
rect 26420 53430 26450 53460
rect 26540 53430 26570 53460
rect 30420 53430 30450 53460
rect 30540 53430 30570 53460
rect 31100 53440 37190 53470
rect 31180 53430 31260 53440
rect 31360 53430 31440 53440
rect 31540 53430 31620 53440
rect 31720 53430 31800 53440
rect 31900 53430 31980 53440
rect 32080 53430 32160 53440
rect 32260 53430 32340 53440
rect 32440 53430 32520 53440
rect 32620 53430 32700 53440
rect 32800 53430 32880 53440
rect 32980 53430 33060 53440
rect 33160 53430 33240 53440
rect 33340 53430 33420 53440
rect 33520 53430 33600 53440
rect 33700 53430 33780 53440
rect 33880 53430 33960 53440
rect 34060 53430 34140 53440
rect 34240 53430 34320 53440
rect 34420 53430 34500 53440
rect 34600 53430 34680 53440
rect 34780 53430 34860 53440
rect 34960 53430 35040 53440
rect 35140 53430 35220 53440
rect 35320 53430 35400 53440
rect 35500 53430 35580 53440
rect 35680 53430 35760 53440
rect 35860 53430 35940 53440
rect 36040 53430 36120 53440
rect 36220 53430 36300 53440
rect 36400 53430 36480 53440
rect 36580 53430 36660 53440
rect 36760 53430 36840 53440
rect 36940 53430 37020 53440
rect 19010 53400 19070 53430
rect 19130 53400 19190 53430
rect 19250 53400 19310 53430
rect 19960 53350 19970 53430
rect 20140 53350 20150 53430
rect 20320 53350 20330 53430
rect 20500 53350 20510 53430
rect 20680 53350 20690 53430
rect 20860 53350 20870 53430
rect 21040 53350 21050 53430
rect 21220 53350 21230 53430
rect 21400 53350 21410 53430
rect 21580 53350 21590 53430
rect 21760 53350 21770 53430
rect 21940 53350 21950 53430
rect 22120 53350 22130 53430
rect 22300 53350 22310 53430
rect 22480 53350 22490 53430
rect 22660 53350 22670 53430
rect 22840 53350 22850 53430
rect 23020 53350 23030 53430
rect 23200 53350 23210 53430
rect 23380 53350 23390 53430
rect 23560 53350 23570 53430
rect 23740 53350 23750 53430
rect 23920 53350 23930 53430
rect 24100 53350 24110 53430
rect 24280 53350 24290 53430
rect 24460 53350 24470 53430
rect 24640 53350 24650 53430
rect 24820 53350 24830 53430
rect 25000 53350 25010 53430
rect 25180 53350 25190 53430
rect 25360 53350 25370 53430
rect 25540 53350 25550 53430
rect 25720 53350 25730 53430
rect 26300 53400 26360 53430
rect 26420 53400 26480 53430
rect 26540 53400 26600 53430
rect 30300 53400 30360 53430
rect 30420 53400 30480 53430
rect 30540 53400 30600 53430
rect 31260 53370 31270 53430
rect 31440 53370 31450 53430
rect 31620 53370 31630 53430
rect 31800 53370 31810 53430
rect 31980 53370 31990 53430
rect 32160 53370 32170 53430
rect 32340 53370 32350 53430
rect 32520 53370 32530 53430
rect 32700 53370 32710 53430
rect 32880 53370 32890 53430
rect 33060 53370 33070 53430
rect 33240 53370 33250 53430
rect 33420 53370 33430 53430
rect 33600 53370 33610 53430
rect 33780 53370 33790 53430
rect 33960 53370 33970 53430
rect 34140 53370 34150 53430
rect 34320 53370 34330 53430
rect 34500 53370 34510 53430
rect 34680 53370 34690 53430
rect 34860 53370 34870 53430
rect 35040 53370 35050 53430
rect 35220 53370 35230 53430
rect 35400 53370 35410 53430
rect 35580 53370 35590 53430
rect 35760 53370 35770 53430
rect 35940 53370 35950 53430
rect 36120 53370 36130 53430
rect 36300 53370 36310 53430
rect 36480 53370 36490 53430
rect 36660 53370 36670 53430
rect 36840 53370 36850 53430
rect 37020 53370 37030 53430
rect 37100 53370 37190 53440
rect 37720 53430 37750 53460
rect 37840 53430 37870 53460
rect 146100 53430 146160 53460
rect 147580 53430 147640 53460
rect 148400 53430 148460 53460
rect 149880 53430 149940 53460
rect 152900 53440 158990 53470
rect 37600 53400 37660 53430
rect 37720 53400 37780 53430
rect 37840 53400 37900 53430
rect 152220 53410 152250 53440
rect 152340 53410 152370 53440
rect 152980 53430 153060 53440
rect 153160 53430 153240 53440
rect 153340 53430 153420 53440
rect 153520 53430 153600 53440
rect 153700 53430 153780 53440
rect 153880 53430 153960 53440
rect 154060 53430 154140 53440
rect 154240 53430 154320 53440
rect 154420 53430 154500 53440
rect 154600 53430 154680 53440
rect 154780 53430 154860 53440
rect 154960 53430 155040 53440
rect 155140 53430 155220 53440
rect 155320 53430 155400 53440
rect 155500 53430 155580 53440
rect 155680 53430 155760 53440
rect 155860 53430 155940 53440
rect 156040 53430 156120 53440
rect 156220 53430 156300 53440
rect 156400 53430 156480 53440
rect 156580 53430 156660 53440
rect 156760 53430 156840 53440
rect 156940 53430 157020 53440
rect 157120 53430 157200 53440
rect 157300 53430 157380 53440
rect 157480 53430 157560 53440
rect 157660 53430 157740 53440
rect 157840 53430 157920 53440
rect 158020 53430 158100 53440
rect 158200 53430 158280 53440
rect 158380 53430 158460 53440
rect 158560 53430 158640 53440
rect 158740 53430 158820 53440
rect 152100 53380 152160 53410
rect 152220 53380 152280 53410
rect 152340 53380 152400 53410
rect 31100 53340 37190 53370
rect 40060 53350 40120 53380
rect 41540 53350 41600 53380
rect 42360 53350 42420 53380
rect 43840 53350 43900 53380
rect 153060 53370 153070 53430
rect 153240 53370 153250 53430
rect 153420 53370 153430 53430
rect 153600 53370 153610 53430
rect 153780 53370 153790 53430
rect 153960 53370 153970 53430
rect 154140 53370 154150 53430
rect 154320 53370 154330 53430
rect 154500 53370 154510 53430
rect 154680 53370 154690 53430
rect 154860 53370 154870 53430
rect 155040 53370 155050 53430
rect 155220 53370 155230 53430
rect 155400 53370 155410 53430
rect 155580 53370 155590 53430
rect 155760 53370 155770 53430
rect 155940 53370 155950 53430
rect 156120 53370 156130 53430
rect 156300 53370 156310 53430
rect 156480 53370 156490 53430
rect 156660 53370 156670 53430
rect 156840 53370 156850 53430
rect 157020 53370 157030 53430
rect 157200 53370 157210 53430
rect 157380 53370 157390 53430
rect 157560 53370 157570 53430
rect 157740 53370 157750 53430
rect 157920 53370 157930 53430
rect 158100 53370 158110 53430
rect 158280 53370 158290 53430
rect 158460 53370 158470 53430
rect 158640 53370 158650 53430
rect 158820 53370 158830 53430
rect 158900 53370 158990 53440
rect 159520 53410 159550 53440
rect 159640 53410 159670 53440
rect 163520 53410 163550 53440
rect 163640 53410 163670 53440
rect 164280 53430 164360 53440
rect 164460 53430 164540 53440
rect 164640 53430 164720 53440
rect 164820 53430 164900 53440
rect 165000 53430 165080 53440
rect 165180 53430 165260 53440
rect 165360 53430 165440 53440
rect 165540 53430 165620 53440
rect 165720 53430 165800 53440
rect 165900 53430 165980 53440
rect 166080 53430 166160 53440
rect 166260 53430 166340 53440
rect 166440 53430 166520 53440
rect 166620 53430 166700 53440
rect 166800 53430 166880 53440
rect 166980 53430 167060 53440
rect 167160 53430 167240 53440
rect 167340 53430 167420 53440
rect 167520 53430 167600 53440
rect 167700 53430 167780 53440
rect 167880 53430 167960 53440
rect 168060 53430 168140 53440
rect 168240 53430 168320 53440
rect 168420 53430 168500 53440
rect 168600 53430 168680 53440
rect 168780 53430 168860 53440
rect 168960 53430 169040 53440
rect 169140 53430 169220 53440
rect 169320 53430 169400 53440
rect 169500 53430 169580 53440
rect 169680 53430 169760 53440
rect 169860 53430 169940 53440
rect 170040 53430 170120 53440
rect 159400 53380 159460 53410
rect 159520 53380 159580 53410
rect 159640 53380 159700 53410
rect 163400 53380 163460 53410
rect 163520 53380 163580 53410
rect 163640 53380 163700 53410
rect 152900 53340 158990 53370
rect 164360 53350 164370 53430
rect 164540 53350 164550 53430
rect 164720 53350 164730 53430
rect 164900 53350 164910 53430
rect 165080 53350 165090 53430
rect 165260 53350 165270 53430
rect 165440 53350 165450 53430
rect 165620 53350 165630 53430
rect 165800 53350 165810 53430
rect 165980 53350 165990 53430
rect 166160 53350 166170 53430
rect 166340 53350 166350 53430
rect 166520 53350 166530 53430
rect 166700 53350 166710 53430
rect 166880 53350 166890 53430
rect 167060 53350 167070 53430
rect 167240 53350 167250 53430
rect 167420 53350 167430 53430
rect 167600 53350 167610 53430
rect 167780 53350 167790 53430
rect 167960 53350 167970 53430
rect 168140 53350 168150 53430
rect 168320 53350 168330 53430
rect 168500 53350 168510 53430
rect 168680 53350 168690 53430
rect 168860 53350 168870 53430
rect 169040 53350 169050 53430
rect 169220 53350 169230 53430
rect 169400 53350 169410 53430
rect 169580 53350 169590 53430
rect 169760 53350 169770 53430
rect 169940 53350 169950 53430
rect 170120 53350 170130 53430
rect 170810 53410 170840 53440
rect 170930 53410 170960 53440
rect 170690 53380 170750 53410
rect 170810 53380 170870 53410
rect 170930 53380 170990 53410
rect 19130 53310 19160 53340
rect 19250 53310 19280 53340
rect 26420 53310 26450 53340
rect 26540 53310 26570 53340
rect 30420 53310 30450 53340
rect 30540 53310 30570 53340
rect 19010 53280 19070 53310
rect 19130 53280 19190 53310
rect 19250 53280 19310 53310
rect 19880 53280 19960 53290
rect 20060 53280 20140 53290
rect 20240 53280 20320 53290
rect 20420 53280 20500 53290
rect 20600 53280 20680 53290
rect 20780 53280 20860 53290
rect 20960 53280 21040 53290
rect 21140 53280 21220 53290
rect 21320 53280 21400 53290
rect 21500 53280 21580 53290
rect 21680 53280 21760 53290
rect 21860 53280 21940 53290
rect 22040 53280 22120 53290
rect 22220 53280 22300 53290
rect 22400 53280 22480 53290
rect 22580 53280 22660 53290
rect 22760 53280 22840 53290
rect 22940 53280 23020 53290
rect 23120 53280 23200 53290
rect 23300 53280 23380 53290
rect 23480 53280 23560 53290
rect 23660 53280 23740 53290
rect 23840 53280 23920 53290
rect 24020 53280 24100 53290
rect 24200 53280 24280 53290
rect 24380 53280 24460 53290
rect 24560 53280 24640 53290
rect 24740 53280 24820 53290
rect 24920 53280 25000 53290
rect 25100 53280 25180 53290
rect 25280 53280 25360 53290
rect 25460 53280 25540 53290
rect 25640 53280 25720 53290
rect 26300 53280 26360 53310
rect 26420 53280 26480 53310
rect 26540 53280 26600 53310
rect 30300 53280 30360 53310
rect 30420 53280 30480 53310
rect 30540 53280 30600 53310
rect 31180 53280 31260 53290
rect 31360 53280 31440 53290
rect 31540 53280 31620 53290
rect 31720 53280 31800 53290
rect 31900 53280 31980 53290
rect 32080 53280 32160 53290
rect 32260 53280 32340 53290
rect 32440 53280 32520 53290
rect 32620 53280 32700 53290
rect 32800 53280 32880 53290
rect 32980 53280 33060 53290
rect 33160 53280 33240 53290
rect 33340 53280 33420 53290
rect 33520 53280 33600 53290
rect 33700 53280 33780 53290
rect 33880 53280 33960 53290
rect 34060 53280 34140 53290
rect 34240 53280 34320 53290
rect 34420 53280 34500 53290
rect 34600 53280 34680 53290
rect 34780 53280 34860 53290
rect 34960 53280 35040 53290
rect 35140 53280 35220 53290
rect 35320 53280 35400 53290
rect 35500 53280 35580 53290
rect 35680 53280 35760 53290
rect 35860 53280 35940 53290
rect 36040 53280 36120 53290
rect 36220 53280 36300 53290
rect 36400 53280 36480 53290
rect 36580 53280 36660 53290
rect 36760 53280 36840 53290
rect 36940 53280 37020 53290
rect 19130 53190 19160 53220
rect 19250 53190 19280 53220
rect 19960 53200 19970 53280
rect 20140 53200 20150 53280
rect 20320 53200 20330 53280
rect 20500 53200 20510 53280
rect 20680 53200 20690 53280
rect 20860 53200 20870 53280
rect 21040 53200 21050 53280
rect 21220 53200 21230 53280
rect 21400 53200 21410 53280
rect 21580 53200 21590 53280
rect 21760 53200 21770 53280
rect 21940 53200 21950 53280
rect 22120 53200 22130 53280
rect 22300 53200 22310 53280
rect 22480 53200 22490 53280
rect 22660 53200 22670 53280
rect 22840 53200 22850 53280
rect 23020 53200 23030 53280
rect 23200 53200 23210 53280
rect 23380 53200 23390 53280
rect 23560 53200 23570 53280
rect 23740 53200 23750 53280
rect 23920 53200 23930 53280
rect 24100 53200 24110 53280
rect 24280 53200 24290 53280
rect 24460 53200 24470 53280
rect 24640 53200 24650 53280
rect 24820 53200 24830 53280
rect 25000 53200 25010 53280
rect 25180 53200 25190 53280
rect 25360 53200 25370 53280
rect 25540 53200 25550 53280
rect 25720 53200 25730 53280
rect 26420 53190 26450 53220
rect 26540 53190 26570 53220
rect 30420 53190 30450 53220
rect 30540 53190 30570 53220
rect 31260 53200 31270 53280
rect 31440 53200 31450 53280
rect 31620 53200 31630 53280
rect 31800 53200 31810 53280
rect 31980 53200 31990 53280
rect 32160 53200 32170 53280
rect 32340 53200 32350 53280
rect 32520 53200 32530 53280
rect 32700 53200 32710 53280
rect 32880 53200 32890 53280
rect 33060 53200 33070 53280
rect 33240 53200 33250 53280
rect 33420 53200 33430 53280
rect 33600 53200 33610 53280
rect 33780 53200 33790 53280
rect 33960 53200 33970 53280
rect 34140 53200 34150 53280
rect 34320 53200 34330 53280
rect 34500 53200 34510 53280
rect 34680 53200 34690 53280
rect 34860 53200 34870 53280
rect 35040 53200 35050 53280
rect 35220 53200 35230 53280
rect 35400 53200 35410 53280
rect 35580 53200 35590 53280
rect 35760 53200 35770 53280
rect 35940 53200 35950 53280
rect 36120 53200 36130 53280
rect 36300 53200 36310 53280
rect 36480 53200 36490 53280
rect 36660 53200 36670 53280
rect 36840 53200 36850 53280
rect 37020 53200 37030 53280
rect 19010 53160 19070 53190
rect 19130 53160 19190 53190
rect 19250 53160 19310 53190
rect 26300 53160 26360 53190
rect 26420 53160 26480 53190
rect 26540 53160 26600 53190
rect 30300 53160 30360 53190
rect 30420 53160 30480 53190
rect 30540 53160 30600 53190
rect 37100 53140 37190 53340
rect 37720 53310 37750 53340
rect 37840 53310 37870 53340
rect 146100 53310 146160 53340
rect 147580 53310 147640 53340
rect 148400 53310 148460 53340
rect 149880 53310 149940 53340
rect 37600 53280 37660 53310
rect 37720 53280 37780 53310
rect 37840 53280 37900 53310
rect 152220 53290 152250 53320
rect 152340 53290 152370 53320
rect 152100 53260 152160 53290
rect 152220 53260 152280 53290
rect 152340 53260 152400 53290
rect 152980 53280 153060 53290
rect 153160 53280 153240 53290
rect 153340 53280 153420 53290
rect 153520 53280 153600 53290
rect 153700 53280 153780 53290
rect 153880 53280 153960 53290
rect 154060 53280 154140 53290
rect 154240 53280 154320 53290
rect 154420 53280 154500 53290
rect 154600 53280 154680 53290
rect 154780 53280 154860 53290
rect 154960 53280 155040 53290
rect 155140 53280 155220 53290
rect 155320 53280 155400 53290
rect 155500 53280 155580 53290
rect 155680 53280 155760 53290
rect 155860 53280 155940 53290
rect 156040 53280 156120 53290
rect 156220 53280 156300 53290
rect 156400 53280 156480 53290
rect 156580 53280 156660 53290
rect 156760 53280 156840 53290
rect 156940 53280 157020 53290
rect 157120 53280 157200 53290
rect 157300 53280 157380 53290
rect 157480 53280 157560 53290
rect 157660 53280 157740 53290
rect 157840 53280 157920 53290
rect 158020 53280 158100 53290
rect 158200 53280 158280 53290
rect 158380 53280 158460 53290
rect 158560 53280 158640 53290
rect 158740 53280 158820 53290
rect 40060 53230 40120 53260
rect 41540 53230 41600 53260
rect 42360 53230 42420 53260
rect 43840 53230 43900 53260
rect 37720 53190 37750 53220
rect 37840 53190 37870 53220
rect 146100 53190 146160 53220
rect 147580 53190 147640 53220
rect 148400 53190 148460 53220
rect 149880 53190 149940 53220
rect 153060 53200 153070 53280
rect 153240 53200 153250 53280
rect 153420 53200 153430 53280
rect 153600 53200 153610 53280
rect 153780 53200 153790 53280
rect 153960 53200 153970 53280
rect 154140 53200 154150 53280
rect 154320 53200 154330 53280
rect 154500 53200 154510 53280
rect 154680 53200 154690 53280
rect 154860 53200 154870 53280
rect 155040 53200 155050 53280
rect 155220 53200 155230 53280
rect 155400 53200 155410 53280
rect 155580 53200 155590 53280
rect 155760 53200 155770 53280
rect 155940 53200 155950 53280
rect 156120 53200 156130 53280
rect 156300 53200 156310 53280
rect 156480 53200 156490 53280
rect 156660 53200 156670 53280
rect 156840 53200 156850 53280
rect 157020 53200 157030 53280
rect 157200 53200 157210 53280
rect 157380 53200 157390 53280
rect 157560 53200 157570 53280
rect 157740 53200 157750 53280
rect 157920 53200 157930 53280
rect 158100 53200 158110 53280
rect 158280 53200 158290 53280
rect 158460 53200 158470 53280
rect 158640 53200 158650 53280
rect 158820 53200 158830 53280
rect 37600 53160 37660 53190
rect 37720 53160 37780 53190
rect 37840 53160 37900 53190
rect 152220 53170 152250 53200
rect 152340 53170 152370 53200
rect 152100 53140 152160 53170
rect 152220 53140 152280 53170
rect 152340 53140 152400 53170
rect 158900 53140 158990 53340
rect 159520 53290 159550 53320
rect 159640 53290 159670 53320
rect 163520 53290 163550 53320
rect 163640 53290 163670 53320
rect 170810 53290 170840 53320
rect 170930 53290 170960 53320
rect 159400 53260 159460 53290
rect 159520 53260 159580 53290
rect 159640 53260 159700 53290
rect 163400 53260 163460 53290
rect 163520 53260 163580 53290
rect 163640 53260 163700 53290
rect 164280 53280 164360 53290
rect 164460 53280 164540 53290
rect 164640 53280 164720 53290
rect 164820 53280 164900 53290
rect 165000 53280 165080 53290
rect 165180 53280 165260 53290
rect 165360 53280 165440 53290
rect 165540 53280 165620 53290
rect 165720 53280 165800 53290
rect 165900 53280 165980 53290
rect 166080 53280 166160 53290
rect 166260 53280 166340 53290
rect 166440 53280 166520 53290
rect 166620 53280 166700 53290
rect 166800 53280 166880 53290
rect 166980 53280 167060 53290
rect 167160 53280 167240 53290
rect 167340 53280 167420 53290
rect 167520 53280 167600 53290
rect 167700 53280 167780 53290
rect 167880 53280 167960 53290
rect 168060 53280 168140 53290
rect 168240 53280 168320 53290
rect 168420 53280 168500 53290
rect 168600 53280 168680 53290
rect 168780 53280 168860 53290
rect 168960 53280 169040 53290
rect 169140 53280 169220 53290
rect 169320 53280 169400 53290
rect 169500 53280 169580 53290
rect 169680 53280 169760 53290
rect 169860 53280 169940 53290
rect 170040 53280 170120 53290
rect 164360 53200 164370 53280
rect 164540 53200 164550 53280
rect 164720 53200 164730 53280
rect 164900 53200 164910 53280
rect 165080 53200 165090 53280
rect 165260 53200 165270 53280
rect 165440 53200 165450 53280
rect 165620 53200 165630 53280
rect 165800 53200 165810 53280
rect 165980 53200 165990 53280
rect 166160 53200 166170 53280
rect 166340 53200 166350 53280
rect 166520 53200 166530 53280
rect 166700 53200 166710 53280
rect 166880 53200 166890 53280
rect 167060 53200 167070 53280
rect 167240 53200 167250 53280
rect 167420 53200 167430 53280
rect 167600 53200 167610 53280
rect 167780 53200 167790 53280
rect 167960 53200 167970 53280
rect 168140 53200 168150 53280
rect 168320 53200 168330 53280
rect 168500 53200 168510 53280
rect 168680 53200 168690 53280
rect 168860 53200 168870 53280
rect 169040 53200 169050 53280
rect 169220 53200 169230 53280
rect 169400 53200 169410 53280
rect 169580 53200 169590 53280
rect 169760 53200 169770 53280
rect 169940 53200 169950 53280
rect 170120 53200 170130 53280
rect 170690 53260 170750 53290
rect 170810 53260 170870 53290
rect 170930 53260 170990 53290
rect 159520 53170 159550 53200
rect 159640 53170 159670 53200
rect 163520 53170 163550 53200
rect 163640 53170 163670 53200
rect 170810 53170 170840 53200
rect 170930 53170 170960 53200
rect 159400 53140 159460 53170
rect 159520 53140 159580 53170
rect 159640 53140 159700 53170
rect 163400 53140 163460 53170
rect 163520 53140 163580 53170
rect 163640 53140 163700 53170
rect 170690 53140 170750 53170
rect 170810 53140 170870 53170
rect 170930 53140 170990 53170
rect 19880 53130 19960 53140
rect 20060 53130 20140 53140
rect 20240 53130 20320 53140
rect 20420 53130 20500 53140
rect 20600 53130 20680 53140
rect 20780 53130 20860 53140
rect 20960 53130 21040 53140
rect 21140 53130 21220 53140
rect 21320 53130 21400 53140
rect 21500 53130 21580 53140
rect 21680 53130 21760 53140
rect 21860 53130 21940 53140
rect 22040 53130 22120 53140
rect 22220 53130 22300 53140
rect 22400 53130 22480 53140
rect 22580 53130 22660 53140
rect 22760 53130 22840 53140
rect 22940 53130 23020 53140
rect 23120 53130 23200 53140
rect 23300 53130 23380 53140
rect 23480 53130 23560 53140
rect 23660 53130 23740 53140
rect 23840 53130 23920 53140
rect 24020 53130 24100 53140
rect 24200 53130 24280 53140
rect 24380 53130 24460 53140
rect 24560 53130 24640 53140
rect 24740 53130 24820 53140
rect 24920 53130 25000 53140
rect 25100 53130 25180 53140
rect 25280 53130 25360 53140
rect 25460 53130 25540 53140
rect 25640 53130 25720 53140
rect 19130 53070 19160 53100
rect 19250 53070 19280 53100
rect 19010 53040 19070 53070
rect 19130 53040 19190 53070
rect 19250 53040 19310 53070
rect 19960 53050 19970 53130
rect 20140 53050 20150 53130
rect 20320 53050 20330 53130
rect 20500 53050 20510 53130
rect 20680 53050 20690 53130
rect 20860 53050 20870 53130
rect 21040 53050 21050 53130
rect 21220 53050 21230 53130
rect 21400 53050 21410 53130
rect 21580 53050 21590 53130
rect 21760 53050 21770 53130
rect 21940 53050 21950 53130
rect 22120 53050 22130 53130
rect 22300 53050 22310 53130
rect 22480 53050 22490 53130
rect 22660 53050 22670 53130
rect 22840 53050 22850 53130
rect 23020 53050 23030 53130
rect 23200 53050 23210 53130
rect 23380 53050 23390 53130
rect 23560 53050 23570 53130
rect 23740 53050 23750 53130
rect 23920 53050 23930 53130
rect 24100 53050 24110 53130
rect 24280 53050 24290 53130
rect 24460 53050 24470 53130
rect 24640 53050 24650 53130
rect 24820 53050 24830 53130
rect 25000 53050 25010 53130
rect 25180 53050 25190 53130
rect 25360 53050 25370 53130
rect 25540 53050 25550 53130
rect 25720 53050 25730 53130
rect 31100 53110 37190 53140
rect 40060 53110 40120 53140
rect 41540 53110 41600 53140
rect 42360 53110 42420 53140
rect 43840 53110 43900 53140
rect 152900 53110 158990 53140
rect 164280 53130 164360 53140
rect 164460 53130 164540 53140
rect 164640 53130 164720 53140
rect 164820 53130 164900 53140
rect 165000 53130 165080 53140
rect 165180 53130 165260 53140
rect 165360 53130 165440 53140
rect 165540 53130 165620 53140
rect 165720 53130 165800 53140
rect 165900 53130 165980 53140
rect 166080 53130 166160 53140
rect 166260 53130 166340 53140
rect 166440 53130 166520 53140
rect 166620 53130 166700 53140
rect 166800 53130 166880 53140
rect 166980 53130 167060 53140
rect 167160 53130 167240 53140
rect 167340 53130 167420 53140
rect 167520 53130 167600 53140
rect 167700 53130 167780 53140
rect 167880 53130 167960 53140
rect 168060 53130 168140 53140
rect 168240 53130 168320 53140
rect 168420 53130 168500 53140
rect 168600 53130 168680 53140
rect 168780 53130 168860 53140
rect 168960 53130 169040 53140
rect 169140 53130 169220 53140
rect 169320 53130 169400 53140
rect 169500 53130 169580 53140
rect 169680 53130 169760 53140
rect 169860 53130 169940 53140
rect 170040 53130 170120 53140
rect 26420 53070 26450 53100
rect 26540 53070 26570 53100
rect 30420 53070 30450 53100
rect 30540 53070 30570 53100
rect 26300 53040 26360 53070
rect 26420 53040 26480 53070
rect 26540 53040 26600 53070
rect 30300 53040 30360 53070
rect 30420 53040 30480 53070
rect 30540 53040 30600 53070
rect 31260 53050 31270 53110
rect 31440 53050 31450 53110
rect 31620 53050 31630 53110
rect 31800 53050 31810 53110
rect 31980 53050 31990 53110
rect 32160 53050 32170 53110
rect 32340 53050 32350 53110
rect 32520 53050 32530 53110
rect 32700 53050 32710 53110
rect 32880 53050 32890 53110
rect 33060 53050 33070 53110
rect 33240 53050 33250 53110
rect 33420 53050 33430 53110
rect 33600 53050 33610 53110
rect 33780 53050 33790 53110
rect 33960 53050 33970 53110
rect 34140 53050 34150 53110
rect 34320 53050 34330 53110
rect 34500 53050 34510 53110
rect 34680 53050 34690 53110
rect 34860 53050 34870 53110
rect 35040 53050 35050 53110
rect 35220 53050 35230 53110
rect 35400 53050 35410 53110
rect 35580 53050 35590 53110
rect 35760 53050 35770 53110
rect 35940 53050 35950 53110
rect 36120 53050 36130 53110
rect 36300 53050 36310 53110
rect 36480 53050 36490 53110
rect 36660 53050 36670 53110
rect 36840 53050 36850 53110
rect 37020 53050 37030 53110
rect 37100 53040 37190 53110
rect 37720 53070 37750 53100
rect 37840 53070 37870 53100
rect 146100 53070 146160 53100
rect 147580 53070 147640 53100
rect 148400 53070 148460 53100
rect 149880 53070 149940 53100
rect 37600 53040 37660 53070
rect 37720 53040 37780 53070
rect 37840 53040 37900 53070
rect 152220 53050 152250 53080
rect 152340 53050 152370 53080
rect 153060 53050 153070 53110
rect 153240 53050 153250 53110
rect 153420 53050 153430 53110
rect 153600 53050 153610 53110
rect 153780 53050 153790 53110
rect 153960 53050 153970 53110
rect 154140 53050 154150 53110
rect 154320 53050 154330 53110
rect 154500 53050 154510 53110
rect 154680 53050 154690 53110
rect 154860 53050 154870 53110
rect 155040 53050 155050 53110
rect 155220 53050 155230 53110
rect 155400 53050 155410 53110
rect 155580 53050 155590 53110
rect 155760 53050 155770 53110
rect 155940 53050 155950 53110
rect 156120 53050 156130 53110
rect 156300 53050 156310 53110
rect 156480 53050 156490 53110
rect 156660 53050 156670 53110
rect 156840 53050 156850 53110
rect 157020 53050 157030 53110
rect 157200 53050 157210 53110
rect 157380 53050 157390 53110
rect 157560 53050 157570 53110
rect 157740 53050 157750 53110
rect 157920 53050 157930 53110
rect 158100 53050 158110 53110
rect 158280 53050 158290 53110
rect 158460 53050 158470 53110
rect 158640 53050 158650 53110
rect 158820 53050 158830 53110
rect 31100 53010 37190 53040
rect 152100 53020 152160 53050
rect 152220 53020 152280 53050
rect 152340 53020 152400 53050
rect 158900 53040 158990 53110
rect 159520 53050 159550 53080
rect 159640 53050 159670 53080
rect 163520 53050 163550 53080
rect 163640 53050 163670 53080
rect 164360 53050 164370 53130
rect 164540 53050 164550 53130
rect 164720 53050 164730 53130
rect 164900 53050 164910 53130
rect 165080 53050 165090 53130
rect 165260 53050 165270 53130
rect 165440 53050 165450 53130
rect 165620 53050 165630 53130
rect 165800 53050 165810 53130
rect 165980 53050 165990 53130
rect 166160 53050 166170 53130
rect 166340 53050 166350 53130
rect 166520 53050 166530 53130
rect 166700 53050 166710 53130
rect 166880 53050 166890 53130
rect 167060 53050 167070 53130
rect 167240 53050 167250 53130
rect 167420 53050 167430 53130
rect 167600 53050 167610 53130
rect 167780 53050 167790 53130
rect 167960 53050 167970 53130
rect 168140 53050 168150 53130
rect 168320 53050 168330 53130
rect 168500 53050 168510 53130
rect 168680 53050 168690 53130
rect 168860 53050 168870 53130
rect 169040 53050 169050 53130
rect 169220 53050 169230 53130
rect 169400 53050 169410 53130
rect 169580 53050 169590 53130
rect 169760 53050 169770 53130
rect 169940 53050 169950 53130
rect 170120 53050 170130 53130
rect 170810 53050 170840 53080
rect 170930 53050 170960 53080
rect 37100 53000 37190 53010
rect 19800 52990 25800 53000
rect 31100 52990 37190 53000
rect 40060 52990 40120 53020
rect 41540 52990 41600 53020
rect 42360 52990 42420 53020
rect 43840 52990 43900 53020
rect 152900 53010 158990 53040
rect 159400 53020 159460 53050
rect 159520 53020 159580 53050
rect 159640 53020 159700 53050
rect 163400 53020 163460 53050
rect 163520 53020 163580 53050
rect 163640 53020 163700 53050
rect 170690 53020 170750 53050
rect 170810 53020 170870 53050
rect 170930 53020 170990 53050
rect 158900 53000 158990 53010
rect 152900 52990 158990 53000
rect 164200 52990 170200 53000
rect 19130 52950 19160 52980
rect 19250 52950 19280 52980
rect 26420 52950 26450 52980
rect 26540 52950 26570 52980
rect 30420 52950 30450 52980
rect 30540 52950 30570 52980
rect 19010 52920 19070 52950
rect 19130 52920 19190 52950
rect 19250 52920 19310 52950
rect 26300 52920 26360 52950
rect 26420 52920 26480 52950
rect 26540 52920 26600 52950
rect 30300 52920 30360 52950
rect 30420 52920 30480 52950
rect 30540 52920 30600 52950
rect 19130 52830 19160 52860
rect 19250 52830 19280 52860
rect 26420 52830 26450 52860
rect 26540 52830 26570 52860
rect 30420 52830 30450 52860
rect 30540 52830 30570 52860
rect 19010 52800 19070 52830
rect 19130 52800 19190 52830
rect 19250 52800 19310 52830
rect 26300 52800 26360 52830
rect 26420 52800 26480 52830
rect 26540 52800 26600 52830
rect 30300 52800 30360 52830
rect 30420 52800 30480 52830
rect 30540 52800 30600 52830
rect 31180 52810 31260 52820
rect 31360 52810 31440 52820
rect 31540 52810 31620 52820
rect 31720 52810 31800 52820
rect 31900 52810 31980 52820
rect 32080 52810 32160 52820
rect 32260 52810 32340 52820
rect 32440 52810 32520 52820
rect 32620 52810 32700 52820
rect 32800 52810 32880 52820
rect 32980 52810 33060 52820
rect 33160 52810 33240 52820
rect 33340 52810 33420 52820
rect 33520 52810 33600 52820
rect 33700 52810 33780 52820
rect 33880 52810 33960 52820
rect 34060 52810 34140 52820
rect 34240 52810 34320 52820
rect 34420 52810 34500 52820
rect 34600 52810 34680 52820
rect 34780 52810 34860 52820
rect 34960 52810 35040 52820
rect 35140 52810 35220 52820
rect 35320 52810 35400 52820
rect 35500 52810 35580 52820
rect 35680 52810 35760 52820
rect 35860 52810 35940 52820
rect 36040 52810 36120 52820
rect 36220 52810 36300 52820
rect 36400 52810 36480 52820
rect 36580 52810 36660 52820
rect 36760 52810 36840 52820
rect 36940 52810 37020 52820
rect 19880 52790 19960 52800
rect 20060 52790 20140 52800
rect 20240 52790 20320 52800
rect 20420 52790 20500 52800
rect 20600 52790 20680 52800
rect 20780 52790 20860 52800
rect 20960 52790 21040 52800
rect 21140 52790 21220 52800
rect 21320 52790 21400 52800
rect 21500 52790 21580 52800
rect 21680 52790 21760 52800
rect 21860 52790 21940 52800
rect 22040 52790 22120 52800
rect 22220 52790 22300 52800
rect 22400 52790 22480 52800
rect 22580 52790 22660 52800
rect 22760 52790 22840 52800
rect 22940 52790 23020 52800
rect 23120 52790 23200 52800
rect 23300 52790 23380 52800
rect 23480 52790 23560 52800
rect 23660 52790 23740 52800
rect 23840 52790 23920 52800
rect 24020 52790 24100 52800
rect 24200 52790 24280 52800
rect 24380 52790 24460 52800
rect 24560 52790 24640 52800
rect 24740 52790 24820 52800
rect 24920 52790 25000 52800
rect 25100 52790 25180 52800
rect 25280 52790 25360 52800
rect 25460 52790 25540 52800
rect 25640 52790 25720 52800
rect 19130 52710 19160 52740
rect 19250 52710 19280 52740
rect 19960 52710 19970 52790
rect 20140 52710 20150 52790
rect 20320 52710 20330 52790
rect 20500 52710 20510 52790
rect 20680 52710 20690 52790
rect 20860 52710 20870 52790
rect 21040 52710 21050 52790
rect 21220 52710 21230 52790
rect 21400 52710 21410 52790
rect 21580 52710 21590 52790
rect 21760 52710 21770 52790
rect 21940 52710 21950 52790
rect 22120 52710 22130 52790
rect 22300 52710 22310 52790
rect 22480 52710 22490 52790
rect 22660 52710 22670 52790
rect 22840 52710 22850 52790
rect 23020 52710 23030 52790
rect 23200 52710 23210 52790
rect 23380 52710 23390 52790
rect 23560 52710 23570 52790
rect 23740 52710 23750 52790
rect 23920 52710 23930 52790
rect 24100 52710 24110 52790
rect 24280 52710 24290 52790
rect 24460 52710 24470 52790
rect 24640 52710 24650 52790
rect 24820 52710 24830 52790
rect 25000 52710 25010 52790
rect 25180 52710 25190 52790
rect 25360 52710 25370 52790
rect 25540 52710 25550 52790
rect 25720 52710 25730 52790
rect 26420 52710 26450 52740
rect 26540 52710 26570 52740
rect 30420 52710 30450 52740
rect 30540 52710 30570 52740
rect 31260 52730 31270 52810
rect 31440 52730 31450 52810
rect 31620 52730 31630 52810
rect 31800 52730 31810 52810
rect 31980 52730 31990 52810
rect 32160 52730 32170 52810
rect 32340 52730 32350 52810
rect 32520 52730 32530 52810
rect 32700 52730 32710 52810
rect 32880 52730 32890 52810
rect 33060 52730 33070 52810
rect 33240 52730 33250 52810
rect 33420 52730 33430 52810
rect 33600 52730 33610 52810
rect 33780 52730 33790 52810
rect 33960 52730 33970 52810
rect 34140 52730 34150 52810
rect 34320 52730 34330 52810
rect 34500 52730 34510 52810
rect 34680 52730 34690 52810
rect 34860 52730 34870 52810
rect 35040 52730 35050 52810
rect 35220 52730 35230 52810
rect 35400 52730 35410 52810
rect 35580 52730 35590 52810
rect 35760 52730 35770 52810
rect 35940 52730 35950 52810
rect 36120 52730 36130 52810
rect 36300 52730 36310 52810
rect 36480 52730 36490 52810
rect 36660 52730 36670 52810
rect 36840 52730 36850 52810
rect 37020 52730 37030 52810
rect 19010 52680 19070 52710
rect 19130 52680 19190 52710
rect 19250 52680 19310 52710
rect 26300 52680 26360 52710
rect 26420 52680 26480 52710
rect 26540 52680 26600 52710
rect 30300 52680 30360 52710
rect 30420 52680 30480 52710
rect 30540 52680 30600 52710
rect 19130 52590 19160 52620
rect 19250 52590 19280 52620
rect 26420 52590 26450 52620
rect 26540 52590 26570 52620
rect 30420 52590 30450 52620
rect 30540 52590 30570 52620
rect 19010 52560 19070 52590
rect 19130 52560 19190 52590
rect 19250 52560 19310 52590
rect 26300 52560 26360 52590
rect 26420 52560 26480 52590
rect 26540 52560 26600 52590
rect 30300 52560 30360 52590
rect 30420 52560 30480 52590
rect 30540 52560 30600 52590
rect 19130 52470 19160 52500
rect 19250 52470 19280 52500
rect 19880 52490 19960 52500
rect 20060 52490 20140 52500
rect 20240 52490 20320 52500
rect 20420 52490 20500 52500
rect 20600 52490 20680 52500
rect 20780 52490 20860 52500
rect 20960 52490 21040 52500
rect 21140 52490 21220 52500
rect 21320 52490 21400 52500
rect 21500 52490 21580 52500
rect 21680 52490 21760 52500
rect 21860 52490 21940 52500
rect 22040 52490 22120 52500
rect 22220 52490 22300 52500
rect 22400 52490 22480 52500
rect 22580 52490 22660 52500
rect 22760 52490 22840 52500
rect 22940 52490 23020 52500
rect 23120 52490 23200 52500
rect 23300 52490 23380 52500
rect 23480 52490 23560 52500
rect 23660 52490 23740 52500
rect 23840 52490 23920 52500
rect 24020 52490 24100 52500
rect 24200 52490 24280 52500
rect 24380 52490 24460 52500
rect 24560 52490 24640 52500
rect 24740 52490 24820 52500
rect 24920 52490 25000 52500
rect 25100 52490 25180 52500
rect 25280 52490 25360 52500
rect 25460 52490 25540 52500
rect 25640 52490 25720 52500
rect 19010 52440 19070 52470
rect 19130 52440 19190 52470
rect 19250 52440 19310 52470
rect 19960 52410 19970 52490
rect 20140 52410 20150 52490
rect 20320 52410 20330 52490
rect 20500 52410 20510 52490
rect 20680 52410 20690 52490
rect 20860 52410 20870 52490
rect 21040 52410 21050 52490
rect 21220 52410 21230 52490
rect 21400 52410 21410 52490
rect 21580 52410 21590 52490
rect 21760 52410 21770 52490
rect 21940 52410 21950 52490
rect 22120 52410 22130 52490
rect 22300 52410 22310 52490
rect 22480 52410 22490 52490
rect 22660 52410 22670 52490
rect 22840 52410 22850 52490
rect 23020 52410 23030 52490
rect 23200 52410 23210 52490
rect 23380 52410 23390 52490
rect 23560 52410 23570 52490
rect 23740 52410 23750 52490
rect 23920 52410 23930 52490
rect 24100 52410 24110 52490
rect 24280 52410 24290 52490
rect 24460 52410 24470 52490
rect 24640 52410 24650 52490
rect 24820 52410 24830 52490
rect 25000 52410 25010 52490
rect 25180 52410 25190 52490
rect 25360 52410 25370 52490
rect 25540 52410 25550 52490
rect 25720 52410 25730 52490
rect 26420 52470 26450 52500
rect 26540 52470 26570 52500
rect 30420 52470 30450 52500
rect 30540 52470 30570 52500
rect 31180 52490 31260 52500
rect 31360 52490 31440 52500
rect 31540 52490 31620 52500
rect 31720 52490 31800 52500
rect 31900 52490 31980 52500
rect 32080 52490 32160 52500
rect 32260 52490 32340 52500
rect 32440 52490 32520 52500
rect 32620 52490 32700 52500
rect 32800 52490 32880 52500
rect 32980 52490 33060 52500
rect 33160 52490 33240 52500
rect 33340 52490 33420 52500
rect 33520 52490 33600 52500
rect 33700 52490 33780 52500
rect 33880 52490 33960 52500
rect 34060 52490 34140 52500
rect 34240 52490 34320 52500
rect 34420 52490 34500 52500
rect 34600 52490 34680 52500
rect 34780 52490 34860 52500
rect 34960 52490 35040 52500
rect 35140 52490 35220 52500
rect 35320 52490 35400 52500
rect 35500 52490 35580 52500
rect 35680 52490 35760 52500
rect 35860 52490 35940 52500
rect 36040 52490 36120 52500
rect 36220 52490 36300 52500
rect 36400 52490 36480 52500
rect 36580 52490 36660 52500
rect 36760 52490 36840 52500
rect 36940 52490 37020 52500
rect 26300 52440 26360 52470
rect 26420 52440 26480 52470
rect 26540 52440 26600 52470
rect 30300 52440 30360 52470
rect 30420 52440 30480 52470
rect 30540 52440 30600 52470
rect 31260 52410 31270 52490
rect 31440 52410 31450 52490
rect 31620 52410 31630 52490
rect 31800 52410 31810 52490
rect 31980 52410 31990 52490
rect 32160 52410 32170 52490
rect 32340 52410 32350 52490
rect 32520 52410 32530 52490
rect 32700 52410 32710 52490
rect 32880 52410 32890 52490
rect 33060 52410 33070 52490
rect 33240 52410 33250 52490
rect 33420 52410 33430 52490
rect 33600 52410 33610 52490
rect 33780 52410 33790 52490
rect 33960 52410 33970 52490
rect 34140 52410 34150 52490
rect 34320 52410 34330 52490
rect 34500 52410 34510 52490
rect 34680 52410 34690 52490
rect 34860 52410 34870 52490
rect 35040 52410 35050 52490
rect 35220 52410 35230 52490
rect 35400 52410 35410 52490
rect 35580 52410 35590 52490
rect 35760 52410 35770 52490
rect 35940 52410 35950 52490
rect 36120 52410 36130 52490
rect 36300 52410 36310 52490
rect 36480 52410 36490 52490
rect 36660 52410 36670 52490
rect 36840 52410 36850 52490
rect 37020 52410 37030 52490
rect 19130 52350 19160 52380
rect 19250 52350 19280 52380
rect 26420 52350 26450 52380
rect 26540 52350 26570 52380
rect 30420 52350 30450 52380
rect 30540 52350 30570 52380
rect 19010 52320 19070 52350
rect 19130 52320 19190 52350
rect 19250 52320 19310 52350
rect 26300 52320 26360 52350
rect 26420 52320 26480 52350
rect 26540 52320 26600 52350
rect 30300 52320 30360 52350
rect 30420 52320 30480 52350
rect 30540 52320 30600 52350
rect 37100 52320 37190 52990
rect 37720 52950 37750 52980
rect 37840 52950 37870 52980
rect 42595 52975 42675 52985
rect 37600 52920 37660 52950
rect 37720 52920 37780 52950
rect 37840 52920 37900 52950
rect 42675 52905 42685 52975
rect 146100 52950 146160 52980
rect 147580 52950 147640 52980
rect 148400 52950 148460 52980
rect 149880 52950 149940 52980
rect 152220 52930 152250 52960
rect 152340 52930 152370 52960
rect 40060 52870 40120 52900
rect 41540 52870 41600 52900
rect 42360 52870 42420 52900
rect 42595 52895 42685 52905
rect 152100 52900 152160 52930
rect 152220 52900 152280 52930
rect 152340 52900 152400 52930
rect 43840 52870 43900 52900
rect 37720 52830 37750 52860
rect 37840 52830 37870 52860
rect 37600 52800 37660 52830
rect 37720 52800 37780 52830
rect 37840 52800 37900 52830
rect 42595 52815 42675 52825
rect 40060 52750 40120 52780
rect 41540 52750 41600 52780
rect 42360 52750 42420 52780
rect 37720 52710 37750 52740
rect 37840 52710 37870 52740
rect 42675 52735 42685 52815
rect 43030 52800 43390 52860
rect 146100 52830 146160 52860
rect 147580 52830 147640 52860
rect 148400 52830 148460 52860
rect 149880 52830 149940 52860
rect 152220 52810 152250 52840
rect 152340 52810 152370 52840
rect 152980 52810 153060 52820
rect 153160 52810 153240 52820
rect 153340 52810 153420 52820
rect 153520 52810 153600 52820
rect 153700 52810 153780 52820
rect 153880 52810 153960 52820
rect 154060 52810 154140 52820
rect 154240 52810 154320 52820
rect 154420 52810 154500 52820
rect 154600 52810 154680 52820
rect 154780 52810 154860 52820
rect 154960 52810 155040 52820
rect 155140 52810 155220 52820
rect 155320 52810 155400 52820
rect 155500 52810 155580 52820
rect 155680 52810 155760 52820
rect 155860 52810 155940 52820
rect 156040 52810 156120 52820
rect 156220 52810 156300 52820
rect 156400 52810 156480 52820
rect 156580 52810 156660 52820
rect 156760 52810 156840 52820
rect 156940 52810 157020 52820
rect 157120 52810 157200 52820
rect 157300 52810 157380 52820
rect 157480 52810 157560 52820
rect 157660 52810 157740 52820
rect 157840 52810 157920 52820
rect 158020 52810 158100 52820
rect 158200 52810 158280 52820
rect 158380 52810 158460 52820
rect 158560 52810 158640 52820
rect 158740 52810 158820 52820
rect 152100 52780 152160 52810
rect 152220 52780 152280 52810
rect 152340 52780 152400 52810
rect 43840 52750 43900 52780
rect 38595 52715 38675 52725
rect 38775 52715 38855 52725
rect 38955 52715 39035 52725
rect 39135 52715 39215 52725
rect 39315 52715 39395 52725
rect 37600 52680 37660 52710
rect 37720 52680 37780 52710
rect 37840 52680 37900 52710
rect 38675 52635 38685 52715
rect 38855 52635 38865 52715
rect 39035 52635 39045 52715
rect 39215 52635 39225 52715
rect 39395 52635 39405 52715
rect 43580 52670 43700 52730
rect 146100 52710 146160 52740
rect 147580 52710 147640 52740
rect 148400 52710 148460 52740
rect 149880 52710 149940 52740
rect 153060 52730 153070 52810
rect 153240 52730 153250 52810
rect 153420 52730 153430 52810
rect 153600 52730 153610 52810
rect 153780 52730 153790 52810
rect 153960 52730 153970 52810
rect 154140 52730 154150 52810
rect 154320 52730 154330 52810
rect 154500 52730 154510 52810
rect 154680 52730 154690 52810
rect 154860 52730 154870 52810
rect 155040 52730 155050 52810
rect 155220 52730 155230 52810
rect 155400 52730 155410 52810
rect 155580 52730 155590 52810
rect 155760 52730 155770 52810
rect 155940 52730 155950 52810
rect 156120 52730 156130 52810
rect 156300 52730 156310 52810
rect 156480 52730 156490 52810
rect 156660 52730 156670 52810
rect 156840 52730 156850 52810
rect 157020 52730 157030 52810
rect 157200 52730 157210 52810
rect 157380 52730 157390 52810
rect 157560 52730 157570 52810
rect 157740 52730 157750 52810
rect 157920 52730 157930 52810
rect 158100 52730 158110 52810
rect 158280 52730 158290 52810
rect 158460 52730 158470 52810
rect 158640 52730 158650 52810
rect 158820 52730 158830 52810
rect 152220 52690 152250 52720
rect 152340 52690 152370 52720
rect 40060 52630 40120 52660
rect 41540 52630 41600 52660
rect 42360 52630 42420 52660
rect 42950 52650 43560 52660
rect 43550 52645 43560 52650
rect 42910 52635 43560 52645
rect 37720 52590 37750 52620
rect 37840 52590 37870 52620
rect 37600 52560 37660 52590
rect 37720 52560 37780 52590
rect 37840 52560 37900 52590
rect 42900 52585 42910 52635
rect 38595 52535 38675 52545
rect 38775 52535 38855 52545
rect 38955 52535 39035 52545
rect 39135 52535 39215 52545
rect 39315 52535 39395 52545
rect 43030 52540 43390 52600
rect 37720 52470 37750 52500
rect 37840 52470 37870 52500
rect 37600 52440 37660 52470
rect 37720 52440 37780 52470
rect 37840 52440 37900 52470
rect 38675 52455 38685 52535
rect 38855 52455 38865 52535
rect 39035 52455 39045 52535
rect 39215 52455 39225 52535
rect 39395 52455 39405 52535
rect 40060 52510 40120 52540
rect 41540 52510 41600 52540
rect 42360 52510 42420 52540
rect 42682 52460 42822 52530
rect 40060 52390 40120 52420
rect 40678 52399 40758 52409
rect 40838 52399 40918 52409
rect 37720 52350 37750 52380
rect 37840 52350 37870 52380
rect 38595 52355 38675 52365
rect 38775 52355 38855 52365
rect 38955 52355 39035 52365
rect 39135 52355 39215 52365
rect 39315 52355 39395 52365
rect 37600 52320 37660 52350
rect 37720 52320 37780 52350
rect 37840 52320 37900 52350
rect 19800 52310 25800 52320
rect 31100 52310 37190 52320
rect 19130 52230 19160 52260
rect 19250 52230 19280 52260
rect 26420 52230 26450 52260
rect 26540 52230 26570 52260
rect 30420 52230 30450 52260
rect 30540 52230 30570 52260
rect 19010 52200 19070 52230
rect 19130 52200 19190 52230
rect 19250 52200 19310 52230
rect 26300 52200 26360 52230
rect 26420 52200 26480 52230
rect 26540 52200 26600 52230
rect 30300 52200 30360 52230
rect 30420 52200 30480 52230
rect 30540 52200 30600 52230
rect 37100 52210 37190 52310
rect 38675 52275 38685 52355
rect 38855 52275 38865 52355
rect 39035 52275 39045 52355
rect 39215 52275 39225 52355
rect 39395 52275 39405 52355
rect 40758 52319 40768 52399
rect 40838 52319 40848 52399
rect 40918 52319 40928 52399
rect 41540 52390 41600 52420
rect 42360 52390 42420 52420
rect 42822 52400 42892 52460
rect 42822 52390 43470 52400
rect 43550 52390 43560 52635
rect 43700 52550 43760 52670
rect 152100 52660 152160 52690
rect 152220 52660 152280 52690
rect 152340 52660 152400 52690
rect 43840 52630 43900 52660
rect 146100 52590 146160 52620
rect 147580 52590 147640 52620
rect 148400 52590 148460 52620
rect 149880 52590 149940 52620
rect 152220 52570 152250 52600
rect 152340 52570 152370 52600
rect 152100 52540 152160 52570
rect 152220 52540 152280 52570
rect 152340 52540 152400 52570
rect 43840 52510 43900 52540
rect 146100 52470 146160 52500
rect 147580 52470 147640 52500
rect 148400 52470 148460 52500
rect 149880 52470 149940 52500
rect 152980 52490 153060 52500
rect 153160 52490 153240 52500
rect 153340 52490 153420 52500
rect 153520 52490 153600 52500
rect 153700 52490 153780 52500
rect 153880 52490 153960 52500
rect 154060 52490 154140 52500
rect 154240 52490 154320 52500
rect 154420 52490 154500 52500
rect 154600 52490 154680 52500
rect 154780 52490 154860 52500
rect 154960 52490 155040 52500
rect 155140 52490 155220 52500
rect 155320 52490 155400 52500
rect 155500 52490 155580 52500
rect 155680 52490 155760 52500
rect 155860 52490 155940 52500
rect 156040 52490 156120 52500
rect 156220 52490 156300 52500
rect 156400 52490 156480 52500
rect 156580 52490 156660 52500
rect 156760 52490 156840 52500
rect 156940 52490 157020 52500
rect 157120 52490 157200 52500
rect 157300 52490 157380 52500
rect 157480 52490 157560 52500
rect 157660 52490 157740 52500
rect 157840 52490 157920 52500
rect 158020 52490 158100 52500
rect 158200 52490 158280 52500
rect 158380 52490 158460 52500
rect 158560 52490 158640 52500
rect 158740 52490 158820 52500
rect 43580 52410 43700 52470
rect 152220 52450 152250 52480
rect 152340 52450 152370 52480
rect 152100 52420 152160 52450
rect 152220 52420 152280 52450
rect 152340 52420 152400 52450
rect 42822 52320 42892 52390
rect 42910 52375 43560 52385
rect 42900 52325 42910 52375
rect 40060 52270 40120 52300
rect 37720 52230 37750 52260
rect 37840 52230 37870 52260
rect 40685 52250 40925 52280
rect 41540 52270 41600 52300
rect 42360 52270 42420 52300
rect 42682 52260 42822 52320
rect 43030 52280 43390 52340
rect 43700 52290 43760 52410
rect 43840 52390 43900 52420
rect 153060 52410 153070 52490
rect 153240 52410 153250 52490
rect 153420 52410 153430 52490
rect 153600 52410 153610 52490
rect 153780 52410 153790 52490
rect 153960 52410 153970 52490
rect 154140 52410 154150 52490
rect 154320 52410 154330 52490
rect 154500 52410 154510 52490
rect 154680 52410 154690 52490
rect 154860 52410 154870 52490
rect 155040 52410 155050 52490
rect 155220 52410 155230 52490
rect 155400 52410 155410 52490
rect 155580 52410 155590 52490
rect 155760 52410 155770 52490
rect 155940 52410 155950 52490
rect 156120 52410 156130 52490
rect 156300 52410 156310 52490
rect 156480 52410 156490 52490
rect 156660 52410 156670 52490
rect 156840 52410 156850 52490
rect 157020 52410 157030 52490
rect 157200 52410 157210 52490
rect 157380 52410 157390 52490
rect 157560 52410 157570 52490
rect 157740 52410 157750 52490
rect 157920 52410 157930 52490
rect 158100 52410 158110 52490
rect 158280 52410 158290 52490
rect 158460 52410 158470 52490
rect 158640 52410 158650 52490
rect 158820 52410 158830 52490
rect 146100 52350 146160 52380
rect 147580 52350 147640 52380
rect 148400 52350 148460 52380
rect 149880 52350 149940 52380
rect 152220 52330 152250 52360
rect 152340 52330 152370 52360
rect 152100 52300 152160 52330
rect 152220 52300 152280 52330
rect 152340 52300 152400 52330
rect 158900 52320 158990 52990
rect 159520 52930 159550 52960
rect 159640 52930 159670 52960
rect 163520 52930 163550 52960
rect 163640 52930 163670 52960
rect 170810 52930 170840 52960
rect 170930 52930 170960 52960
rect 159400 52900 159460 52930
rect 159520 52900 159580 52930
rect 159640 52900 159700 52930
rect 163400 52900 163460 52930
rect 163520 52900 163580 52930
rect 163640 52900 163700 52930
rect 170690 52900 170750 52930
rect 170810 52900 170870 52930
rect 170930 52900 170990 52930
rect 159520 52810 159550 52840
rect 159640 52810 159670 52840
rect 163520 52810 163550 52840
rect 163640 52810 163670 52840
rect 164280 52810 164360 52820
rect 164460 52810 164540 52820
rect 164640 52810 164720 52820
rect 164820 52810 164900 52820
rect 165000 52810 165080 52820
rect 165180 52810 165260 52820
rect 165360 52810 165440 52820
rect 165540 52810 165620 52820
rect 165720 52810 165800 52820
rect 165900 52810 165980 52820
rect 166080 52810 166160 52820
rect 166260 52810 166340 52820
rect 166440 52810 166520 52820
rect 166620 52810 166700 52820
rect 166800 52810 166880 52820
rect 166980 52810 167060 52820
rect 167160 52810 167240 52820
rect 167340 52810 167420 52820
rect 167520 52810 167600 52820
rect 167700 52810 167780 52820
rect 167880 52810 167960 52820
rect 168060 52810 168140 52820
rect 168240 52810 168320 52820
rect 168420 52810 168500 52820
rect 168600 52810 168680 52820
rect 168780 52810 168860 52820
rect 168960 52810 169040 52820
rect 169140 52810 169220 52820
rect 169320 52810 169400 52820
rect 169500 52810 169580 52820
rect 169680 52810 169760 52820
rect 169860 52810 169940 52820
rect 170040 52810 170120 52820
rect 170810 52810 170840 52840
rect 170930 52810 170960 52840
rect 159400 52780 159460 52810
rect 159520 52780 159580 52810
rect 159640 52780 159700 52810
rect 163400 52780 163460 52810
rect 163520 52780 163580 52810
rect 163640 52780 163700 52810
rect 164360 52730 164370 52810
rect 164540 52730 164550 52810
rect 164720 52730 164730 52810
rect 164900 52730 164910 52810
rect 165080 52730 165090 52810
rect 165260 52730 165270 52810
rect 165440 52730 165450 52810
rect 165620 52730 165630 52810
rect 165800 52730 165810 52810
rect 165980 52730 165990 52810
rect 166160 52730 166170 52810
rect 166340 52730 166350 52810
rect 166520 52730 166530 52810
rect 166700 52730 166710 52810
rect 166880 52730 166890 52810
rect 167060 52730 167070 52810
rect 167240 52730 167250 52810
rect 167420 52730 167430 52810
rect 167600 52730 167610 52810
rect 167780 52730 167790 52810
rect 167960 52730 167970 52810
rect 168140 52730 168150 52810
rect 168320 52730 168330 52810
rect 168500 52730 168510 52810
rect 168680 52730 168690 52810
rect 168860 52730 168870 52810
rect 169040 52730 169050 52810
rect 169220 52730 169230 52810
rect 169400 52730 169410 52810
rect 169580 52730 169590 52810
rect 169760 52730 169770 52810
rect 169940 52730 169950 52810
rect 170120 52730 170130 52810
rect 170690 52780 170750 52810
rect 170810 52780 170870 52810
rect 170930 52780 170990 52810
rect 159520 52690 159550 52720
rect 159640 52690 159670 52720
rect 163520 52690 163550 52720
rect 163640 52690 163670 52720
rect 170810 52690 170840 52720
rect 170930 52690 170960 52720
rect 159400 52660 159460 52690
rect 159520 52660 159580 52690
rect 159640 52660 159700 52690
rect 163400 52660 163460 52690
rect 163520 52660 163580 52690
rect 163640 52660 163700 52690
rect 170690 52660 170750 52690
rect 170810 52660 170870 52690
rect 170930 52660 170990 52690
rect 159520 52570 159550 52600
rect 159640 52570 159670 52600
rect 163520 52570 163550 52600
rect 163640 52570 163670 52600
rect 170810 52570 170840 52600
rect 170930 52570 170960 52600
rect 159400 52540 159460 52570
rect 159520 52540 159580 52570
rect 159640 52540 159700 52570
rect 163400 52540 163460 52570
rect 163520 52540 163580 52570
rect 163640 52540 163700 52570
rect 170690 52540 170750 52570
rect 170810 52540 170870 52570
rect 170930 52540 170990 52570
rect 164280 52510 164360 52520
rect 164460 52510 164540 52520
rect 164640 52510 164720 52520
rect 164820 52510 164900 52520
rect 165000 52510 165080 52520
rect 165180 52510 165260 52520
rect 165360 52510 165440 52520
rect 165540 52510 165620 52520
rect 165720 52510 165800 52520
rect 165900 52510 165980 52520
rect 166080 52510 166160 52520
rect 166260 52510 166340 52520
rect 166440 52510 166520 52520
rect 166620 52510 166700 52520
rect 166800 52510 166880 52520
rect 166980 52510 167060 52520
rect 167160 52510 167240 52520
rect 167340 52510 167420 52520
rect 167520 52510 167600 52520
rect 167700 52510 167780 52520
rect 167880 52510 167960 52520
rect 168060 52510 168140 52520
rect 168240 52510 168320 52520
rect 168420 52510 168500 52520
rect 168600 52510 168680 52520
rect 168780 52510 168860 52520
rect 168960 52510 169040 52520
rect 169140 52510 169220 52520
rect 169320 52510 169400 52520
rect 169500 52510 169580 52520
rect 169680 52510 169760 52520
rect 169860 52510 169940 52520
rect 170040 52510 170120 52520
rect 159520 52450 159550 52480
rect 159640 52450 159670 52480
rect 163520 52450 163550 52480
rect 163640 52450 163670 52480
rect 159400 52420 159460 52450
rect 159520 52420 159580 52450
rect 159640 52420 159700 52450
rect 163400 52420 163460 52450
rect 163520 52420 163580 52450
rect 163640 52420 163700 52450
rect 164360 52430 164370 52510
rect 164540 52430 164550 52510
rect 164720 52430 164730 52510
rect 164900 52430 164910 52510
rect 165080 52430 165090 52510
rect 165260 52430 165270 52510
rect 165440 52430 165450 52510
rect 165620 52430 165630 52510
rect 165800 52430 165810 52510
rect 165980 52430 165990 52510
rect 166160 52430 166170 52510
rect 166340 52430 166350 52510
rect 166520 52430 166530 52510
rect 166700 52430 166710 52510
rect 166880 52430 166890 52510
rect 167060 52430 167070 52510
rect 167240 52430 167250 52510
rect 167420 52430 167430 52510
rect 167600 52430 167610 52510
rect 167780 52430 167790 52510
rect 167960 52430 167970 52510
rect 168140 52430 168150 52510
rect 168320 52430 168330 52510
rect 168500 52430 168510 52510
rect 168680 52430 168690 52510
rect 168860 52430 168870 52510
rect 169040 52430 169050 52510
rect 169220 52430 169230 52510
rect 169400 52430 169410 52510
rect 169580 52430 169590 52510
rect 169760 52430 169770 52510
rect 169940 52430 169950 52510
rect 170120 52430 170130 52510
rect 170810 52450 170840 52480
rect 170930 52450 170960 52480
rect 170690 52420 170750 52450
rect 170810 52420 170870 52450
rect 170930 52420 170990 52450
rect 159520 52330 159550 52360
rect 159640 52330 159670 52360
rect 163520 52330 163550 52360
rect 163640 52330 163670 52360
rect 170810 52330 170840 52360
rect 170930 52330 170960 52360
rect 152900 52310 158990 52320
rect 43840 52270 43900 52300
rect 31100 52180 37190 52210
rect 37600 52200 37660 52230
rect 37720 52200 37780 52230
rect 37840 52200 37900 52230
rect 40685 52190 40715 52250
rect 40775 52190 40865 52250
rect 40895 52190 40925 52250
rect 19880 52170 19960 52180
rect 20060 52170 20140 52180
rect 20240 52170 20320 52180
rect 20420 52170 20500 52180
rect 20600 52170 20680 52180
rect 20780 52170 20860 52180
rect 20960 52170 21040 52180
rect 21140 52170 21220 52180
rect 21320 52170 21400 52180
rect 21500 52170 21580 52180
rect 21680 52170 21760 52180
rect 21860 52170 21940 52180
rect 22040 52170 22120 52180
rect 22220 52170 22300 52180
rect 22400 52170 22480 52180
rect 22580 52170 22660 52180
rect 22760 52170 22840 52180
rect 22940 52170 23020 52180
rect 23120 52170 23200 52180
rect 23300 52170 23380 52180
rect 23480 52170 23560 52180
rect 23660 52170 23740 52180
rect 23840 52170 23920 52180
rect 24020 52170 24100 52180
rect 24200 52170 24280 52180
rect 24380 52170 24460 52180
rect 24560 52170 24640 52180
rect 24740 52170 24820 52180
rect 24920 52170 25000 52180
rect 25100 52170 25180 52180
rect 25280 52170 25360 52180
rect 25460 52170 25540 52180
rect 25640 52170 25720 52180
rect 31180 52170 31260 52180
rect 31360 52170 31440 52180
rect 31540 52170 31620 52180
rect 31720 52170 31800 52180
rect 31900 52170 31980 52180
rect 32080 52170 32160 52180
rect 32260 52170 32340 52180
rect 32440 52170 32520 52180
rect 32620 52170 32700 52180
rect 32800 52170 32880 52180
rect 32980 52170 33060 52180
rect 33160 52170 33240 52180
rect 33340 52170 33420 52180
rect 33520 52170 33600 52180
rect 33700 52170 33780 52180
rect 33880 52170 33960 52180
rect 34060 52170 34140 52180
rect 34240 52170 34320 52180
rect 34420 52170 34500 52180
rect 34600 52170 34680 52180
rect 34780 52170 34860 52180
rect 34960 52170 35040 52180
rect 35140 52170 35220 52180
rect 35320 52170 35400 52180
rect 35500 52170 35580 52180
rect 35680 52170 35760 52180
rect 35860 52170 35940 52180
rect 36040 52170 36120 52180
rect 36220 52170 36300 52180
rect 36400 52170 36480 52180
rect 36580 52170 36660 52180
rect 36760 52170 36840 52180
rect 36940 52170 37020 52180
rect 19130 52110 19160 52140
rect 19250 52110 19280 52140
rect 19010 52080 19070 52110
rect 19130 52080 19190 52110
rect 19250 52080 19310 52110
rect 19960 52090 19970 52170
rect 20140 52090 20150 52170
rect 20320 52090 20330 52170
rect 20500 52090 20510 52170
rect 20680 52090 20690 52170
rect 20860 52090 20870 52170
rect 21040 52090 21050 52170
rect 21220 52090 21230 52170
rect 21400 52090 21410 52170
rect 21580 52090 21590 52170
rect 21760 52090 21770 52170
rect 21940 52090 21950 52170
rect 22120 52090 22130 52170
rect 22300 52090 22310 52170
rect 22480 52090 22490 52170
rect 22660 52090 22670 52170
rect 22840 52090 22850 52170
rect 23020 52090 23030 52170
rect 23200 52090 23210 52170
rect 23380 52090 23390 52170
rect 23560 52090 23570 52170
rect 23740 52090 23750 52170
rect 23920 52090 23930 52170
rect 24100 52090 24110 52170
rect 24280 52090 24290 52170
rect 24460 52090 24470 52170
rect 24640 52090 24650 52170
rect 24820 52090 24830 52170
rect 25000 52090 25010 52170
rect 25180 52090 25190 52170
rect 25360 52090 25370 52170
rect 25540 52090 25550 52170
rect 25720 52090 25730 52170
rect 26420 52110 26450 52140
rect 26540 52110 26570 52140
rect 30420 52110 30450 52140
rect 30540 52110 30570 52140
rect 31260 52110 31270 52170
rect 31440 52110 31450 52170
rect 31620 52110 31630 52170
rect 31800 52110 31810 52170
rect 31980 52110 31990 52170
rect 32160 52110 32170 52170
rect 32340 52110 32350 52170
rect 32520 52110 32530 52170
rect 32700 52110 32710 52170
rect 32880 52110 32890 52170
rect 33060 52110 33070 52170
rect 33240 52110 33250 52170
rect 33420 52110 33430 52170
rect 33600 52110 33610 52170
rect 33780 52110 33790 52170
rect 33960 52110 33970 52170
rect 34140 52110 34150 52170
rect 34320 52110 34330 52170
rect 34500 52110 34510 52170
rect 34680 52110 34690 52170
rect 34860 52110 34870 52170
rect 35040 52110 35050 52170
rect 35220 52110 35230 52170
rect 35400 52110 35410 52170
rect 35580 52110 35590 52170
rect 35760 52110 35770 52170
rect 35940 52110 35950 52170
rect 36120 52110 36130 52170
rect 36300 52110 36310 52170
rect 36480 52110 36490 52170
rect 36660 52110 36670 52170
rect 36840 52110 36850 52170
rect 37020 52110 37030 52170
rect 37100 52110 37190 52180
rect 38595 52175 38675 52185
rect 38775 52175 38855 52185
rect 38955 52175 39035 52185
rect 39135 52175 39215 52185
rect 39315 52175 39395 52185
rect 37720 52110 37750 52140
rect 37840 52110 37870 52140
rect 26300 52080 26360 52110
rect 26420 52080 26480 52110
rect 26540 52080 26600 52110
rect 30300 52080 30360 52110
rect 30420 52080 30480 52110
rect 30540 52080 30600 52110
rect 31100 52080 37190 52110
rect 37600 52080 37660 52110
rect 37720 52080 37780 52110
rect 37840 52080 37900 52110
rect 38675 52095 38685 52175
rect 38855 52095 38865 52175
rect 39035 52095 39045 52175
rect 39215 52095 39225 52175
rect 39395 52095 39405 52175
rect 40060 52150 40120 52180
rect 40685 52160 40925 52190
rect 41540 52150 41600 52180
rect 42360 52150 42420 52180
rect 40678 52129 40758 52139
rect 40838 52129 40918 52139
rect 19880 52020 19960 52030
rect 20060 52020 20140 52030
rect 20240 52020 20320 52030
rect 20420 52020 20500 52030
rect 20600 52020 20680 52030
rect 20780 52020 20860 52030
rect 20960 52020 21040 52030
rect 21140 52020 21220 52030
rect 21320 52020 21400 52030
rect 21500 52020 21580 52030
rect 21680 52020 21760 52030
rect 21860 52020 21940 52030
rect 22040 52020 22120 52030
rect 22220 52020 22300 52030
rect 22400 52020 22480 52030
rect 22580 52020 22660 52030
rect 22760 52020 22840 52030
rect 22940 52020 23020 52030
rect 23120 52020 23200 52030
rect 23300 52020 23380 52030
rect 23480 52020 23560 52030
rect 23660 52020 23740 52030
rect 23840 52020 23920 52030
rect 24020 52020 24100 52030
rect 24200 52020 24280 52030
rect 24380 52020 24460 52030
rect 24560 52020 24640 52030
rect 24740 52020 24820 52030
rect 24920 52020 25000 52030
rect 25100 52020 25180 52030
rect 25280 52020 25360 52030
rect 25460 52020 25540 52030
rect 25640 52020 25720 52030
rect 31180 52020 31260 52030
rect 31360 52020 31440 52030
rect 31540 52020 31620 52030
rect 31720 52020 31800 52030
rect 31900 52020 31980 52030
rect 32080 52020 32160 52030
rect 32260 52020 32340 52030
rect 32440 52020 32520 52030
rect 32620 52020 32700 52030
rect 32800 52020 32880 52030
rect 32980 52020 33060 52030
rect 33160 52020 33240 52030
rect 33340 52020 33420 52030
rect 33520 52020 33600 52030
rect 33700 52020 33780 52030
rect 33880 52020 33960 52030
rect 34060 52020 34140 52030
rect 34240 52020 34320 52030
rect 34420 52020 34500 52030
rect 34600 52020 34680 52030
rect 34780 52020 34860 52030
rect 34960 52020 35040 52030
rect 35140 52020 35220 52030
rect 35320 52020 35400 52030
rect 35500 52020 35580 52030
rect 35680 52020 35760 52030
rect 35860 52020 35940 52030
rect 36040 52020 36120 52030
rect 36220 52020 36300 52030
rect 36400 52020 36480 52030
rect 36580 52020 36660 52030
rect 36760 52020 36840 52030
rect 36940 52020 37020 52030
rect 19130 51990 19160 52020
rect 19250 51990 19280 52020
rect 19010 51960 19070 51990
rect 19130 51960 19190 51990
rect 19250 51960 19310 51990
rect 19960 51940 19970 52020
rect 20140 51940 20150 52020
rect 20320 51940 20330 52020
rect 20500 51940 20510 52020
rect 20680 51940 20690 52020
rect 20860 51940 20870 52020
rect 21040 51940 21050 52020
rect 21220 51940 21230 52020
rect 21400 51940 21410 52020
rect 21580 51940 21590 52020
rect 21760 51940 21770 52020
rect 21940 51940 21950 52020
rect 22120 51940 22130 52020
rect 22300 51940 22310 52020
rect 22480 51940 22490 52020
rect 22660 51940 22670 52020
rect 22840 51940 22850 52020
rect 23020 51940 23030 52020
rect 23200 51940 23210 52020
rect 23380 51940 23390 52020
rect 23560 51940 23570 52020
rect 23740 51940 23750 52020
rect 23920 51940 23930 52020
rect 24100 51940 24110 52020
rect 24280 51940 24290 52020
rect 24460 51940 24470 52020
rect 24640 51940 24650 52020
rect 24820 51940 24830 52020
rect 25000 51940 25010 52020
rect 25180 51940 25190 52020
rect 25360 51940 25370 52020
rect 25540 51940 25550 52020
rect 25720 51940 25730 52020
rect 26420 51990 26450 52020
rect 26540 51990 26570 52020
rect 30420 51990 30450 52020
rect 30540 51990 30570 52020
rect 26300 51960 26360 51990
rect 26420 51960 26480 51990
rect 26540 51960 26600 51990
rect 30300 51960 30360 51990
rect 30420 51960 30480 51990
rect 30540 51960 30600 51990
rect 31260 51940 31270 52020
rect 31440 51940 31450 52020
rect 31620 51940 31630 52020
rect 31800 51940 31810 52020
rect 31980 51940 31990 52020
rect 32160 51940 32170 52020
rect 32340 51940 32350 52020
rect 32520 51940 32530 52020
rect 32700 51940 32710 52020
rect 32880 51940 32890 52020
rect 33060 51940 33070 52020
rect 33240 51940 33250 52020
rect 33420 51940 33430 52020
rect 33600 51940 33610 52020
rect 33780 51940 33790 52020
rect 33960 51940 33970 52020
rect 34140 51940 34150 52020
rect 34320 51940 34330 52020
rect 34500 51940 34510 52020
rect 34680 51940 34690 52020
rect 34860 51940 34870 52020
rect 35040 51940 35050 52020
rect 35220 51940 35230 52020
rect 35400 51940 35410 52020
rect 35580 51940 35590 52020
rect 35760 51940 35770 52020
rect 35940 51940 35950 52020
rect 36120 51940 36130 52020
rect 36300 51940 36310 52020
rect 36480 51940 36490 52020
rect 36660 51940 36670 52020
rect 36840 51940 36850 52020
rect 37020 51940 37030 52020
rect 19130 51870 19160 51900
rect 19250 51870 19280 51900
rect 19880 51870 19960 51880
rect 20060 51870 20140 51880
rect 20240 51870 20320 51880
rect 20420 51870 20500 51880
rect 20600 51870 20680 51880
rect 20780 51870 20860 51880
rect 20960 51870 21040 51880
rect 21140 51870 21220 51880
rect 21320 51870 21400 51880
rect 21500 51870 21580 51880
rect 21680 51870 21760 51880
rect 21860 51870 21940 51880
rect 22040 51870 22120 51880
rect 22220 51870 22300 51880
rect 22400 51870 22480 51880
rect 22580 51870 22660 51880
rect 22760 51870 22840 51880
rect 22940 51870 23020 51880
rect 23120 51870 23200 51880
rect 23300 51870 23380 51880
rect 23480 51870 23560 51880
rect 23660 51870 23740 51880
rect 23840 51870 23920 51880
rect 24020 51870 24100 51880
rect 24200 51870 24280 51880
rect 24380 51870 24460 51880
rect 24560 51870 24640 51880
rect 24740 51870 24820 51880
rect 24920 51870 25000 51880
rect 25100 51870 25180 51880
rect 25280 51870 25360 51880
rect 25460 51870 25540 51880
rect 25640 51870 25720 51880
rect 26420 51870 26450 51900
rect 26540 51870 26570 51900
rect 30420 51870 30450 51900
rect 30540 51870 30570 51900
rect 37100 51880 37190 52080
rect 40060 52030 40120 52060
rect 40758 52049 40768 52129
rect 40838 52049 40848 52129
rect 40918 52049 40928 52129
rect 42822 52120 42892 52260
rect 146100 52230 146160 52260
rect 147580 52230 147640 52260
rect 148400 52230 148460 52260
rect 149880 52230 149940 52260
rect 152220 52210 152250 52240
rect 152340 52210 152370 52240
rect 158900 52210 158990 52310
rect 159400 52300 159460 52330
rect 159520 52300 159580 52330
rect 159640 52300 159700 52330
rect 163400 52300 163460 52330
rect 163520 52300 163580 52330
rect 163640 52300 163700 52330
rect 164200 52310 170200 52320
rect 170690 52300 170750 52330
rect 170810 52300 170870 52330
rect 170930 52300 170990 52330
rect 159520 52210 159550 52240
rect 159640 52210 159670 52240
rect 163520 52210 163550 52240
rect 163640 52210 163670 52240
rect 170810 52210 170840 52240
rect 170930 52210 170960 52240
rect 43580 52150 43700 52210
rect 152100 52180 152160 52210
rect 152220 52180 152280 52210
rect 152340 52180 152400 52210
rect 152900 52180 158990 52210
rect 159400 52180 159460 52210
rect 159520 52180 159580 52210
rect 159640 52180 159700 52210
rect 163400 52180 163460 52210
rect 163520 52180 163580 52210
rect 163640 52180 163700 52210
rect 170690 52180 170750 52210
rect 170810 52180 170870 52210
rect 170930 52180 170990 52210
rect 43840 52150 43900 52180
rect 152980 52170 153060 52180
rect 153160 52170 153240 52180
rect 153340 52170 153420 52180
rect 153520 52170 153600 52180
rect 153700 52170 153780 52180
rect 153880 52170 153960 52180
rect 154060 52170 154140 52180
rect 154240 52170 154320 52180
rect 154420 52170 154500 52180
rect 154600 52170 154680 52180
rect 154780 52170 154860 52180
rect 154960 52170 155040 52180
rect 155140 52170 155220 52180
rect 155320 52170 155400 52180
rect 155500 52170 155580 52180
rect 155680 52170 155760 52180
rect 155860 52170 155940 52180
rect 156040 52170 156120 52180
rect 156220 52170 156300 52180
rect 156400 52170 156480 52180
rect 156580 52170 156660 52180
rect 156760 52170 156840 52180
rect 156940 52170 157020 52180
rect 157120 52170 157200 52180
rect 157300 52170 157380 52180
rect 157480 52170 157560 52180
rect 157660 52170 157740 52180
rect 157840 52170 157920 52180
rect 158020 52170 158100 52180
rect 158200 52170 158280 52180
rect 158380 52170 158460 52180
rect 158560 52170 158640 52180
rect 158740 52170 158820 52180
rect 42950 52130 43560 52140
rect 43550 52125 43560 52130
rect 42682 52060 42822 52120
rect 42910 52115 43560 52125
rect 42900 52065 42910 52115
rect 41540 52030 41600 52060
rect 42360 52030 42420 52060
rect 37720 51990 37750 52020
rect 37840 51990 37870 52020
rect 38595 51995 38675 52005
rect 38775 51995 38855 52005
rect 38955 51995 39035 52005
rect 39135 51995 39215 52005
rect 39315 51995 39395 52005
rect 37600 51960 37660 51990
rect 37720 51960 37780 51990
rect 37840 51960 37900 51990
rect 38675 51915 38685 51995
rect 38855 51915 38865 51995
rect 39035 51915 39045 51995
rect 39215 51915 39225 51995
rect 39395 51915 39405 51995
rect 40060 51910 40120 51940
rect 41540 51910 41600 51940
rect 42360 51910 42420 51940
rect 42822 51920 42892 52060
rect 43030 52020 43390 52080
rect 19010 51840 19070 51870
rect 19130 51840 19190 51870
rect 19250 51840 19310 51870
rect 19960 51790 19970 51870
rect 20140 51790 20150 51870
rect 20320 51790 20330 51870
rect 20500 51790 20510 51870
rect 20680 51790 20690 51870
rect 20860 51790 20870 51870
rect 21040 51790 21050 51870
rect 21220 51790 21230 51870
rect 21400 51790 21410 51870
rect 21580 51790 21590 51870
rect 21760 51790 21770 51870
rect 21940 51790 21950 51870
rect 22120 51790 22130 51870
rect 22300 51790 22310 51870
rect 22480 51790 22490 51870
rect 22660 51790 22670 51870
rect 22840 51790 22850 51870
rect 23020 51790 23030 51870
rect 23200 51790 23210 51870
rect 23380 51790 23390 51870
rect 23560 51790 23570 51870
rect 23740 51790 23750 51870
rect 23920 51790 23930 51870
rect 24100 51790 24110 51870
rect 24280 51790 24290 51870
rect 24460 51790 24470 51870
rect 24640 51790 24650 51870
rect 24820 51790 24830 51870
rect 25000 51790 25010 51870
rect 25180 51790 25190 51870
rect 25360 51790 25370 51870
rect 25540 51790 25550 51870
rect 25720 51790 25730 51870
rect 26300 51840 26360 51870
rect 26420 51840 26480 51870
rect 26540 51840 26600 51870
rect 30300 51840 30360 51870
rect 30420 51840 30480 51870
rect 30540 51840 30600 51870
rect 31100 51850 37190 51880
rect 37720 51870 37750 51900
rect 37840 51870 37870 51900
rect 31260 51790 31270 51850
rect 31440 51790 31450 51850
rect 31620 51790 31630 51850
rect 31800 51790 31810 51850
rect 31980 51790 31990 51850
rect 32160 51790 32170 51850
rect 32340 51790 32350 51850
rect 32520 51790 32530 51850
rect 32700 51790 32710 51850
rect 32880 51790 32890 51850
rect 33060 51790 33070 51850
rect 33240 51790 33250 51850
rect 33420 51790 33430 51850
rect 33600 51790 33610 51850
rect 33780 51790 33790 51850
rect 33960 51790 33970 51850
rect 34140 51790 34150 51850
rect 34320 51790 34330 51850
rect 34500 51790 34510 51850
rect 34680 51790 34690 51850
rect 34860 51790 34870 51850
rect 35040 51790 35050 51850
rect 35220 51790 35230 51850
rect 35400 51790 35410 51850
rect 35580 51790 35590 51850
rect 35760 51790 35770 51850
rect 35940 51790 35950 51850
rect 36120 51790 36130 51850
rect 36300 51790 36310 51850
rect 36480 51790 36490 51850
rect 36660 51790 36670 51850
rect 36840 51790 36850 51850
rect 37020 51790 37030 51850
rect 37100 51780 37190 51850
rect 37600 51840 37660 51870
rect 37720 51840 37780 51870
rect 37840 51840 37900 51870
rect 40170 51820 40180 51910
rect 40060 51790 40120 51820
rect 19130 51750 19160 51780
rect 19250 51750 19280 51780
rect 26420 51750 26450 51780
rect 26540 51750 26570 51780
rect 30420 51750 30450 51780
rect 30540 51750 30570 51780
rect 31100 51750 37190 51780
rect 37720 51750 37750 51780
rect 37840 51750 37870 51780
rect 19010 51720 19070 51750
rect 19130 51720 19190 51750
rect 19250 51720 19310 51750
rect 19800 51730 25800 51740
rect 26300 51720 26360 51750
rect 26420 51720 26480 51750
rect 26540 51720 26600 51750
rect 30300 51720 30360 51750
rect 30420 51720 30480 51750
rect 30540 51720 30600 51750
rect 37100 51740 37190 51750
rect 31100 51730 37190 51740
rect 19130 51630 19160 51660
rect 19250 51630 19280 51660
rect 26420 51630 26450 51660
rect 26540 51630 26570 51660
rect 30420 51630 30450 51660
rect 30540 51630 30570 51660
rect 19010 51600 19070 51630
rect 19130 51600 19190 51630
rect 19250 51600 19310 51630
rect 26300 51600 26360 51630
rect 26420 51600 26480 51630
rect 26540 51600 26600 51630
rect 30300 51600 30360 51630
rect 30420 51600 30480 51630
rect 30540 51600 30600 51630
rect 31180 51550 31260 51560
rect 31360 51550 31440 51560
rect 31540 51550 31620 51560
rect 31720 51550 31800 51560
rect 31900 51550 31980 51560
rect 32080 51550 32160 51560
rect 32260 51550 32340 51560
rect 32440 51550 32520 51560
rect 32620 51550 32700 51560
rect 32800 51550 32880 51560
rect 32980 51550 33060 51560
rect 33160 51550 33240 51560
rect 33340 51550 33420 51560
rect 33520 51550 33600 51560
rect 33700 51550 33780 51560
rect 33880 51550 33960 51560
rect 34060 51550 34140 51560
rect 34240 51550 34320 51560
rect 34420 51550 34500 51560
rect 34600 51550 34680 51560
rect 34780 51550 34860 51560
rect 34960 51550 35040 51560
rect 35140 51550 35220 51560
rect 35320 51550 35400 51560
rect 35500 51550 35580 51560
rect 35680 51550 35760 51560
rect 35860 51550 35940 51560
rect 36040 51550 36120 51560
rect 36220 51550 36300 51560
rect 36400 51550 36480 51560
rect 36580 51550 36660 51560
rect 36760 51550 36840 51560
rect 36940 51550 37020 51560
rect 19130 51510 19160 51540
rect 19250 51510 19280 51540
rect 19880 51530 19960 51540
rect 20060 51530 20140 51540
rect 20240 51530 20320 51540
rect 20420 51530 20500 51540
rect 20600 51530 20680 51540
rect 20780 51530 20860 51540
rect 20960 51530 21040 51540
rect 21140 51530 21220 51540
rect 21320 51530 21400 51540
rect 21500 51530 21580 51540
rect 21680 51530 21760 51540
rect 21860 51530 21940 51540
rect 22040 51530 22120 51540
rect 22220 51530 22300 51540
rect 22400 51530 22480 51540
rect 22580 51530 22660 51540
rect 22760 51530 22840 51540
rect 22940 51530 23020 51540
rect 23120 51530 23200 51540
rect 23300 51530 23380 51540
rect 23480 51530 23560 51540
rect 23660 51530 23740 51540
rect 23840 51530 23920 51540
rect 24020 51530 24100 51540
rect 24200 51530 24280 51540
rect 24380 51530 24460 51540
rect 24560 51530 24640 51540
rect 24740 51530 24820 51540
rect 24920 51530 25000 51540
rect 25100 51530 25180 51540
rect 25280 51530 25360 51540
rect 25460 51530 25540 51540
rect 25640 51530 25720 51540
rect 19010 51480 19070 51510
rect 19130 51480 19190 51510
rect 19250 51480 19310 51510
rect 19960 51450 19970 51530
rect 20140 51450 20150 51530
rect 20320 51450 20330 51530
rect 20500 51450 20510 51530
rect 20680 51450 20690 51530
rect 20860 51450 20870 51530
rect 21040 51450 21050 51530
rect 21220 51450 21230 51530
rect 21400 51450 21410 51530
rect 21580 51450 21590 51530
rect 21760 51450 21770 51530
rect 21940 51450 21950 51530
rect 22120 51450 22130 51530
rect 22300 51450 22310 51530
rect 22480 51450 22490 51530
rect 22660 51450 22670 51530
rect 22840 51450 22850 51530
rect 23020 51450 23030 51530
rect 23200 51450 23210 51530
rect 23380 51450 23390 51530
rect 23560 51450 23570 51530
rect 23740 51450 23750 51530
rect 23920 51450 23930 51530
rect 24100 51450 24110 51530
rect 24280 51450 24290 51530
rect 24460 51450 24470 51530
rect 24640 51450 24650 51530
rect 24820 51450 24830 51530
rect 25000 51450 25010 51530
rect 25180 51450 25190 51530
rect 25360 51450 25370 51530
rect 25540 51450 25550 51530
rect 25720 51450 25730 51530
rect 26420 51510 26450 51540
rect 26540 51510 26570 51540
rect 30420 51510 30450 51540
rect 30540 51510 30570 51540
rect 26300 51480 26360 51510
rect 26420 51480 26480 51510
rect 26540 51480 26600 51510
rect 30300 51480 30360 51510
rect 30420 51480 30480 51510
rect 30540 51480 30600 51510
rect 31260 51470 31270 51550
rect 31440 51470 31450 51550
rect 31620 51470 31630 51550
rect 31800 51470 31810 51550
rect 31980 51470 31990 51550
rect 32160 51470 32170 51550
rect 32340 51470 32350 51550
rect 32520 51470 32530 51550
rect 32700 51470 32710 51550
rect 32880 51470 32890 51550
rect 33060 51470 33070 51550
rect 33240 51470 33250 51550
rect 33420 51470 33430 51550
rect 33600 51470 33610 51550
rect 33780 51470 33790 51550
rect 33960 51470 33970 51550
rect 34140 51470 34150 51550
rect 34320 51470 34330 51550
rect 34500 51470 34510 51550
rect 34680 51470 34690 51550
rect 34860 51470 34870 51550
rect 35040 51470 35050 51550
rect 35220 51470 35230 51550
rect 35400 51470 35410 51550
rect 35580 51470 35590 51550
rect 35760 51470 35770 51550
rect 35940 51470 35950 51550
rect 36120 51470 36130 51550
rect 36300 51470 36310 51550
rect 36480 51470 36490 51550
rect 36660 51470 36670 51550
rect 36840 51470 36850 51550
rect 37020 51470 37030 51550
rect 19130 51390 19160 51420
rect 19250 51390 19280 51420
rect 26420 51390 26450 51420
rect 26540 51390 26570 51420
rect 30420 51390 30450 51420
rect 30540 51390 30570 51420
rect 19010 51360 19070 51390
rect 19130 51360 19190 51390
rect 19250 51360 19310 51390
rect 26300 51360 26360 51390
rect 26420 51360 26480 51390
rect 26540 51360 26600 51390
rect 30300 51360 30360 51390
rect 30420 51360 30480 51390
rect 30540 51360 30600 51390
rect 19130 51270 19160 51300
rect 19250 51270 19280 51300
rect 26420 51270 26450 51300
rect 26540 51270 26570 51300
rect 30420 51270 30450 51300
rect 30540 51270 30570 51300
rect 19010 51240 19070 51270
rect 19130 51240 19190 51270
rect 19250 51240 19310 51270
rect 26300 51240 26360 51270
rect 26420 51240 26480 51270
rect 26540 51240 26600 51270
rect 30300 51240 30360 51270
rect 30420 51240 30480 51270
rect 30540 51240 30600 51270
rect 19880 51230 19960 51240
rect 20060 51230 20140 51240
rect 20240 51230 20320 51240
rect 20420 51230 20500 51240
rect 20600 51230 20680 51240
rect 20780 51230 20860 51240
rect 20960 51230 21040 51240
rect 21140 51230 21220 51240
rect 21320 51230 21400 51240
rect 21500 51230 21580 51240
rect 21680 51230 21760 51240
rect 21860 51230 21940 51240
rect 22040 51230 22120 51240
rect 22220 51230 22300 51240
rect 22400 51230 22480 51240
rect 22580 51230 22660 51240
rect 22760 51230 22840 51240
rect 22940 51230 23020 51240
rect 23120 51230 23200 51240
rect 23300 51230 23380 51240
rect 23480 51230 23560 51240
rect 23660 51230 23740 51240
rect 23840 51230 23920 51240
rect 24020 51230 24100 51240
rect 24200 51230 24280 51240
rect 24380 51230 24460 51240
rect 24560 51230 24640 51240
rect 24740 51230 24820 51240
rect 24920 51230 25000 51240
rect 25100 51230 25180 51240
rect 25280 51230 25360 51240
rect 25460 51230 25540 51240
rect 25640 51230 25720 51240
rect 31180 51230 31260 51240
rect 31360 51230 31440 51240
rect 31540 51230 31620 51240
rect 31720 51230 31800 51240
rect 31900 51230 31980 51240
rect 32080 51230 32160 51240
rect 32260 51230 32340 51240
rect 32440 51230 32520 51240
rect 32620 51230 32700 51240
rect 32800 51230 32880 51240
rect 32980 51230 33060 51240
rect 33160 51230 33240 51240
rect 33340 51230 33420 51240
rect 33520 51230 33600 51240
rect 33700 51230 33780 51240
rect 33880 51230 33960 51240
rect 34060 51230 34140 51240
rect 34240 51230 34320 51240
rect 34420 51230 34500 51240
rect 34600 51230 34680 51240
rect 34780 51230 34860 51240
rect 34960 51230 35040 51240
rect 35140 51230 35220 51240
rect 35320 51230 35400 51240
rect 35500 51230 35580 51240
rect 35680 51230 35760 51240
rect 35860 51230 35940 51240
rect 36040 51230 36120 51240
rect 36220 51230 36300 51240
rect 36400 51230 36480 51240
rect 36580 51230 36660 51240
rect 36760 51230 36840 51240
rect 36940 51230 37020 51240
rect 19130 51150 19160 51180
rect 19250 51150 19280 51180
rect 19960 51150 19970 51230
rect 20140 51150 20150 51230
rect 20320 51150 20330 51230
rect 20500 51150 20510 51230
rect 20680 51150 20690 51230
rect 20860 51150 20870 51230
rect 21040 51150 21050 51230
rect 21220 51150 21230 51230
rect 21400 51150 21410 51230
rect 21580 51150 21590 51230
rect 21760 51150 21770 51230
rect 21940 51150 21950 51230
rect 22120 51150 22130 51230
rect 22300 51150 22310 51230
rect 22480 51150 22490 51230
rect 22660 51150 22670 51230
rect 22840 51150 22850 51230
rect 23020 51150 23030 51230
rect 23200 51150 23210 51230
rect 23380 51150 23390 51230
rect 23560 51150 23570 51230
rect 23740 51150 23750 51230
rect 23920 51150 23930 51230
rect 24100 51150 24110 51230
rect 24280 51150 24290 51230
rect 24460 51150 24470 51230
rect 24640 51150 24650 51230
rect 24820 51150 24830 51230
rect 25000 51150 25010 51230
rect 25180 51150 25190 51230
rect 25360 51150 25370 51230
rect 25540 51150 25550 51230
rect 25720 51150 25730 51230
rect 26420 51150 26450 51180
rect 26540 51150 26570 51180
rect 30420 51150 30450 51180
rect 30540 51150 30570 51180
rect 31260 51150 31270 51230
rect 31440 51150 31450 51230
rect 31620 51150 31630 51230
rect 31800 51150 31810 51230
rect 31980 51150 31990 51230
rect 32160 51150 32170 51230
rect 32340 51150 32350 51230
rect 32520 51150 32530 51230
rect 32700 51150 32710 51230
rect 32880 51150 32890 51230
rect 33060 51150 33070 51230
rect 33240 51150 33250 51230
rect 33420 51150 33430 51230
rect 33600 51150 33610 51230
rect 33780 51150 33790 51230
rect 33960 51150 33970 51230
rect 34140 51150 34150 51230
rect 34320 51150 34330 51230
rect 34500 51150 34510 51230
rect 34680 51150 34690 51230
rect 34860 51150 34870 51230
rect 35040 51150 35050 51230
rect 35220 51150 35230 51230
rect 35400 51150 35410 51230
rect 35580 51150 35590 51230
rect 35760 51150 35770 51230
rect 35940 51150 35950 51230
rect 36120 51150 36130 51230
rect 36300 51150 36310 51230
rect 36480 51150 36490 51230
rect 36660 51150 36670 51230
rect 36840 51150 36850 51230
rect 37020 51150 37030 51230
rect 19010 51120 19070 51150
rect 19130 51120 19190 51150
rect 19250 51120 19310 51150
rect 26300 51120 26360 51150
rect 26420 51120 26480 51150
rect 26540 51120 26600 51150
rect 30300 51120 30360 51150
rect 30420 51120 30480 51150
rect 30540 51120 30600 51150
rect 37100 51060 37190 51730
rect 37600 51720 37660 51750
rect 37720 51720 37780 51750
rect 37840 51720 37900 51750
rect 40060 51670 40120 51700
rect 37720 51630 37750 51660
rect 37840 51630 37870 51660
rect 37600 51600 37660 51630
rect 37720 51600 37780 51630
rect 37840 51600 37900 51630
rect 40060 51550 40120 51580
rect 37720 51510 37750 51540
rect 37840 51510 37870 51540
rect 37600 51480 37660 51510
rect 37720 51480 37780 51510
rect 37840 51480 37900 51510
rect 40060 51430 40120 51460
rect 37720 51390 37750 51420
rect 37840 51390 37870 51420
rect 37600 51360 37660 51390
rect 37720 51360 37780 51390
rect 37840 51360 37900 51390
rect 40060 51310 40120 51340
rect 37720 51270 37750 51300
rect 37840 51270 37870 51300
rect 37600 51240 37660 51270
rect 37720 51240 37780 51270
rect 37840 51240 37900 51270
rect 40060 51190 40120 51220
rect 37720 51150 37750 51180
rect 37840 51150 37870 51180
rect 37600 51120 37660 51150
rect 37720 51120 37780 51150
rect 37840 51120 37900 51150
rect 40060 51070 40120 51100
rect 19130 51030 19160 51060
rect 19250 51030 19280 51060
rect 19800 51050 25800 51060
rect 26420 51030 26450 51060
rect 26540 51030 26570 51060
rect 30420 51030 30450 51060
rect 30540 51030 30570 51060
rect 31100 51050 37190 51060
rect 19010 51000 19070 51030
rect 19130 51000 19190 51030
rect 19250 51000 19310 51030
rect 26300 51000 26360 51030
rect 26420 51000 26480 51030
rect 26540 51000 26600 51030
rect 30300 51000 30360 51030
rect 30420 51000 30480 51030
rect 30540 51000 30600 51030
rect 37100 50950 37190 51050
rect 37720 51030 37750 51060
rect 37840 51030 37870 51060
rect 40260 51030 40270 51820
rect 40380 51810 41180 51900
rect 40650 51780 40770 51810
rect 40930 51780 41050 51810
rect 41090 51780 41180 51810
rect 40650 51690 40660 51780
rect 40760 51750 40830 51780
rect 40770 51660 40830 51750
rect 40930 51690 40940 51780
rect 41050 51660 41180 51780
rect 41260 51740 41340 51750
rect 41340 51690 41350 51740
rect 41090 51625 41180 51660
rect 41230 51630 41350 51690
rect 40470 51620 41180 51625
rect 40370 51610 41180 51620
rect 40370 51530 40380 51610
rect 40470 51605 41180 51610
rect 40420 51595 41210 51605
rect 41090 51545 41180 51595
rect 40470 51530 41180 51545
rect 40460 51515 41180 51530
rect 40460 51325 40470 51515
rect 40650 51480 40770 51515
rect 40930 51480 41050 51515
rect 41090 51480 41180 51515
rect 41350 51510 41410 51630
rect 40770 51470 40830 51480
rect 40530 51460 40610 51470
rect 40670 51460 40750 51470
rect 40770 51460 40890 51470
rect 40950 51460 41030 51470
rect 40610 51380 40620 51460
rect 40750 51380 40760 51460
rect 40770 51360 40830 51460
rect 40890 51380 40900 51460
rect 41030 51380 41040 51460
rect 41050 51360 41180 51480
rect 41260 51460 41340 51470
rect 41340 51390 41350 51460
rect 41090 51325 41180 51360
rect 41230 51330 41350 51390
rect 40460 51310 41180 51325
rect 40470 51305 41180 51310
rect 40420 51295 41210 51305
rect 41090 51245 41180 51295
rect 40470 51215 41180 51245
rect 40650 51180 40770 51215
rect 40930 51180 41050 51215
rect 41090 51180 41180 51215
rect 41350 51210 41410 51330
rect 41480 51180 41490 51890
rect 42860 51870 43470 51880
rect 43550 51870 43560 52115
rect 43700 52030 43760 52150
rect 146100 52110 146160 52140
rect 147580 52110 147640 52140
rect 148400 52110 148460 52140
rect 149880 52110 149940 52140
rect 152220 52090 152250 52120
rect 152340 52090 152370 52120
rect 153060 52110 153070 52170
rect 153240 52110 153250 52170
rect 153420 52110 153430 52170
rect 153600 52110 153610 52170
rect 153780 52110 153790 52170
rect 153960 52110 153970 52170
rect 154140 52110 154150 52170
rect 154320 52110 154330 52170
rect 154500 52110 154510 52170
rect 154680 52110 154690 52170
rect 154860 52110 154870 52170
rect 155040 52110 155050 52170
rect 155220 52110 155230 52170
rect 155400 52110 155410 52170
rect 155580 52110 155590 52170
rect 155760 52110 155770 52170
rect 155940 52110 155950 52170
rect 156120 52110 156130 52170
rect 156300 52110 156310 52170
rect 156480 52110 156490 52170
rect 156660 52110 156670 52170
rect 156840 52110 156850 52170
rect 157020 52110 157030 52170
rect 157200 52110 157210 52170
rect 157380 52110 157390 52170
rect 157560 52110 157570 52170
rect 157740 52110 157750 52170
rect 157920 52110 157930 52170
rect 158100 52110 158110 52170
rect 158280 52110 158290 52170
rect 158460 52110 158470 52170
rect 158640 52110 158650 52170
rect 158820 52110 158830 52170
rect 158900 52110 158990 52180
rect 164280 52170 164360 52180
rect 164460 52170 164540 52180
rect 164640 52170 164720 52180
rect 164820 52170 164900 52180
rect 165000 52170 165080 52180
rect 165180 52170 165260 52180
rect 165360 52170 165440 52180
rect 165540 52170 165620 52180
rect 165720 52170 165800 52180
rect 165900 52170 165980 52180
rect 166080 52170 166160 52180
rect 166260 52170 166340 52180
rect 166440 52170 166520 52180
rect 166620 52170 166700 52180
rect 166800 52170 166880 52180
rect 166980 52170 167060 52180
rect 167160 52170 167240 52180
rect 167340 52170 167420 52180
rect 167520 52170 167600 52180
rect 167700 52170 167780 52180
rect 167880 52170 167960 52180
rect 168060 52170 168140 52180
rect 168240 52170 168320 52180
rect 168420 52170 168500 52180
rect 168600 52170 168680 52180
rect 168780 52170 168860 52180
rect 168960 52170 169040 52180
rect 169140 52170 169220 52180
rect 169320 52170 169400 52180
rect 169500 52170 169580 52180
rect 169680 52170 169760 52180
rect 169860 52170 169940 52180
rect 170040 52170 170120 52180
rect 152100 52060 152160 52090
rect 152220 52060 152280 52090
rect 152340 52060 152400 52090
rect 152900 52080 158990 52110
rect 159520 52090 159550 52120
rect 159640 52090 159670 52120
rect 163520 52090 163550 52120
rect 163640 52090 163670 52120
rect 164360 52090 164370 52170
rect 164540 52090 164550 52170
rect 164720 52090 164730 52170
rect 164900 52090 164910 52170
rect 165080 52090 165090 52170
rect 165260 52090 165270 52170
rect 165440 52090 165450 52170
rect 165620 52090 165630 52170
rect 165800 52090 165810 52170
rect 165980 52090 165990 52170
rect 166160 52090 166170 52170
rect 166340 52090 166350 52170
rect 166520 52090 166530 52170
rect 166700 52090 166710 52170
rect 166880 52090 166890 52170
rect 167060 52090 167070 52170
rect 167240 52090 167250 52170
rect 167420 52090 167430 52170
rect 167600 52090 167610 52170
rect 167780 52090 167790 52170
rect 167960 52090 167970 52170
rect 168140 52090 168150 52170
rect 168320 52090 168330 52170
rect 168500 52090 168510 52170
rect 168680 52090 168690 52170
rect 168860 52090 168870 52170
rect 169040 52090 169050 52170
rect 169220 52090 169230 52170
rect 169400 52090 169410 52170
rect 169580 52090 169590 52170
rect 169760 52090 169770 52170
rect 169940 52090 169950 52170
rect 170120 52090 170130 52170
rect 170810 52090 170840 52120
rect 170930 52090 170960 52120
rect 43840 52030 43900 52060
rect 152980 52020 153060 52030
rect 153160 52020 153240 52030
rect 153340 52020 153420 52030
rect 153520 52020 153600 52030
rect 153700 52020 153780 52030
rect 153880 52020 153960 52030
rect 154060 52020 154140 52030
rect 154240 52020 154320 52030
rect 154420 52020 154500 52030
rect 154600 52020 154680 52030
rect 154780 52020 154860 52030
rect 154960 52020 155040 52030
rect 155140 52020 155220 52030
rect 155320 52020 155400 52030
rect 155500 52020 155580 52030
rect 155680 52020 155760 52030
rect 155860 52020 155940 52030
rect 156040 52020 156120 52030
rect 156220 52020 156300 52030
rect 156400 52020 156480 52030
rect 156580 52020 156660 52030
rect 156760 52020 156840 52030
rect 156940 52020 157020 52030
rect 157120 52020 157200 52030
rect 157300 52020 157380 52030
rect 157480 52020 157560 52030
rect 157660 52020 157740 52030
rect 157840 52020 157920 52030
rect 158020 52020 158100 52030
rect 158200 52020 158280 52030
rect 158380 52020 158460 52030
rect 158560 52020 158640 52030
rect 158740 52020 158820 52030
rect 146100 51990 146160 52020
rect 147580 51990 147640 52020
rect 148400 51990 148460 52020
rect 149880 51990 149940 52020
rect 152220 51970 152250 52000
rect 152340 51970 152370 52000
rect 43580 51890 43700 51950
rect 152100 51940 152160 51970
rect 152220 51940 152280 51970
rect 152340 51940 152400 51970
rect 153060 51940 153070 52020
rect 153240 51940 153250 52020
rect 153420 51940 153430 52020
rect 153600 51940 153610 52020
rect 153780 51940 153790 52020
rect 153960 51940 153970 52020
rect 154140 51940 154150 52020
rect 154320 51940 154330 52020
rect 154500 51940 154510 52020
rect 154680 51940 154690 52020
rect 154860 51940 154870 52020
rect 155040 51940 155050 52020
rect 155220 51940 155230 52020
rect 155400 51940 155410 52020
rect 155580 51940 155590 52020
rect 155760 51940 155770 52020
rect 155940 51940 155950 52020
rect 156120 51940 156130 52020
rect 156300 51940 156310 52020
rect 156480 51940 156490 52020
rect 156660 51940 156670 52020
rect 156840 51940 156850 52020
rect 157020 51940 157030 52020
rect 157200 51940 157210 52020
rect 157380 51940 157390 52020
rect 157560 51940 157570 52020
rect 157740 51940 157750 52020
rect 157920 51940 157930 52020
rect 158100 51940 158110 52020
rect 158280 51940 158290 52020
rect 158460 51940 158470 52020
rect 158640 51940 158650 52020
rect 158820 51940 158830 52020
rect 43840 51910 43900 51940
rect 42910 51855 43560 51865
rect 41540 51790 41600 51820
rect 42360 51790 42420 51820
rect 42900 51805 42910 51855
rect 43030 51760 43390 51820
rect 43700 51770 43760 51890
rect 146100 51870 146160 51900
rect 147580 51870 147640 51900
rect 148400 51870 148460 51900
rect 149880 51870 149940 51900
rect 158900 51880 158990 52080
rect 159400 52060 159460 52090
rect 159520 52060 159580 52090
rect 159640 52060 159700 52090
rect 163400 52060 163460 52090
rect 163520 52060 163580 52090
rect 163640 52060 163700 52090
rect 170690 52060 170750 52090
rect 170810 52060 170870 52090
rect 170930 52060 170990 52090
rect 164280 52020 164360 52030
rect 164460 52020 164540 52030
rect 164640 52020 164720 52030
rect 164820 52020 164900 52030
rect 165000 52020 165080 52030
rect 165180 52020 165260 52030
rect 165360 52020 165440 52030
rect 165540 52020 165620 52030
rect 165720 52020 165800 52030
rect 165900 52020 165980 52030
rect 166080 52020 166160 52030
rect 166260 52020 166340 52030
rect 166440 52020 166520 52030
rect 166620 52020 166700 52030
rect 166800 52020 166880 52030
rect 166980 52020 167060 52030
rect 167160 52020 167240 52030
rect 167340 52020 167420 52030
rect 167520 52020 167600 52030
rect 167700 52020 167780 52030
rect 167880 52020 167960 52030
rect 168060 52020 168140 52030
rect 168240 52020 168320 52030
rect 168420 52020 168500 52030
rect 168600 52020 168680 52030
rect 168780 52020 168860 52030
rect 168960 52020 169040 52030
rect 169140 52020 169220 52030
rect 169320 52020 169400 52030
rect 169500 52020 169580 52030
rect 169680 52020 169760 52030
rect 169860 52020 169940 52030
rect 170040 52020 170120 52030
rect 159520 51970 159550 52000
rect 159640 51970 159670 52000
rect 163520 51970 163550 52000
rect 163640 51970 163670 52000
rect 159400 51940 159460 51970
rect 159520 51940 159580 51970
rect 159640 51940 159700 51970
rect 163400 51940 163460 51970
rect 163520 51940 163580 51970
rect 163640 51940 163700 51970
rect 164360 51940 164370 52020
rect 164540 51940 164550 52020
rect 164720 51940 164730 52020
rect 164900 51940 164910 52020
rect 165080 51940 165090 52020
rect 165260 51940 165270 52020
rect 165440 51940 165450 52020
rect 165620 51940 165630 52020
rect 165800 51940 165810 52020
rect 165980 51940 165990 52020
rect 166160 51940 166170 52020
rect 166340 51940 166350 52020
rect 166520 51940 166530 52020
rect 166700 51940 166710 52020
rect 166880 51940 166890 52020
rect 167060 51940 167070 52020
rect 167240 51940 167250 52020
rect 167420 51940 167430 52020
rect 167600 51940 167610 52020
rect 167780 51940 167790 52020
rect 167960 51940 167970 52020
rect 168140 51940 168150 52020
rect 168320 51940 168330 52020
rect 168500 51940 168510 52020
rect 168680 51940 168690 52020
rect 168860 51940 168870 52020
rect 169040 51940 169050 52020
rect 169220 51940 169230 52020
rect 169400 51940 169410 52020
rect 169580 51940 169590 52020
rect 169760 51940 169770 52020
rect 169940 51940 169950 52020
rect 170120 51940 170130 52020
rect 170810 51970 170840 52000
rect 170930 51970 170960 52000
rect 170690 51940 170750 51970
rect 170810 51940 170870 51970
rect 170930 51940 170990 51970
rect 152220 51850 152250 51880
rect 152340 51850 152370 51880
rect 152900 51850 158990 51880
rect 159520 51850 159550 51880
rect 159640 51850 159670 51880
rect 163520 51850 163550 51880
rect 163640 51850 163670 51880
rect 164280 51870 164360 51880
rect 164460 51870 164540 51880
rect 164640 51870 164720 51880
rect 164820 51870 164900 51880
rect 165000 51870 165080 51880
rect 165180 51870 165260 51880
rect 165360 51870 165440 51880
rect 165540 51870 165620 51880
rect 165720 51870 165800 51880
rect 165900 51870 165980 51880
rect 166080 51870 166160 51880
rect 166260 51870 166340 51880
rect 166440 51870 166520 51880
rect 166620 51870 166700 51880
rect 166800 51870 166880 51880
rect 166980 51870 167060 51880
rect 167160 51870 167240 51880
rect 167340 51870 167420 51880
rect 167520 51870 167600 51880
rect 167700 51870 167780 51880
rect 167880 51870 167960 51880
rect 168060 51870 168140 51880
rect 168240 51870 168320 51880
rect 168420 51870 168500 51880
rect 168600 51870 168680 51880
rect 168780 51870 168860 51880
rect 168960 51870 169040 51880
rect 169140 51870 169220 51880
rect 169320 51870 169400 51880
rect 169500 51870 169580 51880
rect 169680 51870 169760 51880
rect 169860 51870 169940 51880
rect 170040 51870 170120 51880
rect 152100 51820 152160 51850
rect 152220 51820 152280 51850
rect 152340 51820 152400 51850
rect 43840 51790 43900 51820
rect 153060 51790 153070 51850
rect 153240 51790 153250 51850
rect 153420 51790 153430 51850
rect 153600 51790 153610 51850
rect 153780 51790 153790 51850
rect 153960 51790 153970 51850
rect 154140 51790 154150 51850
rect 154320 51790 154330 51850
rect 154500 51790 154510 51850
rect 154680 51790 154690 51850
rect 154860 51790 154870 51850
rect 155040 51790 155050 51850
rect 155220 51790 155230 51850
rect 155400 51790 155410 51850
rect 155580 51790 155590 51850
rect 155760 51790 155770 51850
rect 155940 51790 155950 51850
rect 156120 51790 156130 51850
rect 156300 51790 156310 51850
rect 156480 51790 156490 51850
rect 156660 51790 156670 51850
rect 156840 51790 156850 51850
rect 157020 51790 157030 51850
rect 157200 51790 157210 51850
rect 157380 51790 157390 51850
rect 157560 51790 157570 51850
rect 157740 51790 157750 51850
rect 157920 51790 157930 51850
rect 158100 51790 158110 51850
rect 158280 51790 158290 51850
rect 158460 51790 158470 51850
rect 158640 51790 158650 51850
rect 158820 51790 158830 51850
rect 158900 51780 158990 51850
rect 159400 51820 159460 51850
rect 159520 51820 159580 51850
rect 159640 51820 159700 51850
rect 163400 51820 163460 51850
rect 163520 51820 163580 51850
rect 163640 51820 163700 51850
rect 164360 51790 164370 51870
rect 164540 51790 164550 51870
rect 164720 51790 164730 51870
rect 164900 51790 164910 51870
rect 165080 51790 165090 51870
rect 165260 51790 165270 51870
rect 165440 51790 165450 51870
rect 165620 51790 165630 51870
rect 165800 51790 165810 51870
rect 165980 51790 165990 51870
rect 166160 51790 166170 51870
rect 166340 51790 166350 51870
rect 166520 51790 166530 51870
rect 166700 51790 166710 51870
rect 166880 51790 166890 51870
rect 167060 51790 167070 51870
rect 167240 51790 167250 51870
rect 167420 51790 167430 51870
rect 167600 51790 167610 51870
rect 167780 51790 167790 51870
rect 167960 51790 167970 51870
rect 168140 51790 168150 51870
rect 168320 51790 168330 51870
rect 168500 51790 168510 51870
rect 168680 51790 168690 51870
rect 168860 51790 168870 51870
rect 169040 51790 169050 51870
rect 169220 51790 169230 51870
rect 169400 51790 169410 51870
rect 169580 51790 169590 51870
rect 169760 51790 169770 51870
rect 169940 51790 169950 51870
rect 170120 51790 170130 51870
rect 170810 51850 170840 51880
rect 170930 51850 170960 51880
rect 170690 51820 170750 51850
rect 170810 51820 170870 51850
rect 170930 51820 170990 51850
rect 146100 51750 146160 51780
rect 147580 51750 147640 51780
rect 148400 51750 148460 51780
rect 149880 51750 149940 51780
rect 41540 51670 41600 51700
rect 42360 51670 42420 51700
rect 42470 51660 42480 51750
rect 152220 51730 152250 51760
rect 152340 51730 152370 51760
rect 152900 51750 158990 51780
rect 158900 51740 158990 51750
rect 152900 51730 158990 51740
rect 159520 51730 159550 51760
rect 159640 51730 159670 51760
rect 163520 51730 163550 51760
rect 163640 51730 163670 51760
rect 164200 51730 170200 51740
rect 170810 51730 170840 51760
rect 170930 51730 170960 51760
rect 152100 51700 152160 51730
rect 152220 51700 152280 51730
rect 152340 51700 152400 51730
rect 43840 51670 43900 51700
rect 41540 51550 41600 51580
rect 42360 51550 42420 51580
rect 41540 51430 41600 51460
rect 42360 51430 42420 51460
rect 41540 51310 41600 51340
rect 42360 51310 42420 51340
rect 41540 51190 41600 51220
rect 42360 51190 42420 51220
rect 42560 51180 42570 51660
rect 146100 51630 146160 51660
rect 147580 51630 147640 51660
rect 148400 51630 148460 51660
rect 149880 51630 149940 51660
rect 42960 51620 43460 51630
rect 152220 51610 152250 51640
rect 152340 51610 152370 51640
rect 42620 51600 42700 51610
rect 42700 51530 42710 51600
rect 42620 51520 42710 51530
rect 42770 51520 42780 51610
rect 152100 51580 152160 51610
rect 152220 51580 152280 51610
rect 152340 51580 152400 51610
rect 43840 51550 43900 51580
rect 152980 51550 153060 51560
rect 153160 51550 153240 51560
rect 153340 51550 153420 51560
rect 153520 51550 153600 51560
rect 153700 51550 153780 51560
rect 153880 51550 153960 51560
rect 154060 51550 154140 51560
rect 154240 51550 154320 51560
rect 154420 51550 154500 51560
rect 154600 51550 154680 51560
rect 154780 51550 154860 51560
rect 154960 51550 155040 51560
rect 155140 51550 155220 51560
rect 155320 51550 155400 51560
rect 155500 51550 155580 51560
rect 155680 51550 155760 51560
rect 155860 51550 155940 51560
rect 156040 51550 156120 51560
rect 156220 51550 156300 51560
rect 156400 51550 156480 51560
rect 156580 51550 156660 51560
rect 156760 51550 156840 51560
rect 156940 51550 157020 51560
rect 157120 51550 157200 51560
rect 157300 51550 157380 51560
rect 157480 51550 157560 51560
rect 157660 51550 157740 51560
rect 157840 51550 157920 51560
rect 158020 51550 158100 51560
rect 158200 51550 158280 51560
rect 158380 51550 158460 51560
rect 158560 51550 158640 51560
rect 158740 51550 158820 51560
rect 42620 51440 42700 51450
rect 42700 51390 42710 51440
rect 42610 51330 42730 51390
rect 42730 51305 42790 51330
rect 42860 51320 42870 51520
rect 42910 51480 43030 51540
rect 43190 51480 43310 51540
rect 146100 51510 146160 51540
rect 147580 51510 147640 51540
rect 148400 51510 148460 51540
rect 149880 51510 149940 51540
rect 152220 51490 152250 51520
rect 152340 51490 152370 51520
rect 43030 51470 43090 51480
rect 43310 51470 43370 51480
rect 42930 51460 43010 51470
rect 43030 51460 43150 51470
rect 43210 51460 43290 51470
rect 43310 51460 43430 51470
rect 152100 51460 152160 51490
rect 152220 51460 152280 51490
rect 152340 51460 152400 51490
rect 153060 51470 153070 51550
rect 153240 51470 153250 51550
rect 153420 51470 153430 51550
rect 153600 51470 153610 51550
rect 153780 51470 153790 51550
rect 153960 51470 153970 51550
rect 154140 51470 154150 51550
rect 154320 51470 154330 51550
rect 154500 51470 154510 51550
rect 154680 51470 154690 51550
rect 154860 51470 154870 51550
rect 155040 51470 155050 51550
rect 155220 51470 155230 51550
rect 155400 51470 155410 51550
rect 155580 51470 155590 51550
rect 155760 51470 155770 51550
rect 155940 51470 155950 51550
rect 156120 51470 156130 51550
rect 156300 51470 156310 51550
rect 156480 51470 156490 51550
rect 156660 51470 156670 51550
rect 156840 51470 156850 51550
rect 157020 51470 157030 51550
rect 157200 51470 157210 51550
rect 157380 51470 157390 51550
rect 157560 51470 157570 51550
rect 157740 51470 157750 51550
rect 157920 51470 157930 51550
rect 158100 51470 158110 51550
rect 158280 51470 158290 51550
rect 158460 51470 158470 51550
rect 158640 51470 158650 51550
rect 158820 51470 158830 51550
rect 43010 51380 43020 51460
rect 43030 51360 43090 51460
rect 43150 51380 43160 51460
rect 43290 51380 43300 51460
rect 43310 51360 43370 51460
rect 43430 51380 43440 51460
rect 43840 51430 43900 51460
rect 146100 51390 146160 51420
rect 147580 51390 147640 51420
rect 148400 51390 148460 51420
rect 149880 51390 149940 51420
rect 152220 51370 152250 51400
rect 152340 51370 152370 51400
rect 152100 51340 152160 51370
rect 152220 51340 152280 51370
rect 152340 51340 152400 51370
rect 42860 51310 43500 51320
rect 43840 51310 43900 51340
rect 42730 51295 43540 51305
rect 42730 51210 42790 51295
rect 43540 51245 43550 51295
rect 146100 51270 146160 51300
rect 147580 51270 147640 51300
rect 148400 51270 148460 51300
rect 149880 51270 149940 51300
rect 152220 51250 152250 51280
rect 152340 51250 152370 51280
rect 42860 51180 42870 51230
rect 42910 51180 43030 51240
rect 43190 51180 43310 51240
rect 152100 51220 152160 51250
rect 152220 51220 152280 51250
rect 152340 51220 152400 51250
rect 152980 51230 153060 51240
rect 153160 51230 153240 51240
rect 153340 51230 153420 51240
rect 153520 51230 153600 51240
rect 153700 51230 153780 51240
rect 153880 51230 153960 51240
rect 154060 51230 154140 51240
rect 154240 51230 154320 51240
rect 154420 51230 154500 51240
rect 154600 51230 154680 51240
rect 154780 51230 154860 51240
rect 154960 51230 155040 51240
rect 155140 51230 155220 51240
rect 155320 51230 155400 51240
rect 155500 51230 155580 51240
rect 155680 51230 155760 51240
rect 155860 51230 155940 51240
rect 156040 51230 156120 51240
rect 156220 51230 156300 51240
rect 156400 51230 156480 51240
rect 156580 51230 156660 51240
rect 156760 51230 156840 51240
rect 156940 51230 157020 51240
rect 157120 51230 157200 51240
rect 157300 51230 157380 51240
rect 157480 51230 157560 51240
rect 157660 51230 157740 51240
rect 157840 51230 157920 51240
rect 158020 51230 158100 51240
rect 158200 51230 158280 51240
rect 158380 51230 158460 51240
rect 158560 51230 158640 51240
rect 158740 51230 158820 51240
rect 43840 51190 43900 51220
rect 40770 51170 40830 51180
rect 40530 51160 40610 51170
rect 40770 51160 40890 51170
rect 40610 51080 40620 51160
rect 40770 51060 40830 51160
rect 40890 51080 40900 51160
rect 41050 51060 41180 51180
rect 43030 51170 43090 51180
rect 43310 51170 43370 51180
rect 43030 51160 43150 51170
rect 43310 51160 43430 51170
rect 41540 51070 41600 51100
rect 42360 51070 42420 51100
rect 43030 51060 43090 51160
rect 43150 51080 43160 51160
rect 43310 51060 43370 51160
rect 43430 51080 43440 51160
rect 146100 51150 146160 51180
rect 147580 51150 147640 51180
rect 148400 51150 148460 51180
rect 149880 51150 149940 51180
rect 152220 51130 152250 51160
rect 152340 51130 152370 51160
rect 153060 51150 153070 51230
rect 153240 51150 153250 51230
rect 153420 51150 153430 51230
rect 153600 51150 153610 51230
rect 153780 51150 153790 51230
rect 153960 51150 153970 51230
rect 154140 51150 154150 51230
rect 154320 51150 154330 51230
rect 154500 51150 154510 51230
rect 154680 51150 154690 51230
rect 154860 51150 154870 51230
rect 155040 51150 155050 51230
rect 155220 51150 155230 51230
rect 155400 51150 155410 51230
rect 155580 51150 155590 51230
rect 155760 51150 155770 51230
rect 155940 51150 155950 51230
rect 156120 51150 156130 51230
rect 156300 51150 156310 51230
rect 156480 51150 156490 51230
rect 156660 51150 156670 51230
rect 156840 51150 156850 51230
rect 157020 51150 157030 51230
rect 157200 51150 157210 51230
rect 157380 51150 157390 51230
rect 157560 51150 157570 51230
rect 157740 51150 157750 51230
rect 157920 51150 157930 51230
rect 158100 51150 158110 51230
rect 158280 51150 158290 51230
rect 158460 51150 158470 51230
rect 158640 51150 158650 51230
rect 158820 51150 158830 51230
rect 152100 51100 152160 51130
rect 152220 51100 152280 51130
rect 152340 51100 152400 51130
rect 43840 51070 43900 51100
rect 158900 51060 158990 51730
rect 159400 51700 159460 51730
rect 159520 51700 159580 51730
rect 159640 51700 159700 51730
rect 163400 51700 163460 51730
rect 163520 51700 163580 51730
rect 163640 51700 163700 51730
rect 170690 51700 170750 51730
rect 170810 51700 170870 51730
rect 170930 51700 170990 51730
rect 159520 51610 159550 51640
rect 159640 51610 159670 51640
rect 163520 51610 163550 51640
rect 163640 51610 163670 51640
rect 170810 51610 170840 51640
rect 170930 51610 170960 51640
rect 159400 51580 159460 51610
rect 159520 51580 159580 51610
rect 159640 51580 159700 51610
rect 163400 51580 163460 51610
rect 163520 51580 163580 51610
rect 163640 51580 163700 51610
rect 170690 51580 170750 51610
rect 170810 51580 170870 51610
rect 170930 51580 170990 51610
rect 164280 51550 164360 51560
rect 164460 51550 164540 51560
rect 164640 51550 164720 51560
rect 164820 51550 164900 51560
rect 165000 51550 165080 51560
rect 165180 51550 165260 51560
rect 165360 51550 165440 51560
rect 165540 51550 165620 51560
rect 165720 51550 165800 51560
rect 165900 51550 165980 51560
rect 166080 51550 166160 51560
rect 166260 51550 166340 51560
rect 166440 51550 166520 51560
rect 166620 51550 166700 51560
rect 166800 51550 166880 51560
rect 166980 51550 167060 51560
rect 167160 51550 167240 51560
rect 167340 51550 167420 51560
rect 167520 51550 167600 51560
rect 167700 51550 167780 51560
rect 167880 51550 167960 51560
rect 168060 51550 168140 51560
rect 168240 51550 168320 51560
rect 168420 51550 168500 51560
rect 168600 51550 168680 51560
rect 168780 51550 168860 51560
rect 168960 51550 169040 51560
rect 169140 51550 169220 51560
rect 169320 51550 169400 51560
rect 169500 51550 169580 51560
rect 169680 51550 169760 51560
rect 169860 51550 169940 51560
rect 170040 51550 170120 51560
rect 159520 51490 159550 51520
rect 159640 51490 159670 51520
rect 163520 51490 163550 51520
rect 163640 51490 163670 51520
rect 159400 51460 159460 51490
rect 159520 51460 159580 51490
rect 159640 51460 159700 51490
rect 163400 51460 163460 51490
rect 163520 51460 163580 51490
rect 163640 51460 163700 51490
rect 164360 51470 164370 51550
rect 164540 51470 164550 51550
rect 164720 51470 164730 51550
rect 164900 51470 164910 51550
rect 165080 51470 165090 51550
rect 165260 51470 165270 51550
rect 165440 51470 165450 51550
rect 165620 51470 165630 51550
rect 165800 51470 165810 51550
rect 165980 51470 165990 51550
rect 166160 51470 166170 51550
rect 166340 51470 166350 51550
rect 166520 51470 166530 51550
rect 166700 51470 166710 51550
rect 166880 51470 166890 51550
rect 167060 51470 167070 51550
rect 167240 51470 167250 51550
rect 167420 51470 167430 51550
rect 167600 51470 167610 51550
rect 167780 51470 167790 51550
rect 167960 51470 167970 51550
rect 168140 51470 168150 51550
rect 168320 51470 168330 51550
rect 168500 51470 168510 51550
rect 168680 51470 168690 51550
rect 168860 51470 168870 51550
rect 169040 51470 169050 51550
rect 169220 51470 169230 51550
rect 169400 51470 169410 51550
rect 169580 51470 169590 51550
rect 169760 51470 169770 51550
rect 169940 51470 169950 51550
rect 170120 51470 170130 51550
rect 170810 51490 170840 51520
rect 170930 51490 170960 51520
rect 170690 51460 170750 51490
rect 170810 51460 170870 51490
rect 170930 51460 170990 51490
rect 159520 51370 159550 51400
rect 159640 51370 159670 51400
rect 163520 51370 163550 51400
rect 163640 51370 163670 51400
rect 170810 51370 170840 51400
rect 170930 51370 170960 51400
rect 159400 51340 159460 51370
rect 159520 51340 159580 51370
rect 159640 51340 159700 51370
rect 163400 51340 163460 51370
rect 163520 51340 163580 51370
rect 163640 51340 163700 51370
rect 170690 51340 170750 51370
rect 170810 51340 170870 51370
rect 170930 51340 170990 51370
rect 159520 51250 159550 51280
rect 159640 51250 159670 51280
rect 163520 51250 163550 51280
rect 163640 51250 163670 51280
rect 164280 51250 164360 51260
rect 164460 51250 164540 51260
rect 164640 51250 164720 51260
rect 164820 51250 164900 51260
rect 165000 51250 165080 51260
rect 165180 51250 165260 51260
rect 165360 51250 165440 51260
rect 165540 51250 165620 51260
rect 165720 51250 165800 51260
rect 165900 51250 165980 51260
rect 166080 51250 166160 51260
rect 166260 51250 166340 51260
rect 166440 51250 166520 51260
rect 166620 51250 166700 51260
rect 166800 51250 166880 51260
rect 166980 51250 167060 51260
rect 167160 51250 167240 51260
rect 167340 51250 167420 51260
rect 167520 51250 167600 51260
rect 167700 51250 167780 51260
rect 167880 51250 167960 51260
rect 168060 51250 168140 51260
rect 168240 51250 168320 51260
rect 168420 51250 168500 51260
rect 168600 51250 168680 51260
rect 168780 51250 168860 51260
rect 168960 51250 169040 51260
rect 169140 51250 169220 51260
rect 169320 51250 169400 51260
rect 169500 51250 169580 51260
rect 169680 51250 169760 51260
rect 169860 51250 169940 51260
rect 170040 51250 170120 51260
rect 170810 51250 170840 51280
rect 170930 51250 170960 51280
rect 159400 51220 159460 51250
rect 159520 51220 159580 51250
rect 159640 51220 159700 51250
rect 163400 51220 163460 51250
rect 163520 51220 163580 51250
rect 163640 51220 163700 51250
rect 164360 51170 164370 51250
rect 164540 51170 164550 51250
rect 164720 51170 164730 51250
rect 164900 51170 164910 51250
rect 165080 51170 165090 51250
rect 165260 51170 165270 51250
rect 165440 51170 165450 51250
rect 165620 51170 165630 51250
rect 165800 51170 165810 51250
rect 165980 51170 165990 51250
rect 166160 51170 166170 51250
rect 166340 51170 166350 51250
rect 166520 51170 166530 51250
rect 166700 51170 166710 51250
rect 166880 51170 166890 51250
rect 167060 51170 167070 51250
rect 167240 51170 167250 51250
rect 167420 51170 167430 51250
rect 167600 51170 167610 51250
rect 167780 51170 167790 51250
rect 167960 51170 167970 51250
rect 168140 51170 168150 51250
rect 168320 51170 168330 51250
rect 168500 51170 168510 51250
rect 168680 51170 168690 51250
rect 168860 51170 168870 51250
rect 169040 51170 169050 51250
rect 169220 51170 169230 51250
rect 169400 51170 169410 51250
rect 169580 51170 169590 51250
rect 169760 51170 169770 51250
rect 169940 51170 169950 51250
rect 170120 51170 170130 51250
rect 170690 51220 170750 51250
rect 170810 51220 170870 51250
rect 170930 51220 170990 51250
rect 159520 51130 159550 51160
rect 159640 51130 159670 51160
rect 163520 51130 163550 51160
rect 163640 51130 163670 51160
rect 170810 51130 170840 51160
rect 170930 51130 170960 51160
rect 159400 51100 159460 51130
rect 159520 51100 159580 51130
rect 159640 51100 159700 51130
rect 163400 51100 163460 51130
rect 163520 51100 163580 51130
rect 163640 51100 163700 51130
rect 170690 51100 170750 51130
rect 170810 51100 170870 51130
rect 170930 51100 170990 51130
rect 41090 51050 41180 51060
rect 40470 51030 41180 51050
rect 146100 51030 146160 51060
rect 147580 51030 147640 51060
rect 148400 51030 148460 51060
rect 149880 51030 149940 51060
rect 152900 51050 158990 51060
rect 164200 51050 170200 51060
rect 37600 51000 37660 51030
rect 37720 51000 37780 51030
rect 37840 51000 37900 51030
rect 40060 50950 40120 50980
rect 19130 50910 19160 50940
rect 19250 50910 19280 50940
rect 19880 50910 19960 50920
rect 20060 50910 20140 50920
rect 20240 50910 20320 50920
rect 20420 50910 20500 50920
rect 20600 50910 20680 50920
rect 20780 50910 20860 50920
rect 20960 50910 21040 50920
rect 21140 50910 21220 50920
rect 21320 50910 21400 50920
rect 21500 50910 21580 50920
rect 21680 50910 21760 50920
rect 21860 50910 21940 50920
rect 22040 50910 22120 50920
rect 22220 50910 22300 50920
rect 22400 50910 22480 50920
rect 22580 50910 22660 50920
rect 22760 50910 22840 50920
rect 22940 50910 23020 50920
rect 23120 50910 23200 50920
rect 23300 50910 23380 50920
rect 23480 50910 23560 50920
rect 23660 50910 23740 50920
rect 23840 50910 23920 50920
rect 24020 50910 24100 50920
rect 24200 50910 24280 50920
rect 24380 50910 24460 50920
rect 24560 50910 24640 50920
rect 24740 50910 24820 50920
rect 24920 50910 25000 50920
rect 25100 50910 25180 50920
rect 25280 50910 25360 50920
rect 25460 50910 25540 50920
rect 25640 50910 25720 50920
rect 26420 50910 26450 50940
rect 26540 50910 26570 50940
rect 30420 50910 30450 50940
rect 30540 50910 30570 50940
rect 31100 50920 37190 50950
rect 40170 50940 40180 51030
rect 40260 51020 41100 51030
rect 31180 50910 31260 50920
rect 31360 50910 31440 50920
rect 31540 50910 31620 50920
rect 31720 50910 31800 50920
rect 31900 50910 31980 50920
rect 32080 50910 32160 50920
rect 32260 50910 32340 50920
rect 32440 50910 32520 50920
rect 32620 50910 32700 50920
rect 32800 50910 32880 50920
rect 32980 50910 33060 50920
rect 33160 50910 33240 50920
rect 33340 50910 33420 50920
rect 33520 50910 33600 50920
rect 33700 50910 33780 50920
rect 33880 50910 33960 50920
rect 34060 50910 34140 50920
rect 34240 50910 34320 50920
rect 34420 50910 34500 50920
rect 34600 50910 34680 50920
rect 34780 50910 34860 50920
rect 34960 50910 35040 50920
rect 35140 50910 35220 50920
rect 35320 50910 35400 50920
rect 35500 50910 35580 50920
rect 35680 50910 35760 50920
rect 35860 50910 35940 50920
rect 36040 50910 36120 50920
rect 36220 50910 36300 50920
rect 36400 50910 36480 50920
rect 36580 50910 36660 50920
rect 36760 50910 36840 50920
rect 36940 50910 37020 50920
rect 19010 50880 19070 50910
rect 19130 50880 19190 50910
rect 19250 50880 19310 50910
rect 19960 50830 19970 50910
rect 20140 50830 20150 50910
rect 20320 50830 20330 50910
rect 20500 50830 20510 50910
rect 20680 50830 20690 50910
rect 20860 50830 20870 50910
rect 21040 50830 21050 50910
rect 21220 50830 21230 50910
rect 21400 50830 21410 50910
rect 21580 50830 21590 50910
rect 21760 50830 21770 50910
rect 21940 50830 21950 50910
rect 22120 50830 22130 50910
rect 22300 50830 22310 50910
rect 22480 50830 22490 50910
rect 22660 50830 22670 50910
rect 22840 50830 22850 50910
rect 23020 50830 23030 50910
rect 23200 50830 23210 50910
rect 23380 50830 23390 50910
rect 23560 50830 23570 50910
rect 23740 50830 23750 50910
rect 23920 50830 23930 50910
rect 24100 50830 24110 50910
rect 24280 50830 24290 50910
rect 24460 50830 24470 50910
rect 24640 50830 24650 50910
rect 24820 50830 24830 50910
rect 25000 50830 25010 50910
rect 25180 50830 25190 50910
rect 25360 50830 25370 50910
rect 25540 50830 25550 50910
rect 25720 50830 25730 50910
rect 26300 50880 26360 50910
rect 26420 50880 26480 50910
rect 26540 50880 26600 50910
rect 30300 50880 30360 50910
rect 30420 50880 30480 50910
rect 30540 50880 30600 50910
rect 31260 50850 31270 50910
rect 31440 50850 31450 50910
rect 31620 50850 31630 50910
rect 31800 50850 31810 50910
rect 31980 50850 31990 50910
rect 32160 50850 32170 50910
rect 32340 50850 32350 50910
rect 32520 50850 32530 50910
rect 32700 50850 32710 50910
rect 32880 50850 32890 50910
rect 33060 50850 33070 50910
rect 33240 50850 33250 50910
rect 33420 50850 33430 50910
rect 33600 50850 33610 50910
rect 33780 50850 33790 50910
rect 33960 50850 33970 50910
rect 34140 50850 34150 50910
rect 34320 50850 34330 50910
rect 34500 50850 34510 50910
rect 34680 50850 34690 50910
rect 34860 50850 34870 50910
rect 35040 50850 35050 50910
rect 35220 50850 35230 50910
rect 35400 50850 35410 50910
rect 35580 50850 35590 50910
rect 35760 50850 35770 50910
rect 35940 50850 35950 50910
rect 36120 50850 36130 50910
rect 36300 50850 36310 50910
rect 36480 50850 36490 50910
rect 36660 50850 36670 50910
rect 36840 50850 36850 50910
rect 37020 50850 37030 50910
rect 37100 50850 37190 50920
rect 37720 50910 37750 50940
rect 37840 50910 37870 50940
rect 37600 50880 37660 50910
rect 37720 50880 37780 50910
rect 37840 50880 37900 50910
rect 31100 50820 37190 50850
rect 40060 50830 40120 50860
rect 19130 50790 19160 50820
rect 19250 50790 19280 50820
rect 26420 50790 26450 50820
rect 26540 50790 26570 50820
rect 30420 50790 30450 50820
rect 30540 50790 30570 50820
rect 19010 50760 19070 50790
rect 19130 50760 19190 50790
rect 19250 50760 19310 50790
rect 19880 50760 19960 50770
rect 20060 50760 20140 50770
rect 20240 50760 20320 50770
rect 20420 50760 20500 50770
rect 20600 50760 20680 50770
rect 20780 50760 20860 50770
rect 20960 50760 21040 50770
rect 21140 50760 21220 50770
rect 21320 50760 21400 50770
rect 21500 50760 21580 50770
rect 21680 50760 21760 50770
rect 21860 50760 21940 50770
rect 22040 50760 22120 50770
rect 22220 50760 22300 50770
rect 22400 50760 22480 50770
rect 22580 50760 22660 50770
rect 22760 50760 22840 50770
rect 22940 50760 23020 50770
rect 23120 50760 23200 50770
rect 23300 50760 23380 50770
rect 23480 50760 23560 50770
rect 23660 50760 23740 50770
rect 23840 50760 23920 50770
rect 24020 50760 24100 50770
rect 24200 50760 24280 50770
rect 24380 50760 24460 50770
rect 24560 50760 24640 50770
rect 24740 50760 24820 50770
rect 24920 50760 25000 50770
rect 25100 50760 25180 50770
rect 25280 50760 25360 50770
rect 25460 50760 25540 50770
rect 25640 50760 25720 50770
rect 26300 50760 26360 50790
rect 26420 50760 26480 50790
rect 26540 50760 26600 50790
rect 30300 50760 30360 50790
rect 30420 50760 30480 50790
rect 30540 50760 30600 50790
rect 31180 50760 31260 50770
rect 31360 50760 31440 50770
rect 31540 50760 31620 50770
rect 31720 50760 31800 50770
rect 31900 50760 31980 50770
rect 32080 50760 32160 50770
rect 32260 50760 32340 50770
rect 32440 50760 32520 50770
rect 32620 50760 32700 50770
rect 32800 50760 32880 50770
rect 32980 50760 33060 50770
rect 33160 50760 33240 50770
rect 33340 50760 33420 50770
rect 33520 50760 33600 50770
rect 33700 50760 33780 50770
rect 33880 50760 33960 50770
rect 34060 50760 34140 50770
rect 34240 50760 34320 50770
rect 34420 50760 34500 50770
rect 34600 50760 34680 50770
rect 34780 50760 34860 50770
rect 34960 50760 35040 50770
rect 35140 50760 35220 50770
rect 35320 50760 35400 50770
rect 35500 50760 35580 50770
rect 35680 50760 35760 50770
rect 35860 50760 35940 50770
rect 36040 50760 36120 50770
rect 36220 50760 36300 50770
rect 36400 50760 36480 50770
rect 36580 50760 36660 50770
rect 36760 50760 36840 50770
rect 36940 50760 37020 50770
rect 19130 50670 19160 50700
rect 19250 50670 19280 50700
rect 19960 50680 19970 50760
rect 20140 50680 20150 50760
rect 20320 50680 20330 50760
rect 20500 50680 20510 50760
rect 20680 50680 20690 50760
rect 20860 50680 20870 50760
rect 21040 50680 21050 50760
rect 21220 50680 21230 50760
rect 21400 50680 21410 50760
rect 21580 50680 21590 50760
rect 21760 50680 21770 50760
rect 21940 50680 21950 50760
rect 22120 50680 22130 50760
rect 22300 50680 22310 50760
rect 22480 50680 22490 50760
rect 22660 50680 22670 50760
rect 22840 50680 22850 50760
rect 23020 50680 23030 50760
rect 23200 50680 23210 50760
rect 23380 50680 23390 50760
rect 23560 50680 23570 50760
rect 23740 50680 23750 50760
rect 23920 50680 23930 50760
rect 24100 50680 24110 50760
rect 24280 50680 24290 50760
rect 24460 50680 24470 50760
rect 24640 50680 24650 50760
rect 24820 50680 24830 50760
rect 25000 50680 25010 50760
rect 25180 50680 25190 50760
rect 25360 50680 25370 50760
rect 25540 50680 25550 50760
rect 25720 50680 25730 50760
rect 26420 50670 26450 50700
rect 26540 50670 26570 50700
rect 30420 50670 30450 50700
rect 30540 50670 30570 50700
rect 31260 50680 31270 50760
rect 31440 50680 31450 50760
rect 31620 50680 31630 50760
rect 31800 50680 31810 50760
rect 31980 50680 31990 50760
rect 32160 50680 32170 50760
rect 32340 50680 32350 50760
rect 32520 50680 32530 50760
rect 32700 50680 32710 50760
rect 32880 50680 32890 50760
rect 33060 50680 33070 50760
rect 33240 50680 33250 50760
rect 33420 50680 33430 50760
rect 33600 50680 33610 50760
rect 33780 50680 33790 50760
rect 33960 50680 33970 50760
rect 34140 50680 34150 50760
rect 34320 50680 34330 50760
rect 34500 50680 34510 50760
rect 34680 50680 34690 50760
rect 34860 50680 34870 50760
rect 35040 50680 35050 50760
rect 35220 50680 35230 50760
rect 35400 50680 35410 50760
rect 35580 50680 35590 50760
rect 35760 50680 35770 50760
rect 35940 50680 35950 50760
rect 36120 50680 36130 50760
rect 36300 50680 36310 50760
rect 36480 50680 36490 50760
rect 36660 50680 36670 50760
rect 36840 50680 36850 50760
rect 37020 50680 37030 50760
rect 19010 50640 19070 50670
rect 19130 50640 19190 50670
rect 19250 50640 19310 50670
rect 26300 50640 26360 50670
rect 26420 50640 26480 50670
rect 26540 50640 26600 50670
rect 30300 50640 30360 50670
rect 30420 50640 30480 50670
rect 30540 50640 30600 50670
rect 37100 50620 37190 50820
rect 37720 50790 37750 50820
rect 37840 50790 37870 50820
rect 37600 50760 37660 50790
rect 37720 50760 37780 50790
rect 37840 50760 37900 50790
rect 40060 50710 40120 50740
rect 37720 50670 37750 50700
rect 37840 50670 37870 50700
rect 37600 50640 37660 50670
rect 37720 50640 37780 50670
rect 37840 50640 37900 50670
rect 19880 50610 19960 50620
rect 20060 50610 20140 50620
rect 20240 50610 20320 50620
rect 20420 50610 20500 50620
rect 20600 50610 20680 50620
rect 20780 50610 20860 50620
rect 20960 50610 21040 50620
rect 21140 50610 21220 50620
rect 21320 50610 21400 50620
rect 21500 50610 21580 50620
rect 21680 50610 21760 50620
rect 21860 50610 21940 50620
rect 22040 50610 22120 50620
rect 22220 50610 22300 50620
rect 22400 50610 22480 50620
rect 22580 50610 22660 50620
rect 22760 50610 22840 50620
rect 22940 50610 23020 50620
rect 23120 50610 23200 50620
rect 23300 50610 23380 50620
rect 23480 50610 23560 50620
rect 23660 50610 23740 50620
rect 23840 50610 23920 50620
rect 24020 50610 24100 50620
rect 24200 50610 24280 50620
rect 24380 50610 24460 50620
rect 24560 50610 24640 50620
rect 24740 50610 24820 50620
rect 24920 50610 25000 50620
rect 25100 50610 25180 50620
rect 25280 50610 25360 50620
rect 25460 50610 25540 50620
rect 25640 50610 25720 50620
rect 19130 50550 19160 50580
rect 19250 50550 19280 50580
rect 19010 50520 19070 50550
rect 19130 50520 19190 50550
rect 19250 50520 19310 50550
rect 19960 50530 19970 50610
rect 20140 50530 20150 50610
rect 20320 50530 20330 50610
rect 20500 50530 20510 50610
rect 20680 50530 20690 50610
rect 20860 50530 20870 50610
rect 21040 50530 21050 50610
rect 21220 50530 21230 50610
rect 21400 50530 21410 50610
rect 21580 50530 21590 50610
rect 21760 50530 21770 50610
rect 21940 50530 21950 50610
rect 22120 50530 22130 50610
rect 22300 50530 22310 50610
rect 22480 50530 22490 50610
rect 22660 50530 22670 50610
rect 22840 50530 22850 50610
rect 23020 50530 23030 50610
rect 23200 50530 23210 50610
rect 23380 50530 23390 50610
rect 23560 50530 23570 50610
rect 23740 50530 23750 50610
rect 23920 50530 23930 50610
rect 24100 50530 24110 50610
rect 24280 50530 24290 50610
rect 24460 50530 24470 50610
rect 24640 50530 24650 50610
rect 24820 50530 24830 50610
rect 25000 50530 25010 50610
rect 25180 50530 25190 50610
rect 25360 50530 25370 50610
rect 25540 50530 25550 50610
rect 25720 50530 25730 50610
rect 31100 50590 37190 50620
rect 40060 50590 40120 50620
rect 26420 50550 26450 50580
rect 26540 50550 26570 50580
rect 30420 50550 30450 50580
rect 30540 50550 30570 50580
rect 26300 50520 26360 50550
rect 26420 50520 26480 50550
rect 26540 50520 26600 50550
rect 30300 50520 30360 50550
rect 30420 50520 30480 50550
rect 30540 50520 30600 50550
rect 31260 50530 31270 50590
rect 31440 50530 31450 50590
rect 31620 50530 31630 50590
rect 31800 50530 31810 50590
rect 31980 50530 31990 50590
rect 32160 50530 32170 50590
rect 32340 50530 32350 50590
rect 32520 50530 32530 50590
rect 32700 50530 32710 50590
rect 32880 50530 32890 50590
rect 33060 50530 33070 50590
rect 33240 50530 33250 50590
rect 33420 50530 33430 50590
rect 33600 50530 33610 50590
rect 33780 50530 33790 50590
rect 33960 50530 33970 50590
rect 34140 50530 34150 50590
rect 34320 50530 34330 50590
rect 34500 50530 34510 50590
rect 34680 50530 34690 50590
rect 34860 50530 34870 50590
rect 35040 50530 35050 50590
rect 35220 50530 35230 50590
rect 35400 50530 35410 50590
rect 35580 50530 35590 50590
rect 35760 50530 35770 50590
rect 35940 50530 35950 50590
rect 36120 50530 36130 50590
rect 36300 50530 36310 50590
rect 36480 50530 36490 50590
rect 36660 50530 36670 50590
rect 36840 50530 36850 50590
rect 37020 50530 37030 50590
rect 37100 50520 37190 50590
rect 37720 50550 37750 50580
rect 37840 50550 37870 50580
rect 37600 50520 37660 50550
rect 37720 50520 37780 50550
rect 37840 50520 37900 50550
rect 31100 50490 37190 50520
rect 37100 50480 37190 50490
rect 19800 50470 25800 50480
rect 31100 50470 37190 50480
rect 40060 50470 40120 50500
rect 19130 50430 19160 50460
rect 19250 50430 19280 50460
rect 26420 50430 26450 50460
rect 26540 50430 26570 50460
rect 30420 50430 30450 50460
rect 30540 50430 30570 50460
rect 19010 50400 19070 50430
rect 19130 50400 19190 50430
rect 19250 50400 19310 50430
rect 26300 50400 26360 50430
rect 26420 50400 26480 50430
rect 26540 50400 26600 50430
rect 30300 50400 30360 50430
rect 30420 50400 30480 50430
rect 30540 50400 30600 50430
rect 19130 50310 19160 50340
rect 19250 50310 19280 50340
rect 26420 50310 26450 50340
rect 26540 50310 26570 50340
rect 30420 50310 30450 50340
rect 30540 50310 30570 50340
rect 19010 50280 19070 50310
rect 19130 50280 19190 50310
rect 19250 50280 19310 50310
rect 26300 50280 26360 50310
rect 26420 50280 26480 50310
rect 26540 50280 26600 50310
rect 30300 50280 30360 50310
rect 30420 50280 30480 50310
rect 30540 50280 30600 50310
rect 31180 50290 31260 50300
rect 31360 50290 31440 50300
rect 31540 50290 31620 50300
rect 31720 50290 31800 50300
rect 31900 50290 31980 50300
rect 32080 50290 32160 50300
rect 32260 50290 32340 50300
rect 32440 50290 32520 50300
rect 32620 50290 32700 50300
rect 32800 50290 32880 50300
rect 32980 50290 33060 50300
rect 33160 50290 33240 50300
rect 33340 50290 33420 50300
rect 33520 50290 33600 50300
rect 33700 50290 33780 50300
rect 33880 50290 33960 50300
rect 34060 50290 34140 50300
rect 34240 50290 34320 50300
rect 34420 50290 34500 50300
rect 34600 50290 34680 50300
rect 34780 50290 34860 50300
rect 34960 50290 35040 50300
rect 35140 50290 35220 50300
rect 35320 50290 35400 50300
rect 35500 50290 35580 50300
rect 35680 50290 35760 50300
rect 35860 50290 35940 50300
rect 36040 50290 36120 50300
rect 36220 50290 36300 50300
rect 36400 50290 36480 50300
rect 36580 50290 36660 50300
rect 36760 50290 36840 50300
rect 36940 50290 37020 50300
rect 19880 50270 19960 50280
rect 20060 50270 20140 50280
rect 20240 50270 20320 50280
rect 20420 50270 20500 50280
rect 20600 50270 20680 50280
rect 20780 50270 20860 50280
rect 20960 50270 21040 50280
rect 21140 50270 21220 50280
rect 21320 50270 21400 50280
rect 21500 50270 21580 50280
rect 21680 50270 21760 50280
rect 21860 50270 21940 50280
rect 22040 50270 22120 50280
rect 22220 50270 22300 50280
rect 22400 50270 22480 50280
rect 22580 50270 22660 50280
rect 22760 50270 22840 50280
rect 22940 50270 23020 50280
rect 23120 50270 23200 50280
rect 23300 50270 23380 50280
rect 23480 50270 23560 50280
rect 23660 50270 23740 50280
rect 23840 50270 23920 50280
rect 24020 50270 24100 50280
rect 24200 50270 24280 50280
rect 24380 50270 24460 50280
rect 24560 50270 24640 50280
rect 24740 50270 24820 50280
rect 24920 50270 25000 50280
rect 25100 50270 25180 50280
rect 25280 50270 25360 50280
rect 25460 50270 25540 50280
rect 25640 50270 25720 50280
rect 19130 50190 19160 50220
rect 19250 50190 19280 50220
rect 19960 50190 19970 50270
rect 20140 50190 20150 50270
rect 20320 50190 20330 50270
rect 20500 50190 20510 50270
rect 20680 50190 20690 50270
rect 20860 50190 20870 50270
rect 21040 50190 21050 50270
rect 21220 50190 21230 50270
rect 21400 50190 21410 50270
rect 21580 50190 21590 50270
rect 21760 50190 21770 50270
rect 21940 50190 21950 50270
rect 22120 50190 22130 50270
rect 22300 50190 22310 50270
rect 22480 50190 22490 50270
rect 22660 50190 22670 50270
rect 22840 50190 22850 50270
rect 23020 50190 23030 50270
rect 23200 50190 23210 50270
rect 23380 50190 23390 50270
rect 23560 50190 23570 50270
rect 23740 50190 23750 50270
rect 23920 50190 23930 50270
rect 24100 50190 24110 50270
rect 24280 50190 24290 50270
rect 24460 50190 24470 50270
rect 24640 50190 24650 50270
rect 24820 50190 24830 50270
rect 25000 50190 25010 50270
rect 25180 50190 25190 50270
rect 25360 50190 25370 50270
rect 25540 50190 25550 50270
rect 25720 50190 25730 50270
rect 26420 50190 26450 50220
rect 26540 50190 26570 50220
rect 30420 50190 30450 50220
rect 30540 50190 30570 50220
rect 31260 50210 31270 50290
rect 31440 50210 31450 50290
rect 31620 50210 31630 50290
rect 31800 50210 31810 50290
rect 31980 50210 31990 50290
rect 32160 50210 32170 50290
rect 32340 50210 32350 50290
rect 32520 50210 32530 50290
rect 32700 50210 32710 50290
rect 32880 50210 32890 50290
rect 33060 50210 33070 50290
rect 33240 50210 33250 50290
rect 33420 50210 33430 50290
rect 33600 50210 33610 50290
rect 33780 50210 33790 50290
rect 33960 50210 33970 50290
rect 34140 50210 34150 50290
rect 34320 50210 34330 50290
rect 34500 50210 34510 50290
rect 34680 50210 34690 50290
rect 34860 50210 34870 50290
rect 35040 50210 35050 50290
rect 35220 50210 35230 50290
rect 35400 50210 35410 50290
rect 35580 50210 35590 50290
rect 35760 50210 35770 50290
rect 35940 50210 35950 50290
rect 36120 50210 36130 50290
rect 36300 50210 36310 50290
rect 36480 50210 36490 50290
rect 36660 50210 36670 50290
rect 36840 50210 36850 50290
rect 37020 50210 37030 50290
rect 19010 50160 19070 50190
rect 19130 50160 19190 50190
rect 19250 50160 19310 50190
rect 26300 50160 26360 50190
rect 26420 50160 26480 50190
rect 26540 50160 26600 50190
rect 30300 50160 30360 50190
rect 30420 50160 30480 50190
rect 30540 50160 30600 50190
rect 19130 50070 19160 50100
rect 19250 50070 19280 50100
rect 26420 50070 26450 50100
rect 26540 50070 26570 50100
rect 30420 50070 30450 50100
rect 30540 50070 30570 50100
rect 19010 50040 19070 50070
rect 19130 50040 19190 50070
rect 19250 50040 19310 50070
rect 26300 50040 26360 50070
rect 26420 50040 26480 50070
rect 26540 50040 26600 50070
rect 30300 50040 30360 50070
rect 30420 50040 30480 50070
rect 30540 50040 30600 50070
rect 19130 49950 19160 49980
rect 19250 49950 19280 49980
rect 19880 49970 19960 49980
rect 20060 49970 20140 49980
rect 20240 49970 20320 49980
rect 20420 49970 20500 49980
rect 20600 49970 20680 49980
rect 20780 49970 20860 49980
rect 20960 49970 21040 49980
rect 21140 49970 21220 49980
rect 21320 49970 21400 49980
rect 21500 49970 21580 49980
rect 21680 49970 21760 49980
rect 21860 49970 21940 49980
rect 22040 49970 22120 49980
rect 22220 49970 22300 49980
rect 22400 49970 22480 49980
rect 22580 49970 22660 49980
rect 22760 49970 22840 49980
rect 22940 49970 23020 49980
rect 23120 49970 23200 49980
rect 23300 49970 23380 49980
rect 23480 49970 23560 49980
rect 23660 49970 23740 49980
rect 23840 49970 23920 49980
rect 24020 49970 24100 49980
rect 24200 49970 24280 49980
rect 24380 49970 24460 49980
rect 24560 49970 24640 49980
rect 24740 49970 24820 49980
rect 24920 49970 25000 49980
rect 25100 49970 25180 49980
rect 25280 49970 25360 49980
rect 25460 49970 25540 49980
rect 25640 49970 25720 49980
rect 19010 49920 19070 49950
rect 19130 49920 19190 49950
rect 19250 49920 19310 49950
rect 19960 49890 19970 49970
rect 20140 49890 20150 49970
rect 20320 49890 20330 49970
rect 20500 49890 20510 49970
rect 20680 49890 20690 49970
rect 20860 49890 20870 49970
rect 21040 49890 21050 49970
rect 21220 49890 21230 49970
rect 21400 49890 21410 49970
rect 21580 49890 21590 49970
rect 21760 49890 21770 49970
rect 21940 49890 21950 49970
rect 22120 49890 22130 49970
rect 22300 49890 22310 49970
rect 22480 49890 22490 49970
rect 22660 49890 22670 49970
rect 22840 49890 22850 49970
rect 23020 49890 23030 49970
rect 23200 49890 23210 49970
rect 23380 49890 23390 49970
rect 23560 49890 23570 49970
rect 23740 49890 23750 49970
rect 23920 49890 23930 49970
rect 24100 49890 24110 49970
rect 24280 49890 24290 49970
rect 24460 49890 24470 49970
rect 24640 49890 24650 49970
rect 24820 49890 24830 49970
rect 25000 49890 25010 49970
rect 25180 49890 25190 49970
rect 25360 49890 25370 49970
rect 25540 49890 25550 49970
rect 25720 49890 25730 49970
rect 26420 49950 26450 49980
rect 26540 49950 26570 49980
rect 30420 49950 30450 49980
rect 30540 49950 30570 49980
rect 31180 49970 31260 49980
rect 31360 49970 31440 49980
rect 31540 49970 31620 49980
rect 31720 49970 31800 49980
rect 31900 49970 31980 49980
rect 32080 49970 32160 49980
rect 32260 49970 32340 49980
rect 32440 49970 32520 49980
rect 32620 49970 32700 49980
rect 32800 49970 32880 49980
rect 32980 49970 33060 49980
rect 33160 49970 33240 49980
rect 33340 49970 33420 49980
rect 33520 49970 33600 49980
rect 33700 49970 33780 49980
rect 33880 49970 33960 49980
rect 34060 49970 34140 49980
rect 34240 49970 34320 49980
rect 34420 49970 34500 49980
rect 34600 49970 34680 49980
rect 34780 49970 34860 49980
rect 34960 49970 35040 49980
rect 35140 49970 35220 49980
rect 35320 49970 35400 49980
rect 35500 49970 35580 49980
rect 35680 49970 35760 49980
rect 35860 49970 35940 49980
rect 36040 49970 36120 49980
rect 36220 49970 36300 49980
rect 36400 49970 36480 49980
rect 36580 49970 36660 49980
rect 36760 49970 36840 49980
rect 36940 49970 37020 49980
rect 26300 49920 26360 49950
rect 26420 49920 26480 49950
rect 26540 49920 26600 49950
rect 30300 49920 30360 49950
rect 30420 49920 30480 49950
rect 30540 49920 30600 49950
rect 31260 49890 31270 49970
rect 31440 49890 31450 49970
rect 31620 49890 31630 49970
rect 31800 49890 31810 49970
rect 31980 49890 31990 49970
rect 32160 49890 32170 49970
rect 32340 49890 32350 49970
rect 32520 49890 32530 49970
rect 32700 49890 32710 49970
rect 32880 49890 32890 49970
rect 33060 49890 33070 49970
rect 33240 49890 33250 49970
rect 33420 49890 33430 49970
rect 33600 49890 33610 49970
rect 33780 49890 33790 49970
rect 33960 49890 33970 49970
rect 34140 49890 34150 49970
rect 34320 49890 34330 49970
rect 34500 49890 34510 49970
rect 34680 49890 34690 49970
rect 34860 49890 34870 49970
rect 35040 49890 35050 49970
rect 35220 49890 35230 49970
rect 35400 49890 35410 49970
rect 35580 49890 35590 49970
rect 35760 49890 35770 49970
rect 35940 49890 35950 49970
rect 36120 49890 36130 49970
rect 36300 49890 36310 49970
rect 36480 49890 36490 49970
rect 36660 49890 36670 49970
rect 36840 49890 36850 49970
rect 37020 49890 37030 49970
rect 19130 49830 19160 49860
rect 19250 49830 19280 49860
rect 26420 49830 26450 49860
rect 26540 49830 26570 49860
rect 30420 49830 30450 49860
rect 30540 49830 30570 49860
rect 19010 49800 19070 49830
rect 19130 49800 19190 49830
rect 19250 49800 19310 49830
rect 26300 49800 26360 49830
rect 26420 49800 26480 49830
rect 26540 49800 26600 49830
rect 30300 49800 30360 49830
rect 30420 49800 30480 49830
rect 30540 49800 30600 49830
rect 37100 49800 37190 50470
rect 37720 50430 37750 50460
rect 37840 50430 37870 50460
rect 37600 50400 37660 50430
rect 37720 50400 37780 50430
rect 37840 50400 37900 50430
rect 40060 50350 40120 50380
rect 37720 50310 37750 50340
rect 37840 50310 37870 50340
rect 37600 50280 37660 50310
rect 37720 50280 37780 50310
rect 37840 50280 37900 50310
rect 40060 50230 40120 50260
rect 37720 50190 37750 50220
rect 37840 50190 37870 50220
rect 37600 50160 37660 50190
rect 37720 50160 37780 50190
rect 37840 50160 37900 50190
rect 40060 50110 40120 50140
rect 37720 50070 37750 50100
rect 37840 50070 37870 50100
rect 37600 50040 37660 50070
rect 37720 50040 37780 50070
rect 37840 50040 37900 50070
rect 40060 49990 40120 50020
rect 37720 49950 37750 49980
rect 37840 49950 37870 49980
rect 37600 49920 37660 49950
rect 37720 49920 37780 49950
rect 37840 49920 37900 49950
rect 40060 49870 40120 49900
rect 37720 49830 37750 49860
rect 37840 49830 37870 49860
rect 37600 49800 37660 49830
rect 37720 49800 37780 49830
rect 37840 49800 37900 49830
rect 19800 49790 25800 49800
rect 31100 49790 37190 49800
rect 19130 49710 19160 49740
rect 19250 49710 19280 49740
rect 26420 49710 26450 49740
rect 26540 49710 26570 49740
rect 30420 49710 30450 49740
rect 30540 49710 30570 49740
rect 19010 49680 19070 49710
rect 19130 49680 19190 49710
rect 19250 49680 19310 49710
rect 26300 49680 26360 49710
rect 26420 49680 26480 49710
rect 26540 49680 26600 49710
rect 30300 49680 30360 49710
rect 30420 49680 30480 49710
rect 30540 49680 30600 49710
rect 37100 49690 37190 49790
rect 40060 49750 40120 49780
rect 37720 49710 37750 49740
rect 37840 49710 37870 49740
rect 31100 49660 37190 49690
rect 37600 49680 37660 49710
rect 37720 49680 37780 49710
rect 37840 49680 37900 49710
rect 19880 49650 19960 49660
rect 20060 49650 20140 49660
rect 20240 49650 20320 49660
rect 20420 49650 20500 49660
rect 20600 49650 20680 49660
rect 20780 49650 20860 49660
rect 20960 49650 21040 49660
rect 21140 49650 21220 49660
rect 21320 49650 21400 49660
rect 21500 49650 21580 49660
rect 21680 49650 21760 49660
rect 21860 49650 21940 49660
rect 22040 49650 22120 49660
rect 22220 49650 22300 49660
rect 22400 49650 22480 49660
rect 22580 49650 22660 49660
rect 22760 49650 22840 49660
rect 22940 49650 23020 49660
rect 23120 49650 23200 49660
rect 23300 49650 23380 49660
rect 23480 49650 23560 49660
rect 23660 49650 23740 49660
rect 23840 49650 23920 49660
rect 24020 49650 24100 49660
rect 24200 49650 24280 49660
rect 24380 49650 24460 49660
rect 24560 49650 24640 49660
rect 24740 49650 24820 49660
rect 24920 49650 25000 49660
rect 25100 49650 25180 49660
rect 25280 49650 25360 49660
rect 25460 49650 25540 49660
rect 25640 49650 25720 49660
rect 31180 49650 31260 49660
rect 31360 49650 31440 49660
rect 31540 49650 31620 49660
rect 31720 49650 31800 49660
rect 31900 49650 31980 49660
rect 32080 49650 32160 49660
rect 32260 49650 32340 49660
rect 32440 49650 32520 49660
rect 32620 49650 32700 49660
rect 32800 49650 32880 49660
rect 32980 49650 33060 49660
rect 33160 49650 33240 49660
rect 33340 49650 33420 49660
rect 33520 49650 33600 49660
rect 33700 49650 33780 49660
rect 33880 49650 33960 49660
rect 34060 49650 34140 49660
rect 34240 49650 34320 49660
rect 34420 49650 34500 49660
rect 34600 49650 34680 49660
rect 34780 49650 34860 49660
rect 34960 49650 35040 49660
rect 35140 49650 35220 49660
rect 35320 49650 35400 49660
rect 35500 49650 35580 49660
rect 35680 49650 35760 49660
rect 35860 49650 35940 49660
rect 36040 49650 36120 49660
rect 36220 49650 36300 49660
rect 36400 49650 36480 49660
rect 36580 49650 36660 49660
rect 36760 49650 36840 49660
rect 36940 49650 37020 49660
rect 19130 49590 19160 49620
rect 19250 49590 19280 49620
rect 19010 49560 19070 49590
rect 19130 49560 19190 49590
rect 19250 49560 19310 49590
rect 19960 49570 19970 49650
rect 20140 49570 20150 49650
rect 20320 49570 20330 49650
rect 20500 49570 20510 49650
rect 20680 49570 20690 49650
rect 20860 49570 20870 49650
rect 21040 49570 21050 49650
rect 21220 49570 21230 49650
rect 21400 49570 21410 49650
rect 21580 49570 21590 49650
rect 21760 49570 21770 49650
rect 21940 49570 21950 49650
rect 22120 49570 22130 49650
rect 22300 49570 22310 49650
rect 22480 49570 22490 49650
rect 22660 49570 22670 49650
rect 22840 49570 22850 49650
rect 23020 49570 23030 49650
rect 23200 49570 23210 49650
rect 23380 49570 23390 49650
rect 23560 49570 23570 49650
rect 23740 49570 23750 49650
rect 23920 49570 23930 49650
rect 24100 49570 24110 49650
rect 24280 49570 24290 49650
rect 24460 49570 24470 49650
rect 24640 49570 24650 49650
rect 24820 49570 24830 49650
rect 25000 49570 25010 49650
rect 25180 49570 25190 49650
rect 25360 49570 25370 49650
rect 25540 49570 25550 49650
rect 25720 49570 25730 49650
rect 26420 49590 26450 49620
rect 26540 49590 26570 49620
rect 30420 49590 30450 49620
rect 30540 49590 30570 49620
rect 31260 49590 31270 49650
rect 31440 49590 31450 49650
rect 31620 49590 31630 49650
rect 31800 49590 31810 49650
rect 31980 49590 31990 49650
rect 32160 49590 32170 49650
rect 32340 49590 32350 49650
rect 32520 49590 32530 49650
rect 32700 49590 32710 49650
rect 32880 49590 32890 49650
rect 33060 49590 33070 49650
rect 33240 49590 33250 49650
rect 33420 49590 33430 49650
rect 33600 49590 33610 49650
rect 33780 49590 33790 49650
rect 33960 49590 33970 49650
rect 34140 49590 34150 49650
rect 34320 49590 34330 49650
rect 34500 49590 34510 49650
rect 34680 49590 34690 49650
rect 34860 49590 34870 49650
rect 35040 49590 35050 49650
rect 35220 49590 35230 49650
rect 35400 49590 35410 49650
rect 35580 49590 35590 49650
rect 35760 49590 35770 49650
rect 35940 49590 35950 49650
rect 36120 49590 36130 49650
rect 36300 49590 36310 49650
rect 36480 49590 36490 49650
rect 36660 49590 36670 49650
rect 36840 49590 36850 49650
rect 37020 49590 37030 49650
rect 37100 49590 37190 49660
rect 40060 49630 40120 49660
rect 37720 49590 37750 49620
rect 37840 49590 37870 49620
rect 26300 49560 26360 49590
rect 26420 49560 26480 49590
rect 26540 49560 26600 49590
rect 30300 49560 30360 49590
rect 30420 49560 30480 49590
rect 30540 49560 30600 49590
rect 31100 49560 37190 49590
rect 37600 49560 37660 49590
rect 37720 49560 37780 49590
rect 37840 49560 37900 49590
rect 19880 49500 19960 49510
rect 20060 49500 20140 49510
rect 20240 49500 20320 49510
rect 20420 49500 20500 49510
rect 20600 49500 20680 49510
rect 20780 49500 20860 49510
rect 20960 49500 21040 49510
rect 21140 49500 21220 49510
rect 21320 49500 21400 49510
rect 21500 49500 21580 49510
rect 21680 49500 21760 49510
rect 21860 49500 21940 49510
rect 22040 49500 22120 49510
rect 22220 49500 22300 49510
rect 22400 49500 22480 49510
rect 22580 49500 22660 49510
rect 22760 49500 22840 49510
rect 22940 49500 23020 49510
rect 23120 49500 23200 49510
rect 23300 49500 23380 49510
rect 23480 49500 23560 49510
rect 23660 49500 23740 49510
rect 23840 49500 23920 49510
rect 24020 49500 24100 49510
rect 24200 49500 24280 49510
rect 24380 49500 24460 49510
rect 24560 49500 24640 49510
rect 24740 49500 24820 49510
rect 24920 49500 25000 49510
rect 25100 49500 25180 49510
rect 25280 49500 25360 49510
rect 25460 49500 25540 49510
rect 25640 49500 25720 49510
rect 31180 49500 31260 49510
rect 31360 49500 31440 49510
rect 31540 49500 31620 49510
rect 31720 49500 31800 49510
rect 31900 49500 31980 49510
rect 32080 49500 32160 49510
rect 32260 49500 32340 49510
rect 32440 49500 32520 49510
rect 32620 49500 32700 49510
rect 32800 49500 32880 49510
rect 32980 49500 33060 49510
rect 33160 49500 33240 49510
rect 33340 49500 33420 49510
rect 33520 49500 33600 49510
rect 33700 49500 33780 49510
rect 33880 49500 33960 49510
rect 34060 49500 34140 49510
rect 34240 49500 34320 49510
rect 34420 49500 34500 49510
rect 34600 49500 34680 49510
rect 34780 49500 34860 49510
rect 34960 49500 35040 49510
rect 35140 49500 35220 49510
rect 35320 49500 35400 49510
rect 35500 49500 35580 49510
rect 35680 49500 35760 49510
rect 35860 49500 35940 49510
rect 36040 49500 36120 49510
rect 36220 49500 36300 49510
rect 36400 49500 36480 49510
rect 36580 49500 36660 49510
rect 36760 49500 36840 49510
rect 36940 49500 37020 49510
rect 19130 49470 19160 49500
rect 19250 49470 19280 49500
rect 19010 49440 19070 49470
rect 19130 49440 19190 49470
rect 19250 49440 19310 49470
rect 19960 49420 19970 49500
rect 20140 49420 20150 49500
rect 20320 49420 20330 49500
rect 20500 49420 20510 49500
rect 20680 49420 20690 49500
rect 20860 49420 20870 49500
rect 21040 49420 21050 49500
rect 21220 49420 21230 49500
rect 21400 49420 21410 49500
rect 21580 49420 21590 49500
rect 21760 49420 21770 49500
rect 21940 49420 21950 49500
rect 22120 49420 22130 49500
rect 22300 49420 22310 49500
rect 22480 49420 22490 49500
rect 22660 49420 22670 49500
rect 22840 49420 22850 49500
rect 23020 49420 23030 49500
rect 23200 49420 23210 49500
rect 23380 49420 23390 49500
rect 23560 49420 23570 49500
rect 23740 49420 23750 49500
rect 23920 49420 23930 49500
rect 24100 49420 24110 49500
rect 24280 49420 24290 49500
rect 24460 49420 24470 49500
rect 24640 49420 24650 49500
rect 24820 49420 24830 49500
rect 25000 49420 25010 49500
rect 25180 49420 25190 49500
rect 25360 49420 25370 49500
rect 25540 49420 25550 49500
rect 25720 49420 25730 49500
rect 26420 49470 26450 49500
rect 26540 49470 26570 49500
rect 30420 49470 30450 49500
rect 30540 49470 30570 49500
rect 26300 49440 26360 49470
rect 26420 49440 26480 49470
rect 26540 49440 26600 49470
rect 30300 49440 30360 49470
rect 30420 49440 30480 49470
rect 30540 49440 30600 49470
rect 31260 49420 31270 49500
rect 31440 49420 31450 49500
rect 31620 49420 31630 49500
rect 31800 49420 31810 49500
rect 31980 49420 31990 49500
rect 32160 49420 32170 49500
rect 32340 49420 32350 49500
rect 32520 49420 32530 49500
rect 32700 49420 32710 49500
rect 32880 49420 32890 49500
rect 33060 49420 33070 49500
rect 33240 49420 33250 49500
rect 33420 49420 33430 49500
rect 33600 49420 33610 49500
rect 33780 49420 33790 49500
rect 33960 49420 33970 49500
rect 34140 49420 34150 49500
rect 34320 49420 34330 49500
rect 34500 49420 34510 49500
rect 34680 49420 34690 49500
rect 34860 49420 34870 49500
rect 35040 49420 35050 49500
rect 35220 49420 35230 49500
rect 35400 49420 35410 49500
rect 35580 49420 35590 49500
rect 35760 49420 35770 49500
rect 35940 49420 35950 49500
rect 36120 49420 36130 49500
rect 36300 49420 36310 49500
rect 36480 49420 36490 49500
rect 36660 49420 36670 49500
rect 36840 49420 36850 49500
rect 37020 49420 37030 49500
rect 19130 49350 19160 49380
rect 19250 49350 19280 49380
rect 19880 49350 19960 49360
rect 20060 49350 20140 49360
rect 20240 49350 20320 49360
rect 20420 49350 20500 49360
rect 20600 49350 20680 49360
rect 20780 49350 20860 49360
rect 20960 49350 21040 49360
rect 21140 49350 21220 49360
rect 21320 49350 21400 49360
rect 21500 49350 21580 49360
rect 21680 49350 21760 49360
rect 21860 49350 21940 49360
rect 22040 49350 22120 49360
rect 22220 49350 22300 49360
rect 22400 49350 22480 49360
rect 22580 49350 22660 49360
rect 22760 49350 22840 49360
rect 22940 49350 23020 49360
rect 23120 49350 23200 49360
rect 23300 49350 23380 49360
rect 23480 49350 23560 49360
rect 23660 49350 23740 49360
rect 23840 49350 23920 49360
rect 24020 49350 24100 49360
rect 24200 49350 24280 49360
rect 24380 49350 24460 49360
rect 24560 49350 24640 49360
rect 24740 49350 24820 49360
rect 24920 49350 25000 49360
rect 25100 49350 25180 49360
rect 25280 49350 25360 49360
rect 25460 49350 25540 49360
rect 25640 49350 25720 49360
rect 26420 49350 26450 49380
rect 26540 49350 26570 49380
rect 30420 49350 30450 49380
rect 30540 49350 30570 49380
rect 31180 49350 31260 49360
rect 31360 49350 31440 49360
rect 31540 49350 31620 49360
rect 31720 49350 31800 49360
rect 31900 49350 31980 49360
rect 32080 49350 32160 49360
rect 32260 49350 32340 49360
rect 32440 49350 32520 49360
rect 32620 49350 32700 49360
rect 32800 49350 32880 49360
rect 32980 49350 33060 49360
rect 33160 49350 33240 49360
rect 33340 49350 33420 49360
rect 33520 49350 33600 49360
rect 33700 49350 33780 49360
rect 33880 49350 33960 49360
rect 34060 49350 34140 49360
rect 34240 49350 34320 49360
rect 34420 49350 34500 49360
rect 34600 49350 34680 49360
rect 34780 49350 34860 49360
rect 34960 49350 35040 49360
rect 35140 49350 35220 49360
rect 35320 49350 35400 49360
rect 35500 49350 35580 49360
rect 35680 49350 35760 49360
rect 35860 49350 35940 49360
rect 36040 49350 36120 49360
rect 36220 49350 36300 49360
rect 36400 49350 36480 49360
rect 36580 49350 36660 49360
rect 36760 49350 36840 49360
rect 36940 49350 37020 49360
rect 19010 49320 19070 49350
rect 19130 49320 19190 49350
rect 19250 49320 19310 49350
rect 19960 49270 19970 49350
rect 20140 49270 20150 49350
rect 20320 49270 20330 49350
rect 20500 49270 20510 49350
rect 20680 49270 20690 49350
rect 20860 49270 20870 49350
rect 21040 49270 21050 49350
rect 21220 49270 21230 49350
rect 21400 49270 21410 49350
rect 21580 49270 21590 49350
rect 21760 49270 21770 49350
rect 21940 49270 21950 49350
rect 22120 49270 22130 49350
rect 22300 49270 22310 49350
rect 22480 49270 22490 49350
rect 22660 49270 22670 49350
rect 22840 49270 22850 49350
rect 23020 49270 23030 49350
rect 23200 49270 23210 49350
rect 23380 49270 23390 49350
rect 23560 49270 23570 49350
rect 23740 49270 23750 49350
rect 23920 49270 23930 49350
rect 24100 49270 24110 49350
rect 24280 49270 24290 49350
rect 24460 49270 24470 49350
rect 24640 49270 24650 49350
rect 24820 49270 24830 49350
rect 25000 49270 25010 49350
rect 25180 49270 25190 49350
rect 25360 49270 25370 49350
rect 25540 49270 25550 49350
rect 25720 49270 25730 49350
rect 26300 49320 26360 49350
rect 26420 49320 26480 49350
rect 26540 49320 26600 49350
rect 30300 49320 30360 49350
rect 30420 49320 30480 49350
rect 30540 49320 30600 49350
rect 31260 49270 31270 49350
rect 31440 49270 31450 49350
rect 31620 49270 31630 49350
rect 31800 49270 31810 49350
rect 31980 49270 31990 49350
rect 32160 49270 32170 49350
rect 32340 49270 32350 49350
rect 32520 49270 32530 49350
rect 32700 49270 32710 49350
rect 32880 49270 32890 49350
rect 33060 49270 33070 49350
rect 33240 49270 33250 49350
rect 33420 49270 33430 49350
rect 33600 49270 33610 49350
rect 33780 49270 33790 49350
rect 33960 49270 33970 49350
rect 34140 49270 34150 49350
rect 34320 49270 34330 49350
rect 34500 49270 34510 49350
rect 34680 49270 34690 49350
rect 34860 49270 34870 49350
rect 35040 49270 35050 49350
rect 35220 49270 35230 49350
rect 35400 49270 35410 49350
rect 35580 49270 35590 49350
rect 35760 49270 35770 49350
rect 35940 49270 35950 49350
rect 36120 49270 36130 49350
rect 36300 49270 36310 49350
rect 36480 49270 36490 49350
rect 36660 49270 36670 49350
rect 36840 49270 36850 49350
rect 37020 49270 37030 49350
rect 37100 49330 37190 49560
rect 40060 49510 40120 49540
rect 37720 49470 37750 49500
rect 37840 49470 37870 49500
rect 37600 49440 37660 49470
rect 37720 49440 37780 49470
rect 37840 49440 37900 49470
rect 40060 49390 40120 49420
rect 37720 49350 37750 49380
rect 37840 49350 37870 49380
rect 37600 49320 37660 49350
rect 37720 49320 37780 49350
rect 37840 49320 37900 49350
rect 40060 49270 40120 49300
rect 19130 49200 19160 49260
rect 19250 49200 19280 49260
rect 26420 49200 26450 49260
rect 26540 49200 26570 49260
rect 30420 49230 30450 49260
rect 30540 49230 30570 49260
rect 37720 49230 37750 49260
rect 37840 49230 37870 49260
rect 30300 49200 30360 49230
rect 30420 49200 30480 49230
rect 30540 49200 30600 49230
rect 37600 49200 37660 49230
rect 37720 49200 37780 49230
rect 37840 49200 37900 49230
rect 40060 49150 40120 49180
rect 30420 49080 30450 49140
rect 30540 49080 30570 49140
rect 37720 49080 37750 49140
rect 37840 49080 37870 49140
rect 40060 49030 40120 49060
rect 18980 48940 19060 48950
rect 19160 48940 19240 48950
rect 19340 48940 19420 48950
rect 19520 48940 19600 48950
rect 19700 48940 19780 48950
rect 19880 48940 19960 48950
rect 20060 48940 20140 48950
rect 20240 48940 20320 48950
rect 20420 48940 20500 48950
rect 20600 48940 20680 48950
rect 20780 48940 20860 48950
rect 20960 48940 21040 48950
rect 21140 48940 21220 48950
rect 21320 48940 21400 48950
rect 21500 48940 21580 48950
rect 21680 48940 21760 48950
rect 21860 48940 21940 48950
rect 22040 48940 22120 48950
rect 22220 48940 22300 48950
rect 22400 48940 22480 48950
rect 22580 48940 22660 48950
rect 22760 48940 22840 48950
rect 22940 48940 23020 48950
rect 23120 48940 23200 48950
rect 23300 48940 23380 48950
rect 23480 48940 23560 48950
rect 23660 48940 23740 48950
rect 23840 48940 23920 48950
rect 24020 48940 24100 48950
rect 24200 48940 24280 48950
rect 24380 48940 24460 48950
rect 24560 48940 24640 48950
rect 24740 48940 24820 48950
rect 24920 48940 25000 48950
rect 25100 48940 25180 48950
rect 25280 48940 25360 48950
rect 25460 48940 25540 48950
rect 25640 48940 25720 48950
rect 25820 48940 25900 48950
rect 26000 48940 26080 48950
rect 26180 48940 26260 48950
rect 26360 48940 26440 48950
rect 26540 48940 26620 48950
rect 30280 48940 30360 48950
rect 30460 48940 30540 48950
rect 30640 48940 30720 48950
rect 30820 48940 30900 48950
rect 31000 48940 31080 48950
rect 31180 48940 31260 48950
rect 31360 48940 31440 48950
rect 31540 48940 31620 48950
rect 31720 48940 31800 48950
rect 31900 48940 31980 48950
rect 32080 48940 32160 48950
rect 32260 48940 32340 48950
rect 32440 48940 32520 48950
rect 32620 48940 32700 48950
rect 32800 48940 32880 48950
rect 32980 48940 33060 48950
rect 33160 48940 33240 48950
rect 33340 48940 33420 48950
rect 33520 48940 33600 48950
rect 33700 48940 33780 48950
rect 33880 48940 33960 48950
rect 34060 48940 34140 48950
rect 34240 48940 34320 48950
rect 34420 48940 34500 48950
rect 34600 48940 34680 48950
rect 34780 48940 34860 48950
rect 34960 48940 35040 48950
rect 35140 48940 35220 48950
rect 35320 48940 35400 48950
rect 35500 48940 35580 48950
rect 35680 48940 35760 48950
rect 35860 48940 35940 48950
rect 36040 48940 36120 48950
rect 36220 48940 36300 48950
rect 36400 48940 36480 48950
rect 36580 48940 36660 48950
rect 36760 48940 36840 48950
rect 36940 48940 37020 48950
rect 37120 48940 37200 48950
rect 37300 48940 37380 48950
rect 37480 48940 37560 48950
rect 37660 48940 37740 48950
rect 37840 48940 37920 48950
rect 40260 48940 40270 50940
rect 40380 50930 41180 51020
rect 152220 51010 152250 51040
rect 152340 51010 152370 51040
rect 152100 50980 152160 51010
rect 152220 50980 152280 51010
rect 152340 50980 152400 51010
rect 41540 50950 41600 50980
rect 42360 50950 42420 50980
rect 43840 50950 43900 50980
rect 158900 50950 158990 51050
rect 159520 51010 159550 51040
rect 159640 51010 159670 51040
rect 163520 51010 163550 51040
rect 163640 51010 163670 51040
rect 170810 51010 170840 51040
rect 170930 51010 170960 51040
rect 159400 50980 159460 51010
rect 159520 50980 159580 51010
rect 159640 50980 159700 51010
rect 163400 50980 163460 51010
rect 163520 50980 163580 51010
rect 163640 50980 163700 51010
rect 170690 50980 170750 51010
rect 170810 50980 170870 51010
rect 170930 50980 170990 51010
rect 40650 50900 40770 50930
rect 40930 50900 41050 50930
rect 41090 50900 41180 50930
rect 146100 50910 146160 50940
rect 147580 50910 147640 50940
rect 148400 50910 148460 50940
rect 149880 50910 149940 50940
rect 152900 50920 158990 50950
rect 40650 50810 40660 50900
rect 40760 50870 40830 50900
rect 40770 50780 40830 50870
rect 40930 50810 40940 50900
rect 41050 50780 41180 50900
rect 152220 50890 152250 50920
rect 152340 50890 152370 50920
rect 152980 50910 153060 50920
rect 153160 50910 153240 50920
rect 153340 50910 153420 50920
rect 153520 50910 153600 50920
rect 153700 50910 153780 50920
rect 153880 50910 153960 50920
rect 154060 50910 154140 50920
rect 154240 50910 154320 50920
rect 154420 50910 154500 50920
rect 154600 50910 154680 50920
rect 154780 50910 154860 50920
rect 154960 50910 155040 50920
rect 155140 50910 155220 50920
rect 155320 50910 155400 50920
rect 155500 50910 155580 50920
rect 155680 50910 155760 50920
rect 155860 50910 155940 50920
rect 156040 50910 156120 50920
rect 156220 50910 156300 50920
rect 156400 50910 156480 50920
rect 156580 50910 156660 50920
rect 156760 50910 156840 50920
rect 156940 50910 157020 50920
rect 157120 50910 157200 50920
rect 157300 50910 157380 50920
rect 157480 50910 157560 50920
rect 157660 50910 157740 50920
rect 157840 50910 157920 50920
rect 158020 50910 158100 50920
rect 158200 50910 158280 50920
rect 158380 50910 158460 50920
rect 158560 50910 158640 50920
rect 158740 50910 158820 50920
rect 41090 50745 41180 50780
rect 41230 50750 41350 50810
rect 40470 50740 41180 50745
rect 40370 50730 41180 50740
rect 40370 50650 40380 50730
rect 40470 50725 41180 50730
rect 40420 50715 41210 50725
rect 41090 50665 41180 50715
rect 40470 50650 41180 50665
rect 40460 50635 41180 50650
rect 40460 50445 40470 50635
rect 40650 50600 40770 50635
rect 40930 50600 41050 50635
rect 41090 50600 41180 50635
rect 41350 50630 41410 50750
rect 40770 50590 40830 50600
rect 40530 50580 40610 50590
rect 40670 50580 40750 50590
rect 40770 50580 40890 50590
rect 40950 50580 41030 50590
rect 40610 50500 40620 50580
rect 40750 50500 40760 50580
rect 40770 50480 40830 50580
rect 40890 50500 40900 50580
rect 41030 50500 41040 50580
rect 41050 50480 41180 50600
rect 41260 50580 41340 50590
rect 41340 50510 41350 50580
rect 41090 50445 41180 50480
rect 41230 50450 41350 50510
rect 40460 50430 41180 50445
rect 40470 50425 41180 50430
rect 40420 50415 41210 50425
rect 41090 50365 41180 50415
rect 40470 50335 41180 50365
rect 40650 50300 40770 50335
rect 40930 50300 41050 50335
rect 41090 50300 41180 50335
rect 41350 50330 41410 50450
rect 40650 50210 40660 50300
rect 40760 50270 40830 50300
rect 40770 50180 40830 50270
rect 40930 50210 40940 50300
rect 41050 50180 41180 50300
rect 41260 50280 41340 50290
rect 41340 50210 41350 50280
rect 41090 50145 41180 50180
rect 41230 50150 41350 50210
rect 40370 50130 40460 50140
rect 40370 50050 40380 50130
rect 40470 50125 41180 50145
rect 40420 50115 41210 50125
rect 41090 50065 41180 50115
rect 40470 50050 41180 50065
rect 40460 50035 41180 50050
rect 40460 49845 40470 50035
rect 40650 50000 40770 50035
rect 40930 50000 41050 50035
rect 41090 50000 41180 50035
rect 41350 50030 41410 50150
rect 40770 49990 40830 50000
rect 40530 49980 40610 49990
rect 40670 49980 40750 49990
rect 40770 49980 40890 49990
rect 40950 49980 41030 49990
rect 40610 49900 40620 49980
rect 40750 49900 40760 49980
rect 40770 49880 40830 49980
rect 40890 49900 40900 49980
rect 41030 49900 41040 49980
rect 41050 49880 41180 50000
rect 41260 49980 41340 49990
rect 41340 49910 41350 49980
rect 41090 49845 41180 49880
rect 41230 49850 41350 49910
rect 40460 49830 41180 49845
rect 40470 49825 41180 49830
rect 40420 49815 41210 49825
rect 41090 49765 41180 49815
rect 40470 49735 41180 49765
rect 40650 49700 40770 49735
rect 40930 49700 41050 49735
rect 41090 49700 41180 49735
rect 41350 49730 41410 49850
rect 40650 49610 40660 49700
rect 40760 49670 40830 49700
rect 40770 49580 40830 49670
rect 40930 49610 40940 49700
rect 41050 49580 41180 49700
rect 41260 49680 41340 49690
rect 41340 49610 41350 49680
rect 41090 49545 41180 49580
rect 41230 49550 41350 49610
rect 40370 49530 40460 49540
rect 40370 49450 40380 49530
rect 40470 49525 41180 49545
rect 40420 49515 41210 49525
rect 41090 49465 41180 49515
rect 40470 49450 41180 49465
rect 40460 49435 41180 49450
rect 40460 49245 40470 49435
rect 40650 49400 40770 49435
rect 40930 49400 41050 49435
rect 41090 49400 41180 49435
rect 41350 49430 41410 49550
rect 40770 49390 40830 49400
rect 40530 49380 40610 49390
rect 40670 49380 40750 49390
rect 40770 49380 40890 49390
rect 40950 49380 41030 49390
rect 40610 49300 40620 49380
rect 40750 49300 40760 49380
rect 40770 49280 40830 49380
rect 40890 49300 40900 49380
rect 41030 49300 41040 49380
rect 41050 49280 41180 49400
rect 41260 49370 41340 49380
rect 41340 49310 41350 49370
rect 41090 49245 41180 49280
rect 41230 49250 41350 49310
rect 40460 49230 41180 49245
rect 40470 49225 41180 49230
rect 40420 49215 41210 49225
rect 41090 49165 41180 49215
rect 40470 49135 41180 49165
rect 40650 49100 40770 49135
rect 40930 49100 41050 49135
rect 41090 49100 41180 49135
rect 41350 49130 41410 49250
rect 41480 49100 41490 50870
rect 152100 50860 152160 50890
rect 152220 50860 152280 50890
rect 152340 50860 152400 50890
rect 41540 50830 41600 50860
rect 42360 50830 42420 50860
rect 43840 50830 43900 50860
rect 153060 50850 153070 50910
rect 153240 50850 153250 50910
rect 153420 50850 153430 50910
rect 153600 50850 153610 50910
rect 153780 50850 153790 50910
rect 153960 50850 153970 50910
rect 154140 50850 154150 50910
rect 154320 50850 154330 50910
rect 154500 50850 154510 50910
rect 154680 50850 154690 50910
rect 154860 50850 154870 50910
rect 155040 50850 155050 50910
rect 155220 50850 155230 50910
rect 155400 50850 155410 50910
rect 155580 50850 155590 50910
rect 155760 50850 155770 50910
rect 155940 50850 155950 50910
rect 156120 50850 156130 50910
rect 156300 50850 156310 50910
rect 156480 50850 156490 50910
rect 156660 50850 156670 50910
rect 156840 50850 156850 50910
rect 157020 50850 157030 50910
rect 157200 50850 157210 50910
rect 157380 50850 157390 50910
rect 157560 50850 157570 50910
rect 157740 50850 157750 50910
rect 157920 50850 157930 50910
rect 158100 50850 158110 50910
rect 158280 50850 158290 50910
rect 158460 50850 158470 50910
rect 158640 50850 158650 50910
rect 158820 50850 158830 50910
rect 158900 50850 158990 50920
rect 159520 50890 159550 50920
rect 159640 50890 159670 50920
rect 163520 50890 163550 50920
rect 163640 50890 163670 50920
rect 164280 50910 164360 50920
rect 164460 50910 164540 50920
rect 164640 50910 164720 50920
rect 164820 50910 164900 50920
rect 165000 50910 165080 50920
rect 165180 50910 165260 50920
rect 165360 50910 165440 50920
rect 165540 50910 165620 50920
rect 165720 50910 165800 50920
rect 165900 50910 165980 50920
rect 166080 50910 166160 50920
rect 166260 50910 166340 50920
rect 166440 50910 166520 50920
rect 166620 50910 166700 50920
rect 166800 50910 166880 50920
rect 166980 50910 167060 50920
rect 167160 50910 167240 50920
rect 167340 50910 167420 50920
rect 167520 50910 167600 50920
rect 167700 50910 167780 50920
rect 167880 50910 167960 50920
rect 168060 50910 168140 50920
rect 168240 50910 168320 50920
rect 168420 50910 168500 50920
rect 168600 50910 168680 50920
rect 168780 50910 168860 50920
rect 168960 50910 169040 50920
rect 169140 50910 169220 50920
rect 169320 50910 169400 50920
rect 169500 50910 169580 50920
rect 169680 50910 169760 50920
rect 169860 50910 169940 50920
rect 170040 50910 170120 50920
rect 159400 50860 159460 50890
rect 159520 50860 159580 50890
rect 159640 50860 159700 50890
rect 163400 50860 163460 50890
rect 163520 50860 163580 50890
rect 163640 50860 163700 50890
rect 152900 50820 158990 50850
rect 164360 50830 164370 50910
rect 164540 50830 164550 50910
rect 164720 50830 164730 50910
rect 164900 50830 164910 50910
rect 165080 50830 165090 50910
rect 165260 50830 165270 50910
rect 165440 50830 165450 50910
rect 165620 50830 165630 50910
rect 165800 50830 165810 50910
rect 165980 50830 165990 50910
rect 166160 50830 166170 50910
rect 166340 50830 166350 50910
rect 166520 50830 166530 50910
rect 166700 50830 166710 50910
rect 166880 50830 166890 50910
rect 167060 50830 167070 50910
rect 167240 50830 167250 50910
rect 167420 50830 167430 50910
rect 167600 50830 167610 50910
rect 167780 50830 167790 50910
rect 167960 50830 167970 50910
rect 168140 50830 168150 50910
rect 168320 50830 168330 50910
rect 168500 50830 168510 50910
rect 168680 50830 168690 50910
rect 168860 50830 168870 50910
rect 169040 50830 169050 50910
rect 169220 50830 169230 50910
rect 169400 50830 169410 50910
rect 169580 50830 169590 50910
rect 169760 50830 169770 50910
rect 169940 50830 169950 50910
rect 170120 50830 170130 50910
rect 170810 50890 170840 50920
rect 170930 50890 170960 50920
rect 170690 50860 170750 50890
rect 170810 50860 170870 50890
rect 170930 50860 170990 50890
rect 146100 50790 146160 50820
rect 147580 50790 147640 50820
rect 148400 50790 148460 50820
rect 149880 50790 149940 50820
rect 152220 50770 152250 50800
rect 152340 50770 152370 50800
rect 152100 50740 152160 50770
rect 152220 50740 152280 50770
rect 152340 50740 152400 50770
rect 152980 50760 153060 50770
rect 153160 50760 153240 50770
rect 153340 50760 153420 50770
rect 153520 50760 153600 50770
rect 153700 50760 153780 50770
rect 153880 50760 153960 50770
rect 154060 50760 154140 50770
rect 154240 50760 154320 50770
rect 154420 50760 154500 50770
rect 154600 50760 154680 50770
rect 154780 50760 154860 50770
rect 154960 50760 155040 50770
rect 155140 50760 155220 50770
rect 155320 50760 155400 50770
rect 155500 50760 155580 50770
rect 155680 50760 155760 50770
rect 155860 50760 155940 50770
rect 156040 50760 156120 50770
rect 156220 50760 156300 50770
rect 156400 50760 156480 50770
rect 156580 50760 156660 50770
rect 156760 50760 156840 50770
rect 156940 50760 157020 50770
rect 157120 50760 157200 50770
rect 157300 50760 157380 50770
rect 157480 50760 157560 50770
rect 157660 50760 157740 50770
rect 157840 50760 157920 50770
rect 158020 50760 158100 50770
rect 158200 50760 158280 50770
rect 158380 50760 158460 50770
rect 158560 50760 158640 50770
rect 158740 50760 158820 50770
rect 41540 50710 41600 50740
rect 42360 50710 42420 50740
rect 43840 50710 43900 50740
rect 41540 50590 41600 50620
rect 42360 50590 42420 50620
rect 42910 50600 43030 50660
rect 43190 50600 43310 50660
rect 43030 50590 43090 50600
rect 43310 50590 43370 50600
rect 43840 50590 43900 50620
rect 42930 50580 43010 50590
rect 43030 50580 43150 50590
rect 43210 50580 43290 50590
rect 43310 50580 43430 50590
rect 41540 50470 41600 50500
rect 42360 50470 42420 50500
rect 42470 50480 42480 50570
rect 41540 50350 41600 50380
rect 42360 50350 42420 50380
rect 41540 50230 41600 50260
rect 42360 50230 42420 50260
rect 41540 50110 41600 50140
rect 42360 50110 42420 50140
rect 41540 49990 41600 50020
rect 42360 49990 42420 50020
rect 41540 49870 41600 49900
rect 42360 49870 42420 49900
rect 41540 49750 41600 49780
rect 42360 49750 42420 49780
rect 41540 49630 41600 49660
rect 42360 49630 42420 49660
rect 41540 49510 41600 49540
rect 42360 49510 42420 49540
rect 41540 49390 41600 49420
rect 42360 49390 42420 49420
rect 41540 49270 41600 49300
rect 42360 49270 42420 49300
rect 41540 49150 41600 49180
rect 42360 49150 42420 49180
rect 42560 49120 42570 50480
rect 42610 50450 42730 50510
rect 42730 50425 42790 50450
rect 42860 50440 42870 50570
rect 43010 50500 43020 50580
rect 43030 50480 43090 50580
rect 43150 50500 43160 50580
rect 43290 50500 43300 50580
rect 43310 50480 43370 50580
rect 43430 50500 43440 50580
rect 146100 50670 146160 50700
rect 147580 50670 147640 50700
rect 148400 50670 148460 50700
rect 149880 50670 149940 50700
rect 153060 50680 153070 50760
rect 153240 50680 153250 50760
rect 153420 50680 153430 50760
rect 153600 50680 153610 50760
rect 153780 50680 153790 50760
rect 153960 50680 153970 50760
rect 154140 50680 154150 50760
rect 154320 50680 154330 50760
rect 154500 50680 154510 50760
rect 154680 50680 154690 50760
rect 154860 50680 154870 50760
rect 155040 50680 155050 50760
rect 155220 50680 155230 50760
rect 155400 50680 155410 50760
rect 155580 50680 155590 50760
rect 155760 50680 155770 50760
rect 155940 50680 155950 50760
rect 156120 50680 156130 50760
rect 156300 50680 156310 50760
rect 156480 50680 156490 50760
rect 156660 50680 156670 50760
rect 156840 50680 156850 50760
rect 157020 50680 157030 50760
rect 157200 50680 157210 50760
rect 157380 50680 157390 50760
rect 157560 50680 157570 50760
rect 157740 50680 157750 50760
rect 157920 50680 157930 50760
rect 158100 50680 158110 50760
rect 158280 50680 158290 50760
rect 158460 50680 158470 50760
rect 158640 50680 158650 50760
rect 158820 50680 158830 50760
rect 152220 50650 152250 50680
rect 152340 50650 152370 50680
rect 152100 50620 152160 50650
rect 152220 50620 152280 50650
rect 152340 50620 152400 50650
rect 158900 50620 158990 50820
rect 159520 50770 159550 50800
rect 159640 50770 159670 50800
rect 163520 50770 163550 50800
rect 163640 50770 163670 50800
rect 170810 50770 170840 50800
rect 170930 50770 170960 50800
rect 159400 50740 159460 50770
rect 159520 50740 159580 50770
rect 159640 50740 159700 50770
rect 163400 50740 163460 50770
rect 163520 50740 163580 50770
rect 163640 50740 163700 50770
rect 164280 50760 164360 50770
rect 164460 50760 164540 50770
rect 164640 50760 164720 50770
rect 164820 50760 164900 50770
rect 165000 50760 165080 50770
rect 165180 50760 165260 50770
rect 165360 50760 165440 50770
rect 165540 50760 165620 50770
rect 165720 50760 165800 50770
rect 165900 50760 165980 50770
rect 166080 50760 166160 50770
rect 166260 50760 166340 50770
rect 166440 50760 166520 50770
rect 166620 50760 166700 50770
rect 166800 50760 166880 50770
rect 166980 50760 167060 50770
rect 167160 50760 167240 50770
rect 167340 50760 167420 50770
rect 167520 50760 167600 50770
rect 167700 50760 167780 50770
rect 167880 50760 167960 50770
rect 168060 50760 168140 50770
rect 168240 50760 168320 50770
rect 168420 50760 168500 50770
rect 168600 50760 168680 50770
rect 168780 50760 168860 50770
rect 168960 50760 169040 50770
rect 169140 50760 169220 50770
rect 169320 50760 169400 50770
rect 169500 50760 169580 50770
rect 169680 50760 169760 50770
rect 169860 50760 169940 50770
rect 170040 50760 170120 50770
rect 164360 50680 164370 50760
rect 164540 50680 164550 50760
rect 164720 50680 164730 50760
rect 164900 50680 164910 50760
rect 165080 50680 165090 50760
rect 165260 50680 165270 50760
rect 165440 50680 165450 50760
rect 165620 50680 165630 50760
rect 165800 50680 165810 50760
rect 165980 50680 165990 50760
rect 166160 50680 166170 50760
rect 166340 50680 166350 50760
rect 166520 50680 166530 50760
rect 166700 50680 166710 50760
rect 166880 50680 166890 50760
rect 167060 50680 167070 50760
rect 167240 50680 167250 50760
rect 167420 50680 167430 50760
rect 167600 50680 167610 50760
rect 167780 50680 167790 50760
rect 167960 50680 167970 50760
rect 168140 50680 168150 50760
rect 168320 50680 168330 50760
rect 168500 50680 168510 50760
rect 168680 50680 168690 50760
rect 168860 50680 168870 50760
rect 169040 50680 169050 50760
rect 169220 50680 169230 50760
rect 169400 50680 169410 50760
rect 169580 50680 169590 50760
rect 169760 50680 169770 50760
rect 169940 50680 169950 50760
rect 170120 50680 170130 50760
rect 170690 50740 170750 50770
rect 170810 50740 170870 50770
rect 170930 50740 170990 50770
rect 159520 50650 159550 50680
rect 159640 50650 159670 50680
rect 163520 50650 163550 50680
rect 163640 50650 163670 50680
rect 170810 50650 170840 50680
rect 170930 50650 170960 50680
rect 159400 50620 159460 50650
rect 159520 50620 159580 50650
rect 159640 50620 159700 50650
rect 163400 50620 163460 50650
rect 163520 50620 163580 50650
rect 163640 50620 163700 50650
rect 170690 50620 170750 50650
rect 170810 50620 170870 50650
rect 170930 50620 170990 50650
rect 152900 50590 158990 50620
rect 164280 50610 164360 50620
rect 164460 50610 164540 50620
rect 164640 50610 164720 50620
rect 164820 50610 164900 50620
rect 165000 50610 165080 50620
rect 165180 50610 165260 50620
rect 165360 50610 165440 50620
rect 165540 50610 165620 50620
rect 165720 50610 165800 50620
rect 165900 50610 165980 50620
rect 166080 50610 166160 50620
rect 166260 50610 166340 50620
rect 166440 50610 166520 50620
rect 166620 50610 166700 50620
rect 166800 50610 166880 50620
rect 166980 50610 167060 50620
rect 167160 50610 167240 50620
rect 167340 50610 167420 50620
rect 167520 50610 167600 50620
rect 167700 50610 167780 50620
rect 167880 50610 167960 50620
rect 168060 50610 168140 50620
rect 168240 50610 168320 50620
rect 168420 50610 168500 50620
rect 168600 50610 168680 50620
rect 168780 50610 168860 50620
rect 168960 50610 169040 50620
rect 169140 50610 169220 50620
rect 169320 50610 169400 50620
rect 169500 50610 169580 50620
rect 169680 50610 169760 50620
rect 169860 50610 169940 50620
rect 170040 50610 170120 50620
rect 146100 50550 146160 50580
rect 147580 50550 147640 50580
rect 148400 50550 148460 50580
rect 149880 50550 149940 50580
rect 152220 50530 152250 50560
rect 152340 50530 152370 50560
rect 153060 50530 153070 50590
rect 153240 50530 153250 50590
rect 153420 50530 153430 50590
rect 153600 50530 153610 50590
rect 153780 50530 153790 50590
rect 153960 50530 153970 50590
rect 154140 50530 154150 50590
rect 154320 50530 154330 50590
rect 154500 50530 154510 50590
rect 154680 50530 154690 50590
rect 154860 50530 154870 50590
rect 155040 50530 155050 50590
rect 155220 50530 155230 50590
rect 155400 50530 155410 50590
rect 155580 50530 155590 50590
rect 155760 50530 155770 50590
rect 155940 50530 155950 50590
rect 156120 50530 156130 50590
rect 156300 50530 156310 50590
rect 156480 50530 156490 50590
rect 156660 50530 156670 50590
rect 156840 50530 156850 50590
rect 157020 50530 157030 50590
rect 157200 50530 157210 50590
rect 157380 50530 157390 50590
rect 157560 50530 157570 50590
rect 157740 50530 157750 50590
rect 157920 50530 157930 50590
rect 158100 50530 158110 50590
rect 158280 50530 158290 50590
rect 158460 50530 158470 50590
rect 158640 50530 158650 50590
rect 158820 50530 158830 50590
rect 152100 50500 152160 50530
rect 152220 50500 152280 50530
rect 152340 50500 152400 50530
rect 158900 50520 158990 50590
rect 159520 50530 159550 50560
rect 159640 50530 159670 50560
rect 163520 50530 163550 50560
rect 163640 50530 163670 50560
rect 164360 50530 164370 50610
rect 164540 50530 164550 50610
rect 164720 50530 164730 50610
rect 164900 50530 164910 50610
rect 165080 50530 165090 50610
rect 165260 50530 165270 50610
rect 165440 50530 165450 50610
rect 165620 50530 165630 50610
rect 165800 50530 165810 50610
rect 165980 50530 165990 50610
rect 166160 50530 166170 50610
rect 166340 50530 166350 50610
rect 166520 50530 166530 50610
rect 166700 50530 166710 50610
rect 166880 50530 166890 50610
rect 167060 50530 167070 50610
rect 167240 50530 167250 50610
rect 167420 50530 167430 50610
rect 167600 50530 167610 50610
rect 167780 50530 167790 50610
rect 167960 50530 167970 50610
rect 168140 50530 168150 50610
rect 168320 50530 168330 50610
rect 168500 50530 168510 50610
rect 168680 50530 168690 50610
rect 168860 50530 168870 50610
rect 169040 50530 169050 50610
rect 169220 50530 169230 50610
rect 169400 50530 169410 50610
rect 169580 50530 169590 50610
rect 169760 50530 169770 50610
rect 169940 50530 169950 50610
rect 170120 50530 170130 50610
rect 170810 50530 170840 50560
rect 170930 50530 170960 50560
rect 43840 50470 43900 50500
rect 152900 50490 158990 50520
rect 159400 50500 159460 50530
rect 159520 50500 159580 50530
rect 159640 50500 159700 50530
rect 163400 50500 163460 50530
rect 163520 50500 163580 50530
rect 163640 50500 163700 50530
rect 170690 50500 170750 50530
rect 170810 50500 170870 50530
rect 170930 50500 170990 50530
rect 158900 50480 158990 50490
rect 152900 50470 158990 50480
rect 164200 50470 170200 50480
rect 42860 50430 43500 50440
rect 42730 50415 43540 50425
rect 42730 50330 42790 50415
rect 43540 50365 43550 50415
rect 42620 50240 42700 50250
rect 42700 50160 42710 50240
rect 42860 50160 42870 50350
rect 42910 50300 43030 50360
rect 43190 50300 43310 50360
rect 43020 50270 43090 50300
rect 43030 50180 43090 50270
rect 43190 50210 43200 50300
rect 43300 50270 43370 50300
rect 43310 50180 43370 50270
rect 42860 50150 43490 50160
rect 42860 50140 42870 50150
rect 42620 50060 42700 50070
rect 42700 49980 42710 50060
rect 42770 50050 42780 50140
rect 42610 49860 42730 49920
rect 42730 49835 42790 49860
rect 42860 49850 42870 50050
rect 42910 50010 43030 50070
rect 43190 50010 43310 50070
rect 43030 50000 43090 50010
rect 43310 50000 43370 50010
rect 42930 49990 43010 50000
rect 43030 49990 43150 50000
rect 43210 49990 43290 50000
rect 43310 49990 43430 50000
rect 43010 49910 43020 49990
rect 43030 49890 43090 49990
rect 43150 49910 43160 49990
rect 43290 49910 43300 49990
rect 43310 49890 43370 49990
rect 43430 49910 43440 49990
rect 42860 49840 43500 49850
rect 43580 49840 43590 50140
rect 42730 49825 43540 49835
rect 42730 49740 42790 49825
rect 43540 49775 43550 49825
rect 42620 49640 42700 49650
rect 42700 49560 42710 49640
rect 42860 49570 42870 49760
rect 42910 49710 43030 49770
rect 43190 49710 43310 49770
rect 43020 49680 43090 49710
rect 43030 49590 43090 49680
rect 43190 49620 43200 49710
rect 43300 49680 43370 49710
rect 43310 49590 43370 49680
rect 42860 49560 43490 49570
rect 42860 49550 42870 49560
rect 42620 49460 42700 49470
rect 42770 49460 42780 49550
rect 42700 49380 42710 49460
rect 42610 49270 42730 49330
rect 42730 49245 42790 49270
rect 42860 49260 42870 49460
rect 42910 49420 43030 49480
rect 43190 49420 43310 49480
rect 43030 49410 43090 49420
rect 43310 49410 43370 49420
rect 42930 49400 43010 49410
rect 43030 49400 43150 49410
rect 43210 49400 43290 49410
rect 43310 49400 43430 49410
rect 43010 49320 43020 49400
rect 43030 49300 43090 49400
rect 43150 49320 43160 49400
rect 43290 49320 43300 49400
rect 43310 49300 43370 49400
rect 43430 49320 43440 49400
rect 42860 49250 43500 49260
rect 43580 49250 43590 49550
rect 42730 49235 43540 49245
rect 42730 49150 42790 49235
rect 43540 49185 43550 49235
rect 42860 49120 42870 49170
rect 42910 49120 43030 49180
rect 43190 49120 43310 49180
rect 43030 49110 43090 49120
rect 43310 49110 43370 49120
rect 43030 49100 43150 49110
rect 43310 49100 43430 49110
rect 40770 49090 40830 49100
rect 40530 49080 40610 49090
rect 40770 49080 40890 49090
rect 40610 49000 40620 49080
rect 40770 48980 40830 49080
rect 40890 49000 40900 49080
rect 41050 48980 41180 49100
rect 41540 49030 41600 49060
rect 42360 49030 42420 49060
rect 43030 49000 43090 49100
rect 43150 49020 43160 49100
rect 43310 49000 43370 49100
rect 43430 49020 43440 49100
rect 41090 48950 41180 48980
rect 43780 48960 43790 50440
rect 146100 50430 146160 50460
rect 147580 50430 147640 50460
rect 148400 50430 148460 50460
rect 149880 50430 149940 50460
rect 152220 50410 152250 50440
rect 152340 50410 152370 50440
rect 152100 50380 152160 50410
rect 152220 50380 152280 50410
rect 152340 50380 152400 50410
rect 43840 50350 43900 50380
rect 146100 50310 146160 50340
rect 147580 50310 147640 50340
rect 148400 50310 148460 50340
rect 149880 50310 149940 50340
rect 152220 50290 152250 50320
rect 152340 50290 152370 50320
rect 152980 50290 153060 50300
rect 153160 50290 153240 50300
rect 153340 50290 153420 50300
rect 153520 50290 153600 50300
rect 153700 50290 153780 50300
rect 153880 50290 153960 50300
rect 154060 50290 154140 50300
rect 154240 50290 154320 50300
rect 154420 50290 154500 50300
rect 154600 50290 154680 50300
rect 154780 50290 154860 50300
rect 154960 50290 155040 50300
rect 155140 50290 155220 50300
rect 155320 50290 155400 50300
rect 155500 50290 155580 50300
rect 155680 50290 155760 50300
rect 155860 50290 155940 50300
rect 156040 50290 156120 50300
rect 156220 50290 156300 50300
rect 156400 50290 156480 50300
rect 156580 50290 156660 50300
rect 156760 50290 156840 50300
rect 156940 50290 157020 50300
rect 157120 50290 157200 50300
rect 157300 50290 157380 50300
rect 157480 50290 157560 50300
rect 157660 50290 157740 50300
rect 157840 50290 157920 50300
rect 158020 50290 158100 50300
rect 158200 50290 158280 50300
rect 158380 50290 158460 50300
rect 158560 50290 158640 50300
rect 158740 50290 158820 50300
rect 152100 50260 152160 50290
rect 152220 50260 152280 50290
rect 152340 50260 152400 50290
rect 43840 50230 43900 50260
rect 146100 50190 146160 50220
rect 147580 50190 147640 50220
rect 148400 50190 148460 50220
rect 149880 50190 149940 50220
rect 153060 50210 153070 50290
rect 153240 50210 153250 50290
rect 153420 50210 153430 50290
rect 153600 50210 153610 50290
rect 153780 50210 153790 50290
rect 153960 50210 153970 50290
rect 154140 50210 154150 50290
rect 154320 50210 154330 50290
rect 154500 50210 154510 50290
rect 154680 50210 154690 50290
rect 154860 50210 154870 50290
rect 155040 50210 155050 50290
rect 155220 50210 155230 50290
rect 155400 50210 155410 50290
rect 155580 50210 155590 50290
rect 155760 50210 155770 50290
rect 155940 50210 155950 50290
rect 156120 50210 156130 50290
rect 156300 50210 156310 50290
rect 156480 50210 156490 50290
rect 156660 50210 156670 50290
rect 156840 50210 156850 50290
rect 157020 50210 157030 50290
rect 157200 50210 157210 50290
rect 157380 50210 157390 50290
rect 157560 50210 157570 50290
rect 157740 50210 157750 50290
rect 157920 50210 157930 50290
rect 158100 50210 158110 50290
rect 158280 50210 158290 50290
rect 158460 50210 158470 50290
rect 158640 50210 158650 50290
rect 158820 50210 158830 50290
rect 152220 50170 152250 50200
rect 152340 50170 152370 50200
rect 152100 50140 152160 50170
rect 152220 50140 152280 50170
rect 152340 50140 152400 50170
rect 43840 50110 43900 50140
rect 146100 50070 146160 50100
rect 147580 50070 147640 50100
rect 148400 50070 148460 50100
rect 149880 50070 149940 50100
rect 152220 50050 152250 50080
rect 152340 50050 152370 50080
rect 152100 50020 152160 50050
rect 152220 50020 152280 50050
rect 152340 50020 152400 50050
rect 43840 49990 43900 50020
rect 146100 49950 146160 49980
rect 147580 49950 147640 49980
rect 148400 49950 148460 49980
rect 149880 49950 149940 49980
rect 152980 49970 153060 49980
rect 153160 49970 153240 49980
rect 153340 49970 153420 49980
rect 153520 49970 153600 49980
rect 153700 49970 153780 49980
rect 153880 49970 153960 49980
rect 154060 49970 154140 49980
rect 154240 49970 154320 49980
rect 154420 49970 154500 49980
rect 154600 49970 154680 49980
rect 154780 49970 154860 49980
rect 154960 49970 155040 49980
rect 155140 49970 155220 49980
rect 155320 49970 155400 49980
rect 155500 49970 155580 49980
rect 155680 49970 155760 49980
rect 155860 49970 155940 49980
rect 156040 49970 156120 49980
rect 156220 49970 156300 49980
rect 156400 49970 156480 49980
rect 156580 49970 156660 49980
rect 156760 49970 156840 49980
rect 156940 49970 157020 49980
rect 157120 49970 157200 49980
rect 157300 49970 157380 49980
rect 157480 49970 157560 49980
rect 157660 49970 157740 49980
rect 157840 49970 157920 49980
rect 158020 49970 158100 49980
rect 158200 49970 158280 49980
rect 158380 49970 158460 49980
rect 158560 49970 158640 49980
rect 158740 49970 158820 49980
rect 152220 49930 152250 49960
rect 152340 49930 152370 49960
rect 152100 49900 152160 49930
rect 152220 49900 152280 49930
rect 152340 49900 152400 49930
rect 43840 49870 43900 49900
rect 153060 49890 153070 49970
rect 153240 49890 153250 49970
rect 153420 49890 153430 49970
rect 153600 49890 153610 49970
rect 153780 49890 153790 49970
rect 153960 49890 153970 49970
rect 154140 49890 154150 49970
rect 154320 49890 154330 49970
rect 154500 49890 154510 49970
rect 154680 49890 154690 49970
rect 154860 49890 154870 49970
rect 155040 49890 155050 49970
rect 155220 49890 155230 49970
rect 155400 49890 155410 49970
rect 155580 49890 155590 49970
rect 155760 49890 155770 49970
rect 155940 49890 155950 49970
rect 156120 49890 156130 49970
rect 156300 49890 156310 49970
rect 156480 49890 156490 49970
rect 156660 49890 156670 49970
rect 156840 49890 156850 49970
rect 157020 49890 157030 49970
rect 157200 49890 157210 49970
rect 157380 49890 157390 49970
rect 157560 49890 157570 49970
rect 157740 49890 157750 49970
rect 157920 49890 157930 49970
rect 158100 49890 158110 49970
rect 158280 49890 158290 49970
rect 158460 49890 158470 49970
rect 158640 49890 158650 49970
rect 158820 49890 158830 49970
rect 146100 49830 146160 49860
rect 147580 49830 147640 49860
rect 148400 49830 148460 49860
rect 149880 49830 149940 49860
rect 152220 49810 152250 49840
rect 152340 49810 152370 49840
rect 152100 49780 152160 49810
rect 152220 49780 152280 49810
rect 152340 49780 152400 49810
rect 158900 49800 158990 50470
rect 159520 50410 159550 50440
rect 159640 50410 159670 50440
rect 163520 50410 163550 50440
rect 163640 50410 163670 50440
rect 170810 50410 170840 50440
rect 170930 50410 170960 50440
rect 159400 50380 159460 50410
rect 159520 50380 159580 50410
rect 159640 50380 159700 50410
rect 163400 50380 163460 50410
rect 163520 50380 163580 50410
rect 163640 50380 163700 50410
rect 170690 50380 170750 50410
rect 170810 50380 170870 50410
rect 170930 50380 170990 50410
rect 159520 50290 159550 50320
rect 159640 50290 159670 50320
rect 163520 50290 163550 50320
rect 163640 50290 163670 50320
rect 164280 50290 164360 50300
rect 164460 50290 164540 50300
rect 164640 50290 164720 50300
rect 164820 50290 164900 50300
rect 165000 50290 165080 50300
rect 165180 50290 165260 50300
rect 165360 50290 165440 50300
rect 165540 50290 165620 50300
rect 165720 50290 165800 50300
rect 165900 50290 165980 50300
rect 166080 50290 166160 50300
rect 166260 50290 166340 50300
rect 166440 50290 166520 50300
rect 166620 50290 166700 50300
rect 166800 50290 166880 50300
rect 166980 50290 167060 50300
rect 167160 50290 167240 50300
rect 167340 50290 167420 50300
rect 167520 50290 167600 50300
rect 167700 50290 167780 50300
rect 167880 50290 167960 50300
rect 168060 50290 168140 50300
rect 168240 50290 168320 50300
rect 168420 50290 168500 50300
rect 168600 50290 168680 50300
rect 168780 50290 168860 50300
rect 168960 50290 169040 50300
rect 169140 50290 169220 50300
rect 169320 50290 169400 50300
rect 169500 50290 169580 50300
rect 169680 50290 169760 50300
rect 169860 50290 169940 50300
rect 170040 50290 170120 50300
rect 170810 50290 170840 50320
rect 170930 50290 170960 50320
rect 159400 50260 159460 50290
rect 159520 50260 159580 50290
rect 159640 50260 159700 50290
rect 163400 50260 163460 50290
rect 163520 50260 163580 50290
rect 163640 50260 163700 50290
rect 164360 50210 164370 50290
rect 164540 50210 164550 50290
rect 164720 50210 164730 50290
rect 164900 50210 164910 50290
rect 165080 50210 165090 50290
rect 165260 50210 165270 50290
rect 165440 50210 165450 50290
rect 165620 50210 165630 50290
rect 165800 50210 165810 50290
rect 165980 50210 165990 50290
rect 166160 50210 166170 50290
rect 166340 50210 166350 50290
rect 166520 50210 166530 50290
rect 166700 50210 166710 50290
rect 166880 50210 166890 50290
rect 167060 50210 167070 50290
rect 167240 50210 167250 50290
rect 167420 50210 167430 50290
rect 167600 50210 167610 50290
rect 167780 50210 167790 50290
rect 167960 50210 167970 50290
rect 168140 50210 168150 50290
rect 168320 50210 168330 50290
rect 168500 50210 168510 50290
rect 168680 50210 168690 50290
rect 168860 50210 168870 50290
rect 169040 50210 169050 50290
rect 169220 50210 169230 50290
rect 169400 50210 169410 50290
rect 169580 50210 169590 50290
rect 169760 50210 169770 50290
rect 169940 50210 169950 50290
rect 170120 50210 170130 50290
rect 170690 50260 170750 50290
rect 170810 50260 170870 50290
rect 170930 50260 170990 50290
rect 159520 50170 159550 50200
rect 159640 50170 159670 50200
rect 163520 50170 163550 50200
rect 163640 50170 163670 50200
rect 170810 50170 170840 50200
rect 170930 50170 170960 50200
rect 159400 50140 159460 50170
rect 159520 50140 159580 50170
rect 159640 50140 159700 50170
rect 163400 50140 163460 50170
rect 163520 50140 163580 50170
rect 163640 50140 163700 50170
rect 170690 50140 170750 50170
rect 170810 50140 170870 50170
rect 170930 50140 170990 50170
rect 159520 50050 159550 50080
rect 159640 50050 159670 50080
rect 163520 50050 163550 50080
rect 163640 50050 163670 50080
rect 170810 50050 170840 50080
rect 170930 50050 170960 50080
rect 159400 50020 159460 50050
rect 159520 50020 159580 50050
rect 159640 50020 159700 50050
rect 163400 50020 163460 50050
rect 163520 50020 163580 50050
rect 163640 50020 163700 50050
rect 170690 50020 170750 50050
rect 170810 50020 170870 50050
rect 170930 50020 170990 50050
rect 164280 49990 164360 50000
rect 164460 49990 164540 50000
rect 164640 49990 164720 50000
rect 164820 49990 164900 50000
rect 165000 49990 165080 50000
rect 165180 49990 165260 50000
rect 165360 49990 165440 50000
rect 165540 49990 165620 50000
rect 165720 49990 165800 50000
rect 165900 49990 165980 50000
rect 166080 49990 166160 50000
rect 166260 49990 166340 50000
rect 166440 49990 166520 50000
rect 166620 49990 166700 50000
rect 166800 49990 166880 50000
rect 166980 49990 167060 50000
rect 167160 49990 167240 50000
rect 167340 49990 167420 50000
rect 167520 49990 167600 50000
rect 167700 49990 167780 50000
rect 167880 49990 167960 50000
rect 168060 49990 168140 50000
rect 168240 49990 168320 50000
rect 168420 49990 168500 50000
rect 168600 49990 168680 50000
rect 168780 49990 168860 50000
rect 168960 49990 169040 50000
rect 169140 49990 169220 50000
rect 169320 49990 169400 50000
rect 169500 49990 169580 50000
rect 169680 49990 169760 50000
rect 169860 49990 169940 50000
rect 170040 49990 170120 50000
rect 159520 49930 159550 49960
rect 159640 49930 159670 49960
rect 163520 49930 163550 49960
rect 163640 49930 163670 49960
rect 159400 49900 159460 49930
rect 159520 49900 159580 49930
rect 159640 49900 159700 49930
rect 163400 49900 163460 49930
rect 163520 49900 163580 49930
rect 163640 49900 163700 49930
rect 164360 49910 164370 49990
rect 164540 49910 164550 49990
rect 164720 49910 164730 49990
rect 164900 49910 164910 49990
rect 165080 49910 165090 49990
rect 165260 49910 165270 49990
rect 165440 49910 165450 49990
rect 165620 49910 165630 49990
rect 165800 49910 165810 49990
rect 165980 49910 165990 49990
rect 166160 49910 166170 49990
rect 166340 49910 166350 49990
rect 166520 49910 166530 49990
rect 166700 49910 166710 49990
rect 166880 49910 166890 49990
rect 167060 49910 167070 49990
rect 167240 49910 167250 49990
rect 167420 49910 167430 49990
rect 167600 49910 167610 49990
rect 167780 49910 167790 49990
rect 167960 49910 167970 49990
rect 168140 49910 168150 49990
rect 168320 49910 168330 49990
rect 168500 49910 168510 49990
rect 168680 49910 168690 49990
rect 168860 49910 168870 49990
rect 169040 49910 169050 49990
rect 169220 49910 169230 49990
rect 169400 49910 169410 49990
rect 169580 49910 169590 49990
rect 169760 49910 169770 49990
rect 169940 49910 169950 49990
rect 170120 49910 170130 49990
rect 170810 49930 170840 49960
rect 170930 49930 170960 49960
rect 170690 49900 170750 49930
rect 170810 49900 170870 49930
rect 170930 49900 170990 49930
rect 159520 49810 159550 49840
rect 159640 49810 159670 49840
rect 163520 49810 163550 49840
rect 163640 49810 163670 49840
rect 170810 49810 170840 49840
rect 170930 49810 170960 49840
rect 152900 49790 158990 49800
rect 43840 49750 43900 49780
rect 146100 49710 146160 49740
rect 147580 49710 147640 49740
rect 148400 49710 148460 49740
rect 149880 49710 149940 49740
rect 152220 49690 152250 49720
rect 152340 49690 152370 49720
rect 158900 49690 158990 49790
rect 159400 49780 159460 49810
rect 159520 49780 159580 49810
rect 159640 49780 159700 49810
rect 163400 49780 163460 49810
rect 163520 49780 163580 49810
rect 163640 49780 163700 49810
rect 164200 49790 170200 49800
rect 170690 49780 170750 49810
rect 170810 49780 170870 49810
rect 170930 49780 170990 49810
rect 159520 49690 159550 49720
rect 159640 49690 159670 49720
rect 163520 49690 163550 49720
rect 163640 49690 163670 49720
rect 170810 49690 170840 49720
rect 170930 49690 170960 49720
rect 152100 49660 152160 49690
rect 152220 49660 152280 49690
rect 152340 49660 152400 49690
rect 152900 49660 158990 49690
rect 159400 49660 159460 49690
rect 159520 49660 159580 49690
rect 159640 49660 159700 49690
rect 163400 49660 163460 49690
rect 163520 49660 163580 49690
rect 163640 49660 163700 49690
rect 170690 49660 170750 49690
rect 170810 49660 170870 49690
rect 170930 49660 170990 49690
rect 43840 49630 43900 49660
rect 152980 49650 153060 49660
rect 153160 49650 153240 49660
rect 153340 49650 153420 49660
rect 153520 49650 153600 49660
rect 153700 49650 153780 49660
rect 153880 49650 153960 49660
rect 154060 49650 154140 49660
rect 154240 49650 154320 49660
rect 154420 49650 154500 49660
rect 154600 49650 154680 49660
rect 154780 49650 154860 49660
rect 154960 49650 155040 49660
rect 155140 49650 155220 49660
rect 155320 49650 155400 49660
rect 155500 49650 155580 49660
rect 155680 49650 155760 49660
rect 155860 49650 155940 49660
rect 156040 49650 156120 49660
rect 156220 49650 156300 49660
rect 156400 49650 156480 49660
rect 156580 49650 156660 49660
rect 156760 49650 156840 49660
rect 156940 49650 157020 49660
rect 157120 49650 157200 49660
rect 157300 49650 157380 49660
rect 157480 49650 157560 49660
rect 157660 49650 157740 49660
rect 157840 49650 157920 49660
rect 158020 49650 158100 49660
rect 158200 49650 158280 49660
rect 158380 49650 158460 49660
rect 158560 49650 158640 49660
rect 158740 49650 158820 49660
rect 146100 49590 146160 49620
rect 147580 49590 147640 49620
rect 148400 49590 148460 49620
rect 149880 49590 149940 49620
rect 152220 49570 152250 49600
rect 152340 49570 152370 49600
rect 153060 49590 153070 49650
rect 153240 49590 153250 49650
rect 153420 49590 153430 49650
rect 153600 49590 153610 49650
rect 153780 49590 153790 49650
rect 153960 49590 153970 49650
rect 154140 49590 154150 49650
rect 154320 49590 154330 49650
rect 154500 49590 154510 49650
rect 154680 49590 154690 49650
rect 154860 49590 154870 49650
rect 155040 49590 155050 49650
rect 155220 49590 155230 49650
rect 155400 49590 155410 49650
rect 155580 49590 155590 49650
rect 155760 49590 155770 49650
rect 155940 49590 155950 49650
rect 156120 49590 156130 49650
rect 156300 49590 156310 49650
rect 156480 49590 156490 49650
rect 156660 49590 156670 49650
rect 156840 49590 156850 49650
rect 157020 49590 157030 49650
rect 157200 49590 157210 49650
rect 157380 49590 157390 49650
rect 157560 49590 157570 49650
rect 157740 49590 157750 49650
rect 157920 49590 157930 49650
rect 158100 49590 158110 49650
rect 158280 49590 158290 49650
rect 158460 49590 158470 49650
rect 158640 49590 158650 49650
rect 158820 49590 158830 49650
rect 158900 49590 158990 49660
rect 164280 49650 164360 49660
rect 164460 49650 164540 49660
rect 164640 49650 164720 49660
rect 164820 49650 164900 49660
rect 165000 49650 165080 49660
rect 165180 49650 165260 49660
rect 165360 49650 165440 49660
rect 165540 49650 165620 49660
rect 165720 49650 165800 49660
rect 165900 49650 165980 49660
rect 166080 49650 166160 49660
rect 166260 49650 166340 49660
rect 166440 49650 166520 49660
rect 166620 49650 166700 49660
rect 166800 49650 166880 49660
rect 166980 49650 167060 49660
rect 167160 49650 167240 49660
rect 167340 49650 167420 49660
rect 167520 49650 167600 49660
rect 167700 49650 167780 49660
rect 167880 49650 167960 49660
rect 168060 49650 168140 49660
rect 168240 49650 168320 49660
rect 168420 49650 168500 49660
rect 168600 49650 168680 49660
rect 168780 49650 168860 49660
rect 168960 49650 169040 49660
rect 169140 49650 169220 49660
rect 169320 49650 169400 49660
rect 169500 49650 169580 49660
rect 169680 49650 169760 49660
rect 169860 49650 169940 49660
rect 170040 49650 170120 49660
rect 152100 49540 152160 49570
rect 152220 49540 152280 49570
rect 152340 49540 152400 49570
rect 152900 49560 158990 49590
rect 159520 49570 159550 49600
rect 159640 49570 159670 49600
rect 163520 49570 163550 49600
rect 163640 49570 163670 49600
rect 164360 49570 164370 49650
rect 164540 49570 164550 49650
rect 164720 49570 164730 49650
rect 164900 49570 164910 49650
rect 165080 49570 165090 49650
rect 165260 49570 165270 49650
rect 165440 49570 165450 49650
rect 165620 49570 165630 49650
rect 165800 49570 165810 49650
rect 165980 49570 165990 49650
rect 166160 49570 166170 49650
rect 166340 49570 166350 49650
rect 166520 49570 166530 49650
rect 166700 49570 166710 49650
rect 166880 49570 166890 49650
rect 167060 49570 167070 49650
rect 167240 49570 167250 49650
rect 167420 49570 167430 49650
rect 167600 49570 167610 49650
rect 167780 49570 167790 49650
rect 167960 49570 167970 49650
rect 168140 49570 168150 49650
rect 168320 49570 168330 49650
rect 168500 49570 168510 49650
rect 168680 49570 168690 49650
rect 168860 49570 168870 49650
rect 169040 49570 169050 49650
rect 169220 49570 169230 49650
rect 169400 49570 169410 49650
rect 169580 49570 169590 49650
rect 169760 49570 169770 49650
rect 169940 49570 169950 49650
rect 170120 49570 170130 49650
rect 170810 49570 170840 49600
rect 170930 49570 170960 49600
rect 43840 49510 43900 49540
rect 152980 49500 153060 49510
rect 153160 49500 153240 49510
rect 153340 49500 153420 49510
rect 153520 49500 153600 49510
rect 153700 49500 153780 49510
rect 153880 49500 153960 49510
rect 154060 49500 154140 49510
rect 154240 49500 154320 49510
rect 154420 49500 154500 49510
rect 154600 49500 154680 49510
rect 154780 49500 154860 49510
rect 154960 49500 155040 49510
rect 155140 49500 155220 49510
rect 155320 49500 155400 49510
rect 155500 49500 155580 49510
rect 155680 49500 155760 49510
rect 155860 49500 155940 49510
rect 156040 49500 156120 49510
rect 156220 49500 156300 49510
rect 156400 49500 156480 49510
rect 156580 49500 156660 49510
rect 156760 49500 156840 49510
rect 156940 49500 157020 49510
rect 157120 49500 157200 49510
rect 157300 49500 157380 49510
rect 157480 49500 157560 49510
rect 157660 49500 157740 49510
rect 157840 49500 157920 49510
rect 158020 49500 158100 49510
rect 158200 49500 158280 49510
rect 158380 49500 158460 49510
rect 158560 49500 158640 49510
rect 158740 49500 158820 49510
rect 146100 49470 146160 49500
rect 147580 49470 147640 49500
rect 148400 49470 148460 49500
rect 149880 49470 149940 49500
rect 152220 49450 152250 49480
rect 152340 49450 152370 49480
rect 152100 49420 152160 49450
rect 152220 49420 152280 49450
rect 152340 49420 152400 49450
rect 153060 49420 153070 49500
rect 153240 49420 153250 49500
rect 153420 49420 153430 49500
rect 153600 49420 153610 49500
rect 153780 49420 153790 49500
rect 153960 49420 153970 49500
rect 154140 49420 154150 49500
rect 154320 49420 154330 49500
rect 154500 49420 154510 49500
rect 154680 49420 154690 49500
rect 154860 49420 154870 49500
rect 155040 49420 155050 49500
rect 155220 49420 155230 49500
rect 155400 49420 155410 49500
rect 155580 49420 155590 49500
rect 155760 49420 155770 49500
rect 155940 49420 155950 49500
rect 156120 49420 156130 49500
rect 156300 49420 156310 49500
rect 156480 49420 156490 49500
rect 156660 49420 156670 49500
rect 156840 49420 156850 49500
rect 157020 49420 157030 49500
rect 157200 49420 157210 49500
rect 157380 49420 157390 49500
rect 157560 49420 157570 49500
rect 157740 49420 157750 49500
rect 157920 49420 157930 49500
rect 158100 49420 158110 49500
rect 158280 49420 158290 49500
rect 158460 49420 158470 49500
rect 158640 49420 158650 49500
rect 158820 49420 158830 49500
rect 43840 49390 43900 49420
rect 146100 49350 146160 49380
rect 147580 49350 147640 49380
rect 148400 49350 148460 49380
rect 149880 49350 149940 49380
rect 152220 49330 152250 49360
rect 152340 49330 152370 49360
rect 152980 49350 153060 49360
rect 153160 49350 153240 49360
rect 153340 49350 153420 49360
rect 153520 49350 153600 49360
rect 153700 49350 153780 49360
rect 153880 49350 153960 49360
rect 154060 49350 154140 49360
rect 154240 49350 154320 49360
rect 154420 49350 154500 49360
rect 154600 49350 154680 49360
rect 154780 49350 154860 49360
rect 154960 49350 155040 49360
rect 155140 49350 155220 49360
rect 155320 49350 155400 49360
rect 155500 49350 155580 49360
rect 155680 49350 155760 49360
rect 155860 49350 155940 49360
rect 156040 49350 156120 49360
rect 156220 49350 156300 49360
rect 156400 49350 156480 49360
rect 156580 49350 156660 49360
rect 156760 49350 156840 49360
rect 156940 49350 157020 49360
rect 157120 49350 157200 49360
rect 157300 49350 157380 49360
rect 157480 49350 157560 49360
rect 157660 49350 157740 49360
rect 157840 49350 157920 49360
rect 158020 49350 158100 49360
rect 158200 49350 158280 49360
rect 158380 49350 158460 49360
rect 158560 49350 158640 49360
rect 158740 49350 158820 49360
rect 152100 49300 152160 49330
rect 152220 49300 152280 49330
rect 152340 49300 152400 49330
rect 43840 49270 43900 49300
rect 153060 49270 153070 49350
rect 153240 49270 153250 49350
rect 153420 49270 153430 49350
rect 153600 49270 153610 49350
rect 153780 49270 153790 49350
rect 153960 49270 153970 49350
rect 154140 49270 154150 49350
rect 154320 49270 154330 49350
rect 154500 49270 154510 49350
rect 154680 49270 154690 49350
rect 154860 49270 154870 49350
rect 155040 49270 155050 49350
rect 155220 49270 155230 49350
rect 155400 49270 155410 49350
rect 155580 49270 155590 49350
rect 155760 49270 155770 49350
rect 155940 49270 155950 49350
rect 156120 49270 156130 49350
rect 156300 49270 156310 49350
rect 156480 49270 156490 49350
rect 156660 49270 156670 49350
rect 156840 49270 156850 49350
rect 157020 49270 157030 49350
rect 157200 49270 157210 49350
rect 157380 49270 157390 49350
rect 157560 49270 157570 49350
rect 157740 49270 157750 49350
rect 157920 49270 157930 49350
rect 158100 49270 158110 49350
rect 158280 49270 158290 49350
rect 158460 49270 158470 49350
rect 158640 49270 158650 49350
rect 158820 49270 158830 49350
rect 158900 49330 158990 49560
rect 159400 49540 159460 49570
rect 159520 49540 159580 49570
rect 159640 49540 159700 49570
rect 163400 49540 163460 49570
rect 163520 49540 163580 49570
rect 163640 49540 163700 49570
rect 170690 49540 170750 49570
rect 170810 49540 170870 49570
rect 170930 49540 170990 49570
rect 164280 49500 164360 49510
rect 164460 49500 164540 49510
rect 164640 49500 164720 49510
rect 164820 49500 164900 49510
rect 165000 49500 165080 49510
rect 165180 49500 165260 49510
rect 165360 49500 165440 49510
rect 165540 49500 165620 49510
rect 165720 49500 165800 49510
rect 165900 49500 165980 49510
rect 166080 49500 166160 49510
rect 166260 49500 166340 49510
rect 166440 49500 166520 49510
rect 166620 49500 166700 49510
rect 166800 49500 166880 49510
rect 166980 49500 167060 49510
rect 167160 49500 167240 49510
rect 167340 49500 167420 49510
rect 167520 49500 167600 49510
rect 167700 49500 167780 49510
rect 167880 49500 167960 49510
rect 168060 49500 168140 49510
rect 168240 49500 168320 49510
rect 168420 49500 168500 49510
rect 168600 49500 168680 49510
rect 168780 49500 168860 49510
rect 168960 49500 169040 49510
rect 169140 49500 169220 49510
rect 169320 49500 169400 49510
rect 169500 49500 169580 49510
rect 169680 49500 169760 49510
rect 169860 49500 169940 49510
rect 170040 49500 170120 49510
rect 159520 49450 159550 49480
rect 159640 49450 159670 49480
rect 163520 49450 163550 49480
rect 163640 49450 163670 49480
rect 159400 49420 159460 49450
rect 159520 49420 159580 49450
rect 159640 49420 159700 49450
rect 163400 49420 163460 49450
rect 163520 49420 163580 49450
rect 163640 49420 163700 49450
rect 164360 49420 164370 49500
rect 164540 49420 164550 49500
rect 164720 49420 164730 49500
rect 164900 49420 164910 49500
rect 165080 49420 165090 49500
rect 165260 49420 165270 49500
rect 165440 49420 165450 49500
rect 165620 49420 165630 49500
rect 165800 49420 165810 49500
rect 165980 49420 165990 49500
rect 166160 49420 166170 49500
rect 166340 49420 166350 49500
rect 166520 49420 166530 49500
rect 166700 49420 166710 49500
rect 166880 49420 166890 49500
rect 167060 49420 167070 49500
rect 167240 49420 167250 49500
rect 167420 49420 167430 49500
rect 167600 49420 167610 49500
rect 167780 49420 167790 49500
rect 167960 49420 167970 49500
rect 168140 49420 168150 49500
rect 168320 49420 168330 49500
rect 168500 49420 168510 49500
rect 168680 49420 168690 49500
rect 168860 49420 168870 49500
rect 169040 49420 169050 49500
rect 169220 49420 169230 49500
rect 169400 49420 169410 49500
rect 169580 49420 169590 49500
rect 169760 49420 169770 49500
rect 169940 49420 169950 49500
rect 170120 49420 170130 49500
rect 170810 49450 170840 49480
rect 170930 49450 170960 49480
rect 170690 49420 170750 49450
rect 170810 49420 170870 49450
rect 170930 49420 170990 49450
rect 159520 49330 159550 49360
rect 159640 49330 159670 49360
rect 163520 49330 163550 49360
rect 163640 49330 163670 49360
rect 164280 49350 164360 49360
rect 164460 49350 164540 49360
rect 164640 49350 164720 49360
rect 164820 49350 164900 49360
rect 165000 49350 165080 49360
rect 165180 49350 165260 49360
rect 165360 49350 165440 49360
rect 165540 49350 165620 49360
rect 165720 49350 165800 49360
rect 165900 49350 165980 49360
rect 166080 49350 166160 49360
rect 166260 49350 166340 49360
rect 166440 49350 166520 49360
rect 166620 49350 166700 49360
rect 166800 49350 166880 49360
rect 166980 49350 167060 49360
rect 167160 49350 167240 49360
rect 167340 49350 167420 49360
rect 167520 49350 167600 49360
rect 167700 49350 167780 49360
rect 167880 49350 167960 49360
rect 168060 49350 168140 49360
rect 168240 49350 168320 49360
rect 168420 49350 168500 49360
rect 168600 49350 168680 49360
rect 168780 49350 168860 49360
rect 168960 49350 169040 49360
rect 169140 49350 169220 49360
rect 169320 49350 169400 49360
rect 169500 49350 169580 49360
rect 169680 49350 169760 49360
rect 169860 49350 169940 49360
rect 170040 49350 170120 49360
rect 159400 49300 159460 49330
rect 159520 49300 159580 49330
rect 159640 49300 159700 49330
rect 163400 49300 163460 49330
rect 163520 49300 163580 49330
rect 163640 49300 163700 49330
rect 164360 49270 164370 49350
rect 164540 49270 164550 49350
rect 164720 49270 164730 49350
rect 164900 49270 164910 49350
rect 165080 49270 165090 49350
rect 165260 49270 165270 49350
rect 165440 49270 165450 49350
rect 165620 49270 165630 49350
rect 165800 49270 165810 49350
rect 165980 49270 165990 49350
rect 166160 49270 166170 49350
rect 166340 49270 166350 49350
rect 166520 49270 166530 49350
rect 166700 49270 166710 49350
rect 166880 49270 166890 49350
rect 167060 49270 167070 49350
rect 167240 49270 167250 49350
rect 167420 49270 167430 49350
rect 167600 49270 167610 49350
rect 167780 49270 167790 49350
rect 167960 49270 167970 49350
rect 168140 49270 168150 49350
rect 168320 49270 168330 49350
rect 168500 49270 168510 49350
rect 168680 49270 168690 49350
rect 168860 49270 168870 49350
rect 169040 49270 169050 49350
rect 169220 49270 169230 49350
rect 169400 49270 169410 49350
rect 169580 49270 169590 49350
rect 169760 49270 169770 49350
rect 169940 49270 169950 49350
rect 170120 49270 170130 49350
rect 170810 49330 170840 49360
rect 170930 49330 170960 49360
rect 170690 49300 170750 49330
rect 170810 49300 170870 49330
rect 170930 49300 170990 49330
rect 146100 49230 146160 49260
rect 147580 49230 147640 49260
rect 148400 49230 148460 49260
rect 149880 49230 149940 49260
rect 152220 49210 152250 49240
rect 152340 49210 152370 49240
rect 159520 49210 159550 49240
rect 159640 49210 159670 49240
rect 163520 49210 163550 49240
rect 163640 49210 163670 49240
rect 170810 49210 170840 49240
rect 170930 49210 170960 49240
rect 152100 49180 152160 49210
rect 152220 49180 152280 49210
rect 152340 49180 152400 49210
rect 159400 49180 159460 49210
rect 159520 49180 159580 49210
rect 159640 49180 159700 49210
rect 163400 49180 163460 49210
rect 163520 49180 163580 49210
rect 163640 49180 163700 49210
rect 170690 49180 170750 49210
rect 170810 49180 170870 49210
rect 170930 49180 170990 49210
rect 43840 49150 43900 49180
rect 146100 49110 146160 49140
rect 147580 49110 147640 49140
rect 148400 49110 148460 49140
rect 149880 49110 149940 49140
rect 152220 49060 152250 49120
rect 152340 49060 152370 49120
rect 159520 49060 159550 49120
rect 159640 49060 159670 49120
rect 163520 49060 163550 49120
rect 163640 49060 163670 49120
rect 170810 49060 170840 49120
rect 170930 49060 170960 49120
rect 43840 49030 43900 49060
rect 146100 48990 146160 49020
rect 147580 48990 147640 49020
rect 148400 48990 148460 49020
rect 149880 48990 149940 49020
rect 19060 48860 19070 48940
rect 19240 48860 19250 48940
rect 19420 48860 19430 48940
rect 19600 48860 19610 48940
rect 19780 48860 19790 48940
rect 19960 48860 19970 48940
rect 20140 48860 20150 48940
rect 20320 48860 20330 48940
rect 20500 48860 20510 48940
rect 20680 48860 20690 48940
rect 20860 48860 20870 48940
rect 21040 48860 21050 48940
rect 21220 48860 21230 48940
rect 21400 48860 21410 48940
rect 21580 48860 21590 48940
rect 21760 48860 21770 48940
rect 21940 48860 21950 48940
rect 22120 48860 22130 48940
rect 22300 48860 22310 48940
rect 22480 48860 22490 48940
rect 22660 48860 22670 48940
rect 22840 48860 22850 48940
rect 23020 48860 23030 48940
rect 23200 48860 23210 48940
rect 23380 48860 23390 48940
rect 23560 48860 23570 48940
rect 23740 48860 23750 48940
rect 23920 48860 23930 48940
rect 24100 48860 24110 48940
rect 24280 48860 24290 48940
rect 24460 48860 24470 48940
rect 24640 48860 24650 48940
rect 24820 48860 24830 48940
rect 25000 48860 25010 48940
rect 25180 48860 25190 48940
rect 25360 48860 25370 48940
rect 25540 48860 25550 48940
rect 25720 48860 25730 48940
rect 25900 48860 25910 48940
rect 26080 48860 26090 48940
rect 26260 48860 26270 48940
rect 26440 48860 26450 48940
rect 26620 48860 26630 48940
rect 27315 48915 27395 48925
rect 27495 48915 27575 48925
rect 27675 48915 27755 48925
rect 27855 48915 27935 48925
rect 28035 48915 28115 48925
rect 27395 48835 27405 48915
rect 27575 48835 27585 48915
rect 27755 48835 27765 48915
rect 27935 48835 27945 48915
rect 28115 48835 28125 48915
rect 30360 48860 30370 48940
rect 30540 48860 30550 48940
rect 30720 48860 30730 48940
rect 30900 48860 30910 48940
rect 31080 48860 31090 48940
rect 31260 48860 31270 48940
rect 31440 48860 31450 48940
rect 31620 48860 31630 48940
rect 31800 48860 31810 48940
rect 31980 48860 31990 48940
rect 32160 48860 32170 48940
rect 32340 48860 32350 48940
rect 32520 48860 32530 48940
rect 32700 48860 32710 48940
rect 32880 48860 32890 48940
rect 33060 48860 33070 48940
rect 33240 48860 33250 48940
rect 33420 48860 33430 48940
rect 33600 48860 33610 48940
rect 33780 48860 33790 48940
rect 33960 48860 33970 48940
rect 34140 48860 34150 48940
rect 34320 48860 34330 48940
rect 34500 48860 34510 48940
rect 34680 48860 34690 48940
rect 34860 48860 34870 48940
rect 35040 48860 35050 48940
rect 35220 48860 35230 48940
rect 35400 48860 35410 48940
rect 35580 48860 35590 48940
rect 35760 48860 35770 48940
rect 35940 48860 35950 48940
rect 36120 48860 36130 48940
rect 36300 48860 36310 48940
rect 36480 48860 36490 48940
rect 36660 48860 36670 48940
rect 36840 48860 36850 48940
rect 37020 48860 37030 48940
rect 37200 48860 37210 48940
rect 37380 48860 37390 48940
rect 37560 48860 37570 48940
rect 37740 48860 37750 48940
rect 37920 48860 37930 48940
rect 40060 48910 40120 48940
rect 41540 48910 41600 48940
rect 42360 48910 42420 48940
rect 43840 48910 43900 48940
rect 146100 48870 146160 48900
rect 147580 48870 147640 48900
rect 148400 48870 148460 48900
rect 149880 48870 149940 48900
rect 18980 48790 19060 48800
rect 19160 48790 19240 48800
rect 19340 48790 19420 48800
rect 19520 48790 19600 48800
rect 19700 48790 19780 48800
rect 19880 48790 19960 48800
rect 20060 48790 20140 48800
rect 20240 48790 20320 48800
rect 20420 48790 20500 48800
rect 20600 48790 20680 48800
rect 20780 48790 20860 48800
rect 20960 48790 21040 48800
rect 21140 48790 21220 48800
rect 21320 48790 21400 48800
rect 21500 48790 21580 48800
rect 21680 48790 21760 48800
rect 21860 48790 21940 48800
rect 22040 48790 22120 48800
rect 22220 48790 22300 48800
rect 22400 48790 22480 48800
rect 22580 48790 22660 48800
rect 22760 48790 22840 48800
rect 22940 48790 23020 48800
rect 23120 48790 23200 48800
rect 23300 48790 23380 48800
rect 23480 48790 23560 48800
rect 23660 48790 23740 48800
rect 23840 48790 23920 48800
rect 24020 48790 24100 48800
rect 24200 48790 24280 48800
rect 24380 48790 24460 48800
rect 24560 48790 24640 48800
rect 24740 48790 24820 48800
rect 24920 48790 25000 48800
rect 25100 48790 25180 48800
rect 25280 48790 25360 48800
rect 25460 48790 25540 48800
rect 25640 48790 25720 48800
rect 25820 48790 25900 48800
rect 26000 48790 26080 48800
rect 26180 48790 26260 48800
rect 26360 48790 26440 48800
rect 26540 48790 26620 48800
rect 30280 48790 30360 48800
rect 30460 48790 30540 48800
rect 30640 48790 30720 48800
rect 30820 48790 30900 48800
rect 31000 48790 31080 48800
rect 31180 48790 31260 48800
rect 31360 48790 31440 48800
rect 31540 48790 31620 48800
rect 31720 48790 31800 48800
rect 31900 48790 31980 48800
rect 32080 48790 32160 48800
rect 32260 48790 32340 48800
rect 32440 48790 32520 48800
rect 32620 48790 32700 48800
rect 32800 48790 32880 48800
rect 32980 48790 33060 48800
rect 33160 48790 33240 48800
rect 33340 48790 33420 48800
rect 33520 48790 33600 48800
rect 33700 48790 33780 48800
rect 33880 48790 33960 48800
rect 34060 48790 34140 48800
rect 34240 48790 34320 48800
rect 34420 48790 34500 48800
rect 34600 48790 34680 48800
rect 34780 48790 34860 48800
rect 34960 48790 35040 48800
rect 35140 48790 35220 48800
rect 35320 48790 35400 48800
rect 35500 48790 35580 48800
rect 35680 48790 35760 48800
rect 35860 48790 35940 48800
rect 36040 48790 36120 48800
rect 36220 48790 36300 48800
rect 36400 48790 36480 48800
rect 36580 48790 36660 48800
rect 36760 48790 36840 48800
rect 36940 48790 37020 48800
rect 37120 48790 37200 48800
rect 37300 48790 37380 48800
rect 37480 48790 37560 48800
rect 37660 48790 37740 48800
rect 37840 48790 37920 48800
rect 152080 48790 152160 48800
rect 152260 48790 152340 48800
rect 152440 48790 152520 48800
rect 152620 48790 152700 48800
rect 152800 48790 152880 48800
rect 152980 48790 153060 48800
rect 153160 48790 153240 48800
rect 153340 48790 153420 48800
rect 153520 48790 153600 48800
rect 153700 48790 153780 48800
rect 153880 48790 153960 48800
rect 154060 48790 154140 48800
rect 154240 48790 154320 48800
rect 154420 48790 154500 48800
rect 154600 48790 154680 48800
rect 154780 48790 154860 48800
rect 154960 48790 155040 48800
rect 155140 48790 155220 48800
rect 155320 48790 155400 48800
rect 155500 48790 155580 48800
rect 155680 48790 155760 48800
rect 155860 48790 155940 48800
rect 156040 48790 156120 48800
rect 156220 48790 156300 48800
rect 156400 48790 156480 48800
rect 156580 48790 156660 48800
rect 156760 48790 156840 48800
rect 156940 48790 157020 48800
rect 157120 48790 157200 48800
rect 157300 48790 157380 48800
rect 157480 48790 157560 48800
rect 157660 48790 157740 48800
rect 157840 48790 157920 48800
rect 158020 48790 158100 48800
rect 158200 48790 158280 48800
rect 158380 48790 158460 48800
rect 158560 48790 158640 48800
rect 158740 48790 158820 48800
rect 158920 48790 159000 48800
rect 159100 48790 159180 48800
rect 159280 48790 159360 48800
rect 159460 48790 159540 48800
rect 159640 48790 159720 48800
rect 163380 48790 163460 48800
rect 163560 48790 163640 48800
rect 163740 48790 163820 48800
rect 163920 48790 164000 48800
rect 164100 48790 164180 48800
rect 164280 48790 164360 48800
rect 164460 48790 164540 48800
rect 164640 48790 164720 48800
rect 164820 48790 164900 48800
rect 165000 48790 165080 48800
rect 165180 48790 165260 48800
rect 165360 48790 165440 48800
rect 165540 48790 165620 48800
rect 165720 48790 165800 48800
rect 165900 48790 165980 48800
rect 166080 48790 166160 48800
rect 166260 48790 166340 48800
rect 166440 48790 166520 48800
rect 166620 48790 166700 48800
rect 166800 48790 166880 48800
rect 166980 48790 167060 48800
rect 167160 48790 167240 48800
rect 167340 48790 167420 48800
rect 167520 48790 167600 48800
rect 167700 48790 167780 48800
rect 167880 48790 167960 48800
rect 168060 48790 168140 48800
rect 168240 48790 168320 48800
rect 168420 48790 168500 48800
rect 168600 48790 168680 48800
rect 168780 48790 168860 48800
rect 168960 48790 169040 48800
rect 169140 48790 169220 48800
rect 169320 48790 169400 48800
rect 169500 48790 169580 48800
rect 169680 48790 169760 48800
rect 169860 48790 169940 48800
rect 170040 48790 170120 48800
rect 170220 48790 170300 48800
rect 170400 48790 170480 48800
rect 170580 48790 170660 48800
rect 170760 48790 170840 48800
rect 170940 48790 171020 48800
rect 19060 48710 19070 48790
rect 19240 48710 19250 48790
rect 19420 48710 19430 48790
rect 19600 48710 19610 48790
rect 19780 48710 19790 48790
rect 19960 48710 19970 48790
rect 20140 48710 20150 48790
rect 20320 48710 20330 48790
rect 20500 48710 20510 48790
rect 20680 48710 20690 48790
rect 20860 48710 20870 48790
rect 21040 48710 21050 48790
rect 21220 48710 21230 48790
rect 21400 48710 21410 48790
rect 21580 48710 21590 48790
rect 21760 48710 21770 48790
rect 21940 48710 21950 48790
rect 22120 48710 22130 48790
rect 22300 48710 22310 48790
rect 22480 48710 22490 48790
rect 22660 48710 22670 48790
rect 22840 48710 22850 48790
rect 23020 48710 23030 48790
rect 23200 48710 23210 48790
rect 23380 48710 23390 48790
rect 23560 48710 23570 48790
rect 23740 48710 23750 48790
rect 23920 48710 23930 48790
rect 24100 48710 24110 48790
rect 24280 48710 24290 48790
rect 24460 48710 24470 48790
rect 24640 48710 24650 48790
rect 24820 48710 24830 48790
rect 25000 48710 25010 48790
rect 25180 48710 25190 48790
rect 25360 48710 25370 48790
rect 25540 48710 25550 48790
rect 25720 48710 25730 48790
rect 25900 48710 25910 48790
rect 26080 48710 26090 48790
rect 26260 48710 26270 48790
rect 26440 48710 26450 48790
rect 26620 48710 26630 48790
rect 27315 48735 27395 48745
rect 27495 48735 27575 48745
rect 27675 48735 27755 48745
rect 27855 48735 27935 48745
rect 28035 48735 28115 48745
rect 27395 48655 27405 48735
rect 27575 48655 27585 48735
rect 27755 48655 27765 48735
rect 27935 48655 27945 48735
rect 28115 48655 28125 48735
rect 30360 48710 30370 48790
rect 30540 48710 30550 48790
rect 30720 48710 30730 48790
rect 30900 48710 30910 48790
rect 31080 48710 31090 48790
rect 31260 48710 31270 48790
rect 31440 48710 31450 48790
rect 31620 48710 31630 48790
rect 31800 48710 31810 48790
rect 31980 48710 31990 48790
rect 32160 48710 32170 48790
rect 32340 48710 32350 48790
rect 32520 48710 32530 48790
rect 32700 48710 32710 48790
rect 32880 48710 32890 48790
rect 33060 48710 33070 48790
rect 33240 48710 33250 48790
rect 33420 48710 33430 48790
rect 33600 48710 33610 48790
rect 33780 48710 33790 48790
rect 33960 48710 33970 48790
rect 34140 48710 34150 48790
rect 34320 48710 34330 48790
rect 34500 48710 34510 48790
rect 34680 48710 34690 48790
rect 34860 48710 34870 48790
rect 35040 48710 35050 48790
rect 35220 48710 35230 48790
rect 35400 48710 35410 48790
rect 35580 48710 35590 48790
rect 35760 48710 35770 48790
rect 35940 48710 35950 48790
rect 36120 48710 36130 48790
rect 36300 48710 36310 48790
rect 36480 48710 36490 48790
rect 36660 48710 36670 48790
rect 36840 48710 36850 48790
rect 37020 48710 37030 48790
rect 37200 48710 37210 48790
rect 37380 48710 37390 48790
rect 37560 48710 37570 48790
rect 37740 48710 37750 48790
rect 37920 48710 37930 48790
rect 152160 48710 152170 48790
rect 152340 48710 152350 48790
rect 152520 48710 152530 48790
rect 152700 48710 152710 48790
rect 152880 48710 152890 48790
rect 153060 48710 153070 48790
rect 153240 48710 153250 48790
rect 153420 48710 153430 48790
rect 153600 48710 153610 48790
rect 153780 48710 153790 48790
rect 153960 48710 153970 48790
rect 154140 48710 154150 48790
rect 154320 48710 154330 48790
rect 154500 48710 154510 48790
rect 154680 48710 154690 48790
rect 154860 48710 154870 48790
rect 155040 48710 155050 48790
rect 155220 48710 155230 48790
rect 155400 48710 155410 48790
rect 155580 48710 155590 48790
rect 155760 48710 155770 48790
rect 155940 48710 155950 48790
rect 156120 48710 156130 48790
rect 156300 48710 156310 48790
rect 156480 48710 156490 48790
rect 156660 48710 156670 48790
rect 156840 48710 156850 48790
rect 157020 48710 157030 48790
rect 157200 48710 157210 48790
rect 157380 48710 157390 48790
rect 157560 48710 157570 48790
rect 157740 48710 157750 48790
rect 157920 48710 157930 48790
rect 158100 48710 158110 48790
rect 158280 48710 158290 48790
rect 158460 48710 158470 48790
rect 158640 48710 158650 48790
rect 158820 48710 158830 48790
rect 159000 48710 159010 48790
rect 159180 48710 159190 48790
rect 159360 48710 159370 48790
rect 159540 48710 159550 48790
rect 159720 48710 159730 48790
rect 160430 48765 160510 48775
rect 160590 48765 160670 48775
rect 160750 48765 160830 48775
rect 160910 48765 160990 48775
rect 161070 48765 161150 48775
rect 160510 48685 160520 48765
rect 160590 48685 160600 48765
rect 160670 48685 160680 48765
rect 160750 48685 160760 48765
rect 160830 48685 160840 48765
rect 160910 48685 160920 48765
rect 160990 48685 161000 48765
rect 161070 48685 161080 48765
rect 161150 48685 161160 48765
rect 163460 48710 163470 48790
rect 163640 48710 163650 48790
rect 163820 48710 163830 48790
rect 164000 48710 164010 48790
rect 164180 48710 164190 48790
rect 164360 48710 164370 48790
rect 164540 48710 164550 48790
rect 164720 48710 164730 48790
rect 164900 48710 164910 48790
rect 165080 48710 165090 48790
rect 165260 48710 165270 48790
rect 165440 48710 165450 48790
rect 165620 48710 165630 48790
rect 165800 48710 165810 48790
rect 165980 48710 165990 48790
rect 166160 48710 166170 48790
rect 166340 48710 166350 48790
rect 166520 48710 166530 48790
rect 166700 48710 166710 48790
rect 166880 48710 166890 48790
rect 167060 48710 167070 48790
rect 167240 48710 167250 48790
rect 167420 48710 167430 48790
rect 167600 48710 167610 48790
rect 167780 48710 167790 48790
rect 167960 48710 167970 48790
rect 168140 48710 168150 48790
rect 168320 48710 168330 48790
rect 168500 48710 168510 48790
rect 168680 48710 168690 48790
rect 168860 48710 168870 48790
rect 169040 48710 169050 48790
rect 169220 48710 169230 48790
rect 169400 48710 169410 48790
rect 169580 48710 169590 48790
rect 169760 48710 169770 48790
rect 169940 48710 169950 48790
rect 170120 48710 170130 48790
rect 170300 48710 170310 48790
rect 170480 48710 170490 48790
rect 170660 48710 170670 48790
rect 170840 48710 170850 48790
rect 171020 48710 171030 48790
rect 18980 48640 19060 48650
rect 19160 48640 19240 48650
rect 19340 48640 19420 48650
rect 19520 48640 19600 48650
rect 19700 48640 19780 48650
rect 19880 48640 19960 48650
rect 20060 48640 20140 48650
rect 20240 48640 20320 48650
rect 20420 48640 20500 48650
rect 20600 48640 20680 48650
rect 20780 48640 20860 48650
rect 20960 48640 21040 48650
rect 21140 48640 21220 48650
rect 21320 48640 21400 48650
rect 21500 48640 21580 48650
rect 21680 48640 21760 48650
rect 21860 48640 21940 48650
rect 22040 48640 22120 48650
rect 22220 48640 22300 48650
rect 22400 48640 22480 48650
rect 22580 48640 22660 48650
rect 22760 48640 22840 48650
rect 22940 48640 23020 48650
rect 23120 48640 23200 48650
rect 23300 48640 23380 48650
rect 23480 48640 23560 48650
rect 23660 48640 23740 48650
rect 23840 48640 23920 48650
rect 24020 48640 24100 48650
rect 24200 48640 24280 48650
rect 24380 48640 24460 48650
rect 24560 48640 24640 48650
rect 24740 48640 24820 48650
rect 24920 48640 25000 48650
rect 25100 48640 25180 48650
rect 25280 48640 25360 48650
rect 25460 48640 25540 48650
rect 25640 48640 25720 48650
rect 25820 48640 25900 48650
rect 26000 48640 26080 48650
rect 26180 48640 26260 48650
rect 26360 48640 26440 48650
rect 26540 48640 26620 48650
rect 30280 48640 30360 48650
rect 30460 48640 30540 48650
rect 30640 48640 30720 48650
rect 30820 48640 30900 48650
rect 31000 48640 31080 48650
rect 31180 48640 31260 48650
rect 31360 48640 31440 48650
rect 31540 48640 31620 48650
rect 31720 48640 31800 48650
rect 31900 48640 31980 48650
rect 32080 48640 32160 48650
rect 32260 48640 32340 48650
rect 32440 48640 32520 48650
rect 32620 48640 32700 48650
rect 32800 48640 32880 48650
rect 32980 48640 33060 48650
rect 33160 48640 33240 48650
rect 33340 48640 33420 48650
rect 33520 48640 33600 48650
rect 33700 48640 33780 48650
rect 33880 48640 33960 48650
rect 34060 48640 34140 48650
rect 34240 48640 34320 48650
rect 34420 48640 34500 48650
rect 34600 48640 34680 48650
rect 34780 48640 34860 48650
rect 34960 48640 35040 48650
rect 35140 48640 35220 48650
rect 35320 48640 35400 48650
rect 35500 48640 35580 48650
rect 35680 48640 35760 48650
rect 35860 48640 35940 48650
rect 36040 48640 36120 48650
rect 36220 48640 36300 48650
rect 36400 48640 36480 48650
rect 36580 48640 36660 48650
rect 36760 48640 36840 48650
rect 36940 48640 37020 48650
rect 37120 48640 37200 48650
rect 37300 48640 37380 48650
rect 37480 48640 37560 48650
rect 37660 48640 37740 48650
rect 37840 48640 37920 48650
rect 40060 48640 40140 48650
rect 40200 48640 40280 48650
rect 40340 48640 40420 48650
rect 40480 48640 40560 48650
rect 40620 48640 40700 48650
rect 40760 48640 40840 48650
rect 40900 48640 40980 48650
rect 41040 48640 41120 48650
rect 41180 48640 41260 48650
rect 41320 48640 41400 48650
rect 42360 48640 42440 48650
rect 42500 48640 42580 48650
rect 42640 48640 42720 48650
rect 42780 48640 42860 48650
rect 42920 48640 43000 48650
rect 43060 48640 43140 48650
rect 43200 48640 43280 48650
rect 43340 48640 43420 48650
rect 43480 48640 43560 48650
rect 43620 48640 43700 48650
rect 146300 48640 146380 48650
rect 146440 48640 146520 48650
rect 146580 48640 146660 48650
rect 146720 48640 146800 48650
rect 146860 48640 146940 48650
rect 147000 48640 147080 48650
rect 147140 48640 147220 48650
rect 147280 48640 147360 48650
rect 147420 48640 147500 48650
rect 147560 48640 147640 48650
rect 148600 48640 148680 48650
rect 148740 48640 148820 48650
rect 148880 48640 148960 48650
rect 149020 48640 149100 48650
rect 149160 48640 149240 48650
rect 149300 48640 149380 48650
rect 149440 48640 149520 48650
rect 149580 48640 149660 48650
rect 149720 48640 149800 48650
rect 149860 48640 149940 48650
rect 152080 48640 152160 48650
rect 152260 48640 152340 48650
rect 152440 48640 152520 48650
rect 152620 48640 152700 48650
rect 152800 48640 152880 48650
rect 152980 48640 153060 48650
rect 153160 48640 153240 48650
rect 153340 48640 153420 48650
rect 153520 48640 153600 48650
rect 153700 48640 153780 48650
rect 153880 48640 153960 48650
rect 154060 48640 154140 48650
rect 154240 48640 154320 48650
rect 154420 48640 154500 48650
rect 154600 48640 154680 48650
rect 154780 48640 154860 48650
rect 154960 48640 155040 48650
rect 155140 48640 155220 48650
rect 155320 48640 155400 48650
rect 155500 48640 155580 48650
rect 155680 48640 155760 48650
rect 155860 48640 155940 48650
rect 156040 48640 156120 48650
rect 156220 48640 156300 48650
rect 156400 48640 156480 48650
rect 156580 48640 156660 48650
rect 156760 48640 156840 48650
rect 156940 48640 157020 48650
rect 157120 48640 157200 48650
rect 157300 48640 157380 48650
rect 157480 48640 157560 48650
rect 157660 48640 157740 48650
rect 157840 48640 157920 48650
rect 158020 48640 158100 48650
rect 158200 48640 158280 48650
rect 158380 48640 158460 48650
rect 158560 48640 158640 48650
rect 158740 48640 158820 48650
rect 158920 48640 159000 48650
rect 159100 48640 159180 48650
rect 159280 48640 159360 48650
rect 159460 48640 159540 48650
rect 159640 48640 159720 48650
rect 163380 48640 163460 48650
rect 163560 48640 163640 48650
rect 163740 48640 163820 48650
rect 163920 48640 164000 48650
rect 164100 48640 164180 48650
rect 164280 48640 164360 48650
rect 164460 48640 164540 48650
rect 164640 48640 164720 48650
rect 164820 48640 164900 48650
rect 165000 48640 165080 48650
rect 165180 48640 165260 48650
rect 165360 48640 165440 48650
rect 165540 48640 165620 48650
rect 165720 48640 165800 48650
rect 165900 48640 165980 48650
rect 166080 48640 166160 48650
rect 166260 48640 166340 48650
rect 166440 48640 166520 48650
rect 166620 48640 166700 48650
rect 166800 48640 166880 48650
rect 166980 48640 167060 48650
rect 167160 48640 167240 48650
rect 167340 48640 167420 48650
rect 167520 48640 167600 48650
rect 167700 48640 167780 48650
rect 167880 48640 167960 48650
rect 168060 48640 168140 48650
rect 168240 48640 168320 48650
rect 168420 48640 168500 48650
rect 168600 48640 168680 48650
rect 168780 48640 168860 48650
rect 168960 48640 169040 48650
rect 169140 48640 169220 48650
rect 169320 48640 169400 48650
rect 169500 48640 169580 48650
rect 169680 48640 169760 48650
rect 169860 48640 169940 48650
rect 170040 48640 170120 48650
rect 170220 48640 170300 48650
rect 170400 48640 170480 48650
rect 170580 48640 170660 48650
rect 170760 48640 170840 48650
rect 170940 48640 171020 48650
rect 19060 48560 19070 48640
rect 19240 48560 19250 48640
rect 19420 48560 19430 48640
rect 19600 48560 19610 48640
rect 19780 48560 19790 48640
rect 19960 48560 19970 48640
rect 20140 48560 20150 48640
rect 20320 48560 20330 48640
rect 20500 48560 20510 48640
rect 20680 48560 20690 48640
rect 20860 48560 20870 48640
rect 21040 48560 21050 48640
rect 21220 48560 21230 48640
rect 21400 48560 21410 48640
rect 21580 48560 21590 48640
rect 21760 48560 21770 48640
rect 21940 48560 21950 48640
rect 22120 48560 22130 48640
rect 22300 48560 22310 48640
rect 22480 48560 22490 48640
rect 22660 48560 22670 48640
rect 22840 48560 22850 48640
rect 23020 48560 23030 48640
rect 23200 48560 23210 48640
rect 23380 48560 23390 48640
rect 23560 48560 23570 48640
rect 23740 48560 23750 48640
rect 23920 48560 23930 48640
rect 24100 48560 24110 48640
rect 24280 48560 24290 48640
rect 24460 48560 24470 48640
rect 24640 48560 24650 48640
rect 24820 48560 24830 48640
rect 25000 48560 25010 48640
rect 25180 48560 25190 48640
rect 25360 48560 25370 48640
rect 25540 48560 25550 48640
rect 25720 48560 25730 48640
rect 25900 48560 25910 48640
rect 26080 48560 26090 48640
rect 26260 48560 26270 48640
rect 26440 48560 26450 48640
rect 26620 48560 26630 48640
rect 30360 48560 30370 48640
rect 30540 48560 30550 48640
rect 30720 48560 30730 48640
rect 30900 48560 30910 48640
rect 31080 48560 31090 48640
rect 31260 48560 31270 48640
rect 31440 48560 31450 48640
rect 31620 48560 31630 48640
rect 31800 48560 31810 48640
rect 31980 48560 31990 48640
rect 32160 48560 32170 48640
rect 32340 48560 32350 48640
rect 32520 48560 32530 48640
rect 32700 48560 32710 48640
rect 32880 48560 32890 48640
rect 33060 48560 33070 48640
rect 33240 48560 33250 48640
rect 33420 48560 33430 48640
rect 33600 48560 33610 48640
rect 33780 48560 33790 48640
rect 33960 48560 33970 48640
rect 34140 48560 34150 48640
rect 34320 48560 34330 48640
rect 34500 48560 34510 48640
rect 34680 48560 34690 48640
rect 34860 48560 34870 48640
rect 35040 48560 35050 48640
rect 35220 48560 35230 48640
rect 35400 48560 35410 48640
rect 35580 48560 35590 48640
rect 35760 48560 35770 48640
rect 35940 48560 35950 48640
rect 36120 48560 36130 48640
rect 36300 48560 36310 48640
rect 36480 48560 36490 48640
rect 36660 48560 36670 48640
rect 36840 48560 36850 48640
rect 37020 48560 37030 48640
rect 37200 48560 37210 48640
rect 37380 48560 37390 48640
rect 37560 48560 37570 48640
rect 37740 48560 37750 48640
rect 37920 48560 37930 48640
rect 40140 48560 40150 48640
rect 40280 48560 40290 48640
rect 40420 48560 40430 48640
rect 40560 48560 40570 48640
rect 40700 48560 40710 48640
rect 40840 48560 40850 48640
rect 40980 48560 40990 48640
rect 41120 48560 41130 48640
rect 41260 48560 41270 48640
rect 41400 48560 41410 48640
rect 42440 48560 42450 48640
rect 42580 48560 42590 48640
rect 42720 48560 42730 48640
rect 42860 48560 42870 48640
rect 43000 48560 43010 48640
rect 43140 48560 43150 48640
rect 43280 48560 43290 48640
rect 43420 48560 43430 48640
rect 43560 48560 43570 48640
rect 43700 48560 43710 48640
rect 146380 48560 146390 48640
rect 146520 48560 146530 48640
rect 146660 48560 146670 48640
rect 146800 48560 146810 48640
rect 146940 48560 146950 48640
rect 147080 48560 147090 48640
rect 147220 48560 147230 48640
rect 147360 48560 147370 48640
rect 147500 48560 147510 48640
rect 147640 48560 147650 48640
rect 148680 48560 148690 48640
rect 148820 48560 148830 48640
rect 148960 48560 148970 48640
rect 149100 48560 149110 48640
rect 149240 48560 149250 48640
rect 149380 48560 149390 48640
rect 149520 48560 149530 48640
rect 149660 48560 149670 48640
rect 149800 48560 149810 48640
rect 149940 48560 149950 48640
rect 152160 48560 152170 48640
rect 152340 48560 152350 48640
rect 152520 48560 152530 48640
rect 152700 48560 152710 48640
rect 152880 48560 152890 48640
rect 153060 48560 153070 48640
rect 153240 48560 153250 48640
rect 153420 48560 153430 48640
rect 153600 48560 153610 48640
rect 153780 48560 153790 48640
rect 153960 48560 153970 48640
rect 154140 48560 154150 48640
rect 154320 48560 154330 48640
rect 154500 48560 154510 48640
rect 154680 48560 154690 48640
rect 154860 48560 154870 48640
rect 155040 48560 155050 48640
rect 155220 48560 155230 48640
rect 155400 48560 155410 48640
rect 155580 48560 155590 48640
rect 155760 48560 155770 48640
rect 155940 48560 155950 48640
rect 156120 48560 156130 48640
rect 156300 48560 156310 48640
rect 156480 48560 156490 48640
rect 156660 48560 156670 48640
rect 156840 48560 156850 48640
rect 157020 48560 157030 48640
rect 157200 48560 157210 48640
rect 157380 48560 157390 48640
rect 157560 48560 157570 48640
rect 157740 48560 157750 48640
rect 157920 48560 157930 48640
rect 158100 48560 158110 48640
rect 158280 48560 158290 48640
rect 158460 48560 158470 48640
rect 158640 48560 158650 48640
rect 158820 48560 158830 48640
rect 159000 48560 159010 48640
rect 159180 48560 159190 48640
rect 159360 48560 159370 48640
rect 159540 48560 159550 48640
rect 159720 48560 159730 48640
rect 163460 48560 163470 48640
rect 163640 48560 163650 48640
rect 163820 48560 163830 48640
rect 164000 48560 164010 48640
rect 164180 48560 164190 48640
rect 164360 48560 164370 48640
rect 164540 48560 164550 48640
rect 164720 48560 164730 48640
rect 164900 48560 164910 48640
rect 165080 48560 165090 48640
rect 165260 48560 165270 48640
rect 165440 48560 165450 48640
rect 165620 48560 165630 48640
rect 165800 48560 165810 48640
rect 165980 48560 165990 48640
rect 166160 48560 166170 48640
rect 166340 48560 166350 48640
rect 166520 48560 166530 48640
rect 166700 48560 166710 48640
rect 166880 48560 166890 48640
rect 167060 48560 167070 48640
rect 167240 48560 167250 48640
rect 167420 48560 167430 48640
rect 167600 48560 167610 48640
rect 167780 48560 167790 48640
rect 167960 48560 167970 48640
rect 168140 48560 168150 48640
rect 168320 48560 168330 48640
rect 168500 48560 168510 48640
rect 168680 48560 168690 48640
rect 168860 48560 168870 48640
rect 169040 48560 169050 48640
rect 169220 48560 169230 48640
rect 169400 48560 169410 48640
rect 169580 48560 169590 48640
rect 169760 48560 169770 48640
rect 169940 48560 169950 48640
rect 170120 48560 170130 48640
rect 170300 48560 170310 48640
rect 170480 48560 170490 48640
rect 170660 48560 170670 48640
rect 170840 48560 170850 48640
rect 171020 48560 171030 48640
rect 30360 48455 30440 48465
rect 30680 48455 30760 48465
rect 31000 48455 31080 48465
rect 31320 48455 31400 48465
rect 31640 48455 31720 48465
rect 31960 48455 32040 48465
rect 32280 48455 32360 48465
rect 32600 48455 32680 48465
rect 32920 48455 33000 48465
rect 33240 48455 33320 48465
rect 33560 48455 33640 48465
rect 33880 48455 33960 48465
rect 34200 48455 34280 48465
rect 34520 48455 34600 48465
rect 34840 48455 34920 48465
rect 35160 48455 35240 48465
rect 35480 48455 35560 48465
rect 35800 48455 35880 48465
rect 36120 48455 36200 48465
rect 36440 48455 36520 48465
rect 36760 48455 36840 48465
rect 37080 48455 37160 48465
rect 37400 48455 37480 48465
rect 37720 48455 37800 48465
rect 40180 48455 40260 48465
rect 40500 48455 40580 48465
rect 40820 48455 40900 48465
rect 41140 48455 41220 48465
rect 42560 48455 42640 48465
rect 42880 48455 42960 48465
rect 43200 48455 43280 48465
rect 43520 48455 43600 48465
rect 146400 48455 146480 48465
rect 146720 48455 146800 48465
rect 147040 48455 147120 48465
rect 147360 48455 147440 48465
rect 148780 48455 148860 48465
rect 149100 48455 149180 48465
rect 149420 48455 149500 48465
rect 149740 48455 149820 48465
rect 152200 48455 152280 48465
rect 152520 48455 152600 48465
rect 152840 48455 152920 48465
rect 153160 48455 153240 48465
rect 153480 48455 153560 48465
rect 153800 48455 153880 48465
rect 154120 48455 154200 48465
rect 154440 48455 154520 48465
rect 154760 48455 154840 48465
rect 155080 48455 155160 48465
rect 155400 48455 155480 48465
rect 155720 48455 155800 48465
rect 156040 48455 156120 48465
rect 156360 48455 156440 48465
rect 156680 48455 156760 48465
rect 157000 48455 157080 48465
rect 157320 48455 157400 48465
rect 157640 48455 157720 48465
rect 157960 48455 158040 48465
rect 158280 48455 158360 48465
rect 158600 48455 158680 48465
rect 158920 48455 159000 48465
rect 159240 48455 159320 48465
rect 159560 48455 159640 48465
rect 30440 48375 30450 48455
rect 30760 48375 30770 48455
rect 31080 48375 31090 48455
rect 31400 48375 31410 48455
rect 31720 48375 31730 48455
rect 32040 48375 32050 48455
rect 32360 48375 32370 48455
rect 32680 48375 32690 48455
rect 33000 48375 33010 48455
rect 33320 48375 33330 48455
rect 33640 48375 33650 48455
rect 33960 48375 33970 48455
rect 34280 48375 34290 48455
rect 34600 48375 34610 48455
rect 34920 48375 34930 48455
rect 35240 48375 35250 48455
rect 35560 48375 35570 48455
rect 35880 48375 35890 48455
rect 36200 48375 36210 48455
rect 36520 48375 36530 48455
rect 36840 48375 36850 48455
rect 37160 48375 37170 48455
rect 37480 48375 37490 48455
rect 37800 48375 37810 48455
rect 40260 48375 40270 48455
rect 40580 48375 40590 48455
rect 40900 48375 40910 48455
rect 41220 48375 41230 48455
rect 42640 48375 42650 48455
rect 42960 48375 42970 48455
rect 43280 48375 43290 48455
rect 43600 48375 43610 48455
rect 146480 48375 146490 48455
rect 146800 48375 146810 48455
rect 147120 48375 147130 48455
rect 147440 48375 147450 48455
rect 148860 48375 148870 48455
rect 149180 48375 149190 48455
rect 149500 48375 149510 48455
rect 149820 48375 149830 48455
rect 152280 48375 152290 48455
rect 152600 48375 152610 48455
rect 152920 48375 152930 48455
rect 153240 48375 153250 48455
rect 153560 48375 153570 48455
rect 153880 48375 153890 48455
rect 154200 48375 154210 48455
rect 154520 48375 154530 48455
rect 154840 48375 154850 48455
rect 155160 48375 155170 48455
rect 155480 48375 155490 48455
rect 155800 48375 155810 48455
rect 156120 48375 156130 48455
rect 156440 48375 156450 48455
rect 156760 48375 156770 48455
rect 157080 48375 157090 48455
rect 157400 48375 157410 48455
rect 157720 48375 157730 48455
rect 158040 48375 158050 48455
rect 158360 48375 158370 48455
rect 158680 48375 158690 48455
rect 159000 48375 159010 48455
rect 159320 48375 159330 48455
rect 159640 48375 159650 48455
rect 19130 48335 19210 48345
rect 19450 48335 19530 48345
rect 19770 48335 19850 48345
rect 20090 48335 20170 48345
rect 20410 48335 20490 48345
rect 20730 48335 20810 48345
rect 21050 48335 21130 48345
rect 21370 48335 21450 48345
rect 21690 48335 21770 48345
rect 22010 48335 22090 48345
rect 22330 48335 22410 48345
rect 22650 48335 22730 48345
rect 22970 48335 23050 48345
rect 23290 48335 23370 48345
rect 23610 48335 23690 48345
rect 23930 48335 24010 48345
rect 24250 48335 24330 48345
rect 24570 48335 24650 48345
rect 24890 48335 24970 48345
rect 25210 48335 25290 48345
rect 25530 48335 25610 48345
rect 25850 48335 25930 48345
rect 26170 48335 26250 48345
rect 163750 48335 163830 48345
rect 164070 48335 164150 48345
rect 164390 48335 164470 48345
rect 164710 48335 164790 48345
rect 165030 48335 165110 48345
rect 165350 48335 165430 48345
rect 165670 48335 165750 48345
rect 165990 48335 166070 48345
rect 166310 48335 166390 48345
rect 166630 48335 166710 48345
rect 166950 48335 167030 48345
rect 167270 48335 167350 48345
rect 167590 48335 167670 48345
rect 167910 48335 167990 48345
rect 168230 48335 168310 48345
rect 168550 48335 168630 48345
rect 168870 48335 168950 48345
rect 169190 48335 169270 48345
rect 169510 48335 169590 48345
rect 169830 48335 169910 48345
rect 170150 48335 170230 48345
rect 170470 48335 170550 48345
rect 170790 48335 170870 48345
rect 19210 48255 19220 48335
rect 19530 48255 19540 48335
rect 19850 48255 19860 48335
rect 20170 48255 20180 48335
rect 20490 48255 20500 48335
rect 20810 48255 20820 48335
rect 21130 48255 21140 48335
rect 21450 48255 21460 48335
rect 21770 48255 21780 48335
rect 22090 48255 22100 48335
rect 22410 48255 22420 48335
rect 22730 48255 22740 48335
rect 23050 48255 23060 48335
rect 23370 48255 23380 48335
rect 23690 48255 23700 48335
rect 24010 48255 24020 48335
rect 24330 48255 24340 48335
rect 24650 48255 24660 48335
rect 24970 48255 24980 48335
rect 25290 48255 25300 48335
rect 25610 48255 25620 48335
rect 25930 48255 25940 48335
rect 26250 48255 26260 48335
rect 30520 48295 30600 48305
rect 30840 48295 30920 48305
rect 31160 48295 31240 48305
rect 31480 48295 31560 48305
rect 31800 48295 31880 48305
rect 32120 48295 32200 48305
rect 32440 48295 32520 48305
rect 32760 48295 32840 48305
rect 33080 48295 33160 48305
rect 33400 48295 33480 48305
rect 33720 48295 33800 48305
rect 34040 48295 34120 48305
rect 34360 48295 34440 48305
rect 34680 48295 34760 48305
rect 35000 48295 35080 48305
rect 35320 48295 35400 48305
rect 35640 48295 35720 48305
rect 35960 48295 36040 48305
rect 36280 48295 36360 48305
rect 36600 48295 36680 48305
rect 36920 48295 37000 48305
rect 37240 48295 37320 48305
rect 37560 48295 37640 48305
rect 40340 48295 40420 48305
rect 40660 48295 40740 48305
rect 40980 48295 41060 48305
rect 42720 48295 42800 48305
rect 43040 48295 43120 48305
rect 43360 48295 43440 48305
rect 146560 48295 146640 48305
rect 146880 48295 146960 48305
rect 147200 48295 147280 48305
rect 148940 48295 149020 48305
rect 149260 48295 149340 48305
rect 149580 48295 149660 48305
rect 152360 48295 152440 48305
rect 152680 48295 152760 48305
rect 153000 48295 153080 48305
rect 153320 48295 153400 48305
rect 153640 48295 153720 48305
rect 153960 48295 154040 48305
rect 154280 48295 154360 48305
rect 154600 48295 154680 48305
rect 154920 48295 155000 48305
rect 155240 48295 155320 48305
rect 155560 48295 155640 48305
rect 155880 48295 155960 48305
rect 156200 48295 156280 48305
rect 156520 48295 156600 48305
rect 156840 48295 156920 48305
rect 157160 48295 157240 48305
rect 157480 48295 157560 48305
rect 157800 48295 157880 48305
rect 158120 48295 158200 48305
rect 158440 48295 158520 48305
rect 158760 48295 158840 48305
rect 159080 48295 159160 48305
rect 159400 48295 159480 48305
rect 30600 48215 30610 48295
rect 30920 48215 30930 48295
rect 31240 48215 31250 48295
rect 31560 48215 31570 48295
rect 31880 48215 31890 48295
rect 32200 48215 32210 48295
rect 32520 48215 32530 48295
rect 32840 48215 32850 48295
rect 33160 48215 33170 48295
rect 33480 48215 33490 48295
rect 33800 48215 33810 48295
rect 34120 48215 34130 48295
rect 34440 48215 34450 48295
rect 34760 48215 34770 48295
rect 35080 48215 35090 48295
rect 35400 48215 35410 48295
rect 35720 48215 35730 48295
rect 36040 48215 36050 48295
rect 36360 48215 36370 48295
rect 36680 48215 36690 48295
rect 37000 48215 37010 48295
rect 37320 48215 37330 48295
rect 37640 48215 37650 48295
rect 40420 48215 40430 48295
rect 40740 48215 40750 48295
rect 41060 48215 41070 48295
rect 42800 48215 42810 48295
rect 43120 48215 43130 48295
rect 43440 48215 43450 48295
rect 146640 48215 146650 48295
rect 146960 48215 146970 48295
rect 147280 48215 147290 48295
rect 149020 48215 149030 48295
rect 149340 48215 149350 48295
rect 149660 48215 149670 48295
rect 152440 48215 152450 48295
rect 152760 48215 152770 48295
rect 153080 48215 153090 48295
rect 153400 48215 153410 48295
rect 153720 48215 153730 48295
rect 154040 48215 154050 48295
rect 154360 48215 154370 48295
rect 154680 48215 154690 48295
rect 155000 48215 155010 48295
rect 155320 48215 155330 48295
rect 155640 48215 155650 48295
rect 155960 48215 155970 48295
rect 156280 48215 156290 48295
rect 156600 48215 156610 48295
rect 156920 48215 156930 48295
rect 157240 48215 157250 48295
rect 157560 48215 157570 48295
rect 157880 48215 157890 48295
rect 158200 48215 158210 48295
rect 158520 48215 158530 48295
rect 158840 48215 158850 48295
rect 159160 48215 159170 48295
rect 159480 48215 159490 48295
rect 163830 48255 163840 48335
rect 164150 48255 164160 48335
rect 164470 48255 164480 48335
rect 164790 48255 164800 48335
rect 165110 48255 165120 48335
rect 165430 48255 165440 48335
rect 165750 48255 165760 48335
rect 166070 48255 166080 48335
rect 166390 48255 166400 48335
rect 166710 48255 166720 48335
rect 167030 48255 167040 48335
rect 167350 48255 167360 48335
rect 167670 48255 167680 48335
rect 167990 48255 168000 48335
rect 168310 48255 168320 48335
rect 168630 48255 168640 48335
rect 168950 48255 168960 48335
rect 169270 48255 169280 48335
rect 169590 48255 169600 48335
rect 169910 48255 169920 48335
rect 170230 48255 170240 48335
rect 170550 48255 170560 48335
rect 170870 48255 170880 48335
rect 18970 48175 19050 48185
rect 19290 48175 19370 48185
rect 19610 48175 19690 48185
rect 19930 48175 20010 48185
rect 20250 48175 20330 48185
rect 20570 48175 20650 48185
rect 20890 48175 20970 48185
rect 21210 48175 21290 48185
rect 21530 48175 21610 48185
rect 21850 48175 21930 48185
rect 22170 48175 22250 48185
rect 22490 48175 22570 48185
rect 22810 48175 22890 48185
rect 23130 48175 23210 48185
rect 23450 48175 23530 48185
rect 23770 48175 23850 48185
rect 24090 48175 24170 48185
rect 24410 48175 24490 48185
rect 24730 48175 24810 48185
rect 25050 48175 25130 48185
rect 25370 48175 25450 48185
rect 25690 48175 25770 48185
rect 26010 48175 26090 48185
rect 26330 48175 26410 48185
rect 163590 48175 163670 48185
rect 163910 48175 163990 48185
rect 164230 48175 164310 48185
rect 164550 48175 164630 48185
rect 164870 48175 164950 48185
rect 165190 48175 165270 48185
rect 165510 48175 165590 48185
rect 165830 48175 165910 48185
rect 166150 48175 166230 48185
rect 166470 48175 166550 48185
rect 166790 48175 166870 48185
rect 167110 48175 167190 48185
rect 167430 48175 167510 48185
rect 167750 48175 167830 48185
rect 168070 48175 168150 48185
rect 168390 48175 168470 48185
rect 168710 48175 168790 48185
rect 169030 48175 169110 48185
rect 169350 48175 169430 48185
rect 169670 48175 169750 48185
rect 169990 48175 170070 48185
rect 170310 48175 170390 48185
rect 170630 48175 170710 48185
rect 170950 48175 171030 48185
rect 19050 48095 19060 48175
rect 19370 48095 19380 48175
rect 19690 48095 19700 48175
rect 20010 48095 20020 48175
rect 20330 48095 20340 48175
rect 20650 48095 20660 48175
rect 20970 48095 20980 48175
rect 21290 48095 21300 48175
rect 21610 48095 21620 48175
rect 21930 48095 21940 48175
rect 22250 48095 22260 48175
rect 22570 48095 22580 48175
rect 22890 48095 22900 48175
rect 23210 48095 23220 48175
rect 23530 48095 23540 48175
rect 23850 48095 23860 48175
rect 24170 48095 24180 48175
rect 24490 48095 24500 48175
rect 24810 48095 24820 48175
rect 25130 48095 25140 48175
rect 25450 48095 25460 48175
rect 25770 48095 25780 48175
rect 26090 48095 26100 48175
rect 26410 48095 26420 48175
rect 30360 48135 30440 48145
rect 30680 48135 30760 48145
rect 31000 48135 31080 48145
rect 31320 48135 31400 48145
rect 31640 48135 31720 48145
rect 31960 48135 32040 48145
rect 32280 48135 32360 48145
rect 32600 48135 32680 48145
rect 32920 48135 33000 48145
rect 33240 48135 33320 48145
rect 33560 48135 33640 48145
rect 33880 48135 33960 48145
rect 34200 48135 34280 48145
rect 34520 48135 34600 48145
rect 34840 48135 34920 48145
rect 35160 48135 35240 48145
rect 35480 48135 35560 48145
rect 35800 48135 35880 48145
rect 36120 48135 36200 48145
rect 36440 48135 36520 48145
rect 36760 48135 36840 48145
rect 37080 48135 37160 48145
rect 37400 48135 37480 48145
rect 37720 48135 37800 48145
rect 40180 48135 40260 48145
rect 40500 48135 40580 48145
rect 40820 48135 40900 48145
rect 41140 48135 41220 48145
rect 42560 48135 42640 48145
rect 42880 48135 42960 48145
rect 43200 48135 43280 48145
rect 43520 48135 43600 48145
rect 146400 48135 146480 48145
rect 146720 48135 146800 48145
rect 147040 48135 147120 48145
rect 147360 48135 147440 48145
rect 148780 48135 148860 48145
rect 149100 48135 149180 48145
rect 149420 48135 149500 48145
rect 149740 48135 149820 48145
rect 152200 48135 152280 48145
rect 152520 48135 152600 48145
rect 152840 48135 152920 48145
rect 153160 48135 153240 48145
rect 153480 48135 153560 48145
rect 153800 48135 153880 48145
rect 154120 48135 154200 48145
rect 154440 48135 154520 48145
rect 154760 48135 154840 48145
rect 155080 48135 155160 48145
rect 155400 48135 155480 48145
rect 155720 48135 155800 48145
rect 156040 48135 156120 48145
rect 156360 48135 156440 48145
rect 156680 48135 156760 48145
rect 157000 48135 157080 48145
rect 157320 48135 157400 48145
rect 157640 48135 157720 48145
rect 157960 48135 158040 48145
rect 158280 48135 158360 48145
rect 158600 48135 158680 48145
rect 158920 48135 159000 48145
rect 159240 48135 159320 48145
rect 159560 48135 159640 48145
rect 30440 48055 30450 48135
rect 30760 48055 30770 48135
rect 31080 48055 31090 48135
rect 31400 48055 31410 48135
rect 31720 48055 31730 48135
rect 32040 48055 32050 48135
rect 32360 48055 32370 48135
rect 32680 48055 32690 48135
rect 33000 48055 33010 48135
rect 33320 48055 33330 48135
rect 33640 48055 33650 48135
rect 33960 48055 33970 48135
rect 34280 48055 34290 48135
rect 34600 48055 34610 48135
rect 34920 48055 34930 48135
rect 35240 48055 35250 48135
rect 35560 48055 35570 48135
rect 35880 48055 35890 48135
rect 36200 48055 36210 48135
rect 36520 48055 36530 48135
rect 36840 48055 36850 48135
rect 37160 48055 37170 48135
rect 37480 48055 37490 48135
rect 37800 48055 37810 48135
rect 40260 48055 40270 48135
rect 40580 48055 40590 48135
rect 40900 48055 40910 48135
rect 41220 48055 41230 48135
rect 42640 48055 42650 48135
rect 42960 48055 42970 48135
rect 43280 48055 43290 48135
rect 43600 48055 43610 48135
rect 146480 48055 146490 48135
rect 146800 48055 146810 48135
rect 147120 48055 147130 48135
rect 147440 48055 147450 48135
rect 148860 48055 148870 48135
rect 149180 48055 149190 48135
rect 149500 48055 149510 48135
rect 149820 48055 149830 48135
rect 152280 48055 152290 48135
rect 152600 48055 152610 48135
rect 152920 48055 152930 48135
rect 153240 48055 153250 48135
rect 153560 48055 153570 48135
rect 153880 48055 153890 48135
rect 154200 48055 154210 48135
rect 154520 48055 154530 48135
rect 154840 48055 154850 48135
rect 155160 48055 155170 48135
rect 155480 48055 155490 48135
rect 155800 48055 155810 48135
rect 156120 48055 156130 48135
rect 156440 48055 156450 48135
rect 156760 48055 156770 48135
rect 157080 48055 157090 48135
rect 157400 48055 157410 48135
rect 157720 48055 157730 48135
rect 158040 48055 158050 48135
rect 158360 48055 158370 48135
rect 158680 48055 158690 48135
rect 159000 48055 159010 48135
rect 159320 48055 159330 48135
rect 159640 48055 159650 48135
rect 163670 48095 163680 48175
rect 163990 48095 164000 48175
rect 164310 48095 164320 48175
rect 164630 48095 164640 48175
rect 164950 48095 164960 48175
rect 165270 48095 165280 48175
rect 165590 48095 165600 48175
rect 165910 48095 165920 48175
rect 166230 48095 166240 48175
rect 166550 48095 166560 48175
rect 166870 48095 166880 48175
rect 167190 48095 167200 48175
rect 167510 48095 167520 48175
rect 167830 48095 167840 48175
rect 168150 48095 168160 48175
rect 168470 48095 168480 48175
rect 168790 48095 168800 48175
rect 169110 48095 169120 48175
rect 169430 48095 169440 48175
rect 169750 48095 169760 48175
rect 170070 48095 170080 48175
rect 170390 48095 170400 48175
rect 170710 48095 170720 48175
rect 171030 48095 171040 48175
rect 19130 48015 19210 48025
rect 19450 48015 19530 48025
rect 19770 48015 19850 48025
rect 20090 48015 20170 48025
rect 20410 48015 20490 48025
rect 20730 48015 20810 48025
rect 21050 48015 21130 48025
rect 21370 48015 21450 48025
rect 21690 48015 21770 48025
rect 22010 48015 22090 48025
rect 22330 48015 22410 48025
rect 22650 48015 22730 48025
rect 22970 48015 23050 48025
rect 23290 48015 23370 48025
rect 23610 48015 23690 48025
rect 23930 48015 24010 48025
rect 24250 48015 24330 48025
rect 24570 48015 24650 48025
rect 24890 48015 24970 48025
rect 25210 48015 25290 48025
rect 25530 48015 25610 48025
rect 25850 48015 25930 48025
rect 26170 48015 26250 48025
rect 163750 48015 163830 48025
rect 164070 48015 164150 48025
rect 164390 48015 164470 48025
rect 164710 48015 164790 48025
rect 165030 48015 165110 48025
rect 165350 48015 165430 48025
rect 165670 48015 165750 48025
rect 165990 48015 166070 48025
rect 166310 48015 166390 48025
rect 166630 48015 166710 48025
rect 166950 48015 167030 48025
rect 167270 48015 167350 48025
rect 167590 48015 167670 48025
rect 167910 48015 167990 48025
rect 168230 48015 168310 48025
rect 168550 48015 168630 48025
rect 168870 48015 168950 48025
rect 169190 48015 169270 48025
rect 169510 48015 169590 48025
rect 169830 48015 169910 48025
rect 170150 48015 170230 48025
rect 170470 48015 170550 48025
rect 170790 48015 170870 48025
rect 19210 47935 19220 48015
rect 19530 47935 19540 48015
rect 19850 47935 19860 48015
rect 20170 47935 20180 48015
rect 20490 47935 20500 48015
rect 20810 47935 20820 48015
rect 21130 47935 21140 48015
rect 21450 47935 21460 48015
rect 21770 47935 21780 48015
rect 22090 47935 22100 48015
rect 22410 47935 22420 48015
rect 22730 47935 22740 48015
rect 23050 47935 23060 48015
rect 23370 47935 23380 48015
rect 23690 47935 23700 48015
rect 24010 47935 24020 48015
rect 24330 47935 24340 48015
rect 24650 47935 24660 48015
rect 24970 47935 24980 48015
rect 25290 47935 25300 48015
rect 25610 47935 25620 48015
rect 25930 47935 25940 48015
rect 26250 47935 26260 48015
rect 30520 47975 30600 47985
rect 30840 47975 30920 47985
rect 31160 47975 31240 47985
rect 31480 47975 31560 47985
rect 31800 47975 31880 47985
rect 32120 47975 32200 47985
rect 32440 47975 32520 47985
rect 32760 47975 32840 47985
rect 33080 47975 33160 47985
rect 33400 47975 33480 47985
rect 33720 47975 33800 47985
rect 34040 47975 34120 47985
rect 34360 47975 34440 47985
rect 34680 47975 34760 47985
rect 35000 47975 35080 47985
rect 35320 47975 35400 47985
rect 35640 47975 35720 47985
rect 35960 47975 36040 47985
rect 36280 47975 36360 47985
rect 36600 47975 36680 47985
rect 36920 47975 37000 47985
rect 37240 47975 37320 47985
rect 37560 47975 37640 47985
rect 40340 47975 40420 47985
rect 40660 47975 40740 47985
rect 40980 47975 41060 47985
rect 42720 47975 42800 47985
rect 43040 47975 43120 47985
rect 43360 47975 43440 47985
rect 146560 47975 146640 47985
rect 146880 47975 146960 47985
rect 147200 47975 147280 47985
rect 148940 47975 149020 47985
rect 149260 47975 149340 47985
rect 149580 47975 149660 47985
rect 152360 47975 152440 47985
rect 152680 47975 152760 47985
rect 153000 47975 153080 47985
rect 153320 47975 153400 47985
rect 153640 47975 153720 47985
rect 153960 47975 154040 47985
rect 154280 47975 154360 47985
rect 154600 47975 154680 47985
rect 154920 47975 155000 47985
rect 155240 47975 155320 47985
rect 155560 47975 155640 47985
rect 155880 47975 155960 47985
rect 156200 47975 156280 47985
rect 156520 47975 156600 47985
rect 156840 47975 156920 47985
rect 157160 47975 157240 47985
rect 157480 47975 157560 47985
rect 157800 47975 157880 47985
rect 158120 47975 158200 47985
rect 158440 47975 158520 47985
rect 158760 47975 158840 47985
rect 159080 47975 159160 47985
rect 159400 47975 159480 47985
rect 30600 47895 30610 47975
rect 30920 47895 30930 47975
rect 31240 47895 31250 47975
rect 31560 47895 31570 47975
rect 31880 47895 31890 47975
rect 32200 47895 32210 47975
rect 32520 47895 32530 47975
rect 32840 47895 32850 47975
rect 33160 47895 33170 47975
rect 33480 47895 33490 47975
rect 33800 47895 33810 47975
rect 34120 47895 34130 47975
rect 34440 47895 34450 47975
rect 34760 47895 34770 47975
rect 35080 47895 35090 47975
rect 35400 47895 35410 47975
rect 35720 47895 35730 47975
rect 36040 47895 36050 47975
rect 36360 47895 36370 47975
rect 36680 47895 36690 47975
rect 37000 47895 37010 47975
rect 37320 47895 37330 47975
rect 37640 47895 37650 47975
rect 40420 47895 40430 47975
rect 40740 47895 40750 47975
rect 41060 47895 41070 47975
rect 42800 47895 42810 47975
rect 43120 47895 43130 47975
rect 43440 47895 43450 47975
rect 146640 47895 146650 47975
rect 146960 47895 146970 47975
rect 147280 47895 147290 47975
rect 149020 47895 149030 47975
rect 149340 47895 149350 47975
rect 149660 47895 149670 47975
rect 152440 47895 152450 47975
rect 152760 47895 152770 47975
rect 153080 47895 153090 47975
rect 153400 47895 153410 47975
rect 153720 47895 153730 47975
rect 154040 47895 154050 47975
rect 154360 47895 154370 47975
rect 154680 47895 154690 47975
rect 155000 47895 155010 47975
rect 155320 47895 155330 47975
rect 155640 47895 155650 47975
rect 155960 47895 155970 47975
rect 156280 47895 156290 47975
rect 156600 47895 156610 47975
rect 156920 47895 156930 47975
rect 157240 47895 157250 47975
rect 157560 47895 157570 47975
rect 157880 47895 157890 47975
rect 158200 47895 158210 47975
rect 158520 47895 158530 47975
rect 158840 47895 158850 47975
rect 159160 47895 159170 47975
rect 159480 47895 159490 47975
rect 163830 47935 163840 48015
rect 164150 47935 164160 48015
rect 164470 47935 164480 48015
rect 164790 47935 164800 48015
rect 165110 47935 165120 48015
rect 165430 47935 165440 48015
rect 165750 47935 165760 48015
rect 166070 47935 166080 48015
rect 166390 47935 166400 48015
rect 166710 47935 166720 48015
rect 167030 47935 167040 48015
rect 167350 47935 167360 48015
rect 167670 47935 167680 48015
rect 167990 47935 168000 48015
rect 168310 47935 168320 48015
rect 168630 47935 168640 48015
rect 168950 47935 168960 48015
rect 169270 47935 169280 48015
rect 169590 47935 169600 48015
rect 169910 47935 169920 48015
rect 170230 47935 170240 48015
rect 170550 47935 170560 48015
rect 170870 47935 170880 48015
rect 18970 47855 19050 47865
rect 19290 47855 19370 47865
rect 19610 47855 19690 47865
rect 19930 47855 20010 47865
rect 20250 47855 20330 47865
rect 20570 47855 20650 47865
rect 20890 47855 20970 47865
rect 21210 47855 21290 47865
rect 21530 47855 21610 47865
rect 21850 47855 21930 47865
rect 22170 47855 22250 47865
rect 22490 47855 22570 47865
rect 22810 47855 22890 47865
rect 23130 47855 23210 47865
rect 23450 47855 23530 47865
rect 23770 47855 23850 47865
rect 24090 47855 24170 47865
rect 24410 47855 24490 47865
rect 24730 47855 24810 47865
rect 25050 47855 25130 47865
rect 25370 47855 25450 47865
rect 25690 47855 25770 47865
rect 26010 47855 26090 47865
rect 26330 47855 26410 47865
rect 163590 47855 163670 47865
rect 163910 47855 163990 47865
rect 164230 47855 164310 47865
rect 164550 47855 164630 47865
rect 164870 47855 164950 47865
rect 165190 47855 165270 47865
rect 165510 47855 165590 47865
rect 165830 47855 165910 47865
rect 166150 47855 166230 47865
rect 166470 47855 166550 47865
rect 166790 47855 166870 47865
rect 167110 47855 167190 47865
rect 167430 47855 167510 47865
rect 167750 47855 167830 47865
rect 168070 47855 168150 47865
rect 168390 47855 168470 47865
rect 168710 47855 168790 47865
rect 169030 47855 169110 47865
rect 169350 47855 169430 47865
rect 169670 47855 169750 47865
rect 169990 47855 170070 47865
rect 170310 47855 170390 47865
rect 170630 47855 170710 47865
rect 170950 47855 171030 47865
rect 19050 47775 19060 47855
rect 19370 47775 19380 47855
rect 19690 47775 19700 47855
rect 20010 47775 20020 47855
rect 20330 47775 20340 47855
rect 20650 47775 20660 47855
rect 20970 47775 20980 47855
rect 21290 47775 21300 47855
rect 21610 47775 21620 47855
rect 21930 47775 21940 47855
rect 22250 47775 22260 47855
rect 22570 47775 22580 47855
rect 22890 47775 22900 47855
rect 23210 47775 23220 47855
rect 23530 47775 23540 47855
rect 23850 47775 23860 47855
rect 24170 47775 24180 47855
rect 24490 47775 24500 47855
rect 24810 47775 24820 47855
rect 25130 47775 25140 47855
rect 25450 47775 25460 47855
rect 25770 47775 25780 47855
rect 26090 47775 26100 47855
rect 26410 47775 26420 47855
rect 30360 47815 30440 47825
rect 30680 47815 30760 47825
rect 31000 47815 31080 47825
rect 31320 47815 31400 47825
rect 31640 47815 31720 47825
rect 31960 47815 32040 47825
rect 32280 47815 32360 47825
rect 32600 47815 32680 47825
rect 32920 47815 33000 47825
rect 33240 47815 33320 47825
rect 33560 47815 33640 47825
rect 33880 47815 33960 47825
rect 34200 47815 34280 47825
rect 34520 47815 34600 47825
rect 34840 47815 34920 47825
rect 35160 47815 35240 47825
rect 35480 47815 35560 47825
rect 35800 47815 35880 47825
rect 36120 47815 36200 47825
rect 36440 47815 36520 47825
rect 36760 47815 36840 47825
rect 37080 47815 37160 47825
rect 37400 47815 37480 47825
rect 37720 47815 37800 47825
rect 40180 47815 40260 47825
rect 40500 47815 40580 47825
rect 40820 47815 40900 47825
rect 41140 47815 41220 47825
rect 42560 47815 42640 47825
rect 42880 47815 42960 47825
rect 43200 47815 43280 47825
rect 43520 47815 43600 47825
rect 146400 47815 146480 47825
rect 146720 47815 146800 47825
rect 147040 47815 147120 47825
rect 147360 47815 147440 47825
rect 148780 47815 148860 47825
rect 149100 47815 149180 47825
rect 149420 47815 149500 47825
rect 149740 47815 149820 47825
rect 152200 47815 152280 47825
rect 152520 47815 152600 47825
rect 152840 47815 152920 47825
rect 153160 47815 153240 47825
rect 153480 47815 153560 47825
rect 153800 47815 153880 47825
rect 154120 47815 154200 47825
rect 154440 47815 154520 47825
rect 154760 47815 154840 47825
rect 155080 47815 155160 47825
rect 155400 47815 155480 47825
rect 155720 47815 155800 47825
rect 156040 47815 156120 47825
rect 156360 47815 156440 47825
rect 156680 47815 156760 47825
rect 157000 47815 157080 47825
rect 157320 47815 157400 47825
rect 157640 47815 157720 47825
rect 157960 47815 158040 47825
rect 158280 47815 158360 47825
rect 158600 47815 158680 47825
rect 158920 47815 159000 47825
rect 159240 47815 159320 47825
rect 159560 47815 159640 47825
rect 30440 47735 30450 47815
rect 30760 47735 30770 47815
rect 31080 47735 31090 47815
rect 31400 47735 31410 47815
rect 31720 47735 31730 47815
rect 32040 47735 32050 47815
rect 32360 47735 32370 47815
rect 32680 47735 32690 47815
rect 33000 47735 33010 47815
rect 33320 47735 33330 47815
rect 33640 47735 33650 47815
rect 33960 47735 33970 47815
rect 34280 47735 34290 47815
rect 34600 47735 34610 47815
rect 34920 47735 34930 47815
rect 35240 47735 35250 47815
rect 35560 47735 35570 47815
rect 35880 47735 35890 47815
rect 36200 47735 36210 47815
rect 36520 47735 36530 47815
rect 36840 47735 36850 47815
rect 37160 47735 37170 47815
rect 37480 47735 37490 47815
rect 37800 47735 37810 47815
rect 40260 47735 40270 47815
rect 40580 47735 40590 47815
rect 40900 47735 40910 47815
rect 41220 47735 41230 47815
rect 42640 47735 42650 47815
rect 42960 47735 42970 47815
rect 43280 47735 43290 47815
rect 43600 47735 43610 47815
rect 146480 47735 146490 47815
rect 146800 47735 146810 47815
rect 147120 47735 147130 47815
rect 147440 47735 147450 47815
rect 148860 47735 148870 47815
rect 149180 47735 149190 47815
rect 149500 47735 149510 47815
rect 149820 47735 149830 47815
rect 152280 47735 152290 47815
rect 152600 47735 152610 47815
rect 152920 47735 152930 47815
rect 153240 47735 153250 47815
rect 153560 47735 153570 47815
rect 153880 47735 153890 47815
rect 154200 47735 154210 47815
rect 154520 47735 154530 47815
rect 154840 47735 154850 47815
rect 155160 47735 155170 47815
rect 155480 47735 155490 47815
rect 155800 47735 155810 47815
rect 156120 47735 156130 47815
rect 156440 47735 156450 47815
rect 156760 47735 156770 47815
rect 157080 47735 157090 47815
rect 157400 47735 157410 47815
rect 157720 47735 157730 47815
rect 158040 47735 158050 47815
rect 158360 47735 158370 47815
rect 158680 47735 158690 47815
rect 159000 47735 159010 47815
rect 159320 47735 159330 47815
rect 159640 47735 159650 47815
rect 163670 47775 163680 47855
rect 163990 47775 164000 47855
rect 164310 47775 164320 47855
rect 164630 47775 164640 47855
rect 164950 47775 164960 47855
rect 165270 47775 165280 47855
rect 165590 47775 165600 47855
rect 165910 47775 165920 47855
rect 166230 47775 166240 47855
rect 166550 47775 166560 47855
rect 166870 47775 166880 47855
rect 167190 47775 167200 47855
rect 167510 47775 167520 47855
rect 167830 47775 167840 47855
rect 168150 47775 168160 47855
rect 168470 47775 168480 47855
rect 168790 47775 168800 47855
rect 169110 47775 169120 47855
rect 169430 47775 169440 47855
rect 169750 47775 169760 47855
rect 170070 47775 170080 47855
rect 170390 47775 170400 47855
rect 170710 47775 170720 47855
rect 171030 47775 171040 47855
rect 19130 47695 19210 47705
rect 19450 47695 19530 47705
rect 19770 47695 19850 47705
rect 20090 47695 20170 47705
rect 20410 47695 20490 47705
rect 20730 47695 20810 47705
rect 21050 47695 21130 47705
rect 21370 47695 21450 47705
rect 21690 47695 21770 47705
rect 22010 47695 22090 47705
rect 22330 47695 22410 47705
rect 22650 47695 22730 47705
rect 22970 47695 23050 47705
rect 23290 47695 23370 47705
rect 23610 47695 23690 47705
rect 23930 47695 24010 47705
rect 24250 47695 24330 47705
rect 24570 47695 24650 47705
rect 24890 47695 24970 47705
rect 25210 47695 25290 47705
rect 25530 47695 25610 47705
rect 25850 47695 25930 47705
rect 26170 47695 26250 47705
rect 163750 47695 163830 47705
rect 164070 47695 164150 47705
rect 164390 47695 164470 47705
rect 164710 47695 164790 47705
rect 165030 47695 165110 47705
rect 165350 47695 165430 47705
rect 165670 47695 165750 47705
rect 165990 47695 166070 47705
rect 166310 47695 166390 47705
rect 166630 47695 166710 47705
rect 166950 47695 167030 47705
rect 167270 47695 167350 47705
rect 167590 47695 167670 47705
rect 167910 47695 167990 47705
rect 168230 47695 168310 47705
rect 168550 47695 168630 47705
rect 168870 47695 168950 47705
rect 169190 47695 169270 47705
rect 169510 47695 169590 47705
rect 169830 47695 169910 47705
rect 170150 47695 170230 47705
rect 170470 47695 170550 47705
rect 170790 47695 170870 47705
rect 19210 47615 19220 47695
rect 19530 47615 19540 47695
rect 19850 47615 19860 47695
rect 20170 47615 20180 47695
rect 20490 47615 20500 47695
rect 20810 47615 20820 47695
rect 21130 47615 21140 47695
rect 21450 47615 21460 47695
rect 21770 47615 21780 47695
rect 22090 47615 22100 47695
rect 22410 47615 22420 47695
rect 22730 47615 22740 47695
rect 23050 47615 23060 47695
rect 23370 47615 23380 47695
rect 23690 47615 23700 47695
rect 24010 47615 24020 47695
rect 24330 47615 24340 47695
rect 24650 47615 24660 47695
rect 24970 47615 24980 47695
rect 25290 47615 25300 47695
rect 25610 47615 25620 47695
rect 25930 47615 25940 47695
rect 26250 47615 26260 47695
rect 30520 47655 30600 47665
rect 30840 47655 30920 47665
rect 31160 47655 31240 47665
rect 31480 47655 31560 47665
rect 31800 47655 31880 47665
rect 32120 47655 32200 47665
rect 32440 47655 32520 47665
rect 32760 47655 32840 47665
rect 33080 47655 33160 47665
rect 33400 47655 33480 47665
rect 33720 47655 33800 47665
rect 34040 47655 34120 47665
rect 34360 47655 34440 47665
rect 34680 47655 34760 47665
rect 35000 47655 35080 47665
rect 35320 47655 35400 47665
rect 35640 47655 35720 47665
rect 35960 47655 36040 47665
rect 36280 47655 36360 47665
rect 36600 47655 36680 47665
rect 36920 47655 37000 47665
rect 37240 47655 37320 47665
rect 37560 47655 37640 47665
rect 40340 47655 40420 47665
rect 40660 47655 40740 47665
rect 40980 47655 41060 47665
rect 42720 47655 42800 47665
rect 43040 47655 43120 47665
rect 43360 47655 43440 47665
rect 146560 47655 146640 47665
rect 146880 47655 146960 47665
rect 147200 47655 147280 47665
rect 148940 47655 149020 47665
rect 149260 47655 149340 47665
rect 149580 47655 149660 47665
rect 152360 47655 152440 47665
rect 152680 47655 152760 47665
rect 153000 47655 153080 47665
rect 153320 47655 153400 47665
rect 153640 47655 153720 47665
rect 153960 47655 154040 47665
rect 154280 47655 154360 47665
rect 154600 47655 154680 47665
rect 154920 47655 155000 47665
rect 155240 47655 155320 47665
rect 155560 47655 155640 47665
rect 155880 47655 155960 47665
rect 156200 47655 156280 47665
rect 156520 47655 156600 47665
rect 156840 47655 156920 47665
rect 157160 47655 157240 47665
rect 157480 47655 157560 47665
rect 157800 47655 157880 47665
rect 158120 47655 158200 47665
rect 158440 47655 158520 47665
rect 158760 47655 158840 47665
rect 159080 47655 159160 47665
rect 159400 47655 159480 47665
rect 30600 47575 30610 47655
rect 30920 47575 30930 47655
rect 31240 47575 31250 47655
rect 31560 47575 31570 47655
rect 31880 47575 31890 47655
rect 32200 47575 32210 47655
rect 32520 47575 32530 47655
rect 32840 47575 32850 47655
rect 33160 47575 33170 47655
rect 33480 47575 33490 47655
rect 33800 47575 33810 47655
rect 34120 47575 34130 47655
rect 34440 47575 34450 47655
rect 34760 47575 34770 47655
rect 35080 47575 35090 47655
rect 35400 47575 35410 47655
rect 35720 47575 35730 47655
rect 36040 47575 36050 47655
rect 36360 47575 36370 47655
rect 36680 47575 36690 47655
rect 37000 47575 37010 47655
rect 37320 47575 37330 47655
rect 37640 47575 37650 47655
rect 40420 47575 40430 47655
rect 40740 47575 40750 47655
rect 41060 47575 41070 47655
rect 42800 47575 42810 47655
rect 43120 47575 43130 47655
rect 43440 47575 43450 47655
rect 146640 47575 146650 47655
rect 146960 47575 146970 47655
rect 147280 47575 147290 47655
rect 149020 47575 149030 47655
rect 149340 47575 149350 47655
rect 149660 47575 149670 47655
rect 152440 47575 152450 47655
rect 152760 47575 152770 47655
rect 153080 47575 153090 47655
rect 153400 47575 153410 47655
rect 153720 47575 153730 47655
rect 154040 47575 154050 47655
rect 154360 47575 154370 47655
rect 154680 47575 154690 47655
rect 155000 47575 155010 47655
rect 155320 47575 155330 47655
rect 155640 47575 155650 47655
rect 155960 47575 155970 47655
rect 156280 47575 156290 47655
rect 156600 47575 156610 47655
rect 156920 47575 156930 47655
rect 157240 47575 157250 47655
rect 157560 47575 157570 47655
rect 157880 47575 157890 47655
rect 158200 47575 158210 47655
rect 158520 47575 158530 47655
rect 158840 47575 158850 47655
rect 159160 47575 159170 47655
rect 159480 47575 159490 47655
rect 163830 47615 163840 47695
rect 164150 47615 164160 47695
rect 164470 47615 164480 47695
rect 164790 47615 164800 47695
rect 165110 47615 165120 47695
rect 165430 47615 165440 47695
rect 165750 47615 165760 47695
rect 166070 47615 166080 47695
rect 166390 47615 166400 47695
rect 166710 47615 166720 47695
rect 167030 47615 167040 47695
rect 167350 47615 167360 47695
rect 167670 47615 167680 47695
rect 167990 47615 168000 47695
rect 168310 47615 168320 47695
rect 168630 47615 168640 47695
rect 168950 47615 168960 47695
rect 169270 47615 169280 47695
rect 169590 47615 169600 47695
rect 169910 47615 169920 47695
rect 170230 47615 170240 47695
rect 170550 47615 170560 47695
rect 170870 47615 170880 47695
rect 18970 47535 19050 47545
rect 19290 47535 19370 47545
rect 19610 47535 19690 47545
rect 19930 47535 20010 47545
rect 20250 47535 20330 47545
rect 20570 47535 20650 47545
rect 20890 47535 20970 47545
rect 21210 47535 21290 47545
rect 21530 47535 21610 47545
rect 21850 47535 21930 47545
rect 22170 47535 22250 47545
rect 22490 47535 22570 47545
rect 22810 47535 22890 47545
rect 23130 47535 23210 47545
rect 23450 47535 23530 47545
rect 23770 47535 23850 47545
rect 24090 47535 24170 47545
rect 24410 47535 24490 47545
rect 24730 47535 24810 47545
rect 25050 47535 25130 47545
rect 25370 47535 25450 47545
rect 25690 47535 25770 47545
rect 26010 47535 26090 47545
rect 26330 47535 26410 47545
rect 163590 47535 163670 47545
rect 163910 47535 163990 47545
rect 164230 47535 164310 47545
rect 164550 47535 164630 47545
rect 164870 47535 164950 47545
rect 165190 47535 165270 47545
rect 165510 47535 165590 47545
rect 165830 47535 165910 47545
rect 166150 47535 166230 47545
rect 166470 47535 166550 47545
rect 166790 47535 166870 47545
rect 167110 47535 167190 47545
rect 167430 47535 167510 47545
rect 167750 47535 167830 47545
rect 168070 47535 168150 47545
rect 168390 47535 168470 47545
rect 168710 47535 168790 47545
rect 169030 47535 169110 47545
rect 169350 47535 169430 47545
rect 169670 47535 169750 47545
rect 169990 47535 170070 47545
rect 170310 47535 170390 47545
rect 170630 47535 170710 47545
rect 170950 47535 171030 47545
rect 19050 47455 19060 47535
rect 19370 47455 19380 47535
rect 19690 47455 19700 47535
rect 20010 47455 20020 47535
rect 20330 47455 20340 47535
rect 20650 47455 20660 47535
rect 20970 47455 20980 47535
rect 21290 47455 21300 47535
rect 21610 47455 21620 47535
rect 21930 47455 21940 47535
rect 22250 47455 22260 47535
rect 22570 47455 22580 47535
rect 22890 47455 22900 47535
rect 23210 47455 23220 47535
rect 23530 47455 23540 47535
rect 23850 47455 23860 47535
rect 24170 47455 24180 47535
rect 24490 47455 24500 47535
rect 24810 47455 24820 47535
rect 25130 47455 25140 47535
rect 25450 47455 25460 47535
rect 25770 47455 25780 47535
rect 26090 47455 26100 47535
rect 26410 47455 26420 47535
rect 30360 47495 30440 47505
rect 30680 47495 30760 47505
rect 31000 47495 31080 47505
rect 31320 47495 31400 47505
rect 31640 47495 31720 47505
rect 31960 47495 32040 47505
rect 32280 47495 32360 47505
rect 32600 47495 32680 47505
rect 32920 47495 33000 47505
rect 33240 47495 33320 47505
rect 33560 47495 33640 47505
rect 33880 47495 33960 47505
rect 34200 47495 34280 47505
rect 34520 47495 34600 47505
rect 34840 47495 34920 47505
rect 35160 47495 35240 47505
rect 35480 47495 35560 47505
rect 35800 47495 35880 47505
rect 36120 47495 36200 47505
rect 36440 47495 36520 47505
rect 36760 47495 36840 47505
rect 37080 47495 37160 47505
rect 37400 47495 37480 47505
rect 37720 47495 37800 47505
rect 40180 47495 40260 47505
rect 40500 47495 40580 47505
rect 40820 47495 40900 47505
rect 41140 47495 41220 47505
rect 42560 47495 42640 47505
rect 42880 47495 42960 47505
rect 43200 47495 43280 47505
rect 43520 47495 43600 47505
rect 146400 47495 146480 47505
rect 146720 47495 146800 47505
rect 147040 47495 147120 47505
rect 147360 47495 147440 47505
rect 148780 47495 148860 47505
rect 149100 47495 149180 47505
rect 149420 47495 149500 47505
rect 149740 47495 149820 47505
rect 152200 47495 152280 47505
rect 152520 47495 152600 47505
rect 152840 47495 152920 47505
rect 153160 47495 153240 47505
rect 153480 47495 153560 47505
rect 153800 47495 153880 47505
rect 154120 47495 154200 47505
rect 154440 47495 154520 47505
rect 154760 47495 154840 47505
rect 155080 47495 155160 47505
rect 155400 47495 155480 47505
rect 155720 47495 155800 47505
rect 156040 47495 156120 47505
rect 156360 47495 156440 47505
rect 156680 47495 156760 47505
rect 157000 47495 157080 47505
rect 157320 47495 157400 47505
rect 157640 47495 157720 47505
rect 157960 47495 158040 47505
rect 158280 47495 158360 47505
rect 158600 47495 158680 47505
rect 158920 47495 159000 47505
rect 159240 47495 159320 47505
rect 159560 47495 159640 47505
rect 30440 47415 30450 47495
rect 30760 47415 30770 47495
rect 31080 47415 31090 47495
rect 31400 47415 31410 47495
rect 31720 47415 31730 47495
rect 32040 47415 32050 47495
rect 32360 47415 32370 47495
rect 32680 47415 32690 47495
rect 33000 47415 33010 47495
rect 33320 47415 33330 47495
rect 33640 47415 33650 47495
rect 33960 47415 33970 47495
rect 34280 47415 34290 47495
rect 34600 47415 34610 47495
rect 34920 47415 34930 47495
rect 35240 47415 35250 47495
rect 35560 47415 35570 47495
rect 35880 47415 35890 47495
rect 36200 47415 36210 47495
rect 36520 47415 36530 47495
rect 36840 47415 36850 47495
rect 37160 47415 37170 47495
rect 37480 47415 37490 47495
rect 37800 47415 37810 47495
rect 40260 47415 40270 47495
rect 40580 47415 40590 47495
rect 40900 47415 40910 47495
rect 41220 47415 41230 47495
rect 42640 47415 42650 47495
rect 42960 47415 42970 47495
rect 43280 47415 43290 47495
rect 43600 47415 43610 47495
rect 146480 47415 146490 47495
rect 146800 47415 146810 47495
rect 147120 47415 147130 47495
rect 147440 47415 147450 47495
rect 148860 47415 148870 47495
rect 149180 47415 149190 47495
rect 149500 47415 149510 47495
rect 149820 47415 149830 47495
rect 152280 47415 152290 47495
rect 152600 47415 152610 47495
rect 152920 47415 152930 47495
rect 153240 47415 153250 47495
rect 153560 47415 153570 47495
rect 153880 47415 153890 47495
rect 154200 47415 154210 47495
rect 154520 47415 154530 47495
rect 154840 47415 154850 47495
rect 155160 47415 155170 47495
rect 155480 47415 155490 47495
rect 155800 47415 155810 47495
rect 156120 47415 156130 47495
rect 156440 47415 156450 47495
rect 156760 47415 156770 47495
rect 157080 47415 157090 47495
rect 157400 47415 157410 47495
rect 157720 47415 157730 47495
rect 158040 47415 158050 47495
rect 158360 47415 158370 47495
rect 158680 47415 158690 47495
rect 159000 47415 159010 47495
rect 159320 47415 159330 47495
rect 159640 47415 159650 47495
rect 163670 47455 163680 47535
rect 163990 47455 164000 47535
rect 164310 47455 164320 47535
rect 164630 47455 164640 47535
rect 164950 47455 164960 47535
rect 165270 47455 165280 47535
rect 165590 47455 165600 47535
rect 165910 47455 165920 47535
rect 166230 47455 166240 47535
rect 166550 47455 166560 47535
rect 166870 47455 166880 47535
rect 167190 47455 167200 47535
rect 167510 47455 167520 47535
rect 167830 47455 167840 47535
rect 168150 47455 168160 47535
rect 168470 47455 168480 47535
rect 168790 47455 168800 47535
rect 169110 47455 169120 47535
rect 169430 47455 169440 47535
rect 169750 47455 169760 47535
rect 170070 47455 170080 47535
rect 170390 47455 170400 47535
rect 170710 47455 170720 47535
rect 171030 47455 171040 47535
rect 19130 47375 19210 47385
rect 19450 47375 19530 47385
rect 19770 47375 19850 47385
rect 20090 47375 20170 47385
rect 20410 47375 20490 47385
rect 20730 47375 20810 47385
rect 21050 47375 21130 47385
rect 21370 47375 21450 47385
rect 21690 47375 21770 47385
rect 22010 47375 22090 47385
rect 22330 47375 22410 47385
rect 22650 47375 22730 47385
rect 22970 47375 23050 47385
rect 23290 47375 23370 47385
rect 23610 47375 23690 47385
rect 23930 47375 24010 47385
rect 24250 47375 24330 47385
rect 24570 47375 24650 47385
rect 24890 47375 24970 47385
rect 25210 47375 25290 47385
rect 25530 47375 25610 47385
rect 25850 47375 25930 47385
rect 26170 47375 26250 47385
rect 163750 47375 163830 47385
rect 164070 47375 164150 47385
rect 164390 47375 164470 47385
rect 164710 47375 164790 47385
rect 165030 47375 165110 47385
rect 165350 47375 165430 47385
rect 165670 47375 165750 47385
rect 165990 47375 166070 47385
rect 166310 47375 166390 47385
rect 166630 47375 166710 47385
rect 166950 47375 167030 47385
rect 167270 47375 167350 47385
rect 167590 47375 167670 47385
rect 167910 47375 167990 47385
rect 168230 47375 168310 47385
rect 168550 47375 168630 47385
rect 168870 47375 168950 47385
rect 169190 47375 169270 47385
rect 169510 47375 169590 47385
rect 169830 47375 169910 47385
rect 170150 47375 170230 47385
rect 170470 47375 170550 47385
rect 170790 47375 170870 47385
rect 19210 47295 19220 47375
rect 19530 47295 19540 47375
rect 19850 47295 19860 47375
rect 20170 47295 20180 47375
rect 20490 47295 20500 47375
rect 20810 47295 20820 47375
rect 21130 47295 21140 47375
rect 21450 47295 21460 47375
rect 21770 47295 21780 47375
rect 22090 47295 22100 47375
rect 22410 47295 22420 47375
rect 22730 47295 22740 47375
rect 23050 47295 23060 47375
rect 23370 47295 23380 47375
rect 23690 47295 23700 47375
rect 24010 47295 24020 47375
rect 24330 47295 24340 47375
rect 24650 47295 24660 47375
rect 24970 47295 24980 47375
rect 25290 47295 25300 47375
rect 25610 47295 25620 47375
rect 25930 47295 25940 47375
rect 26250 47295 26260 47375
rect 30520 47335 30600 47345
rect 30840 47335 30920 47345
rect 31160 47335 31240 47345
rect 31480 47335 31560 47345
rect 31800 47335 31880 47345
rect 32120 47335 32200 47345
rect 32440 47335 32520 47345
rect 32760 47335 32840 47345
rect 33080 47335 33160 47345
rect 33400 47335 33480 47345
rect 33720 47335 33800 47345
rect 34040 47335 34120 47345
rect 34360 47335 34440 47345
rect 34680 47335 34760 47345
rect 35000 47335 35080 47345
rect 35320 47335 35400 47345
rect 35640 47335 35720 47345
rect 35960 47335 36040 47345
rect 36280 47335 36360 47345
rect 36600 47335 36680 47345
rect 36920 47335 37000 47345
rect 37240 47335 37320 47345
rect 37560 47335 37640 47345
rect 40340 47335 40420 47345
rect 40660 47335 40740 47345
rect 40980 47335 41060 47345
rect 42720 47335 42800 47345
rect 43040 47335 43120 47345
rect 43360 47335 43440 47345
rect 146560 47335 146640 47345
rect 146880 47335 146960 47345
rect 147200 47335 147280 47345
rect 148940 47335 149020 47345
rect 149260 47335 149340 47345
rect 149580 47335 149660 47345
rect 152360 47335 152440 47345
rect 152680 47335 152760 47345
rect 153000 47335 153080 47345
rect 153320 47335 153400 47345
rect 153640 47335 153720 47345
rect 153960 47335 154040 47345
rect 154280 47335 154360 47345
rect 154600 47335 154680 47345
rect 154920 47335 155000 47345
rect 155240 47335 155320 47345
rect 155560 47335 155640 47345
rect 155880 47335 155960 47345
rect 156200 47335 156280 47345
rect 156520 47335 156600 47345
rect 156840 47335 156920 47345
rect 157160 47335 157240 47345
rect 157480 47335 157560 47345
rect 157800 47335 157880 47345
rect 158120 47335 158200 47345
rect 158440 47335 158520 47345
rect 158760 47335 158840 47345
rect 159080 47335 159160 47345
rect 159400 47335 159480 47345
rect 30600 47255 30610 47335
rect 30920 47255 30930 47335
rect 31240 47255 31250 47335
rect 31560 47255 31570 47335
rect 31880 47255 31890 47335
rect 32200 47255 32210 47335
rect 32520 47255 32530 47335
rect 32840 47255 32850 47335
rect 33160 47255 33170 47335
rect 33480 47255 33490 47335
rect 33800 47255 33810 47335
rect 34120 47255 34130 47335
rect 34440 47255 34450 47335
rect 34760 47255 34770 47335
rect 35080 47255 35090 47335
rect 35400 47255 35410 47335
rect 35720 47255 35730 47335
rect 36040 47255 36050 47335
rect 36360 47255 36370 47335
rect 36680 47255 36690 47335
rect 37000 47255 37010 47335
rect 37320 47255 37330 47335
rect 37640 47255 37650 47335
rect 40420 47255 40430 47335
rect 40740 47255 40750 47335
rect 41060 47255 41070 47335
rect 42800 47255 42810 47335
rect 43120 47255 43130 47335
rect 43440 47255 43450 47335
rect 146640 47255 146650 47335
rect 146960 47255 146970 47335
rect 147280 47255 147290 47335
rect 149020 47255 149030 47335
rect 149340 47255 149350 47335
rect 149660 47255 149670 47335
rect 152440 47255 152450 47335
rect 152760 47255 152770 47335
rect 153080 47255 153090 47335
rect 153400 47255 153410 47335
rect 153720 47255 153730 47335
rect 154040 47255 154050 47335
rect 154360 47255 154370 47335
rect 154680 47255 154690 47335
rect 155000 47255 155010 47335
rect 155320 47255 155330 47335
rect 155640 47255 155650 47335
rect 155960 47255 155970 47335
rect 156280 47255 156290 47335
rect 156600 47255 156610 47335
rect 156920 47255 156930 47335
rect 157240 47255 157250 47335
rect 157560 47255 157570 47335
rect 157880 47255 157890 47335
rect 158200 47255 158210 47335
rect 158520 47255 158530 47335
rect 158840 47255 158850 47335
rect 159160 47255 159170 47335
rect 159480 47255 159490 47335
rect 163830 47295 163840 47375
rect 164150 47295 164160 47375
rect 164470 47295 164480 47375
rect 164790 47295 164800 47375
rect 165110 47295 165120 47375
rect 165430 47295 165440 47375
rect 165750 47295 165760 47375
rect 166070 47295 166080 47375
rect 166390 47295 166400 47375
rect 166710 47295 166720 47375
rect 167030 47295 167040 47375
rect 167350 47295 167360 47375
rect 167670 47295 167680 47375
rect 167990 47295 168000 47375
rect 168310 47295 168320 47375
rect 168630 47295 168640 47375
rect 168950 47295 168960 47375
rect 169270 47295 169280 47375
rect 169590 47295 169600 47375
rect 169910 47295 169920 47375
rect 170230 47295 170240 47375
rect 170550 47295 170560 47375
rect 170870 47295 170880 47375
rect 18970 47215 19050 47225
rect 19290 47215 19370 47225
rect 19610 47215 19690 47225
rect 19930 47215 20010 47225
rect 20250 47215 20330 47225
rect 20570 47215 20650 47225
rect 20890 47215 20970 47225
rect 21210 47215 21290 47225
rect 21530 47215 21610 47225
rect 21850 47215 21930 47225
rect 22170 47215 22250 47225
rect 22490 47215 22570 47225
rect 22810 47215 22890 47225
rect 23130 47215 23210 47225
rect 23450 47215 23530 47225
rect 23770 47215 23850 47225
rect 24090 47215 24170 47225
rect 24410 47215 24490 47225
rect 24730 47215 24810 47225
rect 25050 47215 25130 47225
rect 25370 47215 25450 47225
rect 25690 47215 25770 47225
rect 26010 47215 26090 47225
rect 26330 47215 26410 47225
rect 163590 47215 163670 47225
rect 163910 47215 163990 47225
rect 164230 47215 164310 47225
rect 164550 47215 164630 47225
rect 164870 47215 164950 47225
rect 165190 47215 165270 47225
rect 165510 47215 165590 47225
rect 165830 47215 165910 47225
rect 166150 47215 166230 47225
rect 166470 47215 166550 47225
rect 166790 47215 166870 47225
rect 167110 47215 167190 47225
rect 167430 47215 167510 47225
rect 167750 47215 167830 47225
rect 168070 47215 168150 47225
rect 168390 47215 168470 47225
rect 168710 47215 168790 47225
rect 169030 47215 169110 47225
rect 169350 47215 169430 47225
rect 169670 47215 169750 47225
rect 169990 47215 170070 47225
rect 170310 47215 170390 47225
rect 170630 47215 170710 47225
rect 170950 47215 171030 47225
rect 19050 47135 19060 47215
rect 19370 47135 19380 47215
rect 19690 47135 19700 47215
rect 20010 47135 20020 47215
rect 20330 47135 20340 47215
rect 20650 47135 20660 47215
rect 20970 47135 20980 47215
rect 21290 47135 21300 47215
rect 21610 47135 21620 47215
rect 21930 47135 21940 47215
rect 22250 47135 22260 47215
rect 22570 47135 22580 47215
rect 22890 47135 22900 47215
rect 23210 47135 23220 47215
rect 23530 47135 23540 47215
rect 23850 47135 23860 47215
rect 24170 47135 24180 47215
rect 24490 47135 24500 47215
rect 24810 47135 24820 47215
rect 25130 47135 25140 47215
rect 25450 47135 25460 47215
rect 25770 47135 25780 47215
rect 26090 47135 26100 47215
rect 26410 47135 26420 47215
rect 30360 47175 30440 47185
rect 30680 47175 30760 47185
rect 31000 47175 31080 47185
rect 31320 47175 31400 47185
rect 31640 47175 31720 47185
rect 31960 47175 32040 47185
rect 32280 47175 32360 47185
rect 32600 47175 32680 47185
rect 32920 47175 33000 47185
rect 33240 47175 33320 47185
rect 33560 47175 33640 47185
rect 33880 47175 33960 47185
rect 34200 47175 34280 47185
rect 34520 47175 34600 47185
rect 34840 47175 34920 47185
rect 35160 47175 35240 47185
rect 35480 47175 35560 47185
rect 35800 47175 35880 47185
rect 36120 47175 36200 47185
rect 36440 47175 36520 47185
rect 36760 47175 36840 47185
rect 37080 47175 37160 47185
rect 37400 47175 37480 47185
rect 37720 47175 37800 47185
rect 40180 47175 40260 47185
rect 40500 47175 40580 47185
rect 40820 47175 40900 47185
rect 41140 47175 41220 47185
rect 42560 47175 42640 47185
rect 42880 47175 42960 47185
rect 43200 47175 43280 47185
rect 43520 47175 43600 47185
rect 146400 47175 146480 47185
rect 146720 47175 146800 47185
rect 147040 47175 147120 47185
rect 147360 47175 147440 47185
rect 148780 47175 148860 47185
rect 149100 47175 149180 47185
rect 149420 47175 149500 47185
rect 149740 47175 149820 47185
rect 152200 47175 152280 47185
rect 152520 47175 152600 47185
rect 152840 47175 152920 47185
rect 153160 47175 153240 47185
rect 153480 47175 153560 47185
rect 153800 47175 153880 47185
rect 154120 47175 154200 47185
rect 154440 47175 154520 47185
rect 154760 47175 154840 47185
rect 155080 47175 155160 47185
rect 155400 47175 155480 47185
rect 155720 47175 155800 47185
rect 156040 47175 156120 47185
rect 156360 47175 156440 47185
rect 156680 47175 156760 47185
rect 157000 47175 157080 47185
rect 157320 47175 157400 47185
rect 157640 47175 157720 47185
rect 157960 47175 158040 47185
rect 158280 47175 158360 47185
rect 158600 47175 158680 47185
rect 158920 47175 159000 47185
rect 159240 47175 159320 47185
rect 159560 47175 159640 47185
rect 30440 47095 30450 47175
rect 30760 47095 30770 47175
rect 31080 47095 31090 47175
rect 31400 47095 31410 47175
rect 31720 47095 31730 47175
rect 32040 47095 32050 47175
rect 32360 47095 32370 47175
rect 32680 47095 32690 47175
rect 33000 47095 33010 47175
rect 33320 47095 33330 47175
rect 33640 47095 33650 47175
rect 33960 47095 33970 47175
rect 34280 47095 34290 47175
rect 34600 47095 34610 47175
rect 34920 47095 34930 47175
rect 35240 47095 35250 47175
rect 35560 47095 35570 47175
rect 35880 47095 35890 47175
rect 36200 47095 36210 47175
rect 36520 47095 36530 47175
rect 36840 47095 36850 47175
rect 37160 47095 37170 47175
rect 37480 47095 37490 47175
rect 37800 47095 37810 47175
rect 40260 47095 40270 47175
rect 40580 47095 40590 47175
rect 40900 47095 40910 47175
rect 41220 47095 41230 47175
rect 42640 47095 42650 47175
rect 42960 47095 42970 47175
rect 43280 47095 43290 47175
rect 43600 47095 43610 47175
rect 146480 47095 146490 47175
rect 146800 47095 146810 47175
rect 147120 47095 147130 47175
rect 147440 47095 147450 47175
rect 148860 47095 148870 47175
rect 149180 47095 149190 47175
rect 149500 47095 149510 47175
rect 149820 47095 149830 47175
rect 152280 47095 152290 47175
rect 152600 47095 152610 47175
rect 152920 47095 152930 47175
rect 153240 47095 153250 47175
rect 153560 47095 153570 47175
rect 153880 47095 153890 47175
rect 154200 47095 154210 47175
rect 154520 47095 154530 47175
rect 154840 47095 154850 47175
rect 155160 47095 155170 47175
rect 155480 47095 155490 47175
rect 155800 47095 155810 47175
rect 156120 47095 156130 47175
rect 156440 47095 156450 47175
rect 156760 47095 156770 47175
rect 157080 47095 157090 47175
rect 157400 47095 157410 47175
rect 157720 47095 157730 47175
rect 158040 47095 158050 47175
rect 158360 47095 158370 47175
rect 158680 47095 158690 47175
rect 159000 47095 159010 47175
rect 159320 47095 159330 47175
rect 159640 47095 159650 47175
rect 163670 47135 163680 47215
rect 163990 47135 164000 47215
rect 164310 47135 164320 47215
rect 164630 47135 164640 47215
rect 164950 47135 164960 47215
rect 165270 47135 165280 47215
rect 165590 47135 165600 47215
rect 165910 47135 165920 47215
rect 166230 47135 166240 47215
rect 166550 47135 166560 47215
rect 166870 47135 166880 47215
rect 167190 47135 167200 47215
rect 167510 47135 167520 47215
rect 167830 47135 167840 47215
rect 168150 47135 168160 47215
rect 168470 47135 168480 47215
rect 168790 47135 168800 47215
rect 169110 47135 169120 47215
rect 169430 47135 169440 47215
rect 169750 47135 169760 47215
rect 170070 47135 170080 47215
rect 170390 47135 170400 47215
rect 170710 47135 170720 47215
rect 171030 47135 171040 47215
rect 19130 47055 19210 47065
rect 19450 47055 19530 47065
rect 19770 47055 19850 47065
rect 20090 47055 20170 47065
rect 20410 47055 20490 47065
rect 20730 47055 20810 47065
rect 21050 47055 21130 47065
rect 21370 47055 21450 47065
rect 21690 47055 21770 47065
rect 22010 47055 22090 47065
rect 22330 47055 22410 47065
rect 22650 47055 22730 47065
rect 22970 47055 23050 47065
rect 23290 47055 23370 47065
rect 23610 47055 23690 47065
rect 23930 47055 24010 47065
rect 24250 47055 24330 47065
rect 24570 47055 24650 47065
rect 24890 47055 24970 47065
rect 25210 47055 25290 47065
rect 25530 47055 25610 47065
rect 25850 47055 25930 47065
rect 26170 47055 26250 47065
rect 163750 47055 163830 47065
rect 164070 47055 164150 47065
rect 164390 47055 164470 47065
rect 164710 47055 164790 47065
rect 165030 47055 165110 47065
rect 165350 47055 165430 47065
rect 165670 47055 165750 47065
rect 165990 47055 166070 47065
rect 166310 47055 166390 47065
rect 166630 47055 166710 47065
rect 166950 47055 167030 47065
rect 167270 47055 167350 47065
rect 167590 47055 167670 47065
rect 167910 47055 167990 47065
rect 168230 47055 168310 47065
rect 168550 47055 168630 47065
rect 168870 47055 168950 47065
rect 169190 47055 169270 47065
rect 169510 47055 169590 47065
rect 169830 47055 169910 47065
rect 170150 47055 170230 47065
rect 170470 47055 170550 47065
rect 170790 47055 170870 47065
rect 19210 46975 19220 47055
rect 19530 46975 19540 47055
rect 19850 46975 19860 47055
rect 20170 46975 20180 47055
rect 20490 46975 20500 47055
rect 20810 46975 20820 47055
rect 21130 46975 21140 47055
rect 21450 46975 21460 47055
rect 21770 46975 21780 47055
rect 22090 46975 22100 47055
rect 22410 46975 22420 47055
rect 22730 46975 22740 47055
rect 23050 46975 23060 47055
rect 23370 46975 23380 47055
rect 23690 46975 23700 47055
rect 24010 46975 24020 47055
rect 24330 46975 24340 47055
rect 24650 46975 24660 47055
rect 24970 46975 24980 47055
rect 25290 46975 25300 47055
rect 25610 46975 25620 47055
rect 25930 46975 25940 47055
rect 26250 46975 26260 47055
rect 30520 47015 30600 47025
rect 30840 47015 30920 47025
rect 31160 47015 31240 47025
rect 31480 47015 31560 47025
rect 31800 47015 31880 47025
rect 32120 47015 32200 47025
rect 32440 47015 32520 47025
rect 32760 47015 32840 47025
rect 33080 47015 33160 47025
rect 33400 47015 33480 47025
rect 33720 47015 33800 47025
rect 34040 47015 34120 47025
rect 34360 47015 34440 47025
rect 34680 47015 34760 47025
rect 35000 47015 35080 47025
rect 35320 47015 35400 47025
rect 35640 47015 35720 47025
rect 35960 47015 36040 47025
rect 36280 47015 36360 47025
rect 36600 47015 36680 47025
rect 36920 47015 37000 47025
rect 37240 47015 37320 47025
rect 37560 47015 37640 47025
rect 40340 47015 40420 47025
rect 40660 47015 40740 47025
rect 40980 47015 41060 47025
rect 42720 47015 42800 47025
rect 43040 47015 43120 47025
rect 43360 47015 43440 47025
rect 146560 47015 146640 47025
rect 146880 47015 146960 47025
rect 147200 47015 147280 47025
rect 148940 47015 149020 47025
rect 149260 47015 149340 47025
rect 149580 47015 149660 47025
rect 152360 47015 152440 47025
rect 152680 47015 152760 47025
rect 153000 47015 153080 47025
rect 153320 47015 153400 47025
rect 153640 47015 153720 47025
rect 153960 47015 154040 47025
rect 154280 47015 154360 47025
rect 154600 47015 154680 47025
rect 154920 47015 155000 47025
rect 155240 47015 155320 47025
rect 155560 47015 155640 47025
rect 155880 47015 155960 47025
rect 156200 47015 156280 47025
rect 156520 47015 156600 47025
rect 156840 47015 156920 47025
rect 157160 47015 157240 47025
rect 157480 47015 157560 47025
rect 157800 47015 157880 47025
rect 158120 47015 158200 47025
rect 158440 47015 158520 47025
rect 158760 47015 158840 47025
rect 159080 47015 159160 47025
rect 159400 47015 159480 47025
rect 30600 46935 30610 47015
rect 30920 46935 30930 47015
rect 31240 46935 31250 47015
rect 31560 46935 31570 47015
rect 31880 46935 31890 47015
rect 32200 46935 32210 47015
rect 32520 46935 32530 47015
rect 32840 46935 32850 47015
rect 33160 46935 33170 47015
rect 33480 46935 33490 47015
rect 33800 46935 33810 47015
rect 34120 46935 34130 47015
rect 34440 46935 34450 47015
rect 34760 46935 34770 47015
rect 35080 46935 35090 47015
rect 35400 46935 35410 47015
rect 35720 46935 35730 47015
rect 36040 46935 36050 47015
rect 36360 46935 36370 47015
rect 36680 46935 36690 47015
rect 37000 46935 37010 47015
rect 37320 46935 37330 47015
rect 37640 46935 37650 47015
rect 40420 46935 40430 47015
rect 40740 46935 40750 47015
rect 41060 46935 41070 47015
rect 42800 46935 42810 47015
rect 43120 46935 43130 47015
rect 43440 46935 43450 47015
rect 146640 46935 146650 47015
rect 146960 46935 146970 47015
rect 147280 46935 147290 47015
rect 149020 46935 149030 47015
rect 149340 46935 149350 47015
rect 149660 46935 149670 47015
rect 152440 46935 152450 47015
rect 152760 46935 152770 47015
rect 153080 46935 153090 47015
rect 153400 46935 153410 47015
rect 153720 46935 153730 47015
rect 154040 46935 154050 47015
rect 154360 46935 154370 47015
rect 154680 46935 154690 47015
rect 155000 46935 155010 47015
rect 155320 46935 155330 47015
rect 155640 46935 155650 47015
rect 155960 46935 155970 47015
rect 156280 46935 156290 47015
rect 156600 46935 156610 47015
rect 156920 46935 156930 47015
rect 157240 46935 157250 47015
rect 157560 46935 157570 47015
rect 157880 46935 157890 47015
rect 158200 46935 158210 47015
rect 158520 46935 158530 47015
rect 158840 46935 158850 47015
rect 159160 46935 159170 47015
rect 159480 46935 159490 47015
rect 163830 46975 163840 47055
rect 164150 46975 164160 47055
rect 164470 46975 164480 47055
rect 164790 46975 164800 47055
rect 165110 46975 165120 47055
rect 165430 46975 165440 47055
rect 165750 46975 165760 47055
rect 166070 46975 166080 47055
rect 166390 46975 166400 47055
rect 166710 46975 166720 47055
rect 167030 46975 167040 47055
rect 167350 46975 167360 47055
rect 167670 46975 167680 47055
rect 167990 46975 168000 47055
rect 168310 46975 168320 47055
rect 168630 46975 168640 47055
rect 168950 46975 168960 47055
rect 169270 46975 169280 47055
rect 169590 46975 169600 47055
rect 169910 46975 169920 47055
rect 170230 46975 170240 47055
rect 170550 46975 170560 47055
rect 170870 46975 170880 47055
rect 18970 46895 19050 46905
rect 19290 46895 19370 46905
rect 19610 46895 19690 46905
rect 19930 46895 20010 46905
rect 20250 46895 20330 46905
rect 20570 46895 20650 46905
rect 20890 46895 20970 46905
rect 21210 46895 21290 46905
rect 21530 46895 21610 46905
rect 21850 46895 21930 46905
rect 22170 46895 22250 46905
rect 22490 46895 22570 46905
rect 22810 46895 22890 46905
rect 23130 46895 23210 46905
rect 23450 46895 23530 46905
rect 23770 46895 23850 46905
rect 24090 46895 24170 46905
rect 24410 46895 24490 46905
rect 24730 46895 24810 46905
rect 25050 46895 25130 46905
rect 25370 46895 25450 46905
rect 25690 46895 25770 46905
rect 26010 46895 26090 46905
rect 26330 46895 26410 46905
rect 163590 46895 163670 46905
rect 163910 46895 163990 46905
rect 164230 46895 164310 46905
rect 164550 46895 164630 46905
rect 164870 46895 164950 46905
rect 165190 46895 165270 46905
rect 165510 46895 165590 46905
rect 165830 46895 165910 46905
rect 166150 46895 166230 46905
rect 166470 46895 166550 46905
rect 166790 46895 166870 46905
rect 167110 46895 167190 46905
rect 167430 46895 167510 46905
rect 167750 46895 167830 46905
rect 168070 46895 168150 46905
rect 168390 46895 168470 46905
rect 168710 46895 168790 46905
rect 169030 46895 169110 46905
rect 169350 46895 169430 46905
rect 169670 46895 169750 46905
rect 169990 46895 170070 46905
rect 170310 46895 170390 46905
rect 170630 46895 170710 46905
rect 170950 46895 171030 46905
rect 19050 46815 19060 46895
rect 19370 46815 19380 46895
rect 19690 46815 19700 46895
rect 20010 46815 20020 46895
rect 20330 46815 20340 46895
rect 20650 46815 20660 46895
rect 20970 46815 20980 46895
rect 21290 46815 21300 46895
rect 21610 46815 21620 46895
rect 21930 46815 21940 46895
rect 22250 46815 22260 46895
rect 22570 46815 22580 46895
rect 22890 46815 22900 46895
rect 23210 46815 23220 46895
rect 23530 46815 23540 46895
rect 23850 46815 23860 46895
rect 24170 46815 24180 46895
rect 24490 46815 24500 46895
rect 24810 46815 24820 46895
rect 25130 46815 25140 46895
rect 25450 46815 25460 46895
rect 25770 46815 25780 46895
rect 26090 46815 26100 46895
rect 26410 46815 26420 46895
rect 30360 46855 30440 46865
rect 30680 46855 30760 46865
rect 31000 46855 31080 46865
rect 31320 46855 31400 46865
rect 31640 46855 31720 46865
rect 31960 46855 32040 46865
rect 32280 46855 32360 46865
rect 32600 46855 32680 46865
rect 32920 46855 33000 46865
rect 33240 46855 33320 46865
rect 33560 46855 33640 46865
rect 33880 46855 33960 46865
rect 34200 46855 34280 46865
rect 34520 46855 34600 46865
rect 34840 46855 34920 46865
rect 35160 46855 35240 46865
rect 35480 46855 35560 46865
rect 35800 46855 35880 46865
rect 36120 46855 36200 46865
rect 36440 46855 36520 46865
rect 36760 46855 36840 46865
rect 37080 46855 37160 46865
rect 37400 46855 37480 46865
rect 37720 46855 37800 46865
rect 40180 46855 40260 46865
rect 40500 46855 40580 46865
rect 40820 46855 40900 46865
rect 41140 46855 41220 46865
rect 42560 46855 42640 46865
rect 42880 46855 42960 46865
rect 43200 46855 43280 46865
rect 43520 46855 43600 46865
rect 146400 46855 146480 46865
rect 146720 46855 146800 46865
rect 147040 46855 147120 46865
rect 147360 46855 147440 46865
rect 148780 46855 148860 46865
rect 149100 46855 149180 46865
rect 149420 46855 149500 46865
rect 149740 46855 149820 46865
rect 152200 46855 152280 46865
rect 152520 46855 152600 46865
rect 152840 46855 152920 46865
rect 153160 46855 153240 46865
rect 153480 46855 153560 46865
rect 153800 46855 153880 46865
rect 154120 46855 154200 46865
rect 154440 46855 154520 46865
rect 154760 46855 154840 46865
rect 155080 46855 155160 46865
rect 155400 46855 155480 46865
rect 155720 46855 155800 46865
rect 156040 46855 156120 46865
rect 156360 46855 156440 46865
rect 156680 46855 156760 46865
rect 157000 46855 157080 46865
rect 157320 46855 157400 46865
rect 157640 46855 157720 46865
rect 157960 46855 158040 46865
rect 158280 46855 158360 46865
rect 158600 46855 158680 46865
rect 158920 46855 159000 46865
rect 159240 46855 159320 46865
rect 159560 46855 159640 46865
rect 30440 46775 30450 46855
rect 30760 46775 30770 46855
rect 31080 46775 31090 46855
rect 31400 46775 31410 46855
rect 31720 46775 31730 46855
rect 32040 46775 32050 46855
rect 32360 46775 32370 46855
rect 32680 46775 32690 46855
rect 33000 46775 33010 46855
rect 33320 46775 33330 46855
rect 33640 46775 33650 46855
rect 33960 46775 33970 46855
rect 34280 46775 34290 46855
rect 34600 46775 34610 46855
rect 34920 46775 34930 46855
rect 35240 46775 35250 46855
rect 35560 46775 35570 46855
rect 35880 46775 35890 46855
rect 36200 46775 36210 46855
rect 36520 46775 36530 46855
rect 36840 46775 36850 46855
rect 37160 46775 37170 46855
rect 37480 46775 37490 46855
rect 37800 46775 37810 46855
rect 40260 46775 40270 46855
rect 40580 46775 40590 46855
rect 40900 46775 40910 46855
rect 41220 46775 41230 46855
rect 42640 46775 42650 46855
rect 42960 46775 42970 46855
rect 43280 46775 43290 46855
rect 43600 46775 43610 46855
rect 19130 46735 19210 46745
rect 19450 46735 19530 46745
rect 19770 46735 19850 46745
rect 20090 46735 20170 46745
rect 20410 46735 20490 46745
rect 20730 46735 20810 46745
rect 21050 46735 21130 46745
rect 21370 46735 21450 46745
rect 21690 46735 21770 46745
rect 22010 46735 22090 46745
rect 22330 46735 22410 46745
rect 22650 46735 22730 46745
rect 22970 46735 23050 46745
rect 23290 46735 23370 46745
rect 23610 46735 23690 46745
rect 23930 46735 24010 46745
rect 24250 46735 24330 46745
rect 24570 46735 24650 46745
rect 24890 46735 24970 46745
rect 25210 46735 25290 46745
rect 25530 46735 25610 46745
rect 25850 46735 25930 46745
rect 26170 46735 26250 46745
rect 19210 46655 19220 46735
rect 19530 46655 19540 46735
rect 19850 46655 19860 46735
rect 20170 46655 20180 46735
rect 20490 46655 20500 46735
rect 20810 46655 20820 46735
rect 21130 46655 21140 46735
rect 21450 46655 21460 46735
rect 21770 46655 21780 46735
rect 22090 46655 22100 46735
rect 22410 46655 22420 46735
rect 22730 46655 22740 46735
rect 23050 46655 23060 46735
rect 23370 46655 23380 46735
rect 23690 46655 23700 46735
rect 24010 46655 24020 46735
rect 24330 46655 24340 46735
rect 24650 46655 24660 46735
rect 24970 46655 24980 46735
rect 25290 46655 25300 46735
rect 25610 46655 25620 46735
rect 25930 46655 25940 46735
rect 26250 46655 26260 46735
rect 30520 46695 30600 46705
rect 30840 46695 30920 46705
rect 31160 46695 31240 46705
rect 31480 46695 31560 46705
rect 31800 46695 31880 46705
rect 32120 46695 32200 46705
rect 32440 46695 32520 46705
rect 32760 46695 32840 46705
rect 33080 46695 33160 46705
rect 33400 46695 33480 46705
rect 33720 46695 33800 46705
rect 34040 46695 34120 46705
rect 34360 46695 34440 46705
rect 34680 46695 34760 46705
rect 35000 46695 35080 46705
rect 35320 46695 35400 46705
rect 35640 46695 35720 46705
rect 35960 46695 36040 46705
rect 36280 46695 36360 46705
rect 36600 46695 36680 46705
rect 36920 46695 37000 46705
rect 37240 46695 37320 46705
rect 37560 46695 37640 46705
rect 40340 46695 40420 46705
rect 40660 46695 40740 46705
rect 40980 46695 41060 46705
rect 42720 46695 42800 46705
rect 43040 46695 43120 46705
rect 43360 46695 43440 46705
rect 30600 46615 30610 46695
rect 30920 46615 30930 46695
rect 31240 46615 31250 46695
rect 31560 46615 31570 46695
rect 31880 46615 31890 46695
rect 32200 46615 32210 46695
rect 32520 46615 32530 46695
rect 32840 46615 32850 46695
rect 33160 46615 33170 46695
rect 33480 46615 33490 46695
rect 33800 46615 33810 46695
rect 34120 46615 34130 46695
rect 34440 46615 34450 46695
rect 34760 46615 34770 46695
rect 35080 46615 35090 46695
rect 35400 46615 35410 46695
rect 35720 46615 35730 46695
rect 36040 46615 36050 46695
rect 36360 46615 36370 46695
rect 36680 46615 36690 46695
rect 37000 46615 37010 46695
rect 37320 46615 37330 46695
rect 37640 46615 37650 46695
rect 40420 46615 40430 46695
rect 40740 46615 40750 46695
rect 41060 46615 41070 46695
rect 42800 46615 42810 46695
rect 43120 46615 43130 46695
rect 43440 46615 43450 46695
rect 46660 46660 48000 46840
rect 60000 46660 72000 46840
rect 84000 46800 120000 46840
rect 84000 46660 142200 46800
rect 146480 46775 146490 46855
rect 146800 46775 146810 46855
rect 147120 46775 147130 46855
rect 147440 46775 147450 46855
rect 148860 46775 148870 46855
rect 149180 46775 149190 46855
rect 149500 46775 149510 46855
rect 149820 46775 149830 46855
rect 152280 46775 152290 46855
rect 152600 46775 152610 46855
rect 152920 46775 152930 46855
rect 153240 46775 153250 46855
rect 153560 46775 153570 46855
rect 153880 46775 153890 46855
rect 154200 46775 154210 46855
rect 154520 46775 154530 46855
rect 154840 46775 154850 46855
rect 155160 46775 155170 46855
rect 155480 46775 155490 46855
rect 155800 46775 155810 46855
rect 156120 46775 156130 46855
rect 156440 46775 156450 46855
rect 156760 46775 156770 46855
rect 157080 46775 157090 46855
rect 157400 46775 157410 46855
rect 157720 46775 157730 46855
rect 158040 46775 158050 46855
rect 158360 46775 158370 46855
rect 158680 46775 158690 46855
rect 159000 46775 159010 46855
rect 159320 46775 159330 46855
rect 159640 46775 159650 46855
rect 163670 46815 163680 46895
rect 163990 46815 164000 46895
rect 164310 46815 164320 46895
rect 164630 46815 164640 46895
rect 164950 46815 164960 46895
rect 165270 46815 165280 46895
rect 165590 46815 165600 46895
rect 165910 46815 165920 46895
rect 166230 46815 166240 46895
rect 166550 46815 166560 46895
rect 166870 46815 166880 46895
rect 167190 46815 167200 46895
rect 167510 46815 167520 46895
rect 167830 46815 167840 46895
rect 168150 46815 168160 46895
rect 168470 46815 168480 46895
rect 168790 46815 168800 46895
rect 169110 46815 169120 46895
rect 169430 46815 169440 46895
rect 169750 46815 169760 46895
rect 170070 46815 170080 46895
rect 170390 46815 170400 46895
rect 170710 46815 170720 46895
rect 171030 46815 171040 46895
rect 163750 46735 163830 46745
rect 164070 46735 164150 46745
rect 164390 46735 164470 46745
rect 164710 46735 164790 46745
rect 165030 46735 165110 46745
rect 165350 46735 165430 46745
rect 165670 46735 165750 46745
rect 165990 46735 166070 46745
rect 166310 46735 166390 46745
rect 166630 46735 166710 46745
rect 166950 46735 167030 46745
rect 167270 46735 167350 46745
rect 167590 46735 167670 46745
rect 167910 46735 167990 46745
rect 168230 46735 168310 46745
rect 168550 46735 168630 46745
rect 168870 46735 168950 46745
rect 169190 46735 169270 46745
rect 169510 46735 169590 46745
rect 169830 46735 169910 46745
rect 170150 46735 170230 46745
rect 170470 46735 170550 46745
rect 170790 46735 170870 46745
rect 146560 46695 146640 46705
rect 146880 46695 146960 46705
rect 147200 46695 147280 46705
rect 148940 46695 149020 46705
rect 149260 46695 149340 46705
rect 149580 46695 149660 46705
rect 152360 46695 152440 46705
rect 152680 46695 152760 46705
rect 153000 46695 153080 46705
rect 153320 46695 153400 46705
rect 153640 46695 153720 46705
rect 153960 46695 154040 46705
rect 154280 46695 154360 46705
rect 154600 46695 154680 46705
rect 154920 46695 155000 46705
rect 155240 46695 155320 46705
rect 155560 46695 155640 46705
rect 155880 46695 155960 46705
rect 156200 46695 156280 46705
rect 156520 46695 156600 46705
rect 156840 46695 156920 46705
rect 157160 46695 157240 46705
rect 157480 46695 157560 46705
rect 157800 46695 157880 46705
rect 158120 46695 158200 46705
rect 158440 46695 158520 46705
rect 158760 46695 158840 46705
rect 159080 46695 159160 46705
rect 159400 46695 159480 46705
rect 98310 46630 100140 46640
rect 146640 46615 146650 46695
rect 146960 46615 146970 46695
rect 147280 46615 147290 46695
rect 149020 46615 149030 46695
rect 149340 46615 149350 46695
rect 149660 46615 149670 46695
rect 152440 46615 152450 46695
rect 152760 46615 152770 46695
rect 153080 46615 153090 46695
rect 153400 46615 153410 46695
rect 153720 46615 153730 46695
rect 154040 46615 154050 46695
rect 154360 46615 154370 46695
rect 154680 46615 154690 46695
rect 155000 46615 155010 46695
rect 155320 46615 155330 46695
rect 155640 46615 155650 46695
rect 155960 46615 155970 46695
rect 156280 46615 156290 46695
rect 156600 46615 156610 46695
rect 156920 46615 156930 46695
rect 157240 46615 157250 46695
rect 157560 46615 157570 46695
rect 157880 46615 157890 46695
rect 158200 46615 158210 46695
rect 158520 46615 158530 46695
rect 158840 46615 158850 46695
rect 159160 46615 159170 46695
rect 159480 46615 159490 46695
rect 163830 46655 163840 46735
rect 164150 46655 164160 46735
rect 164470 46655 164480 46735
rect 164790 46655 164800 46735
rect 165110 46655 165120 46735
rect 165430 46655 165440 46735
rect 165750 46655 165760 46735
rect 166070 46655 166080 46735
rect 166390 46655 166400 46735
rect 166710 46655 166720 46735
rect 167030 46655 167040 46735
rect 167350 46655 167360 46735
rect 167670 46655 167680 46735
rect 167990 46655 168000 46735
rect 168310 46655 168320 46735
rect 168630 46655 168640 46735
rect 168950 46655 168960 46735
rect 169270 46655 169280 46735
rect 169590 46655 169600 46735
rect 169910 46655 169920 46735
rect 170230 46655 170240 46735
rect 170550 46655 170560 46735
rect 170870 46655 170880 46735
rect 18970 46575 19050 46585
rect 19290 46575 19370 46585
rect 19610 46575 19690 46585
rect 19930 46575 20010 46585
rect 20250 46575 20330 46585
rect 20570 46575 20650 46585
rect 20890 46575 20970 46585
rect 21210 46575 21290 46585
rect 21530 46575 21610 46585
rect 21850 46575 21930 46585
rect 22170 46575 22250 46585
rect 22490 46575 22570 46585
rect 22810 46575 22890 46585
rect 23130 46575 23210 46585
rect 23450 46575 23530 46585
rect 23770 46575 23850 46585
rect 24090 46575 24170 46585
rect 24410 46575 24490 46585
rect 24730 46575 24810 46585
rect 25050 46575 25130 46585
rect 25370 46575 25450 46585
rect 25690 46575 25770 46585
rect 26010 46575 26090 46585
rect 26330 46575 26410 46585
rect 163590 46575 163670 46585
rect 163910 46575 163990 46585
rect 164230 46575 164310 46585
rect 164550 46575 164630 46585
rect 164870 46575 164950 46585
rect 165190 46575 165270 46585
rect 165510 46575 165590 46585
rect 165830 46575 165910 46585
rect 166150 46575 166230 46585
rect 166470 46575 166550 46585
rect 166790 46575 166870 46585
rect 167110 46575 167190 46585
rect 167430 46575 167510 46585
rect 167750 46575 167830 46585
rect 168070 46575 168150 46585
rect 168390 46575 168470 46585
rect 168710 46575 168790 46585
rect 169030 46575 169110 46585
rect 169350 46575 169430 46585
rect 169670 46575 169750 46585
rect 169990 46575 170070 46585
rect 170310 46575 170390 46585
rect 170630 46575 170710 46585
rect 170950 46575 171030 46585
rect 19050 46495 19060 46575
rect 19370 46495 19380 46575
rect 19690 46495 19700 46575
rect 20010 46495 20020 46575
rect 20330 46495 20340 46575
rect 20650 46495 20660 46575
rect 20970 46495 20980 46575
rect 21290 46495 21300 46575
rect 21610 46495 21620 46575
rect 21930 46495 21940 46575
rect 22250 46495 22260 46575
rect 22570 46495 22580 46575
rect 22890 46495 22900 46575
rect 23210 46495 23220 46575
rect 23530 46495 23540 46575
rect 23850 46495 23860 46575
rect 24170 46495 24180 46575
rect 24490 46495 24500 46575
rect 24810 46495 24820 46575
rect 25130 46495 25140 46575
rect 25450 46495 25460 46575
rect 25770 46495 25780 46575
rect 26090 46495 26100 46575
rect 26410 46495 26420 46575
rect 30360 46535 30440 46545
rect 30680 46535 30760 46545
rect 31000 46535 31080 46545
rect 31320 46535 31400 46545
rect 31640 46535 31720 46545
rect 31960 46535 32040 46545
rect 32280 46535 32360 46545
rect 32600 46535 32680 46545
rect 32920 46535 33000 46545
rect 33240 46535 33320 46545
rect 33560 46535 33640 46545
rect 33880 46535 33960 46545
rect 34200 46535 34280 46545
rect 34520 46535 34600 46545
rect 34840 46535 34920 46545
rect 35160 46535 35240 46545
rect 35480 46535 35560 46545
rect 35800 46535 35880 46545
rect 36120 46535 36200 46545
rect 36440 46535 36520 46545
rect 36760 46535 36840 46545
rect 37080 46535 37160 46545
rect 37400 46535 37480 46545
rect 37720 46535 37800 46545
rect 40180 46535 40260 46545
rect 40500 46535 40580 46545
rect 40820 46535 40900 46545
rect 41140 46535 41220 46545
rect 42560 46535 42640 46545
rect 42880 46535 42960 46545
rect 43200 46535 43280 46545
rect 43520 46535 43600 46545
rect 146400 46535 146480 46545
rect 146720 46535 146800 46545
rect 147040 46535 147120 46545
rect 147360 46535 147440 46545
rect 148780 46535 148860 46545
rect 149100 46535 149180 46545
rect 149420 46535 149500 46545
rect 149740 46535 149820 46545
rect 152200 46535 152280 46545
rect 152520 46535 152600 46545
rect 152840 46535 152920 46545
rect 153160 46535 153240 46545
rect 153480 46535 153560 46545
rect 153800 46535 153880 46545
rect 154120 46535 154200 46545
rect 154440 46535 154520 46545
rect 154760 46535 154840 46545
rect 155080 46535 155160 46545
rect 155400 46535 155480 46545
rect 155720 46535 155800 46545
rect 156040 46535 156120 46545
rect 156360 46535 156440 46545
rect 156680 46535 156760 46545
rect 157000 46535 157080 46545
rect 157320 46535 157400 46545
rect 157640 46535 157720 46545
rect 157960 46535 158040 46545
rect 158280 46535 158360 46545
rect 158600 46535 158680 46545
rect 158920 46535 159000 46545
rect 159240 46535 159320 46545
rect 159560 46535 159640 46545
rect 30440 46455 30450 46535
rect 30760 46455 30770 46535
rect 31080 46455 31090 46535
rect 31400 46455 31410 46535
rect 31720 46455 31730 46535
rect 32040 46455 32050 46535
rect 32360 46455 32370 46535
rect 32680 46455 32690 46535
rect 33000 46455 33010 46535
rect 33320 46455 33330 46535
rect 33640 46455 33650 46535
rect 33960 46455 33970 46535
rect 34280 46455 34290 46535
rect 34600 46455 34610 46535
rect 34920 46455 34930 46535
rect 35240 46455 35250 46535
rect 35560 46455 35570 46535
rect 35880 46455 35890 46535
rect 36200 46455 36210 46535
rect 36520 46455 36530 46535
rect 36840 46455 36850 46535
rect 37160 46455 37170 46535
rect 37480 46455 37490 46535
rect 37800 46455 37810 46535
rect 40260 46455 40270 46535
rect 40580 46455 40590 46535
rect 40900 46455 40910 46535
rect 41220 46455 41230 46535
rect 42640 46455 42650 46535
rect 42960 46455 42970 46535
rect 43280 46455 43290 46535
rect 43600 46455 43610 46535
rect 146480 46455 146490 46535
rect 146800 46455 146810 46535
rect 147120 46455 147130 46535
rect 147440 46455 147450 46535
rect 148860 46455 148870 46535
rect 149180 46455 149190 46535
rect 149500 46455 149510 46535
rect 149820 46455 149830 46535
rect 152280 46455 152290 46535
rect 152600 46455 152610 46535
rect 152920 46455 152930 46535
rect 153240 46455 153250 46535
rect 153560 46455 153570 46535
rect 153880 46455 153890 46535
rect 154200 46455 154210 46535
rect 154520 46455 154530 46535
rect 154840 46455 154850 46535
rect 155160 46455 155170 46535
rect 155480 46455 155490 46535
rect 155800 46455 155810 46535
rect 156120 46455 156130 46535
rect 156440 46455 156450 46535
rect 156760 46455 156770 46535
rect 157080 46455 157090 46535
rect 157400 46455 157410 46535
rect 157720 46455 157730 46535
rect 158040 46455 158050 46535
rect 158360 46455 158370 46535
rect 158680 46455 158690 46535
rect 159000 46455 159010 46535
rect 159320 46455 159330 46535
rect 159640 46455 159650 46535
rect 163670 46495 163680 46575
rect 163990 46495 164000 46575
rect 164310 46495 164320 46575
rect 164630 46495 164640 46575
rect 164950 46495 164960 46575
rect 165270 46495 165280 46575
rect 165590 46495 165600 46575
rect 165910 46495 165920 46575
rect 166230 46495 166240 46575
rect 166550 46495 166560 46575
rect 166870 46495 166880 46575
rect 167190 46495 167200 46575
rect 167510 46495 167520 46575
rect 167830 46495 167840 46575
rect 168150 46495 168160 46575
rect 168470 46495 168480 46575
rect 168790 46495 168800 46575
rect 169110 46495 169120 46575
rect 169430 46495 169440 46575
rect 169750 46495 169760 46575
rect 170070 46495 170080 46575
rect 170390 46495 170400 46575
rect 170710 46495 170720 46575
rect 171030 46495 171040 46575
rect 19130 46415 19210 46425
rect 19450 46415 19530 46425
rect 19770 46415 19850 46425
rect 20090 46415 20170 46425
rect 20410 46415 20490 46425
rect 20730 46415 20810 46425
rect 21050 46415 21130 46425
rect 21370 46415 21450 46425
rect 21690 46415 21770 46425
rect 22010 46415 22090 46425
rect 22330 46415 22410 46425
rect 22650 46415 22730 46425
rect 22970 46415 23050 46425
rect 23290 46415 23370 46425
rect 23610 46415 23690 46425
rect 23930 46415 24010 46425
rect 24250 46415 24330 46425
rect 24570 46415 24650 46425
rect 24890 46415 24970 46425
rect 25210 46415 25290 46425
rect 25530 46415 25610 46425
rect 25850 46415 25930 46425
rect 26170 46415 26250 46425
rect 163750 46415 163830 46425
rect 164070 46415 164150 46425
rect 164390 46415 164470 46425
rect 164710 46415 164790 46425
rect 165030 46415 165110 46425
rect 165350 46415 165430 46425
rect 165670 46415 165750 46425
rect 165990 46415 166070 46425
rect 166310 46415 166390 46425
rect 166630 46415 166710 46425
rect 166950 46415 167030 46425
rect 167270 46415 167350 46425
rect 167590 46415 167670 46425
rect 167910 46415 167990 46425
rect 168230 46415 168310 46425
rect 168550 46415 168630 46425
rect 168870 46415 168950 46425
rect 169190 46415 169270 46425
rect 169510 46415 169590 46425
rect 169830 46415 169910 46425
rect 170150 46415 170230 46425
rect 170470 46415 170550 46425
rect 170790 46415 170870 46425
rect 19210 46335 19220 46415
rect 19530 46335 19540 46415
rect 19850 46335 19860 46415
rect 20170 46335 20180 46415
rect 20490 46335 20500 46415
rect 20810 46335 20820 46415
rect 21130 46335 21140 46415
rect 21450 46335 21460 46415
rect 21770 46335 21780 46415
rect 22090 46335 22100 46415
rect 22410 46335 22420 46415
rect 22730 46335 22740 46415
rect 23050 46335 23060 46415
rect 23370 46335 23380 46415
rect 23690 46335 23700 46415
rect 24010 46335 24020 46415
rect 24330 46335 24340 46415
rect 24650 46335 24660 46415
rect 24970 46335 24980 46415
rect 25290 46335 25300 46415
rect 25610 46335 25620 46415
rect 25930 46335 25940 46415
rect 26250 46335 26260 46415
rect 30520 46375 30600 46385
rect 30840 46375 30920 46385
rect 31160 46375 31240 46385
rect 31480 46375 31560 46385
rect 31800 46375 31880 46385
rect 32120 46375 32200 46385
rect 32440 46375 32520 46385
rect 32760 46375 32840 46385
rect 33080 46375 33160 46385
rect 33400 46375 33480 46385
rect 33720 46375 33800 46385
rect 34040 46375 34120 46385
rect 34360 46375 34440 46385
rect 34680 46375 34760 46385
rect 35000 46375 35080 46385
rect 35320 46375 35400 46385
rect 35640 46375 35720 46385
rect 35960 46375 36040 46385
rect 36280 46375 36360 46385
rect 36600 46375 36680 46385
rect 36920 46375 37000 46385
rect 37240 46375 37320 46385
rect 37560 46375 37640 46385
rect 40340 46375 40420 46385
rect 40660 46375 40740 46385
rect 40980 46375 41060 46385
rect 42720 46375 42800 46385
rect 43040 46375 43120 46385
rect 43360 46375 43440 46385
rect 146560 46375 146640 46385
rect 146880 46375 146960 46385
rect 147200 46375 147280 46385
rect 148940 46375 149020 46385
rect 149260 46375 149340 46385
rect 149580 46375 149660 46385
rect 152360 46375 152440 46385
rect 152680 46375 152760 46385
rect 153000 46375 153080 46385
rect 153320 46375 153400 46385
rect 153640 46375 153720 46385
rect 153960 46375 154040 46385
rect 154280 46375 154360 46385
rect 154600 46375 154680 46385
rect 154920 46375 155000 46385
rect 155240 46375 155320 46385
rect 155560 46375 155640 46385
rect 155880 46375 155960 46385
rect 156200 46375 156280 46385
rect 156520 46375 156600 46385
rect 156840 46375 156920 46385
rect 157160 46375 157240 46385
rect 157480 46375 157560 46385
rect 157800 46375 157880 46385
rect 158120 46375 158200 46385
rect 158440 46375 158520 46385
rect 158760 46375 158840 46385
rect 159080 46375 159160 46385
rect 159400 46375 159480 46385
rect 30600 46295 30610 46375
rect 30920 46295 30930 46375
rect 31240 46295 31250 46375
rect 31560 46295 31570 46375
rect 31880 46295 31890 46375
rect 32200 46295 32210 46375
rect 32520 46295 32530 46375
rect 32840 46295 32850 46375
rect 33160 46295 33170 46375
rect 33480 46295 33490 46375
rect 33800 46295 33810 46375
rect 34120 46295 34130 46375
rect 34440 46295 34450 46375
rect 34760 46295 34770 46375
rect 35080 46295 35090 46375
rect 35400 46295 35410 46375
rect 35720 46295 35730 46375
rect 36040 46295 36050 46375
rect 36360 46295 36370 46375
rect 36680 46295 36690 46375
rect 37000 46295 37010 46375
rect 37320 46295 37330 46375
rect 37640 46295 37650 46375
rect 40420 46295 40430 46375
rect 40740 46295 40750 46375
rect 41060 46295 41070 46375
rect 42800 46295 42810 46375
rect 43120 46295 43130 46375
rect 43440 46295 43450 46375
rect 146640 46295 146650 46375
rect 146960 46295 146970 46375
rect 147280 46295 147290 46375
rect 149020 46295 149030 46375
rect 149340 46295 149350 46375
rect 149660 46295 149670 46375
rect 152440 46295 152450 46375
rect 152760 46295 152770 46375
rect 153080 46295 153090 46375
rect 153400 46295 153410 46375
rect 153720 46295 153730 46375
rect 154040 46295 154050 46375
rect 154360 46295 154370 46375
rect 154680 46295 154690 46375
rect 155000 46295 155010 46375
rect 155320 46295 155330 46375
rect 155640 46295 155650 46375
rect 155960 46295 155970 46375
rect 156280 46295 156290 46375
rect 156600 46295 156610 46375
rect 156920 46295 156930 46375
rect 157240 46295 157250 46375
rect 157560 46295 157570 46375
rect 157880 46295 157890 46375
rect 158200 46295 158210 46375
rect 158520 46295 158530 46375
rect 158840 46295 158850 46375
rect 159160 46295 159170 46375
rect 159480 46295 159490 46375
rect 163830 46335 163840 46415
rect 164150 46335 164160 46415
rect 164470 46335 164480 46415
rect 164790 46335 164800 46415
rect 165110 46335 165120 46415
rect 165430 46335 165440 46415
rect 165750 46335 165760 46415
rect 166070 46335 166080 46415
rect 166390 46335 166400 46415
rect 166710 46335 166720 46415
rect 167030 46335 167040 46415
rect 167350 46335 167360 46415
rect 167670 46335 167680 46415
rect 167990 46335 168000 46415
rect 168310 46335 168320 46415
rect 168630 46335 168640 46415
rect 168950 46335 168960 46415
rect 169270 46335 169280 46415
rect 169590 46335 169600 46415
rect 169910 46335 169920 46415
rect 170230 46335 170240 46415
rect 170550 46335 170560 46415
rect 170870 46335 170880 46415
rect 18970 46255 19050 46265
rect 19290 46255 19370 46265
rect 19610 46255 19690 46265
rect 19930 46255 20010 46265
rect 20250 46255 20330 46265
rect 20570 46255 20650 46265
rect 20890 46255 20970 46265
rect 21210 46255 21290 46265
rect 21530 46255 21610 46265
rect 21850 46255 21930 46265
rect 22170 46255 22250 46265
rect 22490 46255 22570 46265
rect 22810 46255 22890 46265
rect 23130 46255 23210 46265
rect 23450 46255 23530 46265
rect 23770 46255 23850 46265
rect 24090 46255 24170 46265
rect 24410 46255 24490 46265
rect 24730 46255 24810 46265
rect 25050 46255 25130 46265
rect 25370 46255 25450 46265
rect 25690 46255 25770 46265
rect 26010 46255 26090 46265
rect 26330 46255 26410 46265
rect 163590 46255 163670 46265
rect 163910 46255 163990 46265
rect 164230 46255 164310 46265
rect 164550 46255 164630 46265
rect 164870 46255 164950 46265
rect 165190 46255 165270 46265
rect 165510 46255 165590 46265
rect 165830 46255 165910 46265
rect 166150 46255 166230 46265
rect 166470 46255 166550 46265
rect 166790 46255 166870 46265
rect 167110 46255 167190 46265
rect 167430 46255 167510 46265
rect 167750 46255 167830 46265
rect 168070 46255 168150 46265
rect 168390 46255 168470 46265
rect 168710 46255 168790 46265
rect 169030 46255 169110 46265
rect 169350 46255 169430 46265
rect 169670 46255 169750 46265
rect 169990 46255 170070 46265
rect 170310 46255 170390 46265
rect 170630 46255 170710 46265
rect 170950 46255 171030 46265
rect 19050 46175 19060 46255
rect 19370 46175 19380 46255
rect 19690 46175 19700 46255
rect 20010 46175 20020 46255
rect 20330 46175 20340 46255
rect 20650 46175 20660 46255
rect 20970 46175 20980 46255
rect 21290 46175 21300 46255
rect 21610 46175 21620 46255
rect 21930 46175 21940 46255
rect 22250 46175 22260 46255
rect 22570 46175 22580 46255
rect 22890 46175 22900 46255
rect 23210 46175 23220 46255
rect 23530 46175 23540 46255
rect 23850 46175 23860 46255
rect 24170 46175 24180 46255
rect 24490 46175 24500 46255
rect 24810 46175 24820 46255
rect 25130 46175 25140 46255
rect 25450 46175 25460 46255
rect 25770 46175 25780 46255
rect 26090 46175 26100 46255
rect 26410 46175 26420 46255
rect 30360 46215 30440 46225
rect 30680 46215 30760 46225
rect 31000 46215 31080 46225
rect 31320 46215 31400 46225
rect 31640 46215 31720 46225
rect 31960 46215 32040 46225
rect 32280 46215 32360 46225
rect 32600 46215 32680 46225
rect 32920 46215 33000 46225
rect 33240 46215 33320 46225
rect 33560 46215 33640 46225
rect 33880 46215 33960 46225
rect 34200 46215 34280 46225
rect 34520 46215 34600 46225
rect 34840 46215 34920 46225
rect 35160 46215 35240 46225
rect 35480 46215 35560 46225
rect 35800 46215 35880 46225
rect 36120 46215 36200 46225
rect 36440 46215 36520 46225
rect 36760 46215 36840 46225
rect 37080 46215 37160 46225
rect 37400 46215 37480 46225
rect 37720 46215 37800 46225
rect 40180 46215 40260 46225
rect 40500 46215 40580 46225
rect 40820 46215 40900 46225
rect 41140 46215 41220 46225
rect 42560 46215 42640 46225
rect 42880 46215 42960 46225
rect 43200 46215 43280 46225
rect 43520 46215 43600 46225
rect 146400 46215 146480 46225
rect 146720 46215 146800 46225
rect 147040 46215 147120 46225
rect 147360 46215 147440 46225
rect 148780 46215 148860 46225
rect 149100 46215 149180 46225
rect 149420 46215 149500 46225
rect 149740 46215 149820 46225
rect 152200 46215 152280 46225
rect 152520 46215 152600 46225
rect 152840 46215 152920 46225
rect 153160 46215 153240 46225
rect 153480 46215 153560 46225
rect 153800 46215 153880 46225
rect 154120 46215 154200 46225
rect 154440 46215 154520 46225
rect 154760 46215 154840 46225
rect 155080 46215 155160 46225
rect 155400 46215 155480 46225
rect 155720 46215 155800 46225
rect 156040 46215 156120 46225
rect 156360 46215 156440 46225
rect 156680 46215 156760 46225
rect 157000 46215 157080 46225
rect 157320 46215 157400 46225
rect 157640 46215 157720 46225
rect 157960 46215 158040 46225
rect 158280 46215 158360 46225
rect 158600 46215 158680 46225
rect 158920 46215 159000 46225
rect 159240 46215 159320 46225
rect 159560 46215 159640 46225
rect 30440 46135 30450 46215
rect 30760 46135 30770 46215
rect 31080 46135 31090 46215
rect 31400 46135 31410 46215
rect 31720 46135 31730 46215
rect 32040 46135 32050 46215
rect 32360 46135 32370 46215
rect 32680 46135 32690 46215
rect 33000 46135 33010 46215
rect 33320 46135 33330 46215
rect 33640 46135 33650 46215
rect 33960 46135 33970 46215
rect 34280 46135 34290 46215
rect 34600 46135 34610 46215
rect 34920 46135 34930 46215
rect 35240 46135 35250 46215
rect 35560 46135 35570 46215
rect 35880 46135 35890 46215
rect 36200 46135 36210 46215
rect 36520 46135 36530 46215
rect 36840 46135 36850 46215
rect 37160 46135 37170 46215
rect 37480 46135 37490 46215
rect 37800 46135 37810 46215
rect 40260 46135 40270 46215
rect 40580 46135 40590 46215
rect 40900 46135 40910 46215
rect 41220 46135 41230 46215
rect 42640 46135 42650 46215
rect 42960 46135 42970 46215
rect 43280 46135 43290 46215
rect 43600 46135 43610 46215
rect 146480 46135 146490 46215
rect 146800 46135 146810 46215
rect 147120 46135 147130 46215
rect 147440 46135 147450 46215
rect 148860 46135 148870 46215
rect 149180 46135 149190 46215
rect 149500 46135 149510 46215
rect 149820 46135 149830 46215
rect 152280 46135 152290 46215
rect 152600 46135 152610 46215
rect 152920 46135 152930 46215
rect 153240 46135 153250 46215
rect 153560 46135 153570 46215
rect 153880 46135 153890 46215
rect 154200 46135 154210 46215
rect 154520 46135 154530 46215
rect 154840 46135 154850 46215
rect 155160 46135 155170 46215
rect 155480 46135 155490 46215
rect 155800 46135 155810 46215
rect 156120 46135 156130 46215
rect 156440 46135 156450 46215
rect 156760 46135 156770 46215
rect 157080 46135 157090 46215
rect 157400 46135 157410 46215
rect 157720 46135 157730 46215
rect 158040 46135 158050 46215
rect 158360 46135 158370 46215
rect 158680 46135 158690 46215
rect 159000 46135 159010 46215
rect 159320 46135 159330 46215
rect 159640 46135 159650 46215
rect 163670 46175 163680 46255
rect 163990 46175 164000 46255
rect 164310 46175 164320 46255
rect 164630 46175 164640 46255
rect 164950 46175 164960 46255
rect 165270 46175 165280 46255
rect 165590 46175 165600 46255
rect 165910 46175 165920 46255
rect 166230 46175 166240 46255
rect 166550 46175 166560 46255
rect 166870 46175 166880 46255
rect 167190 46175 167200 46255
rect 167510 46175 167520 46255
rect 167830 46175 167840 46255
rect 168150 46175 168160 46255
rect 168470 46175 168480 46255
rect 168790 46175 168800 46255
rect 169110 46175 169120 46255
rect 169430 46175 169440 46255
rect 169750 46175 169760 46255
rect 170070 46175 170080 46255
rect 170390 46175 170400 46255
rect 170710 46175 170720 46255
rect 171030 46175 171040 46255
rect 19130 46095 19210 46105
rect 19450 46095 19530 46105
rect 19770 46095 19850 46105
rect 20090 46095 20170 46105
rect 20410 46095 20490 46105
rect 20730 46095 20810 46105
rect 21050 46095 21130 46105
rect 21370 46095 21450 46105
rect 21690 46095 21770 46105
rect 22010 46095 22090 46105
rect 22330 46095 22410 46105
rect 22650 46095 22730 46105
rect 22970 46095 23050 46105
rect 23290 46095 23370 46105
rect 23610 46095 23690 46105
rect 23930 46095 24010 46105
rect 24250 46095 24330 46105
rect 24570 46095 24650 46105
rect 24890 46095 24970 46105
rect 25210 46095 25290 46105
rect 25530 46095 25610 46105
rect 25850 46095 25930 46105
rect 26170 46095 26250 46105
rect 163750 46095 163830 46105
rect 164070 46095 164150 46105
rect 164390 46095 164470 46105
rect 164710 46095 164790 46105
rect 165030 46095 165110 46105
rect 165350 46095 165430 46105
rect 165670 46095 165750 46105
rect 165990 46095 166070 46105
rect 166310 46095 166390 46105
rect 166630 46095 166710 46105
rect 166950 46095 167030 46105
rect 167270 46095 167350 46105
rect 167590 46095 167670 46105
rect 167910 46095 167990 46105
rect 168230 46095 168310 46105
rect 168550 46095 168630 46105
rect 168870 46095 168950 46105
rect 169190 46095 169270 46105
rect 169510 46095 169590 46105
rect 169830 46095 169910 46105
rect 170150 46095 170230 46105
rect 170470 46095 170550 46105
rect 170790 46095 170870 46105
rect 19210 46015 19220 46095
rect 19530 46015 19540 46095
rect 19850 46015 19860 46095
rect 20170 46015 20180 46095
rect 20490 46015 20500 46095
rect 20810 46015 20820 46095
rect 21130 46015 21140 46095
rect 21450 46015 21460 46095
rect 21770 46015 21780 46095
rect 22090 46015 22100 46095
rect 22410 46015 22420 46095
rect 22730 46015 22740 46095
rect 23050 46015 23060 46095
rect 23370 46015 23380 46095
rect 23690 46015 23700 46095
rect 24010 46015 24020 46095
rect 24330 46015 24340 46095
rect 24650 46015 24660 46095
rect 24970 46015 24980 46095
rect 25290 46015 25300 46095
rect 25610 46015 25620 46095
rect 25930 46015 25940 46095
rect 26250 46015 26260 46095
rect 30520 46055 30600 46065
rect 30840 46055 30920 46065
rect 31160 46055 31240 46065
rect 31480 46055 31560 46065
rect 31800 46055 31880 46065
rect 32120 46055 32200 46065
rect 32440 46055 32520 46065
rect 32760 46055 32840 46065
rect 33080 46055 33160 46065
rect 33400 46055 33480 46065
rect 33720 46055 33800 46065
rect 34040 46055 34120 46065
rect 34360 46055 34440 46065
rect 34680 46055 34760 46065
rect 35000 46055 35080 46065
rect 35320 46055 35400 46065
rect 35640 46055 35720 46065
rect 35960 46055 36040 46065
rect 36280 46055 36360 46065
rect 36600 46055 36680 46065
rect 36920 46055 37000 46065
rect 37240 46055 37320 46065
rect 37560 46055 37640 46065
rect 40340 46055 40420 46065
rect 40660 46055 40740 46065
rect 40980 46055 41060 46065
rect 42720 46055 42800 46065
rect 43040 46055 43120 46065
rect 43360 46055 43440 46065
rect 146560 46055 146640 46065
rect 146880 46055 146960 46065
rect 147200 46055 147280 46065
rect 148940 46055 149020 46065
rect 149260 46055 149340 46065
rect 149580 46055 149660 46065
rect 152360 46055 152440 46065
rect 152680 46055 152760 46065
rect 153000 46055 153080 46065
rect 153320 46055 153400 46065
rect 153640 46055 153720 46065
rect 153960 46055 154040 46065
rect 154280 46055 154360 46065
rect 154600 46055 154680 46065
rect 154920 46055 155000 46065
rect 155240 46055 155320 46065
rect 155560 46055 155640 46065
rect 155880 46055 155960 46065
rect 156200 46055 156280 46065
rect 156520 46055 156600 46065
rect 156840 46055 156920 46065
rect 157160 46055 157240 46065
rect 157480 46055 157560 46065
rect 157800 46055 157880 46065
rect 158120 46055 158200 46065
rect 158440 46055 158520 46065
rect 158760 46055 158840 46065
rect 159080 46055 159160 46065
rect 159400 46055 159480 46065
rect 30600 45975 30610 46055
rect 30920 45975 30930 46055
rect 31240 45975 31250 46055
rect 31560 45975 31570 46055
rect 31880 45975 31890 46055
rect 32200 45975 32210 46055
rect 32520 45975 32530 46055
rect 32840 45975 32850 46055
rect 33160 45975 33170 46055
rect 33480 45975 33490 46055
rect 33800 45975 33810 46055
rect 34120 45975 34130 46055
rect 34440 45975 34450 46055
rect 34760 45975 34770 46055
rect 35080 45975 35090 46055
rect 35400 45975 35410 46055
rect 35720 45975 35730 46055
rect 36040 45975 36050 46055
rect 36360 45975 36370 46055
rect 36680 45975 36690 46055
rect 37000 45975 37010 46055
rect 37320 45975 37330 46055
rect 37640 45975 37650 46055
rect 40420 45975 40430 46055
rect 40740 45975 40750 46055
rect 41060 45975 41070 46055
rect 42800 45975 42810 46055
rect 43120 45975 43130 46055
rect 43440 45975 43450 46055
rect 146640 45975 146650 46055
rect 146960 45975 146970 46055
rect 147280 45975 147290 46055
rect 149020 45975 149030 46055
rect 149340 45975 149350 46055
rect 149660 45975 149670 46055
rect 152440 45975 152450 46055
rect 152760 45975 152770 46055
rect 153080 45975 153090 46055
rect 153400 45975 153410 46055
rect 153720 45975 153730 46055
rect 154040 45975 154050 46055
rect 154360 45975 154370 46055
rect 154680 45975 154690 46055
rect 155000 45975 155010 46055
rect 155320 45975 155330 46055
rect 155640 45975 155650 46055
rect 155960 45975 155970 46055
rect 156280 45975 156290 46055
rect 156600 45975 156610 46055
rect 156920 45975 156930 46055
rect 157240 45975 157250 46055
rect 157560 45975 157570 46055
rect 157880 45975 157890 46055
rect 158200 45975 158210 46055
rect 158520 45975 158530 46055
rect 158840 45975 158850 46055
rect 159160 45975 159170 46055
rect 159480 45975 159490 46055
rect 163830 46015 163840 46095
rect 164150 46015 164160 46095
rect 164470 46015 164480 46095
rect 164790 46015 164800 46095
rect 165110 46015 165120 46095
rect 165430 46015 165440 46095
rect 165750 46015 165760 46095
rect 166070 46015 166080 46095
rect 166390 46015 166400 46095
rect 166710 46015 166720 46095
rect 167030 46015 167040 46095
rect 167350 46015 167360 46095
rect 167670 46015 167680 46095
rect 167990 46015 168000 46095
rect 168310 46015 168320 46095
rect 168630 46015 168640 46095
rect 168950 46015 168960 46095
rect 169270 46015 169280 46095
rect 169590 46015 169600 46095
rect 169910 46015 169920 46095
rect 170230 46015 170240 46095
rect 170550 46015 170560 46095
rect 170870 46015 170880 46095
rect 18970 45935 19050 45945
rect 19290 45935 19370 45945
rect 19610 45935 19690 45945
rect 19930 45935 20010 45945
rect 20250 45935 20330 45945
rect 20570 45935 20650 45945
rect 20890 45935 20970 45945
rect 21210 45935 21290 45945
rect 21530 45935 21610 45945
rect 21850 45935 21930 45945
rect 22170 45935 22250 45945
rect 22490 45935 22570 45945
rect 22810 45935 22890 45945
rect 23130 45935 23210 45945
rect 23450 45935 23530 45945
rect 23770 45935 23850 45945
rect 24090 45935 24170 45945
rect 24410 45935 24490 45945
rect 24730 45935 24810 45945
rect 25050 45935 25130 45945
rect 25370 45935 25450 45945
rect 25690 45935 25770 45945
rect 26010 45935 26090 45945
rect 26330 45935 26410 45945
rect 163590 45935 163670 45945
rect 163910 45935 163990 45945
rect 164230 45935 164310 45945
rect 164550 45935 164630 45945
rect 164870 45935 164950 45945
rect 165190 45935 165270 45945
rect 165510 45935 165590 45945
rect 165830 45935 165910 45945
rect 166150 45935 166230 45945
rect 166470 45935 166550 45945
rect 166790 45935 166870 45945
rect 167110 45935 167190 45945
rect 167430 45935 167510 45945
rect 167750 45935 167830 45945
rect 168070 45935 168150 45945
rect 168390 45935 168470 45945
rect 168710 45935 168790 45945
rect 169030 45935 169110 45945
rect 169350 45935 169430 45945
rect 169670 45935 169750 45945
rect 169990 45935 170070 45945
rect 170310 45935 170390 45945
rect 170630 45935 170710 45945
rect 170950 45935 171030 45945
rect 19050 45855 19060 45935
rect 19370 45855 19380 45935
rect 19690 45855 19700 45935
rect 20010 45855 20020 45935
rect 20330 45855 20340 45935
rect 20650 45855 20660 45935
rect 20970 45855 20980 45935
rect 21290 45855 21300 45935
rect 21610 45855 21620 45935
rect 21930 45855 21940 45935
rect 22250 45855 22260 45935
rect 22570 45855 22580 45935
rect 22890 45855 22900 45935
rect 23210 45855 23220 45935
rect 23530 45855 23540 45935
rect 23850 45855 23860 45935
rect 24170 45855 24180 45935
rect 24490 45855 24500 45935
rect 24810 45855 24820 45935
rect 25130 45855 25140 45935
rect 25450 45855 25460 45935
rect 25770 45855 25780 45935
rect 26090 45855 26100 45935
rect 26410 45855 26420 45935
rect 30360 45895 30440 45905
rect 30680 45895 30760 45905
rect 31000 45895 31080 45905
rect 31320 45895 31400 45905
rect 31640 45895 31720 45905
rect 31960 45895 32040 45905
rect 32280 45895 32360 45905
rect 32600 45895 32680 45905
rect 32920 45895 33000 45905
rect 33240 45895 33320 45905
rect 33560 45895 33640 45905
rect 33880 45895 33960 45905
rect 34200 45895 34280 45905
rect 34520 45895 34600 45905
rect 34840 45895 34920 45905
rect 35160 45895 35240 45905
rect 35480 45895 35560 45905
rect 35800 45895 35880 45905
rect 36120 45895 36200 45905
rect 36440 45895 36520 45905
rect 36760 45895 36840 45905
rect 37080 45895 37160 45905
rect 37400 45895 37480 45905
rect 37720 45895 37800 45905
rect 40180 45895 40260 45905
rect 40500 45895 40580 45905
rect 40820 45895 40900 45905
rect 41140 45895 41220 45905
rect 42560 45895 42640 45905
rect 42880 45895 42960 45905
rect 43200 45895 43280 45905
rect 43520 45895 43600 45905
rect 146400 45895 146480 45905
rect 146720 45895 146800 45905
rect 147040 45895 147120 45905
rect 147360 45895 147440 45905
rect 148780 45895 148860 45905
rect 149100 45895 149180 45905
rect 149420 45895 149500 45905
rect 149740 45895 149820 45905
rect 152200 45895 152280 45905
rect 152520 45895 152600 45905
rect 152840 45895 152920 45905
rect 153160 45895 153240 45905
rect 153480 45895 153560 45905
rect 153800 45895 153880 45905
rect 154120 45895 154200 45905
rect 154440 45895 154520 45905
rect 154760 45895 154840 45905
rect 155080 45895 155160 45905
rect 155400 45895 155480 45905
rect 155720 45895 155800 45905
rect 156040 45895 156120 45905
rect 156360 45895 156440 45905
rect 156680 45895 156760 45905
rect 157000 45895 157080 45905
rect 157320 45895 157400 45905
rect 157640 45895 157720 45905
rect 157960 45895 158040 45905
rect 158280 45895 158360 45905
rect 158600 45895 158680 45905
rect 158920 45895 159000 45905
rect 159240 45895 159320 45905
rect 159560 45895 159640 45905
rect 30440 45815 30450 45895
rect 30760 45815 30770 45895
rect 31080 45815 31090 45895
rect 31400 45815 31410 45895
rect 31720 45815 31730 45895
rect 32040 45815 32050 45895
rect 32360 45815 32370 45895
rect 32680 45815 32690 45895
rect 33000 45815 33010 45895
rect 33320 45815 33330 45895
rect 33640 45815 33650 45895
rect 33960 45815 33970 45895
rect 34280 45815 34290 45895
rect 34600 45815 34610 45895
rect 34920 45815 34930 45895
rect 35240 45815 35250 45895
rect 35560 45815 35570 45895
rect 35880 45815 35890 45895
rect 36200 45815 36210 45895
rect 36520 45815 36530 45895
rect 36840 45815 36850 45895
rect 37160 45815 37170 45895
rect 37480 45815 37490 45895
rect 37800 45815 37810 45895
rect 40260 45815 40270 45895
rect 40580 45815 40590 45895
rect 40900 45815 40910 45895
rect 41220 45815 41230 45895
rect 42640 45815 42650 45895
rect 42960 45815 42970 45895
rect 43280 45815 43290 45895
rect 43600 45815 43610 45895
rect 146480 45815 146490 45895
rect 146800 45815 146810 45895
rect 147120 45815 147130 45895
rect 147440 45815 147450 45895
rect 148860 45815 148870 45895
rect 149180 45815 149190 45895
rect 149500 45815 149510 45895
rect 149820 45815 149830 45895
rect 152280 45815 152290 45895
rect 152600 45815 152610 45895
rect 152920 45815 152930 45895
rect 153240 45815 153250 45895
rect 153560 45815 153570 45895
rect 153880 45815 153890 45895
rect 154200 45815 154210 45895
rect 154520 45815 154530 45895
rect 154840 45815 154850 45895
rect 155160 45815 155170 45895
rect 155480 45815 155490 45895
rect 155800 45815 155810 45895
rect 156120 45815 156130 45895
rect 156440 45815 156450 45895
rect 156760 45815 156770 45895
rect 157080 45815 157090 45895
rect 157400 45815 157410 45895
rect 157720 45815 157730 45895
rect 158040 45815 158050 45895
rect 158360 45815 158370 45895
rect 158680 45815 158690 45895
rect 159000 45815 159010 45895
rect 159320 45815 159330 45895
rect 159640 45815 159650 45895
rect 163670 45855 163680 45935
rect 163990 45855 164000 45935
rect 164310 45855 164320 45935
rect 164630 45855 164640 45935
rect 164950 45855 164960 45935
rect 165270 45855 165280 45935
rect 165590 45855 165600 45935
rect 165910 45855 165920 45935
rect 166230 45855 166240 45935
rect 166550 45855 166560 45935
rect 166870 45855 166880 45935
rect 167190 45855 167200 45935
rect 167510 45855 167520 45935
rect 167830 45855 167840 45935
rect 168150 45855 168160 45935
rect 168470 45855 168480 45935
rect 168790 45855 168800 45935
rect 169110 45855 169120 45935
rect 169430 45855 169440 45935
rect 169750 45855 169760 45935
rect 170070 45855 170080 45935
rect 170390 45855 170400 45935
rect 170710 45855 170720 45935
rect 171030 45855 171040 45935
rect 19130 45775 19210 45785
rect 19450 45775 19530 45785
rect 19770 45775 19850 45785
rect 20090 45775 20170 45785
rect 20410 45775 20490 45785
rect 20730 45775 20810 45785
rect 21050 45775 21130 45785
rect 21370 45775 21450 45785
rect 21690 45775 21770 45785
rect 22010 45775 22090 45785
rect 22330 45775 22410 45785
rect 22650 45775 22730 45785
rect 22970 45775 23050 45785
rect 23290 45775 23370 45785
rect 23610 45775 23690 45785
rect 23930 45775 24010 45785
rect 24250 45775 24330 45785
rect 24570 45775 24650 45785
rect 24890 45775 24970 45785
rect 25210 45775 25290 45785
rect 25530 45775 25610 45785
rect 25850 45775 25930 45785
rect 26170 45775 26250 45785
rect 163750 45775 163830 45785
rect 164070 45775 164150 45785
rect 164390 45775 164470 45785
rect 164710 45775 164790 45785
rect 165030 45775 165110 45785
rect 165350 45775 165430 45785
rect 165670 45775 165750 45785
rect 165990 45775 166070 45785
rect 166310 45775 166390 45785
rect 166630 45775 166710 45785
rect 166950 45775 167030 45785
rect 167270 45775 167350 45785
rect 167590 45775 167670 45785
rect 167910 45775 167990 45785
rect 168230 45775 168310 45785
rect 168550 45775 168630 45785
rect 168870 45775 168950 45785
rect 169190 45775 169270 45785
rect 169510 45775 169590 45785
rect 169830 45775 169910 45785
rect 170150 45775 170230 45785
rect 170470 45775 170550 45785
rect 170790 45775 170870 45785
rect 19210 45695 19220 45775
rect 19530 45695 19540 45775
rect 19850 45695 19860 45775
rect 20170 45695 20180 45775
rect 20490 45695 20500 45775
rect 20810 45695 20820 45775
rect 21130 45695 21140 45775
rect 21450 45695 21460 45775
rect 21770 45695 21780 45775
rect 22090 45695 22100 45775
rect 22410 45695 22420 45775
rect 22730 45695 22740 45775
rect 23050 45695 23060 45775
rect 23370 45695 23380 45775
rect 23690 45695 23700 45775
rect 24010 45695 24020 45775
rect 24330 45695 24340 45775
rect 24650 45695 24660 45775
rect 24970 45695 24980 45775
rect 25290 45695 25300 45775
rect 25610 45695 25620 45775
rect 25930 45695 25940 45775
rect 26250 45695 26260 45775
rect 30520 45735 30600 45745
rect 30840 45735 30920 45745
rect 31160 45735 31240 45745
rect 31480 45735 31560 45745
rect 31800 45735 31880 45745
rect 32120 45735 32200 45745
rect 32440 45735 32520 45745
rect 32760 45735 32840 45745
rect 33080 45735 33160 45745
rect 33400 45735 33480 45745
rect 33720 45735 33800 45745
rect 34040 45735 34120 45745
rect 34360 45735 34440 45745
rect 34680 45735 34760 45745
rect 35000 45735 35080 45745
rect 35320 45735 35400 45745
rect 35640 45735 35720 45745
rect 35960 45735 36040 45745
rect 36280 45735 36360 45745
rect 36600 45735 36680 45745
rect 36920 45735 37000 45745
rect 37240 45735 37320 45745
rect 37560 45735 37640 45745
rect 40340 45735 40420 45745
rect 40660 45735 40740 45745
rect 40980 45735 41060 45745
rect 42720 45735 42800 45745
rect 43040 45735 43120 45745
rect 43360 45735 43440 45745
rect 146560 45735 146640 45745
rect 146880 45735 146960 45745
rect 147200 45735 147280 45745
rect 148940 45735 149020 45745
rect 149260 45735 149340 45745
rect 149580 45735 149660 45745
rect 152360 45735 152440 45745
rect 152680 45735 152760 45745
rect 153000 45735 153080 45745
rect 153320 45735 153400 45745
rect 153640 45735 153720 45745
rect 153960 45735 154040 45745
rect 154280 45735 154360 45745
rect 154600 45735 154680 45745
rect 154920 45735 155000 45745
rect 155240 45735 155320 45745
rect 155560 45735 155640 45745
rect 155880 45735 155960 45745
rect 156200 45735 156280 45745
rect 156520 45735 156600 45745
rect 156840 45735 156920 45745
rect 157160 45735 157240 45745
rect 157480 45735 157560 45745
rect 157800 45735 157880 45745
rect 158120 45735 158200 45745
rect 158440 45735 158520 45745
rect 158760 45735 158840 45745
rect 159080 45735 159160 45745
rect 159400 45735 159480 45745
rect 30600 45655 30610 45735
rect 30920 45655 30930 45735
rect 31240 45655 31250 45735
rect 31560 45655 31570 45735
rect 31880 45655 31890 45735
rect 32200 45655 32210 45735
rect 32520 45655 32530 45735
rect 32840 45655 32850 45735
rect 33160 45655 33170 45735
rect 33480 45655 33490 45735
rect 33800 45655 33810 45735
rect 34120 45655 34130 45735
rect 34440 45655 34450 45735
rect 34760 45655 34770 45735
rect 35080 45655 35090 45735
rect 35400 45655 35410 45735
rect 35720 45655 35730 45735
rect 36040 45655 36050 45735
rect 36360 45655 36370 45735
rect 36680 45655 36690 45735
rect 37000 45655 37010 45735
rect 37320 45655 37330 45735
rect 37640 45655 37650 45735
rect 40420 45655 40430 45735
rect 40740 45655 40750 45735
rect 41060 45655 41070 45735
rect 42800 45655 42810 45735
rect 43120 45655 43130 45735
rect 43440 45655 43450 45735
rect 146640 45655 146650 45735
rect 146960 45655 146970 45735
rect 147280 45655 147290 45735
rect 149020 45655 149030 45735
rect 149340 45655 149350 45735
rect 149660 45655 149670 45735
rect 152440 45655 152450 45735
rect 152760 45655 152770 45735
rect 153080 45655 153090 45735
rect 153400 45655 153410 45735
rect 153720 45655 153730 45735
rect 154040 45655 154050 45735
rect 154360 45655 154370 45735
rect 154680 45655 154690 45735
rect 155000 45655 155010 45735
rect 155320 45655 155330 45735
rect 155640 45655 155650 45735
rect 155960 45655 155970 45735
rect 156280 45655 156290 45735
rect 156600 45655 156610 45735
rect 156920 45655 156930 45735
rect 157240 45655 157250 45735
rect 157560 45655 157570 45735
rect 157880 45655 157890 45735
rect 158200 45655 158210 45735
rect 158520 45655 158530 45735
rect 158840 45655 158850 45735
rect 159160 45655 159170 45735
rect 159480 45655 159490 45735
rect 163830 45695 163840 45775
rect 164150 45695 164160 45775
rect 164470 45695 164480 45775
rect 164790 45695 164800 45775
rect 165110 45695 165120 45775
rect 165430 45695 165440 45775
rect 165750 45695 165760 45775
rect 166070 45695 166080 45775
rect 166390 45695 166400 45775
rect 166710 45695 166720 45775
rect 167030 45695 167040 45775
rect 167350 45695 167360 45775
rect 167670 45695 167680 45775
rect 167990 45695 168000 45775
rect 168310 45695 168320 45775
rect 168630 45695 168640 45775
rect 168950 45695 168960 45775
rect 169270 45695 169280 45775
rect 169590 45695 169600 45775
rect 169910 45695 169920 45775
rect 170230 45695 170240 45775
rect 170550 45695 170560 45775
rect 170870 45695 170880 45775
rect 18970 45615 19050 45625
rect 19290 45615 19370 45625
rect 19610 45615 19690 45625
rect 19930 45615 20010 45625
rect 20250 45615 20330 45625
rect 20570 45615 20650 45625
rect 20890 45615 20970 45625
rect 21210 45615 21290 45625
rect 21530 45615 21610 45625
rect 21850 45615 21930 45625
rect 22170 45615 22250 45625
rect 22490 45615 22570 45625
rect 22810 45615 22890 45625
rect 23130 45615 23210 45625
rect 23450 45615 23530 45625
rect 23770 45615 23850 45625
rect 24090 45615 24170 45625
rect 24410 45615 24490 45625
rect 24730 45615 24810 45625
rect 25050 45615 25130 45625
rect 25370 45615 25450 45625
rect 25690 45615 25770 45625
rect 26010 45615 26090 45625
rect 26330 45615 26410 45625
rect 163590 45615 163670 45625
rect 163910 45615 163990 45625
rect 164230 45615 164310 45625
rect 164550 45615 164630 45625
rect 164870 45615 164950 45625
rect 165190 45615 165270 45625
rect 165510 45615 165590 45625
rect 165830 45615 165910 45625
rect 166150 45615 166230 45625
rect 166470 45615 166550 45625
rect 166790 45615 166870 45625
rect 167110 45615 167190 45625
rect 167430 45615 167510 45625
rect 167750 45615 167830 45625
rect 168070 45615 168150 45625
rect 168390 45615 168470 45625
rect 168710 45615 168790 45625
rect 169030 45615 169110 45625
rect 169350 45615 169430 45625
rect 169670 45615 169750 45625
rect 169990 45615 170070 45625
rect 170310 45615 170390 45625
rect 170630 45615 170710 45625
rect 170950 45615 171030 45625
rect 19050 45535 19060 45615
rect 19370 45535 19380 45615
rect 19690 45535 19700 45615
rect 20010 45535 20020 45615
rect 20330 45535 20340 45615
rect 20650 45535 20660 45615
rect 20970 45535 20980 45615
rect 21290 45535 21300 45615
rect 21610 45535 21620 45615
rect 21930 45535 21940 45615
rect 22250 45535 22260 45615
rect 22570 45535 22580 45615
rect 22890 45535 22900 45615
rect 23210 45535 23220 45615
rect 23530 45535 23540 45615
rect 23850 45535 23860 45615
rect 24170 45535 24180 45615
rect 24490 45535 24500 45615
rect 24810 45535 24820 45615
rect 25130 45535 25140 45615
rect 25450 45535 25460 45615
rect 25770 45535 25780 45615
rect 26090 45535 26100 45615
rect 26410 45535 26420 45615
rect 30360 45575 30440 45585
rect 30680 45575 30760 45585
rect 31000 45575 31080 45585
rect 31320 45575 31400 45585
rect 31640 45575 31720 45585
rect 31960 45575 32040 45585
rect 32280 45575 32360 45585
rect 32600 45575 32680 45585
rect 32920 45575 33000 45585
rect 33240 45575 33320 45585
rect 33560 45575 33640 45585
rect 33880 45575 33960 45585
rect 34200 45575 34280 45585
rect 34520 45575 34600 45585
rect 34840 45575 34920 45585
rect 35160 45575 35240 45585
rect 35480 45575 35560 45585
rect 35800 45575 35880 45585
rect 36120 45575 36200 45585
rect 36440 45575 36520 45585
rect 36760 45575 36840 45585
rect 37080 45575 37160 45585
rect 37400 45575 37480 45585
rect 37720 45575 37800 45585
rect 40180 45575 40260 45585
rect 40500 45575 40580 45585
rect 40820 45575 40900 45585
rect 41140 45575 41220 45585
rect 42560 45575 42640 45585
rect 42880 45575 42960 45585
rect 43200 45575 43280 45585
rect 43520 45575 43600 45585
rect 146400 45575 146480 45585
rect 146720 45575 146800 45585
rect 147040 45575 147120 45585
rect 147360 45575 147440 45585
rect 148780 45575 148860 45585
rect 149100 45575 149180 45585
rect 149420 45575 149500 45585
rect 149740 45575 149820 45585
rect 152200 45575 152280 45585
rect 152520 45575 152600 45585
rect 152840 45575 152920 45585
rect 153160 45575 153240 45585
rect 153480 45575 153560 45585
rect 153800 45575 153880 45585
rect 154120 45575 154200 45585
rect 154440 45575 154520 45585
rect 154760 45575 154840 45585
rect 155080 45575 155160 45585
rect 155400 45575 155480 45585
rect 155720 45575 155800 45585
rect 156040 45575 156120 45585
rect 156360 45575 156440 45585
rect 156680 45575 156760 45585
rect 157000 45575 157080 45585
rect 157320 45575 157400 45585
rect 157640 45575 157720 45585
rect 157960 45575 158040 45585
rect 158280 45575 158360 45585
rect 158600 45575 158680 45585
rect 158920 45575 159000 45585
rect 159240 45575 159320 45585
rect 159560 45575 159640 45585
rect 30440 45495 30450 45575
rect 30760 45495 30770 45575
rect 31080 45495 31090 45575
rect 31400 45495 31410 45575
rect 31720 45495 31730 45575
rect 32040 45495 32050 45575
rect 32360 45495 32370 45575
rect 32680 45495 32690 45575
rect 33000 45495 33010 45575
rect 33320 45495 33330 45575
rect 33640 45495 33650 45575
rect 33960 45495 33970 45575
rect 34280 45495 34290 45575
rect 34600 45495 34610 45575
rect 34920 45495 34930 45575
rect 35240 45495 35250 45575
rect 35560 45495 35570 45575
rect 35880 45495 35890 45575
rect 36200 45495 36210 45575
rect 36520 45495 36530 45575
rect 36840 45495 36850 45575
rect 37160 45495 37170 45575
rect 37480 45495 37490 45575
rect 37800 45495 37810 45575
rect 40260 45495 40270 45575
rect 40580 45495 40590 45575
rect 40900 45495 40910 45575
rect 41220 45495 41230 45575
rect 42640 45495 42650 45575
rect 42960 45495 42970 45575
rect 43280 45495 43290 45575
rect 43600 45495 43610 45575
rect 146480 45495 146490 45575
rect 146800 45495 146810 45575
rect 147120 45495 147130 45575
rect 147440 45495 147450 45575
rect 148860 45495 148870 45575
rect 149180 45495 149190 45575
rect 149500 45495 149510 45575
rect 149820 45495 149830 45575
rect 152280 45495 152290 45575
rect 152600 45495 152610 45575
rect 152920 45495 152930 45575
rect 153240 45495 153250 45575
rect 153560 45495 153570 45575
rect 153880 45495 153890 45575
rect 154200 45495 154210 45575
rect 154520 45495 154530 45575
rect 154840 45495 154850 45575
rect 155160 45495 155170 45575
rect 155480 45495 155490 45575
rect 155800 45495 155810 45575
rect 156120 45495 156130 45575
rect 156440 45495 156450 45575
rect 156760 45495 156770 45575
rect 157080 45495 157090 45575
rect 157400 45495 157410 45575
rect 157720 45495 157730 45575
rect 158040 45495 158050 45575
rect 158360 45495 158370 45575
rect 158680 45495 158690 45575
rect 159000 45495 159010 45575
rect 159320 45495 159330 45575
rect 159640 45495 159650 45575
rect 163670 45535 163680 45615
rect 163990 45535 164000 45615
rect 164310 45535 164320 45615
rect 164630 45535 164640 45615
rect 164950 45535 164960 45615
rect 165270 45535 165280 45615
rect 165590 45535 165600 45615
rect 165910 45535 165920 45615
rect 166230 45535 166240 45615
rect 166550 45535 166560 45615
rect 166870 45535 166880 45615
rect 167190 45535 167200 45615
rect 167510 45535 167520 45615
rect 167830 45535 167840 45615
rect 168150 45535 168160 45615
rect 168470 45535 168480 45615
rect 168790 45535 168800 45615
rect 169110 45535 169120 45615
rect 169430 45535 169440 45615
rect 169750 45535 169760 45615
rect 170070 45535 170080 45615
rect 170390 45535 170400 45615
rect 170710 45535 170720 45615
rect 171030 45535 171040 45615
rect 19130 45455 19210 45465
rect 19450 45455 19530 45465
rect 19770 45455 19850 45465
rect 20090 45455 20170 45465
rect 20410 45455 20490 45465
rect 20730 45455 20810 45465
rect 21050 45455 21130 45465
rect 21370 45455 21450 45465
rect 21690 45455 21770 45465
rect 22010 45455 22090 45465
rect 22330 45455 22410 45465
rect 22650 45455 22730 45465
rect 22970 45455 23050 45465
rect 23290 45455 23370 45465
rect 23610 45455 23690 45465
rect 23930 45455 24010 45465
rect 24250 45455 24330 45465
rect 24570 45455 24650 45465
rect 24890 45455 24970 45465
rect 25210 45455 25290 45465
rect 25530 45455 25610 45465
rect 25850 45455 25930 45465
rect 26170 45455 26250 45465
rect 163750 45455 163830 45465
rect 164070 45455 164150 45465
rect 164390 45455 164470 45465
rect 164710 45455 164790 45465
rect 165030 45455 165110 45465
rect 165350 45455 165430 45465
rect 165670 45455 165750 45465
rect 165990 45455 166070 45465
rect 166310 45455 166390 45465
rect 166630 45455 166710 45465
rect 166950 45455 167030 45465
rect 167270 45455 167350 45465
rect 167590 45455 167670 45465
rect 167910 45455 167990 45465
rect 168230 45455 168310 45465
rect 168550 45455 168630 45465
rect 168870 45455 168950 45465
rect 169190 45455 169270 45465
rect 169510 45455 169590 45465
rect 169830 45455 169910 45465
rect 170150 45455 170230 45465
rect 170470 45455 170550 45465
rect 170790 45455 170870 45465
rect 19210 45375 19220 45455
rect 19530 45375 19540 45455
rect 19850 45375 19860 45455
rect 20170 45375 20180 45455
rect 20490 45375 20500 45455
rect 20810 45375 20820 45455
rect 21130 45375 21140 45455
rect 21450 45375 21460 45455
rect 21770 45375 21780 45455
rect 22090 45375 22100 45455
rect 22410 45375 22420 45455
rect 22730 45375 22740 45455
rect 23050 45375 23060 45455
rect 23370 45375 23380 45455
rect 23690 45375 23700 45455
rect 24010 45375 24020 45455
rect 24330 45375 24340 45455
rect 24650 45375 24660 45455
rect 24970 45375 24980 45455
rect 25290 45375 25300 45455
rect 25610 45375 25620 45455
rect 25930 45375 25940 45455
rect 26250 45375 26260 45455
rect 30520 45415 30600 45425
rect 30840 45415 30920 45425
rect 31160 45415 31240 45425
rect 31480 45415 31560 45425
rect 31800 45415 31880 45425
rect 32120 45415 32200 45425
rect 32440 45415 32520 45425
rect 32760 45415 32840 45425
rect 33080 45415 33160 45425
rect 33400 45415 33480 45425
rect 33720 45415 33800 45425
rect 34040 45415 34120 45425
rect 34360 45415 34440 45425
rect 34680 45415 34760 45425
rect 35000 45415 35080 45425
rect 35320 45415 35400 45425
rect 35640 45415 35720 45425
rect 35960 45415 36040 45425
rect 36280 45415 36360 45425
rect 36600 45415 36680 45425
rect 36920 45415 37000 45425
rect 37240 45415 37320 45425
rect 37560 45415 37640 45425
rect 40340 45415 40420 45425
rect 40660 45415 40740 45425
rect 40980 45415 41060 45425
rect 42720 45415 42800 45425
rect 43040 45415 43120 45425
rect 43360 45415 43440 45425
rect 146560 45415 146640 45425
rect 146880 45415 146960 45425
rect 147200 45415 147280 45425
rect 148940 45415 149020 45425
rect 149260 45415 149340 45425
rect 149580 45415 149660 45425
rect 152360 45415 152440 45425
rect 152680 45415 152760 45425
rect 153000 45415 153080 45425
rect 153320 45415 153400 45425
rect 153640 45415 153720 45425
rect 153960 45415 154040 45425
rect 154280 45415 154360 45425
rect 154600 45415 154680 45425
rect 154920 45415 155000 45425
rect 155240 45415 155320 45425
rect 155560 45415 155640 45425
rect 155880 45415 155960 45425
rect 156200 45415 156280 45425
rect 156520 45415 156600 45425
rect 156840 45415 156920 45425
rect 157160 45415 157240 45425
rect 157480 45415 157560 45425
rect 157800 45415 157880 45425
rect 158120 45415 158200 45425
rect 158440 45415 158520 45425
rect 158760 45415 158840 45425
rect 159080 45415 159160 45425
rect 159400 45415 159480 45425
rect 30600 45335 30610 45415
rect 30920 45335 30930 45415
rect 31240 45335 31250 45415
rect 31560 45335 31570 45415
rect 31880 45335 31890 45415
rect 32200 45335 32210 45415
rect 32520 45335 32530 45415
rect 32840 45335 32850 45415
rect 33160 45335 33170 45415
rect 33480 45335 33490 45415
rect 33800 45335 33810 45415
rect 34120 45335 34130 45415
rect 34440 45335 34450 45415
rect 34760 45335 34770 45415
rect 35080 45335 35090 45415
rect 35400 45335 35410 45415
rect 35720 45335 35730 45415
rect 36040 45335 36050 45415
rect 36360 45335 36370 45415
rect 36680 45335 36690 45415
rect 37000 45335 37010 45415
rect 37320 45335 37330 45415
rect 37640 45335 37650 45415
rect 40420 45335 40430 45415
rect 40740 45335 40750 45415
rect 41060 45335 41070 45415
rect 42800 45335 42810 45415
rect 43120 45335 43130 45415
rect 43440 45335 43450 45415
rect 146640 45335 146650 45415
rect 146960 45335 146970 45415
rect 147280 45335 147290 45415
rect 149020 45335 149030 45415
rect 149340 45335 149350 45415
rect 149660 45335 149670 45415
rect 152440 45335 152450 45415
rect 152760 45335 152770 45415
rect 153080 45335 153090 45415
rect 153400 45335 153410 45415
rect 153720 45335 153730 45415
rect 154040 45335 154050 45415
rect 154360 45335 154370 45415
rect 154680 45335 154690 45415
rect 155000 45335 155010 45415
rect 155320 45335 155330 45415
rect 155640 45335 155650 45415
rect 155960 45335 155970 45415
rect 156280 45335 156290 45415
rect 156600 45335 156610 45415
rect 156920 45335 156930 45415
rect 157240 45335 157250 45415
rect 157560 45335 157570 45415
rect 157880 45335 157890 45415
rect 158200 45335 158210 45415
rect 158520 45335 158530 45415
rect 158840 45335 158850 45415
rect 159160 45335 159170 45415
rect 159480 45335 159490 45415
rect 163830 45375 163840 45455
rect 164150 45375 164160 45455
rect 164470 45375 164480 45455
rect 164790 45375 164800 45455
rect 165110 45375 165120 45455
rect 165430 45375 165440 45455
rect 165750 45375 165760 45455
rect 166070 45375 166080 45455
rect 166390 45375 166400 45455
rect 166710 45375 166720 45455
rect 167030 45375 167040 45455
rect 167350 45375 167360 45455
rect 167670 45375 167680 45455
rect 167990 45375 168000 45455
rect 168310 45375 168320 45455
rect 168630 45375 168640 45455
rect 168950 45375 168960 45455
rect 169270 45375 169280 45455
rect 169590 45375 169600 45455
rect 169910 45375 169920 45455
rect 170230 45375 170240 45455
rect 170550 45375 170560 45455
rect 170870 45375 170880 45455
rect 18970 45295 19050 45305
rect 19290 45295 19370 45305
rect 19610 45295 19690 45305
rect 19930 45295 20010 45305
rect 20250 45295 20330 45305
rect 20570 45295 20650 45305
rect 20890 45295 20970 45305
rect 21210 45295 21290 45305
rect 21530 45295 21610 45305
rect 21850 45295 21930 45305
rect 22170 45295 22250 45305
rect 22490 45295 22570 45305
rect 22810 45295 22890 45305
rect 23130 45295 23210 45305
rect 23450 45295 23530 45305
rect 23770 45295 23850 45305
rect 24090 45295 24170 45305
rect 24410 45295 24490 45305
rect 24730 45295 24810 45305
rect 25050 45295 25130 45305
rect 25370 45295 25450 45305
rect 25690 45295 25770 45305
rect 26010 45295 26090 45305
rect 26330 45295 26410 45305
rect 163590 45295 163670 45305
rect 163910 45295 163990 45305
rect 164230 45295 164310 45305
rect 164550 45295 164630 45305
rect 164870 45295 164950 45305
rect 165190 45295 165270 45305
rect 165510 45295 165590 45305
rect 165830 45295 165910 45305
rect 166150 45295 166230 45305
rect 166470 45295 166550 45305
rect 166790 45295 166870 45305
rect 167110 45295 167190 45305
rect 167430 45295 167510 45305
rect 167750 45295 167830 45305
rect 168070 45295 168150 45305
rect 168390 45295 168470 45305
rect 168710 45295 168790 45305
rect 169030 45295 169110 45305
rect 169350 45295 169430 45305
rect 169670 45295 169750 45305
rect 169990 45295 170070 45305
rect 170310 45295 170390 45305
rect 170630 45295 170710 45305
rect 170950 45295 171030 45305
rect 19050 45215 19060 45295
rect 19370 45215 19380 45295
rect 19690 45215 19700 45295
rect 20010 45215 20020 45295
rect 20330 45215 20340 45295
rect 20650 45215 20660 45295
rect 20970 45215 20980 45295
rect 21290 45215 21300 45295
rect 21610 45215 21620 45295
rect 21930 45215 21940 45295
rect 22250 45215 22260 45295
rect 22570 45215 22580 45295
rect 22890 45215 22900 45295
rect 23210 45215 23220 45295
rect 23530 45215 23540 45295
rect 23850 45215 23860 45295
rect 24170 45215 24180 45295
rect 24490 45215 24500 45295
rect 24810 45215 24820 45295
rect 25130 45215 25140 45295
rect 25450 45215 25460 45295
rect 25770 45215 25780 45295
rect 26090 45215 26100 45295
rect 26410 45215 26420 45295
rect 30360 45255 30440 45265
rect 30680 45255 30760 45265
rect 31000 45255 31080 45265
rect 31320 45255 31400 45265
rect 31640 45255 31720 45265
rect 31960 45255 32040 45265
rect 32280 45255 32360 45265
rect 32600 45255 32680 45265
rect 32920 45255 33000 45265
rect 33240 45255 33320 45265
rect 33560 45255 33640 45265
rect 33880 45255 33960 45265
rect 34200 45255 34280 45265
rect 34520 45255 34600 45265
rect 34840 45255 34920 45265
rect 35160 45255 35240 45265
rect 35480 45255 35560 45265
rect 35800 45255 35880 45265
rect 36120 45255 36200 45265
rect 36440 45255 36520 45265
rect 36760 45255 36840 45265
rect 37080 45255 37160 45265
rect 37400 45255 37480 45265
rect 37720 45255 37800 45265
rect 40180 45255 40260 45265
rect 40500 45255 40580 45265
rect 40820 45255 40900 45265
rect 41140 45255 41220 45265
rect 42560 45255 42640 45265
rect 42880 45255 42960 45265
rect 43200 45255 43280 45265
rect 43520 45255 43600 45265
rect 146400 45255 146480 45265
rect 146720 45255 146800 45265
rect 147040 45255 147120 45265
rect 147360 45255 147440 45265
rect 148780 45255 148860 45265
rect 149100 45255 149180 45265
rect 149420 45255 149500 45265
rect 149740 45255 149820 45265
rect 152200 45255 152280 45265
rect 152520 45255 152600 45265
rect 152840 45255 152920 45265
rect 153160 45255 153240 45265
rect 153480 45255 153560 45265
rect 153800 45255 153880 45265
rect 154120 45255 154200 45265
rect 154440 45255 154520 45265
rect 154760 45255 154840 45265
rect 155080 45255 155160 45265
rect 155400 45255 155480 45265
rect 155720 45255 155800 45265
rect 156040 45255 156120 45265
rect 156360 45255 156440 45265
rect 156680 45255 156760 45265
rect 157000 45255 157080 45265
rect 157320 45255 157400 45265
rect 157640 45255 157720 45265
rect 157960 45255 158040 45265
rect 158280 45255 158360 45265
rect 158600 45255 158680 45265
rect 158920 45255 159000 45265
rect 159240 45255 159320 45265
rect 159560 45255 159640 45265
rect 30440 45175 30450 45255
rect 30760 45175 30770 45255
rect 31080 45175 31090 45255
rect 31400 45175 31410 45255
rect 31720 45175 31730 45255
rect 32040 45175 32050 45255
rect 32360 45175 32370 45255
rect 32680 45175 32690 45255
rect 33000 45175 33010 45255
rect 33320 45175 33330 45255
rect 33640 45175 33650 45255
rect 33960 45175 33970 45255
rect 34280 45175 34290 45255
rect 34600 45175 34610 45255
rect 34920 45175 34930 45255
rect 35240 45175 35250 45255
rect 35560 45175 35570 45255
rect 35880 45175 35890 45255
rect 36200 45175 36210 45255
rect 36520 45175 36530 45255
rect 36840 45175 36850 45255
rect 37160 45175 37170 45255
rect 37480 45175 37490 45255
rect 37800 45175 37810 45255
rect 40260 45175 40270 45255
rect 40580 45175 40590 45255
rect 40900 45175 40910 45255
rect 41220 45175 41230 45255
rect 42640 45175 42650 45255
rect 42960 45175 42970 45255
rect 43280 45175 43290 45255
rect 43600 45175 43610 45255
rect 146480 45175 146490 45255
rect 146800 45175 146810 45255
rect 147120 45175 147130 45255
rect 147440 45175 147450 45255
rect 148860 45175 148870 45255
rect 149180 45175 149190 45255
rect 149500 45175 149510 45255
rect 149820 45175 149830 45255
rect 152280 45175 152290 45255
rect 152600 45175 152610 45255
rect 152920 45175 152930 45255
rect 153240 45175 153250 45255
rect 153560 45175 153570 45255
rect 153880 45175 153890 45255
rect 154200 45175 154210 45255
rect 154520 45175 154530 45255
rect 154840 45175 154850 45255
rect 155160 45175 155170 45255
rect 155480 45175 155490 45255
rect 155800 45175 155810 45255
rect 156120 45175 156130 45255
rect 156440 45175 156450 45255
rect 156760 45175 156770 45255
rect 157080 45175 157090 45255
rect 157400 45175 157410 45255
rect 157720 45175 157730 45255
rect 158040 45175 158050 45255
rect 158360 45175 158370 45255
rect 158680 45175 158690 45255
rect 159000 45175 159010 45255
rect 159320 45175 159330 45255
rect 159640 45175 159650 45255
rect 163670 45215 163680 45295
rect 163990 45215 164000 45295
rect 164310 45215 164320 45295
rect 164630 45215 164640 45295
rect 164950 45215 164960 45295
rect 165270 45215 165280 45295
rect 165590 45215 165600 45295
rect 165910 45215 165920 45295
rect 166230 45215 166240 45295
rect 166550 45215 166560 45295
rect 166870 45215 166880 45295
rect 167190 45215 167200 45295
rect 167510 45215 167520 45295
rect 167830 45215 167840 45295
rect 168150 45215 168160 45295
rect 168470 45215 168480 45295
rect 168790 45215 168800 45295
rect 169110 45215 169120 45295
rect 169430 45215 169440 45295
rect 169750 45215 169760 45295
rect 170070 45215 170080 45295
rect 170390 45215 170400 45295
rect 170710 45215 170720 45295
rect 171030 45215 171040 45295
rect 19130 45135 19210 45145
rect 19450 45135 19530 45145
rect 19770 45135 19850 45145
rect 20090 45135 20170 45145
rect 20410 45135 20490 45145
rect 20730 45135 20810 45145
rect 21050 45135 21130 45145
rect 21370 45135 21450 45145
rect 21690 45135 21770 45145
rect 22010 45135 22090 45145
rect 22330 45135 22410 45145
rect 22650 45135 22730 45145
rect 22970 45135 23050 45145
rect 23290 45135 23370 45145
rect 23610 45135 23690 45145
rect 23930 45135 24010 45145
rect 24250 45135 24330 45145
rect 24570 45135 24650 45145
rect 24890 45135 24970 45145
rect 25210 45135 25290 45145
rect 25530 45135 25610 45145
rect 25850 45135 25930 45145
rect 26170 45135 26250 45145
rect 163750 45135 163830 45145
rect 164070 45135 164150 45145
rect 164390 45135 164470 45145
rect 164710 45135 164790 45145
rect 165030 45135 165110 45145
rect 165350 45135 165430 45145
rect 165670 45135 165750 45145
rect 165990 45135 166070 45145
rect 166310 45135 166390 45145
rect 166630 45135 166710 45145
rect 166950 45135 167030 45145
rect 167270 45135 167350 45145
rect 167590 45135 167670 45145
rect 167910 45135 167990 45145
rect 168230 45135 168310 45145
rect 168550 45135 168630 45145
rect 168870 45135 168950 45145
rect 169190 45135 169270 45145
rect 169510 45135 169590 45145
rect 169830 45135 169910 45145
rect 170150 45135 170230 45145
rect 170470 45135 170550 45145
rect 170790 45135 170870 45145
rect 19210 45055 19220 45135
rect 19530 45055 19540 45135
rect 19850 45055 19860 45135
rect 20170 45055 20180 45135
rect 20490 45055 20500 45135
rect 20810 45055 20820 45135
rect 21130 45055 21140 45135
rect 21450 45055 21460 45135
rect 21770 45055 21780 45135
rect 22090 45055 22100 45135
rect 22410 45055 22420 45135
rect 22730 45055 22740 45135
rect 23050 45055 23060 45135
rect 23370 45055 23380 45135
rect 23690 45055 23700 45135
rect 24010 45055 24020 45135
rect 24330 45055 24340 45135
rect 24650 45055 24660 45135
rect 24970 45055 24980 45135
rect 25290 45055 25300 45135
rect 25610 45055 25620 45135
rect 25930 45055 25940 45135
rect 26250 45055 26260 45135
rect 30520 45095 30600 45105
rect 30840 45095 30920 45105
rect 31160 45095 31240 45105
rect 31480 45095 31560 45105
rect 31800 45095 31880 45105
rect 32120 45095 32200 45105
rect 32440 45095 32520 45105
rect 32760 45095 32840 45105
rect 33080 45095 33160 45105
rect 33400 45095 33480 45105
rect 33720 45095 33800 45105
rect 34040 45095 34120 45105
rect 34360 45095 34440 45105
rect 34680 45095 34760 45105
rect 35000 45095 35080 45105
rect 35320 45095 35400 45105
rect 35640 45095 35720 45105
rect 35960 45095 36040 45105
rect 36280 45095 36360 45105
rect 36600 45095 36680 45105
rect 36920 45095 37000 45105
rect 37240 45095 37320 45105
rect 37560 45095 37640 45105
rect 40340 45095 40420 45105
rect 40660 45095 40740 45105
rect 40980 45095 41060 45105
rect 42720 45095 42800 45105
rect 43040 45095 43120 45105
rect 43360 45095 43440 45105
rect 146560 45095 146640 45105
rect 146880 45095 146960 45105
rect 147200 45095 147280 45105
rect 148940 45095 149020 45105
rect 149260 45095 149340 45105
rect 149580 45095 149660 45105
rect 152360 45095 152440 45105
rect 152680 45095 152760 45105
rect 153000 45095 153080 45105
rect 153320 45095 153400 45105
rect 153640 45095 153720 45105
rect 153960 45095 154040 45105
rect 154280 45095 154360 45105
rect 154600 45095 154680 45105
rect 154920 45095 155000 45105
rect 155240 45095 155320 45105
rect 155560 45095 155640 45105
rect 155880 45095 155960 45105
rect 156200 45095 156280 45105
rect 156520 45095 156600 45105
rect 156840 45095 156920 45105
rect 157160 45095 157240 45105
rect 157480 45095 157560 45105
rect 157800 45095 157880 45105
rect 158120 45095 158200 45105
rect 158440 45095 158520 45105
rect 158760 45095 158840 45105
rect 159080 45095 159160 45105
rect 159400 45095 159480 45105
rect 30600 45015 30610 45095
rect 30920 45015 30930 45095
rect 31240 45015 31250 45095
rect 31560 45015 31570 45095
rect 31880 45015 31890 45095
rect 32200 45015 32210 45095
rect 32520 45015 32530 45095
rect 32840 45015 32850 45095
rect 33160 45015 33170 45095
rect 33480 45015 33490 45095
rect 33800 45015 33810 45095
rect 34120 45015 34130 45095
rect 34440 45015 34450 45095
rect 34760 45015 34770 45095
rect 35080 45015 35090 45095
rect 35400 45015 35410 45095
rect 35720 45015 35730 45095
rect 36040 45015 36050 45095
rect 36360 45015 36370 45095
rect 36680 45015 36690 45095
rect 37000 45015 37010 45095
rect 37320 45015 37330 45095
rect 37640 45015 37650 45095
rect 40420 45015 40430 45095
rect 40740 45015 40750 45095
rect 41060 45015 41070 45095
rect 42800 45015 42810 45095
rect 43120 45015 43130 45095
rect 43440 45015 43450 45095
rect 146640 45015 146650 45095
rect 146960 45015 146970 45095
rect 147280 45015 147290 45095
rect 149020 45015 149030 45095
rect 149340 45015 149350 45095
rect 149660 45015 149670 45095
rect 152440 45015 152450 45095
rect 152760 45015 152770 45095
rect 153080 45015 153090 45095
rect 153400 45015 153410 45095
rect 153720 45015 153730 45095
rect 154040 45015 154050 45095
rect 154360 45015 154370 45095
rect 154680 45015 154690 45095
rect 155000 45015 155010 45095
rect 155320 45015 155330 45095
rect 155640 45015 155650 45095
rect 155960 45015 155970 45095
rect 156280 45015 156290 45095
rect 156600 45015 156610 45095
rect 156920 45015 156930 45095
rect 157240 45015 157250 45095
rect 157560 45015 157570 45095
rect 157880 45015 157890 45095
rect 158200 45015 158210 45095
rect 158520 45015 158530 45095
rect 158840 45015 158850 45095
rect 159160 45015 159170 45095
rect 159480 45015 159490 45095
rect 163830 45055 163840 45135
rect 164150 45055 164160 45135
rect 164470 45055 164480 45135
rect 164790 45055 164800 45135
rect 165110 45055 165120 45135
rect 165430 45055 165440 45135
rect 165750 45055 165760 45135
rect 166070 45055 166080 45135
rect 166390 45055 166400 45135
rect 166710 45055 166720 45135
rect 167030 45055 167040 45135
rect 167350 45055 167360 45135
rect 167670 45055 167680 45135
rect 167990 45055 168000 45135
rect 168310 45055 168320 45135
rect 168630 45055 168640 45135
rect 168950 45055 168960 45135
rect 169270 45055 169280 45135
rect 169590 45055 169600 45135
rect 169910 45055 169920 45135
rect 170230 45055 170240 45135
rect 170550 45055 170560 45135
rect 170870 45055 170880 45135
rect 18970 44975 19050 44985
rect 19290 44975 19370 44985
rect 19610 44975 19690 44985
rect 19930 44975 20010 44985
rect 20250 44975 20330 44985
rect 20570 44975 20650 44985
rect 20890 44975 20970 44985
rect 21210 44975 21290 44985
rect 21530 44975 21610 44985
rect 21850 44975 21930 44985
rect 22170 44975 22250 44985
rect 22490 44975 22570 44985
rect 22810 44975 22890 44985
rect 23130 44975 23210 44985
rect 23450 44975 23530 44985
rect 23770 44975 23850 44985
rect 24090 44975 24170 44985
rect 24410 44975 24490 44985
rect 24730 44975 24810 44985
rect 25050 44975 25130 44985
rect 25370 44975 25450 44985
rect 25690 44975 25770 44985
rect 26010 44975 26090 44985
rect 26330 44975 26410 44985
rect 163590 44975 163670 44985
rect 163910 44975 163990 44985
rect 164230 44975 164310 44985
rect 164550 44975 164630 44985
rect 164870 44975 164950 44985
rect 165190 44975 165270 44985
rect 165510 44975 165590 44985
rect 165830 44975 165910 44985
rect 166150 44975 166230 44985
rect 166470 44975 166550 44985
rect 166790 44975 166870 44985
rect 167110 44975 167190 44985
rect 167430 44975 167510 44985
rect 167750 44975 167830 44985
rect 168070 44975 168150 44985
rect 168390 44975 168470 44985
rect 168710 44975 168790 44985
rect 169030 44975 169110 44985
rect 169350 44975 169430 44985
rect 169670 44975 169750 44985
rect 169990 44975 170070 44985
rect 170310 44975 170390 44985
rect 170630 44975 170710 44985
rect 170950 44975 171030 44985
rect 19050 44895 19060 44975
rect 19370 44895 19380 44975
rect 19690 44895 19700 44975
rect 20010 44895 20020 44975
rect 20330 44895 20340 44975
rect 20650 44895 20660 44975
rect 20970 44895 20980 44975
rect 21290 44895 21300 44975
rect 21610 44895 21620 44975
rect 21930 44895 21940 44975
rect 22250 44895 22260 44975
rect 22570 44895 22580 44975
rect 22890 44895 22900 44975
rect 23210 44895 23220 44975
rect 23530 44895 23540 44975
rect 23850 44895 23860 44975
rect 24170 44895 24180 44975
rect 24490 44895 24500 44975
rect 24810 44895 24820 44975
rect 25130 44895 25140 44975
rect 25450 44895 25460 44975
rect 25770 44895 25780 44975
rect 26090 44895 26100 44975
rect 26410 44895 26420 44975
rect 30360 44935 30440 44945
rect 30680 44935 30760 44945
rect 31000 44935 31080 44945
rect 31320 44935 31400 44945
rect 31640 44935 31720 44945
rect 31960 44935 32040 44945
rect 32280 44935 32360 44945
rect 32600 44935 32680 44945
rect 32920 44935 33000 44945
rect 33240 44935 33320 44945
rect 33560 44935 33640 44945
rect 33880 44935 33960 44945
rect 34200 44935 34280 44945
rect 34520 44935 34600 44945
rect 34840 44935 34920 44945
rect 35160 44935 35240 44945
rect 35480 44935 35560 44945
rect 35800 44935 35880 44945
rect 36120 44935 36200 44945
rect 36440 44935 36520 44945
rect 36760 44935 36840 44945
rect 37080 44935 37160 44945
rect 37400 44935 37480 44945
rect 37720 44935 37800 44945
rect 40180 44935 40260 44945
rect 40500 44935 40580 44945
rect 40820 44935 40900 44945
rect 41140 44935 41220 44945
rect 42560 44935 42640 44945
rect 42880 44935 42960 44945
rect 43200 44935 43280 44945
rect 43520 44935 43600 44945
rect 146400 44935 146480 44945
rect 146720 44935 146800 44945
rect 147040 44935 147120 44945
rect 147360 44935 147440 44945
rect 148780 44935 148860 44945
rect 149100 44935 149180 44945
rect 149420 44935 149500 44945
rect 149740 44935 149820 44945
rect 152200 44935 152280 44945
rect 152520 44935 152600 44945
rect 152840 44935 152920 44945
rect 153160 44935 153240 44945
rect 153480 44935 153560 44945
rect 153800 44935 153880 44945
rect 154120 44935 154200 44945
rect 154440 44935 154520 44945
rect 154760 44935 154840 44945
rect 155080 44935 155160 44945
rect 155400 44935 155480 44945
rect 155720 44935 155800 44945
rect 156040 44935 156120 44945
rect 156360 44935 156440 44945
rect 156680 44935 156760 44945
rect 157000 44935 157080 44945
rect 157320 44935 157400 44945
rect 157640 44935 157720 44945
rect 157960 44935 158040 44945
rect 158280 44935 158360 44945
rect 158600 44935 158680 44945
rect 158920 44935 159000 44945
rect 159240 44935 159320 44945
rect 159560 44935 159640 44945
rect 30440 44855 30450 44935
rect 30760 44855 30770 44935
rect 31080 44855 31090 44935
rect 31400 44855 31410 44935
rect 31720 44855 31730 44935
rect 32040 44855 32050 44935
rect 32360 44855 32370 44935
rect 32680 44855 32690 44935
rect 33000 44855 33010 44935
rect 33320 44855 33330 44935
rect 33640 44855 33650 44935
rect 33960 44855 33970 44935
rect 34280 44855 34290 44935
rect 34600 44855 34610 44935
rect 34920 44855 34930 44935
rect 35240 44855 35250 44935
rect 35560 44855 35570 44935
rect 35880 44855 35890 44935
rect 36200 44855 36210 44935
rect 36520 44855 36530 44935
rect 36840 44855 36850 44935
rect 37160 44855 37170 44935
rect 37480 44855 37490 44935
rect 37800 44855 37810 44935
rect 40260 44855 40270 44935
rect 40580 44855 40590 44935
rect 40900 44855 40910 44935
rect 41220 44855 41230 44935
rect 42640 44855 42650 44935
rect 42960 44855 42970 44935
rect 43280 44855 43290 44935
rect 43600 44855 43610 44935
rect 146480 44855 146490 44935
rect 146800 44855 146810 44935
rect 147120 44855 147130 44935
rect 147440 44855 147450 44935
rect 148860 44855 148870 44935
rect 149180 44855 149190 44935
rect 149500 44855 149510 44935
rect 149820 44855 149830 44935
rect 152280 44855 152290 44935
rect 152600 44855 152610 44935
rect 152920 44855 152930 44935
rect 153240 44855 153250 44935
rect 153560 44855 153570 44935
rect 153880 44855 153890 44935
rect 154200 44855 154210 44935
rect 154520 44855 154530 44935
rect 154840 44855 154850 44935
rect 155160 44855 155170 44935
rect 155480 44855 155490 44935
rect 155800 44855 155810 44935
rect 156120 44855 156130 44935
rect 156440 44855 156450 44935
rect 156760 44855 156770 44935
rect 157080 44855 157090 44935
rect 157400 44855 157410 44935
rect 157720 44855 157730 44935
rect 158040 44855 158050 44935
rect 158360 44855 158370 44935
rect 158680 44855 158690 44935
rect 159000 44855 159010 44935
rect 159320 44855 159330 44935
rect 159640 44855 159650 44935
rect 163670 44895 163680 44975
rect 163990 44895 164000 44975
rect 164310 44895 164320 44975
rect 164630 44895 164640 44975
rect 164950 44895 164960 44975
rect 165270 44895 165280 44975
rect 165590 44895 165600 44975
rect 165910 44895 165920 44975
rect 166230 44895 166240 44975
rect 166550 44895 166560 44975
rect 166870 44895 166880 44975
rect 167190 44895 167200 44975
rect 167510 44895 167520 44975
rect 167830 44895 167840 44975
rect 168150 44895 168160 44975
rect 168470 44895 168480 44975
rect 168790 44895 168800 44975
rect 169110 44895 169120 44975
rect 169430 44895 169440 44975
rect 169750 44895 169760 44975
rect 170070 44895 170080 44975
rect 170390 44895 170400 44975
rect 170710 44895 170720 44975
rect 171030 44895 171040 44975
rect 19130 44815 19210 44825
rect 19450 44815 19530 44825
rect 19770 44815 19850 44825
rect 20090 44815 20170 44825
rect 20410 44815 20490 44825
rect 20730 44815 20810 44825
rect 21050 44815 21130 44825
rect 21370 44815 21450 44825
rect 21690 44815 21770 44825
rect 22010 44815 22090 44825
rect 22330 44815 22410 44825
rect 22650 44815 22730 44825
rect 22970 44815 23050 44825
rect 23290 44815 23370 44825
rect 23610 44815 23690 44825
rect 23930 44815 24010 44825
rect 24250 44815 24330 44825
rect 24570 44815 24650 44825
rect 24890 44815 24970 44825
rect 25210 44815 25290 44825
rect 25530 44815 25610 44825
rect 25850 44815 25930 44825
rect 26170 44815 26250 44825
rect 163750 44815 163830 44825
rect 164070 44815 164150 44825
rect 164390 44815 164470 44825
rect 164710 44815 164790 44825
rect 165030 44815 165110 44825
rect 165350 44815 165430 44825
rect 165670 44815 165750 44825
rect 165990 44815 166070 44825
rect 166310 44815 166390 44825
rect 166630 44815 166710 44825
rect 166950 44815 167030 44825
rect 167270 44815 167350 44825
rect 167590 44815 167670 44825
rect 167910 44815 167990 44825
rect 168230 44815 168310 44825
rect 168550 44815 168630 44825
rect 168870 44815 168950 44825
rect 169190 44815 169270 44825
rect 169510 44815 169590 44825
rect 169830 44815 169910 44825
rect 170150 44815 170230 44825
rect 170470 44815 170550 44825
rect 170790 44815 170870 44825
rect 19210 44735 19220 44815
rect 19530 44735 19540 44815
rect 19850 44735 19860 44815
rect 20170 44735 20180 44815
rect 20490 44735 20500 44815
rect 20810 44735 20820 44815
rect 21130 44735 21140 44815
rect 21450 44735 21460 44815
rect 21770 44735 21780 44815
rect 22090 44735 22100 44815
rect 22410 44735 22420 44815
rect 22730 44735 22740 44815
rect 23050 44735 23060 44815
rect 23370 44735 23380 44815
rect 23690 44735 23700 44815
rect 24010 44735 24020 44815
rect 24330 44735 24340 44815
rect 24650 44735 24660 44815
rect 24970 44735 24980 44815
rect 25290 44735 25300 44815
rect 25610 44735 25620 44815
rect 25930 44735 25940 44815
rect 26250 44735 26260 44815
rect 30520 44775 30600 44785
rect 30840 44775 30920 44785
rect 31160 44775 31240 44785
rect 31480 44775 31560 44785
rect 31800 44775 31880 44785
rect 32120 44775 32200 44785
rect 32440 44775 32520 44785
rect 32760 44775 32840 44785
rect 33080 44775 33160 44785
rect 33400 44775 33480 44785
rect 33720 44775 33800 44785
rect 34040 44775 34120 44785
rect 34360 44775 34440 44785
rect 34680 44775 34760 44785
rect 35000 44775 35080 44785
rect 35320 44775 35400 44785
rect 35640 44775 35720 44785
rect 35960 44775 36040 44785
rect 36280 44775 36360 44785
rect 36600 44775 36680 44785
rect 36920 44775 37000 44785
rect 37240 44775 37320 44785
rect 37560 44775 37640 44785
rect 40340 44775 40420 44785
rect 40660 44775 40740 44785
rect 40980 44775 41060 44785
rect 42720 44775 42800 44785
rect 43040 44775 43120 44785
rect 43360 44775 43440 44785
rect 146560 44775 146640 44785
rect 146880 44775 146960 44785
rect 147200 44775 147280 44785
rect 148940 44775 149020 44785
rect 149260 44775 149340 44785
rect 149580 44775 149660 44785
rect 152360 44775 152440 44785
rect 152680 44775 152760 44785
rect 153000 44775 153080 44785
rect 153320 44775 153400 44785
rect 153640 44775 153720 44785
rect 153960 44775 154040 44785
rect 154280 44775 154360 44785
rect 154600 44775 154680 44785
rect 154920 44775 155000 44785
rect 155240 44775 155320 44785
rect 155560 44775 155640 44785
rect 155880 44775 155960 44785
rect 156200 44775 156280 44785
rect 156520 44775 156600 44785
rect 156840 44775 156920 44785
rect 157160 44775 157240 44785
rect 157480 44775 157560 44785
rect 157800 44775 157880 44785
rect 158120 44775 158200 44785
rect 158440 44775 158520 44785
rect 158760 44775 158840 44785
rect 159080 44775 159160 44785
rect 159400 44775 159480 44785
rect 30600 44695 30610 44775
rect 30920 44695 30930 44775
rect 31240 44695 31250 44775
rect 31560 44695 31570 44775
rect 31880 44695 31890 44775
rect 32200 44695 32210 44775
rect 32520 44695 32530 44775
rect 32840 44695 32850 44775
rect 33160 44695 33170 44775
rect 33480 44695 33490 44775
rect 33800 44695 33810 44775
rect 34120 44695 34130 44775
rect 34440 44695 34450 44775
rect 34760 44695 34770 44775
rect 35080 44695 35090 44775
rect 35400 44695 35410 44775
rect 35720 44695 35730 44775
rect 36040 44695 36050 44775
rect 36360 44695 36370 44775
rect 36680 44695 36690 44775
rect 37000 44695 37010 44775
rect 37320 44695 37330 44775
rect 37640 44695 37650 44775
rect 40420 44695 40430 44775
rect 40740 44695 40750 44775
rect 41060 44695 41070 44775
rect 42800 44695 42810 44775
rect 43120 44695 43130 44775
rect 43440 44695 43450 44775
rect 146640 44695 146650 44775
rect 146960 44695 146970 44775
rect 147280 44695 147290 44775
rect 149020 44695 149030 44775
rect 149340 44695 149350 44775
rect 149660 44695 149670 44775
rect 152440 44695 152450 44775
rect 152760 44695 152770 44775
rect 153080 44695 153090 44775
rect 153400 44695 153410 44775
rect 153720 44695 153730 44775
rect 154040 44695 154050 44775
rect 154360 44695 154370 44775
rect 154680 44695 154690 44775
rect 155000 44695 155010 44775
rect 155320 44695 155330 44775
rect 155640 44695 155650 44775
rect 155960 44695 155970 44775
rect 156280 44695 156290 44775
rect 156600 44695 156610 44775
rect 156920 44695 156930 44775
rect 157240 44695 157250 44775
rect 157560 44695 157570 44775
rect 157880 44695 157890 44775
rect 158200 44695 158210 44775
rect 158520 44695 158530 44775
rect 158840 44695 158850 44775
rect 159160 44695 159170 44775
rect 159480 44695 159490 44775
rect 163830 44735 163840 44815
rect 164150 44735 164160 44815
rect 164470 44735 164480 44815
rect 164790 44735 164800 44815
rect 165110 44735 165120 44815
rect 165430 44735 165440 44815
rect 165750 44735 165760 44815
rect 166070 44735 166080 44815
rect 166390 44735 166400 44815
rect 166710 44735 166720 44815
rect 167030 44735 167040 44815
rect 167350 44735 167360 44815
rect 167670 44735 167680 44815
rect 167990 44735 168000 44815
rect 168310 44735 168320 44815
rect 168630 44735 168640 44815
rect 168950 44735 168960 44815
rect 169270 44735 169280 44815
rect 169590 44735 169600 44815
rect 169910 44735 169920 44815
rect 170230 44735 170240 44815
rect 170550 44735 170560 44815
rect 170870 44735 170880 44815
rect 18970 44655 19050 44665
rect 19290 44655 19370 44665
rect 19610 44655 19690 44665
rect 19930 44655 20010 44665
rect 20250 44655 20330 44665
rect 20570 44655 20650 44665
rect 20890 44655 20970 44665
rect 21210 44655 21290 44665
rect 21530 44655 21610 44665
rect 21850 44655 21930 44665
rect 22170 44655 22250 44665
rect 22490 44655 22570 44665
rect 22810 44655 22890 44665
rect 23130 44655 23210 44665
rect 23450 44655 23530 44665
rect 23770 44655 23850 44665
rect 24090 44655 24170 44665
rect 24410 44655 24490 44665
rect 24730 44655 24810 44665
rect 25050 44655 25130 44665
rect 25370 44655 25450 44665
rect 25690 44655 25770 44665
rect 26010 44655 26090 44665
rect 26330 44655 26410 44665
rect 163590 44655 163670 44665
rect 163910 44655 163990 44665
rect 164230 44655 164310 44665
rect 164550 44655 164630 44665
rect 164870 44655 164950 44665
rect 165190 44655 165270 44665
rect 165510 44655 165590 44665
rect 165830 44655 165910 44665
rect 166150 44655 166230 44665
rect 166470 44655 166550 44665
rect 166790 44655 166870 44665
rect 167110 44655 167190 44665
rect 167430 44655 167510 44665
rect 167750 44655 167830 44665
rect 168070 44655 168150 44665
rect 168390 44655 168470 44665
rect 168710 44655 168790 44665
rect 169030 44655 169110 44665
rect 169350 44655 169430 44665
rect 169670 44655 169750 44665
rect 169990 44655 170070 44665
rect 170310 44655 170390 44665
rect 170630 44655 170710 44665
rect 170950 44655 171030 44665
rect 19050 44575 19060 44655
rect 19370 44575 19380 44655
rect 19690 44575 19700 44655
rect 20010 44575 20020 44655
rect 20330 44575 20340 44655
rect 20650 44575 20660 44655
rect 20970 44575 20980 44655
rect 21290 44575 21300 44655
rect 21610 44575 21620 44655
rect 21930 44575 21940 44655
rect 22250 44575 22260 44655
rect 22570 44575 22580 44655
rect 22890 44575 22900 44655
rect 23210 44575 23220 44655
rect 23530 44575 23540 44655
rect 23850 44575 23860 44655
rect 24170 44575 24180 44655
rect 24490 44575 24500 44655
rect 24810 44575 24820 44655
rect 25130 44575 25140 44655
rect 25450 44575 25460 44655
rect 25770 44575 25780 44655
rect 26090 44575 26100 44655
rect 26410 44575 26420 44655
rect 30360 44615 30440 44625
rect 30680 44615 30760 44625
rect 31000 44615 31080 44625
rect 31320 44615 31400 44625
rect 31640 44615 31720 44625
rect 31960 44615 32040 44625
rect 32280 44615 32360 44625
rect 32600 44615 32680 44625
rect 32920 44615 33000 44625
rect 33240 44615 33320 44625
rect 33560 44615 33640 44625
rect 33880 44615 33960 44625
rect 34200 44615 34280 44625
rect 34520 44615 34600 44625
rect 34840 44615 34920 44625
rect 35160 44615 35240 44625
rect 35480 44615 35560 44625
rect 35800 44615 35880 44625
rect 36120 44615 36200 44625
rect 36440 44615 36520 44625
rect 36760 44615 36840 44625
rect 37080 44615 37160 44625
rect 37400 44615 37480 44625
rect 37720 44615 37800 44625
rect 40180 44615 40260 44625
rect 40500 44615 40580 44625
rect 40820 44615 40900 44625
rect 41140 44615 41220 44625
rect 42560 44615 42640 44625
rect 42880 44615 42960 44625
rect 43200 44615 43280 44625
rect 43520 44615 43600 44625
rect 146400 44615 146480 44625
rect 146720 44615 146800 44625
rect 147040 44615 147120 44625
rect 147360 44615 147440 44625
rect 148780 44615 148860 44625
rect 149100 44615 149180 44625
rect 149420 44615 149500 44625
rect 149740 44615 149820 44625
rect 152200 44615 152280 44625
rect 152520 44615 152600 44625
rect 152840 44615 152920 44625
rect 153160 44615 153240 44625
rect 153480 44615 153560 44625
rect 153800 44615 153880 44625
rect 154120 44615 154200 44625
rect 154440 44615 154520 44625
rect 154760 44615 154840 44625
rect 155080 44615 155160 44625
rect 155400 44615 155480 44625
rect 155720 44615 155800 44625
rect 156040 44615 156120 44625
rect 156360 44615 156440 44625
rect 156680 44615 156760 44625
rect 157000 44615 157080 44625
rect 157320 44615 157400 44625
rect 157640 44615 157720 44625
rect 157960 44615 158040 44625
rect 158280 44615 158360 44625
rect 158600 44615 158680 44625
rect 158920 44615 159000 44625
rect 159240 44615 159320 44625
rect 159560 44615 159640 44625
rect 30440 44535 30450 44615
rect 30760 44535 30770 44615
rect 31080 44535 31090 44615
rect 31400 44535 31410 44615
rect 31720 44535 31730 44615
rect 32040 44535 32050 44615
rect 32360 44535 32370 44615
rect 32680 44535 32690 44615
rect 33000 44535 33010 44615
rect 33320 44535 33330 44615
rect 33640 44535 33650 44615
rect 33960 44535 33970 44615
rect 34280 44535 34290 44615
rect 34600 44535 34610 44615
rect 34920 44535 34930 44615
rect 35240 44535 35250 44615
rect 35560 44535 35570 44615
rect 35880 44535 35890 44615
rect 36200 44535 36210 44615
rect 36520 44535 36530 44615
rect 36840 44535 36850 44615
rect 37160 44535 37170 44615
rect 37480 44535 37490 44615
rect 37800 44535 37810 44615
rect 40260 44535 40270 44615
rect 40580 44535 40590 44615
rect 40900 44535 40910 44615
rect 41220 44535 41230 44615
rect 42640 44535 42650 44615
rect 42960 44535 42970 44615
rect 43280 44535 43290 44615
rect 43600 44535 43610 44615
rect 146480 44535 146490 44615
rect 146800 44535 146810 44615
rect 147120 44535 147130 44615
rect 147440 44535 147450 44615
rect 148860 44535 148870 44615
rect 149180 44535 149190 44615
rect 149500 44535 149510 44615
rect 149820 44535 149830 44615
rect 152280 44535 152290 44615
rect 152600 44535 152610 44615
rect 152920 44535 152930 44615
rect 153240 44535 153250 44615
rect 153560 44535 153570 44615
rect 153880 44535 153890 44615
rect 154200 44535 154210 44615
rect 154520 44535 154530 44615
rect 154840 44535 154850 44615
rect 155160 44535 155170 44615
rect 155480 44535 155490 44615
rect 155800 44535 155810 44615
rect 156120 44535 156130 44615
rect 156440 44535 156450 44615
rect 156760 44535 156770 44615
rect 157080 44535 157090 44615
rect 157400 44535 157410 44615
rect 157720 44535 157730 44615
rect 158040 44535 158050 44615
rect 158360 44535 158370 44615
rect 158680 44535 158690 44615
rect 159000 44535 159010 44615
rect 159320 44535 159330 44615
rect 159640 44535 159650 44615
rect 163670 44575 163680 44655
rect 163990 44575 164000 44655
rect 164310 44575 164320 44655
rect 164630 44575 164640 44655
rect 164950 44575 164960 44655
rect 165270 44575 165280 44655
rect 165590 44575 165600 44655
rect 165910 44575 165920 44655
rect 166230 44575 166240 44655
rect 166550 44575 166560 44655
rect 166870 44575 166880 44655
rect 167190 44575 167200 44655
rect 167510 44575 167520 44655
rect 167830 44575 167840 44655
rect 168150 44575 168160 44655
rect 168470 44575 168480 44655
rect 168790 44575 168800 44655
rect 169110 44575 169120 44655
rect 169430 44575 169440 44655
rect 169750 44575 169760 44655
rect 170070 44575 170080 44655
rect 170390 44575 170400 44655
rect 170710 44575 170720 44655
rect 171030 44575 171040 44655
rect 19130 44495 19210 44505
rect 19450 44495 19530 44505
rect 19770 44495 19850 44505
rect 20090 44495 20170 44505
rect 20410 44495 20490 44505
rect 20730 44495 20810 44505
rect 21050 44495 21130 44505
rect 21370 44495 21450 44505
rect 21690 44495 21770 44505
rect 22010 44495 22090 44505
rect 22330 44495 22410 44505
rect 22650 44495 22730 44505
rect 22970 44495 23050 44505
rect 23290 44495 23370 44505
rect 23610 44495 23690 44505
rect 23930 44495 24010 44505
rect 24250 44495 24330 44505
rect 24570 44495 24650 44505
rect 24890 44495 24970 44505
rect 25210 44495 25290 44505
rect 25530 44495 25610 44505
rect 25850 44495 25930 44505
rect 26170 44495 26250 44505
rect 163750 44495 163830 44505
rect 164070 44495 164150 44505
rect 164390 44495 164470 44505
rect 164710 44495 164790 44505
rect 165030 44495 165110 44505
rect 165350 44495 165430 44505
rect 165670 44495 165750 44505
rect 165990 44495 166070 44505
rect 166310 44495 166390 44505
rect 166630 44495 166710 44505
rect 166950 44495 167030 44505
rect 167270 44495 167350 44505
rect 167590 44495 167670 44505
rect 167910 44495 167990 44505
rect 168230 44495 168310 44505
rect 168550 44495 168630 44505
rect 168870 44495 168950 44505
rect 169190 44495 169270 44505
rect 169510 44495 169590 44505
rect 169830 44495 169910 44505
rect 170150 44495 170230 44505
rect 170470 44495 170550 44505
rect 170790 44495 170870 44505
rect 19210 44415 19220 44495
rect 19530 44415 19540 44495
rect 19850 44415 19860 44495
rect 20170 44415 20180 44495
rect 20490 44415 20500 44495
rect 20810 44415 20820 44495
rect 21130 44415 21140 44495
rect 21450 44415 21460 44495
rect 21770 44415 21780 44495
rect 22090 44415 22100 44495
rect 22410 44415 22420 44495
rect 22730 44415 22740 44495
rect 23050 44415 23060 44495
rect 23370 44415 23380 44495
rect 23690 44415 23700 44495
rect 24010 44415 24020 44495
rect 24330 44415 24340 44495
rect 24650 44415 24660 44495
rect 24970 44415 24980 44495
rect 25290 44415 25300 44495
rect 25610 44415 25620 44495
rect 25930 44415 25940 44495
rect 26250 44415 26260 44495
rect 30520 44455 30600 44465
rect 30840 44455 30920 44465
rect 31160 44455 31240 44465
rect 31480 44455 31560 44465
rect 31800 44455 31880 44465
rect 32120 44455 32200 44465
rect 32440 44455 32520 44465
rect 32760 44455 32840 44465
rect 33080 44455 33160 44465
rect 33400 44455 33480 44465
rect 33720 44455 33800 44465
rect 34040 44455 34120 44465
rect 34360 44455 34440 44465
rect 34680 44455 34760 44465
rect 35000 44455 35080 44465
rect 35320 44455 35400 44465
rect 35640 44455 35720 44465
rect 35960 44455 36040 44465
rect 36280 44455 36360 44465
rect 36600 44455 36680 44465
rect 36920 44455 37000 44465
rect 37240 44455 37320 44465
rect 37560 44455 37640 44465
rect 40340 44455 40420 44465
rect 40660 44455 40740 44465
rect 40980 44455 41060 44465
rect 42720 44455 42800 44465
rect 43040 44455 43120 44465
rect 43360 44455 43440 44465
rect 146560 44455 146640 44465
rect 146880 44455 146960 44465
rect 147200 44455 147280 44465
rect 148940 44455 149020 44465
rect 149260 44455 149340 44465
rect 149580 44455 149660 44465
rect 152360 44455 152440 44465
rect 152680 44455 152760 44465
rect 153000 44455 153080 44465
rect 153320 44455 153400 44465
rect 153640 44455 153720 44465
rect 153960 44455 154040 44465
rect 154280 44455 154360 44465
rect 154600 44455 154680 44465
rect 154920 44455 155000 44465
rect 155240 44455 155320 44465
rect 155560 44455 155640 44465
rect 155880 44455 155960 44465
rect 156200 44455 156280 44465
rect 156520 44455 156600 44465
rect 156840 44455 156920 44465
rect 157160 44455 157240 44465
rect 157480 44455 157560 44465
rect 157800 44455 157880 44465
rect 158120 44455 158200 44465
rect 158440 44455 158520 44465
rect 158760 44455 158840 44465
rect 159080 44455 159160 44465
rect 159400 44455 159480 44465
rect 30600 44375 30610 44455
rect 30920 44375 30930 44455
rect 31240 44375 31250 44455
rect 31560 44375 31570 44455
rect 31880 44375 31890 44455
rect 32200 44375 32210 44455
rect 32520 44375 32530 44455
rect 32840 44375 32850 44455
rect 33160 44375 33170 44455
rect 33480 44375 33490 44455
rect 33800 44375 33810 44455
rect 34120 44375 34130 44455
rect 34440 44375 34450 44455
rect 34760 44375 34770 44455
rect 35080 44375 35090 44455
rect 35400 44375 35410 44455
rect 35720 44375 35730 44455
rect 36040 44375 36050 44455
rect 36360 44375 36370 44455
rect 36680 44375 36690 44455
rect 37000 44375 37010 44455
rect 37320 44375 37330 44455
rect 37640 44375 37650 44455
rect 40420 44375 40430 44455
rect 40740 44375 40750 44455
rect 41060 44375 41070 44455
rect 42800 44375 42810 44455
rect 43120 44375 43130 44455
rect 43440 44375 43450 44455
rect 146640 44375 146650 44455
rect 146960 44375 146970 44455
rect 147280 44375 147290 44455
rect 149020 44375 149030 44455
rect 149340 44375 149350 44455
rect 149660 44375 149670 44455
rect 152440 44375 152450 44455
rect 152760 44375 152770 44455
rect 153080 44375 153090 44455
rect 153400 44375 153410 44455
rect 153720 44375 153730 44455
rect 154040 44375 154050 44455
rect 154360 44375 154370 44455
rect 154680 44375 154690 44455
rect 155000 44375 155010 44455
rect 155320 44375 155330 44455
rect 155640 44375 155650 44455
rect 155960 44375 155970 44455
rect 156280 44375 156290 44455
rect 156600 44375 156610 44455
rect 156920 44375 156930 44455
rect 157240 44375 157250 44455
rect 157560 44375 157570 44455
rect 157880 44375 157890 44455
rect 158200 44375 158210 44455
rect 158520 44375 158530 44455
rect 158840 44375 158850 44455
rect 159160 44375 159170 44455
rect 159480 44375 159490 44455
rect 163830 44415 163840 44495
rect 164150 44415 164160 44495
rect 164470 44415 164480 44495
rect 164790 44415 164800 44495
rect 165110 44415 165120 44495
rect 165430 44415 165440 44495
rect 165750 44415 165760 44495
rect 166070 44415 166080 44495
rect 166390 44415 166400 44495
rect 166710 44415 166720 44495
rect 167030 44415 167040 44495
rect 167350 44415 167360 44495
rect 167670 44415 167680 44495
rect 167990 44415 168000 44495
rect 168310 44415 168320 44495
rect 168630 44415 168640 44495
rect 168950 44415 168960 44495
rect 169270 44415 169280 44495
rect 169590 44415 169600 44495
rect 169910 44415 169920 44495
rect 170230 44415 170240 44495
rect 170550 44415 170560 44495
rect 170870 44415 170880 44495
rect 18970 44335 19050 44345
rect 19290 44335 19370 44345
rect 19610 44335 19690 44345
rect 19930 44335 20010 44345
rect 20250 44335 20330 44345
rect 20570 44335 20650 44345
rect 20890 44335 20970 44345
rect 21210 44335 21290 44345
rect 21530 44335 21610 44345
rect 21850 44335 21930 44345
rect 22170 44335 22250 44345
rect 22490 44335 22570 44345
rect 22810 44335 22890 44345
rect 23130 44335 23210 44345
rect 23450 44335 23530 44345
rect 23770 44335 23850 44345
rect 24090 44335 24170 44345
rect 24410 44335 24490 44345
rect 24730 44335 24810 44345
rect 25050 44335 25130 44345
rect 25370 44335 25450 44345
rect 25690 44335 25770 44345
rect 26010 44335 26090 44345
rect 26330 44335 26410 44345
rect 163590 44335 163670 44345
rect 163910 44335 163990 44345
rect 164230 44335 164310 44345
rect 164550 44335 164630 44345
rect 164870 44335 164950 44345
rect 165190 44335 165270 44345
rect 165510 44335 165590 44345
rect 165830 44335 165910 44345
rect 166150 44335 166230 44345
rect 166470 44335 166550 44345
rect 166790 44335 166870 44345
rect 167110 44335 167190 44345
rect 167430 44335 167510 44345
rect 167750 44335 167830 44345
rect 168070 44335 168150 44345
rect 168390 44335 168470 44345
rect 168710 44335 168790 44345
rect 169030 44335 169110 44345
rect 169350 44335 169430 44345
rect 169670 44335 169750 44345
rect 169990 44335 170070 44345
rect 170310 44335 170390 44345
rect 170630 44335 170710 44345
rect 170950 44335 171030 44345
rect 19050 44255 19060 44335
rect 19370 44255 19380 44335
rect 19690 44255 19700 44335
rect 20010 44255 20020 44335
rect 20330 44255 20340 44335
rect 20650 44255 20660 44335
rect 20970 44255 20980 44335
rect 21290 44255 21300 44335
rect 21610 44255 21620 44335
rect 21930 44255 21940 44335
rect 22250 44255 22260 44335
rect 22570 44255 22580 44335
rect 22890 44255 22900 44335
rect 23210 44255 23220 44335
rect 23530 44255 23540 44335
rect 23850 44255 23860 44335
rect 24170 44255 24180 44335
rect 24490 44255 24500 44335
rect 24810 44255 24820 44335
rect 25130 44255 25140 44335
rect 25450 44255 25460 44335
rect 25770 44255 25780 44335
rect 26090 44255 26100 44335
rect 26410 44255 26420 44335
rect 30360 44295 30440 44305
rect 30680 44295 30760 44305
rect 31000 44295 31080 44305
rect 31320 44295 31400 44305
rect 31640 44295 31720 44305
rect 31960 44295 32040 44305
rect 32280 44295 32360 44305
rect 32600 44295 32680 44305
rect 32920 44295 33000 44305
rect 33240 44295 33320 44305
rect 33560 44295 33640 44305
rect 33880 44295 33960 44305
rect 34200 44295 34280 44305
rect 34520 44295 34600 44305
rect 34840 44295 34920 44305
rect 35160 44295 35240 44305
rect 35480 44295 35560 44305
rect 35800 44295 35880 44305
rect 36120 44295 36200 44305
rect 36440 44295 36520 44305
rect 36760 44295 36840 44305
rect 37080 44295 37160 44305
rect 37400 44295 37480 44305
rect 37720 44295 37800 44305
rect 40180 44295 40260 44305
rect 40500 44295 40580 44305
rect 40820 44295 40900 44305
rect 41140 44295 41220 44305
rect 42560 44295 42640 44305
rect 42880 44295 42960 44305
rect 43200 44295 43280 44305
rect 43520 44295 43600 44305
rect 146400 44295 146480 44305
rect 146720 44295 146800 44305
rect 147040 44295 147120 44305
rect 147360 44295 147440 44305
rect 148780 44295 148860 44305
rect 149100 44295 149180 44305
rect 149420 44295 149500 44305
rect 149740 44295 149820 44305
rect 152200 44295 152280 44305
rect 152520 44295 152600 44305
rect 152840 44295 152920 44305
rect 153160 44295 153240 44305
rect 153480 44295 153560 44305
rect 153800 44295 153880 44305
rect 154120 44295 154200 44305
rect 154440 44295 154520 44305
rect 154760 44295 154840 44305
rect 155080 44295 155160 44305
rect 155400 44295 155480 44305
rect 155720 44295 155800 44305
rect 156040 44295 156120 44305
rect 156360 44295 156440 44305
rect 156680 44295 156760 44305
rect 157000 44295 157080 44305
rect 157320 44295 157400 44305
rect 157640 44295 157720 44305
rect 157960 44295 158040 44305
rect 158280 44295 158360 44305
rect 158600 44295 158680 44305
rect 158920 44295 159000 44305
rect 159240 44295 159320 44305
rect 159560 44295 159640 44305
rect 30440 44215 30450 44295
rect 30760 44215 30770 44295
rect 31080 44215 31090 44295
rect 31400 44215 31410 44295
rect 31720 44215 31730 44295
rect 32040 44215 32050 44295
rect 32360 44215 32370 44295
rect 32680 44215 32690 44295
rect 33000 44215 33010 44295
rect 33320 44215 33330 44295
rect 33640 44215 33650 44295
rect 33960 44215 33970 44295
rect 34280 44215 34290 44295
rect 34600 44215 34610 44295
rect 34920 44215 34930 44295
rect 35240 44215 35250 44295
rect 35560 44215 35570 44295
rect 35880 44215 35890 44295
rect 36200 44215 36210 44295
rect 36520 44215 36530 44295
rect 36840 44215 36850 44295
rect 37160 44215 37170 44295
rect 37480 44215 37490 44295
rect 37800 44215 37810 44295
rect 40260 44215 40270 44295
rect 40580 44215 40590 44295
rect 40900 44215 40910 44295
rect 41220 44215 41230 44295
rect 42640 44215 42650 44295
rect 42960 44215 42970 44295
rect 43280 44215 43290 44295
rect 43600 44215 43610 44295
rect 146480 44215 146490 44295
rect 146800 44215 146810 44295
rect 147120 44215 147130 44295
rect 147440 44215 147450 44295
rect 148860 44215 148870 44295
rect 149180 44215 149190 44295
rect 149500 44215 149510 44295
rect 149820 44215 149830 44295
rect 152280 44215 152290 44295
rect 152600 44215 152610 44295
rect 152920 44215 152930 44295
rect 153240 44215 153250 44295
rect 153560 44215 153570 44295
rect 153880 44215 153890 44295
rect 154200 44215 154210 44295
rect 154520 44215 154530 44295
rect 154840 44215 154850 44295
rect 155160 44215 155170 44295
rect 155480 44215 155490 44295
rect 155800 44215 155810 44295
rect 156120 44215 156130 44295
rect 156440 44215 156450 44295
rect 156760 44215 156770 44295
rect 157080 44215 157090 44295
rect 157400 44215 157410 44295
rect 157720 44215 157730 44295
rect 158040 44215 158050 44295
rect 158360 44215 158370 44295
rect 158680 44215 158690 44295
rect 159000 44215 159010 44295
rect 159320 44215 159330 44295
rect 159640 44215 159650 44295
rect 163670 44255 163680 44335
rect 163990 44255 164000 44335
rect 164310 44255 164320 44335
rect 164630 44255 164640 44335
rect 164950 44255 164960 44335
rect 165270 44255 165280 44335
rect 165590 44255 165600 44335
rect 165910 44255 165920 44335
rect 166230 44255 166240 44335
rect 166550 44255 166560 44335
rect 166870 44255 166880 44335
rect 167190 44255 167200 44335
rect 167510 44255 167520 44335
rect 167830 44255 167840 44335
rect 168150 44255 168160 44335
rect 168470 44255 168480 44335
rect 168790 44255 168800 44335
rect 169110 44255 169120 44335
rect 169430 44255 169440 44335
rect 169750 44255 169760 44335
rect 170070 44255 170080 44335
rect 170390 44255 170400 44335
rect 170710 44255 170720 44335
rect 171030 44255 171040 44335
rect 19130 44175 19210 44185
rect 19450 44175 19530 44185
rect 19770 44175 19850 44185
rect 20090 44175 20170 44185
rect 20410 44175 20490 44185
rect 20730 44175 20810 44185
rect 21050 44175 21130 44185
rect 21370 44175 21450 44185
rect 21690 44175 21770 44185
rect 22010 44175 22090 44185
rect 22330 44175 22410 44185
rect 22650 44175 22730 44185
rect 22970 44175 23050 44185
rect 23290 44175 23370 44185
rect 23610 44175 23690 44185
rect 23930 44175 24010 44185
rect 24250 44175 24330 44185
rect 24570 44175 24650 44185
rect 24890 44175 24970 44185
rect 25210 44175 25290 44185
rect 25530 44175 25610 44185
rect 25850 44175 25930 44185
rect 26170 44175 26250 44185
rect 163750 44175 163830 44185
rect 164070 44175 164150 44185
rect 164390 44175 164470 44185
rect 164710 44175 164790 44185
rect 165030 44175 165110 44185
rect 165350 44175 165430 44185
rect 165670 44175 165750 44185
rect 165990 44175 166070 44185
rect 166310 44175 166390 44185
rect 166630 44175 166710 44185
rect 166950 44175 167030 44185
rect 167270 44175 167350 44185
rect 167590 44175 167670 44185
rect 167910 44175 167990 44185
rect 168230 44175 168310 44185
rect 168550 44175 168630 44185
rect 168870 44175 168950 44185
rect 169190 44175 169270 44185
rect 169510 44175 169590 44185
rect 169830 44175 169910 44185
rect 170150 44175 170230 44185
rect 170470 44175 170550 44185
rect 170790 44175 170870 44185
rect 19210 44095 19220 44175
rect 19530 44095 19540 44175
rect 19850 44095 19860 44175
rect 20170 44095 20180 44175
rect 20490 44095 20500 44175
rect 20810 44095 20820 44175
rect 21130 44095 21140 44175
rect 21450 44095 21460 44175
rect 21770 44095 21780 44175
rect 22090 44095 22100 44175
rect 22410 44095 22420 44175
rect 22730 44095 22740 44175
rect 23050 44095 23060 44175
rect 23370 44095 23380 44175
rect 23690 44095 23700 44175
rect 24010 44095 24020 44175
rect 24330 44095 24340 44175
rect 24650 44095 24660 44175
rect 24970 44095 24980 44175
rect 25290 44095 25300 44175
rect 25610 44095 25620 44175
rect 25930 44095 25940 44175
rect 26250 44095 26260 44175
rect 30520 44135 30600 44145
rect 30840 44135 30920 44145
rect 31160 44135 31240 44145
rect 31480 44135 31560 44145
rect 31800 44135 31880 44145
rect 32120 44135 32200 44145
rect 32440 44135 32520 44145
rect 32760 44135 32840 44145
rect 33080 44135 33160 44145
rect 33400 44135 33480 44145
rect 33720 44135 33800 44145
rect 34040 44135 34120 44145
rect 34360 44135 34440 44145
rect 34680 44135 34760 44145
rect 35000 44135 35080 44145
rect 35320 44135 35400 44145
rect 35640 44135 35720 44145
rect 35960 44135 36040 44145
rect 36280 44135 36360 44145
rect 36600 44135 36680 44145
rect 36920 44135 37000 44145
rect 37240 44135 37320 44145
rect 37560 44135 37640 44145
rect 40340 44135 40420 44145
rect 40660 44135 40740 44145
rect 40980 44135 41060 44145
rect 42720 44135 42800 44145
rect 43040 44135 43120 44145
rect 43360 44135 43440 44145
rect 146560 44135 146640 44145
rect 146880 44135 146960 44145
rect 147200 44135 147280 44145
rect 148940 44135 149020 44145
rect 149260 44135 149340 44145
rect 149580 44135 149660 44145
rect 152360 44135 152440 44145
rect 152680 44135 152760 44145
rect 153000 44135 153080 44145
rect 153320 44135 153400 44145
rect 153640 44135 153720 44145
rect 153960 44135 154040 44145
rect 154280 44135 154360 44145
rect 154600 44135 154680 44145
rect 154920 44135 155000 44145
rect 155240 44135 155320 44145
rect 155560 44135 155640 44145
rect 155880 44135 155960 44145
rect 156200 44135 156280 44145
rect 156520 44135 156600 44145
rect 156840 44135 156920 44145
rect 157160 44135 157240 44145
rect 157480 44135 157560 44145
rect 157800 44135 157880 44145
rect 158120 44135 158200 44145
rect 158440 44135 158520 44145
rect 158760 44135 158840 44145
rect 159080 44135 159160 44145
rect 159400 44135 159480 44145
rect 30600 44055 30610 44135
rect 30920 44055 30930 44135
rect 31240 44055 31250 44135
rect 31560 44055 31570 44135
rect 31880 44055 31890 44135
rect 32200 44055 32210 44135
rect 32520 44055 32530 44135
rect 32840 44055 32850 44135
rect 33160 44055 33170 44135
rect 33480 44055 33490 44135
rect 33800 44055 33810 44135
rect 34120 44055 34130 44135
rect 34440 44055 34450 44135
rect 34760 44055 34770 44135
rect 35080 44055 35090 44135
rect 35400 44055 35410 44135
rect 35720 44055 35730 44135
rect 36040 44055 36050 44135
rect 36360 44055 36370 44135
rect 36680 44055 36690 44135
rect 37000 44055 37010 44135
rect 37320 44055 37330 44135
rect 37640 44055 37650 44135
rect 40420 44055 40430 44135
rect 40740 44055 40750 44135
rect 41060 44055 41070 44135
rect 42800 44055 42810 44135
rect 43120 44055 43130 44135
rect 43440 44055 43450 44135
rect 146640 44055 146650 44135
rect 146960 44055 146970 44135
rect 147280 44055 147290 44135
rect 149020 44055 149030 44135
rect 149340 44055 149350 44135
rect 149660 44055 149670 44135
rect 152440 44055 152450 44135
rect 152760 44055 152770 44135
rect 153080 44055 153090 44135
rect 153400 44055 153410 44135
rect 153720 44055 153730 44135
rect 154040 44055 154050 44135
rect 154360 44055 154370 44135
rect 154680 44055 154690 44135
rect 155000 44055 155010 44135
rect 155320 44055 155330 44135
rect 155640 44055 155650 44135
rect 155960 44055 155970 44135
rect 156280 44055 156290 44135
rect 156600 44055 156610 44135
rect 156920 44055 156930 44135
rect 157240 44055 157250 44135
rect 157560 44055 157570 44135
rect 157880 44055 157890 44135
rect 158200 44055 158210 44135
rect 158520 44055 158530 44135
rect 158840 44055 158850 44135
rect 159160 44055 159170 44135
rect 159480 44055 159490 44135
rect 163830 44095 163840 44175
rect 164150 44095 164160 44175
rect 164470 44095 164480 44175
rect 164790 44095 164800 44175
rect 165110 44095 165120 44175
rect 165430 44095 165440 44175
rect 165750 44095 165760 44175
rect 166070 44095 166080 44175
rect 166390 44095 166400 44175
rect 166710 44095 166720 44175
rect 167030 44095 167040 44175
rect 167350 44095 167360 44175
rect 167670 44095 167680 44175
rect 167990 44095 168000 44175
rect 168310 44095 168320 44175
rect 168630 44095 168640 44175
rect 168950 44095 168960 44175
rect 169270 44095 169280 44175
rect 169590 44095 169600 44175
rect 169910 44095 169920 44175
rect 170230 44095 170240 44175
rect 170550 44095 170560 44175
rect 170870 44095 170880 44175
rect 18970 44015 19050 44025
rect 19290 44015 19370 44025
rect 19610 44015 19690 44025
rect 19930 44015 20010 44025
rect 20250 44015 20330 44025
rect 20570 44015 20650 44025
rect 20890 44015 20970 44025
rect 21210 44015 21290 44025
rect 21530 44015 21610 44025
rect 21850 44015 21930 44025
rect 22170 44015 22250 44025
rect 22490 44015 22570 44025
rect 22810 44015 22890 44025
rect 23130 44015 23210 44025
rect 23450 44015 23530 44025
rect 23770 44015 23850 44025
rect 24090 44015 24170 44025
rect 24410 44015 24490 44025
rect 24730 44015 24810 44025
rect 25050 44015 25130 44025
rect 25370 44015 25450 44025
rect 25690 44015 25770 44025
rect 26010 44015 26090 44025
rect 26330 44015 26410 44025
rect 163590 44015 163670 44025
rect 163910 44015 163990 44025
rect 164230 44015 164310 44025
rect 164550 44015 164630 44025
rect 164870 44015 164950 44025
rect 165190 44015 165270 44025
rect 165510 44015 165590 44025
rect 165830 44015 165910 44025
rect 166150 44015 166230 44025
rect 166470 44015 166550 44025
rect 166790 44015 166870 44025
rect 167110 44015 167190 44025
rect 167430 44015 167510 44025
rect 167750 44015 167830 44025
rect 168070 44015 168150 44025
rect 168390 44015 168470 44025
rect 168710 44015 168790 44025
rect 169030 44015 169110 44025
rect 169350 44015 169430 44025
rect 169670 44015 169750 44025
rect 169990 44015 170070 44025
rect 170310 44015 170390 44025
rect 170630 44015 170710 44025
rect 170950 44015 171030 44025
rect 19050 43935 19060 44015
rect 19370 43935 19380 44015
rect 19690 43935 19700 44015
rect 20010 43935 20020 44015
rect 20330 43935 20340 44015
rect 20650 43935 20660 44015
rect 20970 43935 20980 44015
rect 21290 43935 21300 44015
rect 21610 43935 21620 44015
rect 21930 43935 21940 44015
rect 22250 43935 22260 44015
rect 22570 43935 22580 44015
rect 22890 43935 22900 44015
rect 23210 43935 23220 44015
rect 23530 43935 23540 44015
rect 23850 43935 23860 44015
rect 24170 43935 24180 44015
rect 24490 43935 24500 44015
rect 24810 43935 24820 44015
rect 25130 43935 25140 44015
rect 25450 43935 25460 44015
rect 25770 43935 25780 44015
rect 26090 43935 26100 44015
rect 26410 43935 26420 44015
rect 30360 43975 30440 43985
rect 30680 43975 30760 43985
rect 31000 43975 31080 43985
rect 31320 43975 31400 43985
rect 31640 43975 31720 43985
rect 31960 43975 32040 43985
rect 32280 43975 32360 43985
rect 32600 43975 32680 43985
rect 32920 43975 33000 43985
rect 33240 43975 33320 43985
rect 33560 43975 33640 43985
rect 33880 43975 33960 43985
rect 34200 43975 34280 43985
rect 34520 43975 34600 43985
rect 34840 43975 34920 43985
rect 35160 43975 35240 43985
rect 35480 43975 35560 43985
rect 35800 43975 35880 43985
rect 36120 43975 36200 43985
rect 36440 43975 36520 43985
rect 36760 43975 36840 43985
rect 37080 43975 37160 43985
rect 37400 43975 37480 43985
rect 37720 43975 37800 43985
rect 40180 43975 40260 43985
rect 40500 43975 40580 43985
rect 40820 43975 40900 43985
rect 41140 43975 41220 43985
rect 42560 43975 42640 43985
rect 42880 43975 42960 43985
rect 43200 43975 43280 43985
rect 43520 43975 43600 43985
rect 146400 43975 146480 43985
rect 146720 43975 146800 43985
rect 147040 43975 147120 43985
rect 147360 43975 147440 43985
rect 148780 43975 148860 43985
rect 149100 43975 149180 43985
rect 149420 43975 149500 43985
rect 149740 43975 149820 43985
rect 152200 43975 152280 43985
rect 152520 43975 152600 43985
rect 152840 43975 152920 43985
rect 153160 43975 153240 43985
rect 153480 43975 153560 43985
rect 153800 43975 153880 43985
rect 154120 43975 154200 43985
rect 154440 43975 154520 43985
rect 154760 43975 154840 43985
rect 155080 43975 155160 43985
rect 155400 43975 155480 43985
rect 155720 43975 155800 43985
rect 156040 43975 156120 43985
rect 156360 43975 156440 43985
rect 156680 43975 156760 43985
rect 157000 43975 157080 43985
rect 157320 43975 157400 43985
rect 157640 43975 157720 43985
rect 157960 43975 158040 43985
rect 158280 43975 158360 43985
rect 158600 43975 158680 43985
rect 158920 43975 159000 43985
rect 159240 43975 159320 43985
rect 159560 43975 159640 43985
rect 30440 43895 30450 43975
rect 30760 43895 30770 43975
rect 31080 43895 31090 43975
rect 31400 43895 31410 43975
rect 31720 43895 31730 43975
rect 32040 43895 32050 43975
rect 32360 43895 32370 43975
rect 32680 43895 32690 43975
rect 33000 43895 33010 43975
rect 33320 43895 33330 43975
rect 33640 43895 33650 43975
rect 33960 43895 33970 43975
rect 34280 43895 34290 43975
rect 34600 43895 34610 43975
rect 34920 43895 34930 43975
rect 35240 43895 35250 43975
rect 35560 43895 35570 43975
rect 35880 43895 35890 43975
rect 36200 43895 36210 43975
rect 36520 43895 36530 43975
rect 36840 43895 36850 43975
rect 37160 43895 37170 43975
rect 37480 43895 37490 43975
rect 37800 43895 37810 43975
rect 40260 43895 40270 43975
rect 40580 43895 40590 43975
rect 40900 43895 40910 43975
rect 41220 43895 41230 43975
rect 42640 43895 42650 43975
rect 42960 43895 42970 43975
rect 43280 43895 43290 43975
rect 43600 43895 43610 43975
rect 42420 43780 42500 43790
rect 42740 43780 42820 43790
rect 43060 43780 43140 43790
rect 43380 43780 43460 43790
rect 43700 43780 43780 43790
rect 42500 43700 42510 43780
rect 42820 43700 42830 43780
rect 43140 43700 43150 43780
rect 43460 43700 43470 43780
rect 43780 43700 43790 43780
rect 48500 43710 48605 43960
rect 48870 43840 48900 43900
rect 48990 43840 49020 43900
rect 49110 43840 49140 43900
rect 49230 43840 49260 43900
rect 49350 43840 49380 43900
rect 49470 43840 49500 43900
rect 49590 43840 49620 43900
rect 49710 43840 49740 43900
rect 49830 43840 49860 43900
rect 49950 43840 49980 43900
rect 50070 43840 50100 43900
rect 50190 43840 50220 43900
rect 50310 43840 50340 43900
rect 50430 43840 50460 43900
rect 50550 43840 50580 43900
rect 50670 43840 50700 43900
rect 50790 43840 50820 43900
rect 50910 43840 50940 43900
rect 51030 43840 51060 43900
rect 51150 43840 51180 43900
rect 51270 43840 51300 43900
rect 51390 43840 51420 43900
rect 51510 43840 51540 43900
rect 51630 43840 51660 43900
rect 51750 43840 51780 43900
rect 51870 43840 51900 43900
rect 51990 43840 52020 43900
rect 52110 43840 52140 43900
rect 52230 43840 52260 43900
rect 52350 43840 52380 43900
rect 52470 43840 52500 43900
rect 52590 43840 52620 43900
rect 52710 43840 52740 43900
rect 52830 43840 52860 43900
rect 52950 43840 52980 43900
rect 53070 43840 53100 43900
rect 53190 43840 53220 43900
rect 53310 43840 53340 43900
rect 53430 43840 53460 43900
rect 53550 43840 53580 43900
rect 53670 43840 53700 43900
rect 53790 43840 53820 43900
rect 53910 43840 53940 43900
rect 54030 43840 54060 43900
rect 54150 43840 54180 43900
rect 54270 43840 54300 43900
rect 54390 43840 54420 43900
rect 54510 43840 54540 43900
rect 54630 43840 54660 43900
rect 54750 43840 54780 43900
rect 54870 43840 54900 43900
rect 54990 43840 55020 43900
rect 55110 43840 55140 43900
rect 55230 43840 55260 43900
rect 55350 43840 55380 43900
rect 55470 43840 55500 43900
rect 55590 43840 55620 43900
rect 55710 43840 55740 43900
rect 55830 43840 55860 43900
rect 55950 43840 55980 43900
rect 56070 43840 56100 43900
rect 56190 43840 56220 43900
rect 56310 43840 56340 43900
rect 56430 43840 56460 43900
rect 56550 43840 56580 43900
rect 56670 43840 56700 43900
rect 56790 43840 56820 43900
rect 56910 43840 56940 43900
rect 57030 43840 57060 43900
rect 57150 43840 57180 43900
rect 57270 43840 57300 43900
rect 57390 43840 57420 43900
rect 57510 43840 57540 43900
rect 57630 43840 57660 43900
rect 57750 43840 57780 43900
rect 57870 43840 57900 43900
rect 57990 43840 58020 43900
rect 58110 43840 58140 43900
rect 58230 43840 58260 43900
rect 58350 43840 58380 43900
rect 58470 43840 58500 43900
rect 58590 43840 58620 43900
rect 58710 43840 58740 43900
rect 58830 43840 58860 43900
rect 58950 43840 58980 43900
rect 59070 43840 59100 43900
rect 59190 43840 59220 43900
rect 59310 43840 59340 43900
rect 59430 43840 59460 43900
rect 59550 43840 59580 43900
rect 59670 43840 59700 43900
rect 59790 43840 59820 43900
rect 59910 43840 59940 43900
rect 60030 43840 60060 43900
rect 60150 43840 60180 43900
rect 62370 43840 62400 43900
rect 62490 43840 62520 43900
rect 62610 43840 62640 43900
rect 62730 43840 62760 43900
rect 62850 43840 62880 43900
rect 62970 43840 63000 43900
rect 63090 43840 63120 43900
rect 63210 43840 63240 43900
rect 63330 43840 63360 43900
rect 63450 43840 63480 43900
rect 63570 43840 63600 43900
rect 63690 43840 63720 43900
rect 63810 43840 63840 43900
rect 63930 43840 63960 43900
rect 64050 43840 64080 43900
rect 64170 43840 64200 43900
rect 64290 43840 64320 43900
rect 64410 43840 64440 43900
rect 64530 43840 64560 43900
rect 64650 43840 64680 43900
rect 64770 43840 64800 43900
rect 64890 43840 64920 43900
rect 65010 43840 65040 43900
rect 65130 43840 65160 43900
rect 65250 43840 65280 43900
rect 65370 43840 65400 43900
rect 65490 43840 65520 43900
rect 65610 43840 65640 43900
rect 65730 43840 65760 43900
rect 65850 43840 65880 43900
rect 65970 43840 66000 43900
rect 66090 43840 66120 43900
rect 66210 43840 66240 43900
rect 66330 43840 66360 43900
rect 66450 43840 66480 43900
rect 66570 43840 66600 43900
rect 66690 43840 66720 43900
rect 66810 43840 66840 43900
rect 66930 43840 66960 43900
rect 67050 43840 67080 43900
rect 67170 43840 67200 43900
rect 67290 43840 67320 43900
rect 67410 43840 67440 43900
rect 67530 43840 67560 43900
rect 67650 43840 67680 43900
rect 67770 43840 67800 43900
rect 67890 43840 67920 43900
rect 68010 43840 68040 43900
rect 68130 43840 68160 43900
rect 68250 43840 68280 43900
rect 68370 43840 68400 43900
rect 68490 43840 68520 43900
rect 68610 43840 68640 43900
rect 68730 43840 68760 43900
rect 68850 43840 68880 43900
rect 68970 43840 69000 43900
rect 69090 43840 69120 43900
rect 69210 43840 69240 43900
rect 69330 43840 69360 43900
rect 69450 43840 69480 43900
rect 69570 43840 69600 43900
rect 69690 43840 69720 43900
rect 69810 43840 69840 43900
rect 69930 43840 69960 43900
rect 70050 43840 70080 43900
rect 70170 43840 70200 43900
rect 70290 43840 70320 43900
rect 70410 43840 70440 43900
rect 70530 43840 70560 43900
rect 70650 43840 70680 43900
rect 70770 43840 70800 43900
rect 70890 43840 70920 43900
rect 71010 43840 71040 43900
rect 71130 43840 71160 43900
rect 71250 43840 71280 43900
rect 71370 43840 71400 43900
rect 71490 43840 71520 43900
rect 71610 43840 71640 43900
rect 71730 43840 71760 43900
rect 71850 43840 71880 43900
rect 71970 43840 72000 43900
rect 72090 43840 72120 43900
rect 72210 43840 72240 43900
rect 72330 43840 72360 43900
rect 72450 43840 72480 43900
rect 72570 43840 72600 43900
rect 72690 43840 72720 43900
rect 72810 43840 72840 43900
rect 72930 43840 72960 43900
rect 73050 43840 73080 43900
rect 73170 43840 73200 43900
rect 73290 43840 73320 43900
rect 73410 43840 73440 43900
rect 73530 43840 73560 43900
rect 73650 43840 73680 43900
rect 75870 43840 75900 43900
rect 75990 43840 76020 43900
rect 76110 43840 76140 43900
rect 76230 43840 76260 43900
rect 76350 43840 76380 43900
rect 76470 43840 76500 43900
rect 76590 43840 76620 43900
rect 76710 43840 76740 43900
rect 76830 43840 76860 43900
rect 76950 43840 76980 43900
rect 77070 43840 77100 43900
rect 77190 43840 77220 43900
rect 77310 43840 77340 43900
rect 77430 43840 77460 43900
rect 77550 43840 77580 43900
rect 77670 43840 77700 43900
rect 77790 43840 77820 43900
rect 77910 43840 77940 43900
rect 78030 43840 78060 43900
rect 78150 43840 78180 43900
rect 78270 43840 78300 43900
rect 78390 43840 78420 43900
rect 78510 43840 78540 43900
rect 78630 43840 78660 43900
rect 78750 43840 78780 43900
rect 78870 43840 78900 43900
rect 78990 43840 79020 43900
rect 79110 43840 79140 43900
rect 79230 43840 79260 43900
rect 79350 43840 79380 43900
rect 79470 43840 79500 43900
rect 79590 43840 79620 43900
rect 79710 43840 79740 43900
rect 79830 43840 79860 43900
rect 79950 43840 79980 43900
rect 80070 43840 80100 43900
rect 80190 43840 80220 43900
rect 80310 43840 80340 43900
rect 80430 43840 80460 43900
rect 80550 43840 80580 43900
rect 80670 43840 80700 43900
rect 80790 43840 80820 43900
rect 80910 43840 80940 43900
rect 81030 43840 81060 43900
rect 81150 43840 81180 43900
rect 81270 43840 81300 43900
rect 81390 43840 81420 43900
rect 81510 43840 81540 43900
rect 81630 43840 81660 43900
rect 81750 43840 81780 43900
rect 81870 43840 81900 43900
rect 81990 43840 82020 43900
rect 82110 43840 82140 43900
rect 82230 43840 82260 43900
rect 82350 43840 82380 43900
rect 82470 43840 82500 43900
rect 82590 43840 82620 43900
rect 82710 43840 82740 43900
rect 82830 43840 82860 43900
rect 82950 43840 82980 43900
rect 83070 43840 83100 43900
rect 83190 43840 83220 43900
rect 83310 43840 83340 43900
rect 83430 43840 83460 43900
rect 83550 43840 83580 43900
rect 83670 43840 83700 43900
rect 83790 43840 83820 43900
rect 83910 43840 83940 43900
rect 84030 43840 84060 43900
rect 84150 43840 84180 43900
rect 84270 43840 84300 43900
rect 84390 43840 84420 43900
rect 84510 43840 84540 43900
rect 84630 43840 84660 43900
rect 84750 43840 84780 43900
rect 84870 43840 84900 43900
rect 84990 43840 85020 43900
rect 85110 43840 85140 43900
rect 85230 43840 85260 43900
rect 85350 43840 85380 43900
rect 85470 43840 85500 43900
rect 85590 43840 85620 43900
rect 85710 43840 85740 43900
rect 85830 43840 85860 43900
rect 85950 43840 85980 43900
rect 86070 43840 86100 43900
rect 86190 43840 86220 43900
rect 86310 43840 86340 43900
rect 86430 43840 86460 43900
rect 86550 43840 86580 43900
rect 86670 43840 86700 43900
rect 86790 43840 86820 43900
rect 86910 43840 86940 43900
rect 87030 43840 87060 43900
rect 87150 43840 87180 43900
rect 89370 43840 89400 43900
rect 89490 43840 89520 43900
rect 89610 43840 89640 43900
rect 89730 43840 89760 43900
rect 89850 43840 89880 43900
rect 89970 43840 90000 43900
rect 90090 43840 90120 43900
rect 90210 43840 90240 43900
rect 90330 43840 90360 43900
rect 90450 43840 90480 43900
rect 90570 43840 90600 43900
rect 90690 43840 90720 43900
rect 90810 43840 90840 43900
rect 90930 43840 90960 43900
rect 91050 43840 91080 43900
rect 91170 43840 91200 43900
rect 91290 43840 91320 43900
rect 91410 43840 91440 43900
rect 91530 43840 91560 43900
rect 91650 43840 91680 43900
rect 91770 43840 91800 43900
rect 91890 43840 91920 43900
rect 92010 43840 92040 43900
rect 92130 43840 92160 43900
rect 92250 43840 92280 43900
rect 92370 43840 92400 43900
rect 92490 43840 92520 43900
rect 92610 43840 92640 43900
rect 92730 43840 92760 43900
rect 92850 43840 92880 43900
rect 92970 43840 93000 43900
rect 93090 43840 93120 43900
rect 93210 43840 93240 43900
rect 93330 43840 93360 43900
rect 93450 43840 93480 43900
rect 93570 43840 93600 43900
rect 93690 43840 93720 43900
rect 93810 43840 93840 43900
rect 93930 43840 93960 43900
rect 94050 43840 94080 43900
rect 94170 43840 94200 43900
rect 94290 43840 94320 43900
rect 94410 43840 94440 43900
rect 94530 43840 94560 43900
rect 94650 43840 94680 43900
rect 94770 43840 94800 43900
rect 94890 43840 94920 43900
rect 95010 43840 95040 43900
rect 95130 43840 95160 43900
rect 95250 43840 95280 43900
rect 95370 43840 95400 43900
rect 95490 43840 95520 43900
rect 95610 43840 95640 43900
rect 95730 43840 95760 43900
rect 95850 43840 95880 43900
rect 95970 43840 96000 43900
rect 96090 43840 96120 43900
rect 96210 43840 96240 43900
rect 96330 43840 96360 43900
rect 96450 43840 96480 43900
rect 96570 43840 96600 43900
rect 96690 43840 96720 43900
rect 96810 43840 96840 43900
rect 96930 43840 96960 43900
rect 97050 43840 97080 43900
rect 97170 43840 97200 43900
rect 97290 43840 97320 43900
rect 97410 43840 97440 43900
rect 97530 43840 97560 43900
rect 97650 43840 97680 43900
rect 97770 43840 97800 43900
rect 97890 43840 97920 43900
rect 98010 43840 98040 43900
rect 98130 43840 98160 43900
rect 98250 43840 98280 43900
rect 98370 43840 98400 43900
rect 98490 43840 98520 43900
rect 98610 43840 98640 43900
rect 98730 43840 98760 43900
rect 98850 43840 98880 43900
rect 98970 43840 99000 43900
rect 99090 43840 99120 43900
rect 99210 43840 99240 43900
rect 99330 43840 99360 43900
rect 99450 43840 99480 43900
rect 99570 43840 99600 43900
rect 99690 43840 99720 43900
rect 99810 43840 99840 43900
rect 99930 43840 99960 43900
rect 100050 43840 100080 43900
rect 100170 43840 100200 43900
rect 100290 43840 100320 43900
rect 100410 43840 100440 43900
rect 100530 43840 100560 43900
rect 100650 43840 100680 43900
rect 102870 43840 102900 43900
rect 102990 43840 103020 43900
rect 103110 43840 103140 43900
rect 103230 43840 103260 43900
rect 103350 43840 103380 43900
rect 103470 43840 103500 43900
rect 103590 43840 103620 43900
rect 103710 43840 103740 43900
rect 103830 43840 103860 43900
rect 103950 43840 103980 43900
rect 104070 43840 104100 43900
rect 104190 43840 104220 43900
rect 104310 43840 104340 43900
rect 104430 43840 104460 43900
rect 104550 43840 104580 43900
rect 104670 43840 104700 43900
rect 104790 43840 104820 43900
rect 104910 43840 104940 43900
rect 105030 43840 105060 43900
rect 105150 43840 105180 43900
rect 105270 43840 105300 43900
rect 105390 43840 105420 43900
rect 105510 43840 105540 43900
rect 105630 43840 105660 43900
rect 105750 43840 105780 43900
rect 105870 43840 105900 43900
rect 105990 43840 106020 43900
rect 106110 43840 106140 43900
rect 106230 43840 106260 43900
rect 106350 43840 106380 43900
rect 106470 43840 106500 43900
rect 106590 43840 106620 43900
rect 106710 43840 106740 43900
rect 106830 43840 106860 43900
rect 106950 43840 106980 43900
rect 107070 43840 107100 43900
rect 107190 43840 107220 43900
rect 107310 43840 107340 43900
rect 107430 43840 107460 43900
rect 107550 43840 107580 43900
rect 107670 43840 107700 43900
rect 107790 43840 107820 43900
rect 107910 43840 107940 43900
rect 108030 43840 108060 43900
rect 108150 43840 108180 43900
rect 108270 43840 108300 43900
rect 108390 43840 108420 43900
rect 108510 43840 108540 43900
rect 108630 43840 108660 43900
rect 108750 43840 108780 43900
rect 108870 43840 108900 43900
rect 108990 43840 109020 43900
rect 109110 43840 109140 43900
rect 109230 43840 109260 43900
rect 109350 43840 109380 43900
rect 109470 43840 109500 43900
rect 109590 43840 109620 43900
rect 109710 43840 109740 43900
rect 109830 43840 109860 43900
rect 109950 43840 109980 43900
rect 110070 43840 110100 43900
rect 110190 43840 110220 43900
rect 110310 43840 110340 43900
rect 110430 43840 110460 43900
rect 110550 43840 110580 43900
rect 110670 43840 110700 43900
rect 110790 43840 110820 43900
rect 110910 43840 110940 43900
rect 111030 43840 111060 43900
rect 111150 43840 111180 43900
rect 111270 43840 111300 43900
rect 111390 43840 111420 43900
rect 111510 43840 111540 43900
rect 111630 43840 111660 43900
rect 111750 43840 111780 43900
rect 111870 43840 111900 43900
rect 111990 43840 112020 43900
rect 112110 43840 112140 43900
rect 112230 43840 112260 43900
rect 112350 43840 112380 43900
rect 112470 43840 112500 43900
rect 112590 43840 112620 43900
rect 112710 43840 112740 43900
rect 112830 43840 112860 43900
rect 112950 43840 112980 43900
rect 113070 43840 113100 43900
rect 113190 43840 113220 43900
rect 113310 43840 113340 43900
rect 113430 43840 113460 43900
rect 113550 43840 113580 43900
rect 113670 43840 113700 43900
rect 113790 43840 113820 43900
rect 113910 43840 113940 43900
rect 114030 43840 114060 43900
rect 114150 43840 114180 43900
rect 116370 43840 116400 43900
rect 116490 43840 116520 43900
rect 116610 43840 116640 43900
rect 116730 43840 116760 43900
rect 116850 43840 116880 43900
rect 116970 43840 117000 43900
rect 117090 43840 117120 43900
rect 117210 43840 117240 43900
rect 117330 43840 117360 43900
rect 117450 43840 117480 43900
rect 117570 43840 117600 43900
rect 117690 43840 117720 43900
rect 117810 43840 117840 43900
rect 117930 43840 117960 43900
rect 118050 43840 118080 43900
rect 118170 43840 118200 43900
rect 118290 43840 118320 43900
rect 118410 43840 118440 43900
rect 118530 43840 118560 43900
rect 118650 43840 118680 43900
rect 118770 43840 118800 43900
rect 118890 43840 118920 43900
rect 119010 43840 119040 43900
rect 119130 43840 119160 43900
rect 119250 43840 119280 43900
rect 119370 43840 119400 43900
rect 119490 43840 119520 43900
rect 119610 43840 119640 43900
rect 119730 43840 119760 43900
rect 119850 43840 119880 43900
rect 119970 43840 120000 43900
rect 120090 43840 120120 43900
rect 120210 43840 120240 43900
rect 120330 43840 120360 43900
rect 120450 43840 120480 43900
rect 120570 43840 120600 43900
rect 120690 43840 120720 43900
rect 120810 43840 120840 43900
rect 120930 43840 120960 43900
rect 121050 43840 121080 43900
rect 121170 43840 121200 43900
rect 121290 43840 121320 43900
rect 121410 43840 121440 43900
rect 121530 43840 121560 43900
rect 121650 43840 121680 43900
rect 121770 43840 121800 43900
rect 121890 43840 121920 43900
rect 122010 43840 122040 43900
rect 122130 43840 122160 43900
rect 122250 43840 122280 43900
rect 122370 43840 122400 43900
rect 122490 43840 122520 43900
rect 122610 43840 122640 43900
rect 122730 43840 122760 43900
rect 122850 43840 122880 43900
rect 122970 43840 123000 43900
rect 123090 43840 123120 43900
rect 123210 43840 123240 43900
rect 123330 43840 123360 43900
rect 123450 43840 123480 43900
rect 123570 43840 123600 43900
rect 123690 43840 123720 43900
rect 123810 43840 123840 43900
rect 123930 43840 123960 43900
rect 124050 43840 124080 43900
rect 124170 43840 124200 43900
rect 124290 43840 124320 43900
rect 124410 43840 124440 43900
rect 124530 43840 124560 43900
rect 124650 43840 124680 43900
rect 124770 43840 124800 43900
rect 124890 43840 124920 43900
rect 125010 43840 125040 43900
rect 125130 43840 125160 43900
rect 125250 43840 125280 43900
rect 125370 43840 125400 43900
rect 125490 43840 125520 43900
rect 125610 43840 125640 43900
rect 125730 43840 125760 43900
rect 125850 43840 125880 43900
rect 125970 43840 126000 43900
rect 126090 43840 126120 43900
rect 126210 43840 126240 43900
rect 126330 43840 126360 43900
rect 126450 43840 126480 43900
rect 126570 43840 126600 43900
rect 126690 43840 126720 43900
rect 126810 43840 126840 43900
rect 126930 43840 126960 43900
rect 127050 43840 127080 43900
rect 127170 43840 127200 43900
rect 127290 43840 127320 43900
rect 127410 43840 127440 43900
rect 127530 43840 127560 43900
rect 127650 43840 127680 43900
rect 129870 43840 129900 43900
rect 129990 43840 130020 43900
rect 130110 43840 130140 43900
rect 130230 43840 130260 43900
rect 130350 43840 130380 43900
rect 130470 43840 130500 43900
rect 130590 43840 130620 43900
rect 130710 43840 130740 43900
rect 130830 43840 130860 43900
rect 130950 43840 130980 43900
rect 131070 43840 131100 43900
rect 131190 43840 131220 43900
rect 131310 43840 131340 43900
rect 131430 43840 131460 43900
rect 131550 43840 131580 43900
rect 131670 43840 131700 43900
rect 131790 43840 131820 43900
rect 131910 43840 131940 43900
rect 132030 43840 132060 43900
rect 132150 43840 132180 43900
rect 132270 43840 132300 43900
rect 132390 43840 132420 43900
rect 132510 43840 132540 43900
rect 132630 43840 132660 43900
rect 132750 43840 132780 43900
rect 132870 43840 132900 43900
rect 132990 43840 133020 43900
rect 133110 43840 133140 43900
rect 133230 43840 133260 43900
rect 133350 43840 133380 43900
rect 133470 43840 133500 43900
rect 133590 43840 133620 43900
rect 133710 43840 133740 43900
rect 133830 43840 133860 43900
rect 133950 43840 133980 43900
rect 134070 43840 134100 43900
rect 134190 43840 134220 43900
rect 134310 43840 134340 43900
rect 134430 43840 134460 43900
rect 134550 43840 134580 43900
rect 134670 43840 134700 43900
rect 134790 43840 134820 43900
rect 134910 43840 134940 43900
rect 135030 43840 135060 43900
rect 135150 43840 135180 43900
rect 135270 43840 135300 43900
rect 135390 43840 135420 43900
rect 135510 43840 135540 43900
rect 135630 43840 135660 43900
rect 135750 43840 135780 43900
rect 135870 43840 135900 43900
rect 135990 43840 136020 43900
rect 136110 43840 136140 43900
rect 136230 43840 136260 43900
rect 136350 43840 136380 43900
rect 136470 43840 136500 43900
rect 136590 43840 136620 43900
rect 136710 43840 136740 43900
rect 136830 43840 136860 43900
rect 136950 43840 136980 43900
rect 137070 43840 137100 43900
rect 137190 43840 137220 43900
rect 137310 43840 137340 43900
rect 137430 43840 137460 43900
rect 137550 43840 137580 43900
rect 137670 43840 137700 43900
rect 137790 43840 137820 43900
rect 137910 43840 137940 43900
rect 138030 43840 138060 43900
rect 138150 43840 138180 43900
rect 138270 43840 138300 43900
rect 138390 43840 138420 43900
rect 138510 43840 138540 43900
rect 138630 43840 138660 43900
rect 138750 43840 138780 43900
rect 138870 43840 138900 43900
rect 138990 43840 139020 43900
rect 139110 43840 139140 43900
rect 139230 43840 139260 43900
rect 139350 43840 139380 43900
rect 139470 43840 139500 43900
rect 139590 43840 139620 43900
rect 139710 43840 139740 43900
rect 139830 43840 139860 43900
rect 139950 43840 139980 43900
rect 140070 43840 140100 43900
rect 140190 43840 140220 43900
rect 140310 43840 140340 43900
rect 140430 43840 140460 43900
rect 140550 43840 140580 43900
rect 140670 43840 140700 43900
rect 140790 43840 140820 43900
rect 140910 43840 140940 43900
rect 141030 43840 141060 43900
rect 141150 43840 141180 43900
rect 58560 43780 60130 43790
rect 72060 43780 73630 43790
rect 85560 43780 87130 43790
rect 99060 43780 100630 43790
rect 112560 43780 114130 43790
rect 126060 43780 127630 43790
rect 139560 43780 141130 43790
rect 48500 43700 48640 43710
rect 56330 43700 56450 43760
rect 56590 43700 56710 43760
rect 56850 43700 56970 43760
rect 57110 43700 57230 43760
rect 60360 43700 60440 43710
rect 62060 43700 62140 43710
rect 69830 43700 69950 43760
rect 70090 43700 70210 43760
rect 70350 43700 70470 43760
rect 70610 43700 70730 43760
rect 73860 43700 73940 43710
rect 75560 43700 75640 43710
rect 83330 43700 83450 43760
rect 83590 43700 83710 43760
rect 83850 43700 83970 43760
rect 84110 43700 84230 43760
rect 87360 43700 87440 43710
rect 89060 43700 89140 43710
rect 96830 43700 96950 43760
rect 97090 43700 97210 43760
rect 97350 43700 97470 43760
rect 97610 43700 97730 43760
rect 100860 43700 100940 43710
rect 102560 43700 102640 43710
rect 110330 43700 110450 43760
rect 110590 43700 110710 43760
rect 110850 43700 110970 43760
rect 111110 43700 111230 43760
rect 114360 43700 114440 43710
rect 116060 43700 116140 43710
rect 123830 43700 123950 43760
rect 124090 43700 124210 43760
rect 124350 43700 124470 43760
rect 124610 43700 124730 43760
rect 127860 43700 127940 43710
rect 129560 43700 129640 43710
rect 137330 43700 137450 43760
rect 137590 43700 137710 43760
rect 137850 43700 137970 43760
rect 138110 43700 138230 43760
rect 141360 43700 141440 43710
rect 42580 43620 42660 43630
rect 42900 43620 42980 43630
rect 43220 43620 43300 43630
rect 43540 43620 43620 43630
rect 42660 43540 42670 43620
rect 42980 43540 42990 43620
rect 43300 43540 43310 43620
rect 43620 43540 43630 43620
rect 43785 43600 43865 43610
rect 44105 43600 44185 43610
rect 44425 43600 44505 43610
rect 44745 43600 44825 43610
rect 45065 43600 45145 43610
rect 45385 43600 45465 43610
rect 45705 43600 45785 43610
rect 46025 43600 46105 43610
rect 46345 43600 46425 43610
rect 46665 43600 46745 43610
rect 46985 43600 47065 43610
rect 47305 43600 47385 43610
rect 47625 43600 47705 43610
rect 47945 43600 48025 43610
rect 48265 43600 48345 43610
rect 43865 43550 43875 43600
rect 43785 43520 43875 43550
rect 44185 43520 44195 43600
rect 44505 43520 44515 43600
rect 44825 43520 44835 43600
rect 45145 43520 45155 43600
rect 45465 43520 45475 43600
rect 45785 43520 45795 43600
rect 46105 43520 46115 43600
rect 46425 43520 46435 43600
rect 46745 43520 46755 43600
rect 47065 43520 47075 43600
rect 47385 43520 47395 43600
rect 47705 43520 47715 43600
rect 48025 43520 48035 43600
rect 48345 43520 48355 43600
rect 48500 43570 48605 43700
rect 48640 43620 48650 43700
rect 56450 43580 56510 43700
rect 56710 43580 56770 43700
rect 56970 43580 57030 43700
rect 57230 43580 57290 43700
rect 60440 43620 60450 43700
rect 62140 43620 62150 43700
rect 60580 43600 60660 43610
rect 60900 43600 60980 43610
rect 61320 43600 61400 43610
rect 61640 43600 61720 43610
rect 58860 43580 59250 43590
rect 59450 43580 59840 43590
rect 48500 43560 48640 43570
rect 19060 43460 19140 43470
rect 19380 43460 19460 43470
rect 19700 43460 19780 43470
rect 20020 43460 20100 43470
rect 20340 43460 20420 43470
rect 20660 43460 20740 43470
rect 20980 43460 21060 43470
rect 21300 43460 21380 43470
rect 21620 43460 21700 43470
rect 21940 43460 22020 43470
rect 22260 43460 22340 43470
rect 22580 43460 22660 43470
rect 22900 43460 22980 43470
rect 23220 43460 23300 43470
rect 23540 43460 23620 43470
rect 23860 43460 23940 43470
rect 24180 43460 24260 43470
rect 24500 43460 24580 43470
rect 24820 43460 24900 43470
rect 25140 43460 25220 43470
rect 25460 43460 25540 43470
rect 25780 43460 25860 43470
rect 26100 43460 26180 43470
rect 26420 43460 26500 43470
rect 30580 43460 30660 43470
rect 30900 43460 30980 43470
rect 31220 43460 31300 43470
rect 31540 43460 31620 43470
rect 31860 43460 31940 43470
rect 32180 43460 32260 43470
rect 32500 43460 32580 43470
rect 32820 43460 32900 43470
rect 33140 43460 33220 43470
rect 33460 43460 33540 43470
rect 33780 43460 33860 43470
rect 34100 43460 34180 43470
rect 34420 43460 34500 43470
rect 34740 43460 34820 43470
rect 35060 43460 35140 43470
rect 35380 43460 35460 43470
rect 35700 43460 35780 43470
rect 36020 43460 36100 43470
rect 36340 43460 36420 43470
rect 36660 43460 36740 43470
rect 36980 43460 37060 43470
rect 37300 43460 37380 43470
rect 37620 43460 37700 43470
rect 40180 43460 40260 43470
rect 40500 43460 40580 43470
rect 40820 43460 40900 43470
rect 41140 43460 41220 43470
rect 42420 43460 42500 43470
rect 42740 43460 42820 43470
rect 43060 43460 43140 43470
rect 43380 43460 43460 43470
rect 43700 43460 43780 43470
rect 19140 43380 19150 43460
rect 19460 43380 19470 43460
rect 19780 43380 19790 43460
rect 20100 43380 20110 43460
rect 20420 43380 20430 43460
rect 20740 43380 20750 43460
rect 21060 43380 21070 43460
rect 21380 43380 21390 43460
rect 21700 43380 21710 43460
rect 22020 43380 22030 43460
rect 22340 43380 22350 43460
rect 22660 43380 22670 43460
rect 22980 43380 22990 43460
rect 23300 43380 23310 43460
rect 23620 43380 23630 43460
rect 23940 43380 23950 43460
rect 24260 43380 24270 43460
rect 24580 43380 24590 43460
rect 24900 43380 24910 43460
rect 25220 43380 25230 43460
rect 25540 43380 25550 43460
rect 25860 43380 25870 43460
rect 26180 43380 26190 43460
rect 26500 43380 26510 43460
rect 30660 43380 30670 43460
rect 30980 43380 30990 43460
rect 31300 43380 31310 43460
rect 31620 43380 31630 43460
rect 31940 43380 31950 43460
rect 32260 43380 32270 43460
rect 32580 43380 32590 43460
rect 32900 43380 32910 43460
rect 33220 43380 33230 43460
rect 33540 43380 33550 43460
rect 33860 43380 33870 43460
rect 34180 43380 34190 43460
rect 34500 43380 34510 43460
rect 34820 43380 34830 43460
rect 35140 43380 35150 43460
rect 35460 43380 35470 43460
rect 35780 43380 35790 43460
rect 36100 43380 36110 43460
rect 36420 43380 36430 43460
rect 36740 43380 36750 43460
rect 37060 43380 37070 43460
rect 37380 43380 37390 43460
rect 37700 43380 37710 43460
rect 40260 43380 40270 43460
rect 40580 43380 40590 43460
rect 40900 43380 40910 43460
rect 41220 43380 41230 43460
rect 42500 43380 42510 43460
rect 42820 43380 42830 43460
rect 43140 43380 43150 43460
rect 43460 43380 43470 43460
rect 43780 43380 43790 43460
rect 43945 43440 44025 43450
rect 44265 43440 44345 43450
rect 44585 43440 44665 43450
rect 44905 43440 44985 43450
rect 45225 43440 45305 43450
rect 45545 43440 45625 43450
rect 45865 43440 45945 43450
rect 46185 43440 46265 43450
rect 46505 43440 46585 43450
rect 46825 43440 46905 43450
rect 47145 43440 47225 43450
rect 47465 43440 47545 43450
rect 47785 43440 47865 43450
rect 48105 43440 48185 43450
rect 44025 43360 44035 43440
rect 44345 43360 44355 43440
rect 44665 43360 44675 43440
rect 44985 43360 44995 43440
rect 45305 43360 45315 43440
rect 45625 43360 45635 43440
rect 45945 43360 45955 43440
rect 46265 43360 46275 43440
rect 46585 43360 46595 43440
rect 46905 43360 46915 43440
rect 47225 43360 47235 43440
rect 47545 43360 47555 43440
rect 47865 43360 47875 43440
rect 48185 43360 48195 43440
rect 48500 43430 48605 43560
rect 48640 43480 48650 43560
rect 56340 43550 56700 43560
rect 56340 43470 56350 43550
rect 48500 43420 48640 43430
rect 19220 43300 19300 43310
rect 19540 43300 19620 43310
rect 19860 43300 19940 43310
rect 20180 43300 20260 43310
rect 20500 43300 20580 43310
rect 20820 43300 20900 43310
rect 21140 43300 21220 43310
rect 21460 43300 21540 43310
rect 21780 43300 21860 43310
rect 22100 43300 22180 43310
rect 22420 43300 22500 43310
rect 22740 43300 22820 43310
rect 23060 43300 23140 43310
rect 23380 43300 23460 43310
rect 23700 43300 23780 43310
rect 24020 43300 24100 43310
rect 24340 43300 24420 43310
rect 24660 43300 24740 43310
rect 24980 43300 25060 43310
rect 25300 43300 25380 43310
rect 25620 43300 25700 43310
rect 25940 43300 26020 43310
rect 26260 43300 26340 43310
rect 30420 43300 30500 43310
rect 30740 43300 30820 43310
rect 31060 43300 31140 43310
rect 31380 43300 31460 43310
rect 31700 43300 31780 43310
rect 32020 43300 32100 43310
rect 32340 43300 32420 43310
rect 32660 43300 32740 43310
rect 32980 43300 33060 43310
rect 33300 43300 33380 43310
rect 33620 43300 33700 43310
rect 33940 43300 34020 43310
rect 34260 43300 34340 43310
rect 34580 43300 34660 43310
rect 34900 43300 34980 43310
rect 35220 43300 35300 43310
rect 35540 43300 35620 43310
rect 35860 43300 35940 43310
rect 36180 43300 36260 43310
rect 36500 43300 36580 43310
rect 36820 43300 36900 43310
rect 37140 43300 37220 43310
rect 37460 43300 37540 43310
rect 40340 43300 40420 43310
rect 40660 43300 40740 43310
rect 40980 43300 41060 43310
rect 42580 43300 42660 43310
rect 42900 43300 42980 43310
rect 43220 43300 43300 43310
rect 43540 43300 43620 43310
rect 19300 43220 19310 43300
rect 19620 43220 19630 43300
rect 19940 43220 19950 43300
rect 20260 43220 20270 43300
rect 20580 43220 20590 43300
rect 20900 43220 20910 43300
rect 21220 43220 21230 43300
rect 21540 43220 21550 43300
rect 21860 43220 21870 43300
rect 22180 43220 22190 43300
rect 22500 43220 22510 43300
rect 22820 43220 22830 43300
rect 23140 43220 23150 43300
rect 23460 43220 23470 43300
rect 23780 43220 23790 43300
rect 24100 43220 24110 43300
rect 24420 43220 24430 43300
rect 24740 43220 24750 43300
rect 25060 43220 25070 43300
rect 25380 43220 25390 43300
rect 25700 43220 25710 43300
rect 26020 43220 26030 43300
rect 26340 43220 26350 43300
rect 30500 43220 30510 43300
rect 30820 43220 30830 43300
rect 31140 43220 31150 43300
rect 31460 43220 31470 43300
rect 31780 43220 31790 43300
rect 32100 43220 32110 43300
rect 32420 43220 32430 43300
rect 32740 43220 32750 43300
rect 33060 43220 33070 43300
rect 33380 43220 33390 43300
rect 33700 43220 33710 43300
rect 34020 43220 34030 43300
rect 34340 43220 34350 43300
rect 34660 43220 34670 43300
rect 34980 43220 34990 43300
rect 35300 43220 35310 43300
rect 35620 43220 35630 43300
rect 35940 43220 35950 43300
rect 36260 43220 36270 43300
rect 36580 43220 36590 43300
rect 36900 43220 36910 43300
rect 37220 43220 37230 43300
rect 37540 43220 37550 43300
rect 40420 43220 40430 43300
rect 40740 43220 40750 43300
rect 41060 43220 41070 43300
rect 42660 43220 42670 43300
rect 42980 43220 42990 43300
rect 43300 43220 43310 43300
rect 43620 43220 43630 43300
rect 48500 43290 48605 43420
rect 48640 43340 48650 43420
rect 43785 43280 43865 43290
rect 44105 43280 44185 43290
rect 44425 43280 44505 43290
rect 44745 43280 44825 43290
rect 45065 43280 45145 43290
rect 45385 43280 45465 43290
rect 45705 43280 45785 43290
rect 46025 43280 46105 43290
rect 46345 43280 46425 43290
rect 46665 43280 46745 43290
rect 46985 43280 47065 43290
rect 47305 43280 47385 43290
rect 47625 43280 47705 43290
rect 47945 43280 48025 43290
rect 48265 43280 48345 43290
rect 48500 43280 48640 43290
rect 43865 43230 43875 43280
rect 43785 43200 43875 43230
rect 44185 43200 44195 43280
rect 44505 43200 44515 43280
rect 44825 43200 44835 43280
rect 45145 43200 45155 43280
rect 45465 43200 45475 43280
rect 45785 43200 45795 43280
rect 46105 43200 46115 43280
rect 46425 43200 46435 43280
rect 46745 43200 46755 43280
rect 47065 43200 47075 43280
rect 47385 43200 47395 43280
rect 47705 43200 47715 43280
rect 48025 43200 48035 43280
rect 48345 43200 48355 43280
rect 48500 43150 48605 43280
rect 48640 43200 48650 43280
rect 19060 43140 19140 43150
rect 19380 43140 19460 43150
rect 19700 43140 19780 43150
rect 20020 43140 20100 43150
rect 20340 43140 20420 43150
rect 20660 43140 20740 43150
rect 20980 43140 21060 43150
rect 21300 43140 21380 43150
rect 21620 43140 21700 43150
rect 21940 43140 22020 43150
rect 22260 43140 22340 43150
rect 22580 43140 22660 43150
rect 22900 43140 22980 43150
rect 23220 43140 23300 43150
rect 23540 43140 23620 43150
rect 23860 43140 23940 43150
rect 24180 43140 24260 43150
rect 24500 43140 24580 43150
rect 24820 43140 24900 43150
rect 25140 43140 25220 43150
rect 25460 43140 25540 43150
rect 25780 43140 25860 43150
rect 26100 43140 26180 43150
rect 26420 43140 26500 43150
rect 30580 43140 30660 43150
rect 30900 43140 30980 43150
rect 31220 43140 31300 43150
rect 31540 43140 31620 43150
rect 31860 43140 31940 43150
rect 32180 43140 32260 43150
rect 32500 43140 32580 43150
rect 32820 43140 32900 43150
rect 33140 43140 33220 43150
rect 33460 43140 33540 43150
rect 33780 43140 33860 43150
rect 34100 43140 34180 43150
rect 34420 43140 34500 43150
rect 34740 43140 34820 43150
rect 35060 43140 35140 43150
rect 35380 43140 35460 43150
rect 35700 43140 35780 43150
rect 36020 43140 36100 43150
rect 36340 43140 36420 43150
rect 36660 43140 36740 43150
rect 36980 43140 37060 43150
rect 37300 43140 37380 43150
rect 37620 43140 37700 43150
rect 40180 43140 40260 43150
rect 40500 43140 40580 43150
rect 40820 43140 40900 43150
rect 41140 43140 41220 43150
rect 42420 43140 42500 43150
rect 42740 43140 42820 43150
rect 43060 43140 43140 43150
rect 43380 43140 43460 43150
rect 43700 43140 43780 43150
rect 48500 43140 48640 43150
rect 19140 43060 19150 43140
rect 19460 43060 19470 43140
rect 19780 43060 19790 43140
rect 20100 43060 20110 43140
rect 20420 43060 20430 43140
rect 20740 43060 20750 43140
rect 21060 43060 21070 43140
rect 21380 43060 21390 43140
rect 21700 43060 21710 43140
rect 22020 43060 22030 43140
rect 22340 43060 22350 43140
rect 22660 43060 22670 43140
rect 22980 43060 22990 43140
rect 23300 43060 23310 43140
rect 23620 43060 23630 43140
rect 23940 43060 23950 43140
rect 24260 43060 24270 43140
rect 24580 43060 24590 43140
rect 24900 43060 24910 43140
rect 25220 43060 25230 43140
rect 25540 43060 25550 43140
rect 25860 43060 25870 43140
rect 26180 43060 26190 43140
rect 26500 43060 26510 43140
rect 30660 43060 30670 43140
rect 30980 43060 30990 43140
rect 31300 43060 31310 43140
rect 31620 43060 31630 43140
rect 31940 43060 31950 43140
rect 32260 43060 32270 43140
rect 32580 43060 32590 43140
rect 32900 43060 32910 43140
rect 33220 43060 33230 43140
rect 33540 43060 33550 43140
rect 33860 43060 33870 43140
rect 34180 43060 34190 43140
rect 34500 43060 34510 43140
rect 34820 43060 34830 43140
rect 35140 43060 35150 43140
rect 35460 43060 35470 43140
rect 35780 43060 35790 43140
rect 36100 43060 36110 43140
rect 36420 43060 36430 43140
rect 36740 43060 36750 43140
rect 37060 43060 37070 43140
rect 37380 43060 37390 43140
rect 37700 43060 37710 43140
rect 40260 43060 40270 43140
rect 40580 43060 40590 43140
rect 40900 43060 40910 43140
rect 41220 43060 41230 43140
rect 42500 43060 42510 43140
rect 42820 43060 42830 43140
rect 43140 43060 43150 43140
rect 43460 43060 43470 43140
rect 43780 43060 43790 43140
rect 43945 43120 44025 43130
rect 44265 43120 44345 43130
rect 44585 43120 44665 43130
rect 44905 43120 44985 43130
rect 45225 43120 45305 43130
rect 45545 43120 45625 43130
rect 45865 43120 45945 43130
rect 46185 43120 46265 43130
rect 46505 43120 46585 43130
rect 46825 43120 46905 43130
rect 47145 43120 47225 43130
rect 47465 43120 47545 43130
rect 47785 43120 47865 43130
rect 48105 43120 48185 43130
rect 44025 43040 44035 43120
rect 44345 43040 44355 43120
rect 44665 43040 44675 43120
rect 44985 43040 44995 43120
rect 45305 43040 45315 43120
rect 45625 43040 45635 43120
rect 45945 43040 45955 43120
rect 46265 43040 46275 43120
rect 46585 43040 46595 43120
rect 46905 43040 46915 43120
rect 47225 43040 47235 43120
rect 47545 43040 47555 43120
rect 47865 43040 47875 43120
rect 48185 43040 48195 43120
rect 48500 43010 48605 43140
rect 48640 43060 48650 43140
rect 56320 43030 56380 43390
rect 48500 43000 48640 43010
rect 36180 42980 36260 42990
rect 36500 42980 36580 42990
rect 36820 42980 36900 42990
rect 37140 42980 37220 42990
rect 37460 42980 37540 42990
rect 40340 42980 40420 42990
rect 40660 42980 40740 42990
rect 40980 42980 41060 42990
rect 42580 42980 42660 42990
rect 42900 42980 42980 42990
rect 43220 42980 43300 42990
rect 43540 42980 43620 42990
rect 36260 42900 36270 42980
rect 36580 42900 36590 42980
rect 36900 42900 36910 42980
rect 37220 42900 37230 42980
rect 37540 42900 37550 42980
rect 40420 42900 40430 42980
rect 40740 42900 40750 42980
rect 41060 42900 41070 42980
rect 42660 42900 42670 42980
rect 42980 42900 42990 42980
rect 43300 42900 43310 42980
rect 43620 42900 43630 42980
rect 43785 42960 43865 42970
rect 44105 42960 44185 42970
rect 44425 42960 44505 42970
rect 44745 42960 44825 42970
rect 45065 42960 45145 42970
rect 45385 42960 45465 42970
rect 45705 42960 45785 42970
rect 46025 42960 46105 42970
rect 46345 42960 46425 42970
rect 46665 42960 46745 42970
rect 46985 42960 47065 42970
rect 47305 42960 47385 42970
rect 47625 42960 47705 42970
rect 47945 42960 48025 42970
rect 48265 42960 48345 42970
rect 43865 42910 43875 42960
rect 43785 42880 43875 42910
rect 44185 42880 44195 42960
rect 44505 42880 44515 42960
rect 44825 42880 44835 42960
rect 45145 42880 45155 42960
rect 45465 42880 45475 42960
rect 45785 42880 45795 42960
rect 46105 42880 46115 42960
rect 46425 42880 46435 42960
rect 46745 42880 46755 42960
rect 47065 42880 47075 42960
rect 47385 42880 47395 42960
rect 47705 42880 47715 42960
rect 48025 42880 48035 42960
rect 48345 42880 48355 42960
rect 48500 42870 48605 43000
rect 48640 42920 48650 43000
rect 56415 42910 56425 43550
rect 56430 42950 56440 43470
rect 56580 43030 56640 43390
rect 56675 42910 56685 43550
rect 56690 42950 56700 43550
rect 56860 43550 57220 43560
rect 56860 43470 56870 43550
rect 56840 43030 56900 43390
rect 56935 42910 56945 43550
rect 56950 42950 56960 43470
rect 57100 43030 57160 43390
rect 57195 42910 57205 43550
rect 57210 42950 57220 43550
rect 57705 43540 57755 43550
rect 58585 43540 58635 43550
rect 57360 43030 57420 43390
rect 57490 42960 57500 43490
rect 57540 43430 57620 43440
rect 57620 43370 57630 43430
rect 57520 43310 57640 43370
rect 57540 43290 57620 43300
rect 57620 43210 57630 43290
rect 57640 43190 57700 43310
rect 57540 43150 57620 43160
rect 57620 43090 57630 43150
rect 57520 43030 57640 43090
rect 57540 43010 57620 43020
rect 57620 42930 57630 43010
rect 57640 42910 57700 43030
rect 56365 42900 56415 42910
rect 56625 42900 56675 42910
rect 56885 42900 56935 42910
rect 57145 42900 57195 42910
rect 48500 42860 48640 42870
rect 36020 42820 36100 42830
rect 36340 42820 36420 42830
rect 36660 42820 36740 42830
rect 36980 42820 37060 42830
rect 37300 42820 37380 42830
rect 37620 42820 37700 42830
rect 40180 42820 40260 42830
rect 40500 42820 40580 42830
rect 40820 42820 40900 42830
rect 41140 42820 41220 42830
rect 42740 42820 42820 42830
rect 43060 42820 43140 42830
rect 43380 42820 43460 42830
rect 43700 42820 43780 42830
rect 36100 42740 36110 42820
rect 36420 42740 36430 42820
rect 36740 42740 36750 42820
rect 37060 42740 37070 42820
rect 37380 42740 37390 42820
rect 37700 42740 37710 42820
rect 40260 42740 40270 42820
rect 40580 42740 40590 42820
rect 40900 42740 40910 42820
rect 41220 42740 41230 42820
rect 42820 42740 42830 42820
rect 43140 42740 43150 42820
rect 43460 42740 43470 42820
rect 43780 42740 43790 42820
rect 43945 42800 44025 42810
rect 44265 42800 44345 42810
rect 44585 42800 44665 42810
rect 44905 42800 44985 42810
rect 45225 42800 45305 42810
rect 45545 42800 45625 42810
rect 45865 42800 45945 42810
rect 46185 42800 46265 42810
rect 46505 42800 46585 42810
rect 46825 42800 46905 42810
rect 47145 42800 47225 42810
rect 47465 42800 47545 42810
rect 47785 42800 47865 42810
rect 48105 42800 48185 42810
rect 44025 42720 44035 42800
rect 44345 42720 44355 42800
rect 44665 42720 44675 42800
rect 44985 42720 44995 42800
rect 45305 42720 45315 42800
rect 45625 42720 45635 42800
rect 45945 42720 45955 42800
rect 46265 42720 46275 42800
rect 46585 42720 46595 42800
rect 46905 42720 46915 42800
rect 47225 42720 47235 42800
rect 47545 42720 47555 42800
rect 47865 42720 47875 42800
rect 48185 42720 48195 42800
rect 48500 42730 48605 42860
rect 48640 42780 48650 42860
rect 56540 42822 56680 42892
rect 56740 42822 56880 42892
rect 56940 42822 57080 42892
rect 57480 42860 57690 42870
rect 48500 42720 48640 42730
rect 36180 42660 36260 42670
rect 36500 42660 36580 42670
rect 36820 42660 36900 42670
rect 37140 42660 37220 42670
rect 37460 42660 37540 42670
rect 40340 42660 40420 42670
rect 40660 42660 40740 42670
rect 40980 42660 41060 42670
rect 42900 42660 42980 42670
rect 43220 42660 43300 42670
rect 43540 42660 43620 42670
rect 36260 42580 36270 42660
rect 36580 42580 36590 42660
rect 36900 42580 36910 42660
rect 37220 42580 37230 42660
rect 37540 42580 37550 42660
rect 40420 42580 40430 42660
rect 40740 42580 40750 42660
rect 41060 42580 41070 42660
rect 42980 42580 42990 42660
rect 43300 42580 43310 42660
rect 43620 42580 43630 42660
rect 43785 42640 43865 42650
rect 44105 42640 44185 42650
rect 44425 42640 44505 42650
rect 44745 42640 44825 42650
rect 45065 42640 45145 42650
rect 45385 42640 45465 42650
rect 45705 42640 45785 42650
rect 46025 42640 46105 42650
rect 46345 42640 46425 42650
rect 46665 42640 46745 42650
rect 46985 42640 47065 42650
rect 47305 42640 47385 42650
rect 47625 42640 47705 42650
rect 47945 42640 48025 42650
rect 48265 42640 48345 42650
rect 43865 42590 43875 42640
rect 43785 42560 43875 42590
rect 44185 42560 44195 42640
rect 44505 42560 44515 42640
rect 44825 42560 44835 42640
rect 45145 42560 45155 42640
rect 45465 42560 45475 42640
rect 45785 42560 45795 42640
rect 46105 42560 46115 42640
rect 46425 42560 46435 42640
rect 46745 42560 46755 42640
rect 47065 42560 47075 42640
rect 47385 42560 47395 42640
rect 47705 42560 47715 42640
rect 48025 42560 48035 42640
rect 48345 42560 48355 42640
rect 48500 42590 48605 42720
rect 48640 42640 48650 42720
rect 56025 42675 56105 42685
rect 56185 42675 56265 42685
rect 56680 42682 56740 42822
rect 56880 42682 56940 42822
rect 57080 42682 57150 42822
rect 57755 42790 57765 43540
rect 57770 42870 57780 43500
rect 57840 43430 57920 43440
rect 58420 43430 58500 43440
rect 57920 43370 57930 43430
rect 58500 43370 58510 43430
rect 57820 43310 57940 43370
rect 58400 43310 58520 43370
rect 57940 43190 58000 43310
rect 58420 43290 58500 43300
rect 58500 43210 58510 43290
rect 58520 43190 58580 43310
rect 57840 43150 57920 43160
rect 58420 43150 58500 43160
rect 57920 43090 57930 43150
rect 58500 43090 58510 43150
rect 57820 43030 57940 43090
rect 58400 43030 58520 43090
rect 57940 42910 58000 43030
rect 58420 43010 58500 43020
rect 58500 42930 58510 43010
rect 58520 42910 58580 43030
rect 57770 42860 57910 42870
rect 58430 42860 58570 42870
rect 58635 42790 58645 43540
rect 58650 42870 58660 43580
rect 59175 43540 59225 43550
rect 58700 43310 58820 43370
rect 58820 43200 58880 43310
rect 58700 43190 58880 43200
rect 58700 43030 58820 43090
rect 58820 42910 58880 43030
rect 58960 42870 58970 43490
rect 59010 43430 59090 43440
rect 59090 43370 59100 43430
rect 58990 43310 59110 43370
rect 59010 43290 59090 43300
rect 59090 43210 59100 43290
rect 59110 43190 59170 43310
rect 59010 43150 59090 43160
rect 59090 43090 59100 43150
rect 58990 43030 59110 43090
rect 59010 43010 59090 43020
rect 59090 42930 59100 43010
rect 59110 42910 59170 43030
rect 58650 42860 58860 42870
rect 58950 42860 59160 42870
rect 59225 42790 59235 43540
rect 59240 42870 59250 43580
rect 59765 43540 59815 43550
rect 59290 43310 59410 43370
rect 59410 43200 59470 43310
rect 59290 43190 59470 43200
rect 59290 43030 59410 43090
rect 59410 42910 59470 43030
rect 59550 42870 59560 43490
rect 59600 43430 59680 43440
rect 59680 43370 59690 43430
rect 59580 43310 59700 43370
rect 59600 43290 59680 43300
rect 59680 43210 59690 43290
rect 59700 43190 59760 43310
rect 59600 43150 59680 43160
rect 59680 43090 59690 43150
rect 59580 43030 59700 43090
rect 59600 43010 59680 43020
rect 59680 42930 59690 43010
rect 59700 42910 59760 43030
rect 59240 42860 59450 42870
rect 59540 42860 59750 42870
rect 59815 42790 59825 43540
rect 59830 42870 59840 43580
rect 60360 43560 60440 43570
rect 60440 43480 60450 43560
rect 60660 43520 60670 43600
rect 60980 43520 60990 43600
rect 61400 43520 61410 43600
rect 61720 43520 61730 43600
rect 69950 43580 70010 43700
rect 70210 43580 70270 43700
rect 70470 43580 70530 43700
rect 70730 43580 70790 43700
rect 73940 43620 73950 43700
rect 75640 43620 75650 43700
rect 74080 43600 74160 43610
rect 74400 43600 74480 43610
rect 74820 43600 74900 43610
rect 75140 43600 75220 43610
rect 72360 43580 72750 43590
rect 72950 43580 73340 43590
rect 62060 43560 62140 43570
rect 62140 43480 62150 43560
rect 69840 43550 70200 43560
rect 69840 43470 69850 43550
rect 60740 43440 60820 43450
rect 61060 43440 61140 43450
rect 61480 43440 61560 43450
rect 61800 43440 61880 43450
rect 59900 43430 59980 43440
rect 59980 43370 59990 43430
rect 60360 43420 60440 43430
rect 59880 43310 60000 43370
rect 60440 43340 60450 43420
rect 60820 43360 60830 43440
rect 61140 43360 61150 43440
rect 61560 43360 61570 43440
rect 61880 43360 61890 43440
rect 62060 43420 62140 43430
rect 62140 43340 62150 43420
rect 60000 43190 60060 43310
rect 60360 43280 60440 43290
rect 60580 43280 60660 43290
rect 60900 43280 60980 43290
rect 61320 43280 61400 43290
rect 61640 43280 61720 43290
rect 62060 43280 62140 43290
rect 60440 43200 60450 43280
rect 60660 43200 60670 43280
rect 60980 43200 60990 43280
rect 61400 43200 61410 43280
rect 61720 43200 61730 43280
rect 62140 43200 62150 43280
rect 59900 43150 59980 43160
rect 59980 43090 59990 43150
rect 60360 43140 60440 43150
rect 62060 43140 62140 43150
rect 59880 43030 60000 43090
rect 60440 43060 60450 43140
rect 60740 43120 60820 43130
rect 61060 43120 61140 43130
rect 61480 43120 61560 43130
rect 61800 43120 61880 43130
rect 60820 43040 60830 43120
rect 61140 43040 61150 43120
rect 61560 43040 61570 43120
rect 61880 43040 61890 43120
rect 62140 43060 62150 43140
rect 69820 43030 69880 43390
rect 60000 42910 60060 43030
rect 60360 43000 60440 43010
rect 62060 43000 62140 43010
rect 60440 42920 60450 43000
rect 60580 42960 60660 42970
rect 60900 42960 60980 42970
rect 61320 42960 61400 42970
rect 61640 42960 61720 42970
rect 60660 42880 60670 42960
rect 60980 42880 60990 42960
rect 61400 42880 61410 42960
rect 61720 42880 61730 42960
rect 62140 42920 62150 43000
rect 69915 42910 69925 43550
rect 69930 42950 69940 43470
rect 70080 43030 70140 43390
rect 70175 42910 70185 43550
rect 70190 42950 70200 43550
rect 70360 43550 70720 43560
rect 70360 43470 70370 43550
rect 70340 43030 70400 43390
rect 70435 42910 70445 43550
rect 70450 42950 70460 43470
rect 70600 43030 70660 43390
rect 70695 42910 70705 43550
rect 70710 42950 70720 43550
rect 71205 43540 71255 43550
rect 72085 43540 72135 43550
rect 70860 43030 70920 43390
rect 70990 42960 71000 43490
rect 71040 43430 71120 43440
rect 71120 43370 71130 43430
rect 71020 43310 71140 43370
rect 71040 43290 71120 43300
rect 71120 43210 71130 43290
rect 71140 43190 71200 43310
rect 71040 43150 71120 43160
rect 71120 43090 71130 43150
rect 71020 43030 71140 43090
rect 71040 43010 71120 43020
rect 71120 42930 71130 43010
rect 71140 42910 71200 43030
rect 69865 42900 69915 42910
rect 70125 42900 70175 42910
rect 70385 42900 70435 42910
rect 70645 42900 70695 42910
rect 59830 42860 59970 42870
rect 60360 42860 60440 42870
rect 62060 42860 62140 42870
rect 70040 42860 70180 42892
rect 70240 42860 70380 42892
rect 70440 42860 70580 42892
rect 70980 42860 71190 42870
rect 71255 42860 71265 43540
rect 71270 42870 71280 43500
rect 71340 43430 71420 43440
rect 71920 43430 72000 43440
rect 71420 43370 71430 43430
rect 72000 43370 72010 43430
rect 71320 43310 71440 43370
rect 71900 43310 72020 43370
rect 71440 43190 71500 43310
rect 71920 43290 72000 43300
rect 72000 43210 72010 43290
rect 72020 43190 72080 43310
rect 71340 43150 71420 43160
rect 71920 43150 72000 43160
rect 71420 43090 71430 43150
rect 72000 43090 72010 43150
rect 71320 43030 71440 43090
rect 71900 43030 72020 43090
rect 71440 42910 71500 43030
rect 71920 43010 72000 43020
rect 72000 42935 72010 43010
rect 72020 42935 72080 43030
rect 72135 42935 72145 43540
rect 72150 42935 72160 43580
rect 72675 43540 72725 43550
rect 72200 43310 72320 43370
rect 72320 43200 72380 43310
rect 72200 43190 72380 43200
rect 72200 43030 72320 43090
rect 72320 42935 72380 43030
rect 72460 42935 72470 43490
rect 72510 43430 72590 43440
rect 72590 43370 72600 43430
rect 72490 43310 72610 43370
rect 72510 43290 72590 43300
rect 72590 43210 72600 43290
rect 72610 43190 72670 43310
rect 72510 43150 72590 43160
rect 72590 43090 72600 43150
rect 72490 43030 72610 43090
rect 72510 43010 72590 43020
rect 72590 42935 72600 43010
rect 72610 42935 72670 43030
rect 72725 42935 72735 43540
rect 72740 42935 72750 43580
rect 73265 43540 73315 43550
rect 72790 43310 72910 43370
rect 72910 43200 72970 43310
rect 72790 43190 72970 43200
rect 72790 43030 72910 43090
rect 72910 42935 72970 43030
rect 73050 42935 73060 43490
rect 73100 43430 73180 43440
rect 73180 43370 73190 43430
rect 73080 43310 73200 43370
rect 73100 43290 73180 43300
rect 73180 43210 73190 43290
rect 73200 43190 73260 43310
rect 73100 43150 73180 43160
rect 73180 43090 73190 43150
rect 73080 43030 73200 43090
rect 73100 43010 73180 43020
rect 73180 42935 73190 43010
rect 73200 42935 73260 43030
rect 73245 42910 73260 42935
rect 71270 42860 71410 42870
rect 71930 42860 72000 42870
rect 73245 42860 73250 42870
rect 57670 42730 57790 42790
rect 58550 42730 58670 42790
rect 59140 42730 59260 42790
rect 59730 42730 59850 42790
rect 60440 42780 60450 42860
rect 60740 42800 60820 42810
rect 61060 42800 61140 42810
rect 61480 42800 61560 42810
rect 61800 42800 61880 42810
rect 57400 42700 57480 42710
rect 57560 42700 57640 42710
rect 56105 42595 56115 42675
rect 56185 42595 56195 42675
rect 56265 42595 56275 42675
rect 57480 42620 57490 42700
rect 57560 42620 57570 42700
rect 57640 42620 57650 42700
rect 57790 42610 57850 42730
rect 58670 42610 58730 42730
rect 58760 42700 58840 42710
rect 58940 42700 59020 42710
rect 58840 42620 58850 42700
rect 59020 42620 59030 42700
rect 59260 42610 59320 42730
rect 59360 42700 59440 42710
rect 59540 42700 59620 42710
rect 59440 42620 59450 42700
rect 59620 42620 59630 42700
rect 59850 42610 59910 42730
rect 60360 42720 60440 42730
rect 60820 42720 60830 42800
rect 61140 42720 61150 42800
rect 61560 42720 61570 42800
rect 61880 42720 61890 42800
rect 62140 42780 62150 42860
rect 73315 42790 73325 43540
rect 73330 42870 73340 43580
rect 73860 43560 73940 43570
rect 73940 43480 73950 43560
rect 74160 43520 74170 43600
rect 74480 43520 74490 43600
rect 74900 43520 74910 43600
rect 75220 43520 75230 43600
rect 83450 43580 83510 43700
rect 83710 43580 83770 43700
rect 83970 43580 84030 43700
rect 84230 43580 84290 43700
rect 87440 43620 87450 43700
rect 89140 43620 89150 43700
rect 87580 43600 87660 43610
rect 87900 43600 87980 43610
rect 88320 43600 88400 43610
rect 88640 43600 88720 43610
rect 85860 43580 86250 43590
rect 86450 43580 86840 43590
rect 75560 43560 75640 43570
rect 75640 43480 75650 43560
rect 83340 43550 83700 43560
rect 83340 43470 83350 43550
rect 74240 43440 74320 43450
rect 74560 43440 74640 43450
rect 74980 43440 75060 43450
rect 75300 43440 75380 43450
rect 73400 43430 73480 43440
rect 73480 43370 73490 43430
rect 73860 43420 73940 43430
rect 73380 43310 73500 43370
rect 73940 43340 73950 43420
rect 74320 43360 74330 43440
rect 74640 43360 74650 43440
rect 75060 43360 75070 43440
rect 75380 43360 75390 43440
rect 75560 43420 75640 43430
rect 75640 43340 75650 43420
rect 73500 43190 73560 43310
rect 73860 43280 73940 43290
rect 74080 43280 74160 43290
rect 74400 43280 74480 43290
rect 74820 43280 74900 43290
rect 75140 43280 75220 43290
rect 75560 43280 75640 43290
rect 73940 43200 73950 43280
rect 74160 43200 74170 43280
rect 74480 43200 74490 43280
rect 74900 43200 74910 43280
rect 75220 43200 75230 43280
rect 75640 43200 75650 43280
rect 73400 43150 73480 43160
rect 73480 43090 73490 43150
rect 73860 43140 73940 43150
rect 75560 43140 75640 43150
rect 73380 43030 73500 43090
rect 73940 43060 73950 43140
rect 74240 43120 74320 43130
rect 74560 43120 74640 43130
rect 74980 43120 75060 43130
rect 75300 43120 75380 43130
rect 74320 43040 74330 43120
rect 74640 43040 74650 43120
rect 75060 43040 75070 43120
rect 75380 43040 75390 43120
rect 75640 43060 75650 43140
rect 83320 43030 83380 43390
rect 73500 42910 73560 43030
rect 73860 43000 73940 43010
rect 75560 43000 75640 43010
rect 73940 42920 73950 43000
rect 74080 42960 74160 42970
rect 74400 42960 74480 42970
rect 74820 42960 74900 42970
rect 75140 42960 75220 42970
rect 74160 42880 74170 42960
rect 74480 42880 74490 42960
rect 74900 42880 74910 42960
rect 75220 42880 75230 42960
rect 75640 42920 75650 43000
rect 83415 42935 83425 43550
rect 83430 42950 83440 43470
rect 83580 43030 83640 43390
rect 83675 42935 83685 43550
rect 83690 42950 83700 43550
rect 83860 43550 84220 43560
rect 83860 43470 83870 43550
rect 83840 43030 83900 43390
rect 83935 42935 83945 43550
rect 83950 42950 83960 43470
rect 84100 43030 84160 43390
rect 84195 42910 84205 43550
rect 84210 42950 84220 43550
rect 84705 43540 84755 43550
rect 85585 43540 85635 43550
rect 84360 43030 84420 43390
rect 84490 42960 84500 43490
rect 84540 43430 84620 43440
rect 84620 43370 84630 43430
rect 84520 43310 84640 43370
rect 84540 43290 84620 43300
rect 84620 43210 84630 43290
rect 84640 43190 84700 43310
rect 84540 43150 84620 43160
rect 84620 43090 84630 43150
rect 84520 43030 84640 43090
rect 84540 43010 84620 43020
rect 84620 42930 84630 43010
rect 84640 42910 84700 43030
rect 84145 42900 84195 42910
rect 73330 42860 73470 42870
rect 73860 42860 73940 42870
rect 75560 42860 75640 42870
rect 84000 42860 84080 42892
rect 84480 42860 84690 42870
rect 84755 42860 84765 43540
rect 84770 42870 84780 43500
rect 84840 43430 84920 43440
rect 85420 43430 85500 43440
rect 84920 43370 84930 43430
rect 85500 43370 85510 43430
rect 84820 43310 84940 43370
rect 85400 43310 85520 43370
rect 84940 43190 85000 43310
rect 85420 43290 85500 43300
rect 85500 43210 85510 43290
rect 85520 43190 85580 43310
rect 84840 43150 84920 43160
rect 85420 43150 85500 43160
rect 84920 43090 84930 43150
rect 85500 43090 85510 43150
rect 84820 43030 84940 43090
rect 85400 43030 85520 43090
rect 84940 42910 85000 43030
rect 85420 43010 85500 43020
rect 85500 42930 85510 43010
rect 85520 42910 85580 43030
rect 84770 42860 84910 42870
rect 85430 42860 85570 42870
rect 85635 42860 85645 43540
rect 85650 42870 85660 43580
rect 86175 43540 86225 43550
rect 85700 43310 85820 43370
rect 85820 43200 85880 43310
rect 85700 43190 85880 43200
rect 85700 43030 85820 43090
rect 85820 42910 85880 43030
rect 85960 42870 85970 43490
rect 86010 43430 86090 43440
rect 86090 43370 86100 43430
rect 85990 43310 86110 43370
rect 86010 43290 86090 43300
rect 86090 43210 86100 43290
rect 86110 43190 86170 43310
rect 86010 43150 86090 43160
rect 86090 43090 86100 43150
rect 85990 43030 86110 43090
rect 86010 43010 86090 43020
rect 86090 42930 86100 43010
rect 86110 42910 86170 43030
rect 85650 42860 85860 42870
rect 85950 42860 86160 42870
rect 86225 42860 86235 43540
rect 86240 42870 86250 43580
rect 86765 43540 86815 43550
rect 86290 43310 86410 43370
rect 86410 43200 86470 43310
rect 86290 43190 86470 43200
rect 86290 43030 86410 43090
rect 86410 42910 86470 43030
rect 86550 42870 86560 43490
rect 86600 43430 86680 43440
rect 86680 43370 86690 43430
rect 86580 43310 86700 43370
rect 86600 43290 86680 43300
rect 86680 43210 86690 43290
rect 86700 43190 86760 43310
rect 86600 43150 86680 43160
rect 86680 43090 86690 43150
rect 86580 43030 86700 43090
rect 86600 43010 86680 43020
rect 86680 42930 86690 43010
rect 86700 42910 86760 43030
rect 86240 42860 86450 42870
rect 86540 42860 86750 42870
rect 73245 42730 73350 42790
rect 73940 42780 73950 42860
rect 74240 42800 74320 42810
rect 74560 42800 74640 42810
rect 74980 42800 75060 42810
rect 75300 42800 75380 42810
rect 62060 42720 62140 42730
rect 60440 42640 60450 42720
rect 60580 42640 60660 42650
rect 60900 42640 60980 42650
rect 61320 42640 61400 42650
rect 61640 42640 61720 42650
rect 62140 42640 62150 42720
rect 48500 42580 48640 42590
rect 60360 42580 60440 42590
rect 36020 42500 36100 42510
rect 36340 42500 36420 42510
rect 36660 42500 36740 42510
rect 36980 42500 37060 42510
rect 37300 42500 37380 42510
rect 37620 42500 37700 42510
rect 40180 42500 40260 42510
rect 40500 42500 40580 42510
rect 40820 42500 40900 42510
rect 41140 42500 41220 42510
rect 43060 42500 43140 42510
rect 43380 42500 43460 42510
rect 43700 42500 43780 42510
rect 36100 42420 36110 42500
rect 36420 42420 36430 42500
rect 36740 42420 36750 42500
rect 37060 42420 37070 42500
rect 37380 42420 37390 42500
rect 37700 42420 37710 42500
rect 40260 42420 40270 42500
rect 40580 42420 40590 42500
rect 40900 42420 40910 42500
rect 41220 42420 41230 42500
rect 43140 42420 43150 42500
rect 43460 42420 43470 42500
rect 43780 42420 43790 42500
rect 48500 42450 48605 42580
rect 48640 42500 48650 42580
rect 57340 42560 57820 42570
rect 58520 42560 59880 42570
rect 60440 42500 60450 42580
rect 60660 42560 60670 42640
rect 60980 42560 60990 42640
rect 61400 42560 61410 42640
rect 61720 42560 61730 42640
rect 73350 42610 73410 42730
rect 73860 42720 73940 42730
rect 74320 42720 74330 42800
rect 74640 42720 74650 42800
rect 75060 42720 75070 42800
rect 75380 42720 75390 42800
rect 75640 42780 75650 42860
rect 86815 42790 86825 43540
rect 86830 42870 86840 43580
rect 87360 43560 87440 43570
rect 87440 43480 87450 43560
rect 87660 43520 87670 43600
rect 87980 43520 87990 43600
rect 88400 43520 88410 43600
rect 88720 43520 88730 43600
rect 96950 43580 97010 43700
rect 97210 43580 97270 43700
rect 97470 43580 97530 43700
rect 97730 43580 97790 43700
rect 100940 43620 100950 43700
rect 102640 43620 102650 43700
rect 101080 43600 101160 43610
rect 101400 43600 101480 43610
rect 101820 43600 101900 43610
rect 102140 43600 102220 43610
rect 99360 43580 99750 43590
rect 99950 43580 100340 43590
rect 89060 43560 89140 43570
rect 89140 43480 89150 43560
rect 96840 43550 97200 43560
rect 96840 43470 96850 43550
rect 87740 43440 87820 43450
rect 88060 43440 88140 43450
rect 88480 43440 88560 43450
rect 88800 43440 88880 43450
rect 86900 43430 86980 43440
rect 86980 43370 86990 43430
rect 87360 43420 87440 43430
rect 86880 43310 87000 43370
rect 87440 43340 87450 43420
rect 87820 43360 87830 43440
rect 88140 43360 88150 43440
rect 88560 43360 88570 43440
rect 88880 43360 88890 43440
rect 89060 43420 89140 43430
rect 89140 43340 89150 43420
rect 87000 43190 87060 43310
rect 87360 43280 87440 43290
rect 87580 43280 87660 43290
rect 87900 43280 87980 43290
rect 88320 43280 88400 43290
rect 88640 43280 88720 43290
rect 89060 43280 89140 43290
rect 87440 43200 87450 43280
rect 87660 43200 87670 43280
rect 87980 43200 87990 43280
rect 88400 43200 88410 43280
rect 88720 43200 88730 43280
rect 89140 43200 89150 43280
rect 86900 43150 86980 43160
rect 86980 43090 86990 43150
rect 87360 43140 87440 43150
rect 89060 43140 89140 43150
rect 86880 43030 87000 43090
rect 87440 43060 87450 43140
rect 87740 43120 87820 43130
rect 88060 43120 88140 43130
rect 88480 43120 88560 43130
rect 88800 43120 88880 43130
rect 87820 43040 87830 43120
rect 88140 43040 88150 43120
rect 88560 43040 88570 43120
rect 88880 43040 88890 43120
rect 89140 43060 89150 43140
rect 96820 43030 96880 43390
rect 87000 42910 87060 43030
rect 87360 43000 87440 43010
rect 89060 43000 89140 43010
rect 87440 42920 87450 43000
rect 87580 42960 87660 42970
rect 87900 42960 87980 42970
rect 88320 42960 88400 42970
rect 88640 42960 88720 42970
rect 87660 42880 87670 42960
rect 87980 42880 87990 42960
rect 88400 42880 88410 42960
rect 88720 42880 88730 42960
rect 89140 42920 89150 43000
rect 96915 42910 96925 43550
rect 96930 42950 96940 43470
rect 97080 43030 97140 43390
rect 97175 42910 97185 43550
rect 97190 42950 97200 43550
rect 97360 43550 97720 43560
rect 97360 43470 97370 43550
rect 97340 43030 97400 43390
rect 97435 42910 97445 43550
rect 97450 42950 97460 43470
rect 97600 43030 97660 43390
rect 97695 42910 97705 43550
rect 97710 42950 97720 43550
rect 98205 43540 98255 43550
rect 99085 43540 99135 43550
rect 97860 43030 97920 43390
rect 97990 42960 98000 43490
rect 98040 43430 98120 43440
rect 98120 43370 98130 43430
rect 98020 43310 98140 43370
rect 98040 43290 98120 43300
rect 98120 43210 98130 43290
rect 98140 43190 98200 43310
rect 98040 43150 98120 43160
rect 98120 43090 98130 43150
rect 98020 43030 98140 43090
rect 98040 43010 98120 43020
rect 98120 42930 98130 43010
rect 98140 42910 98200 43030
rect 96865 42900 96915 42910
rect 97125 42900 97175 42910
rect 97385 42900 97435 42910
rect 97645 42900 97695 42910
rect 98255 42900 98265 43540
rect 98270 42900 98280 43500
rect 98340 43430 98420 43440
rect 98920 43430 99000 43440
rect 98420 43370 98430 43430
rect 99000 43370 99010 43430
rect 98320 43310 98440 43370
rect 98900 43310 99020 43370
rect 98440 43190 98500 43310
rect 98920 43290 99000 43300
rect 99000 43210 99010 43290
rect 99020 43190 99080 43310
rect 98340 43150 98420 43160
rect 98920 43150 99000 43160
rect 98420 43090 98430 43150
rect 99000 43090 99010 43150
rect 98320 43030 98440 43090
rect 98900 43030 99020 43090
rect 98440 42910 98500 43030
rect 98920 43010 99000 43020
rect 99000 42930 99010 43010
rect 99020 42910 99080 43030
rect 99135 42900 99145 43540
rect 99150 42900 99160 43580
rect 99675 43540 99725 43550
rect 99200 43310 99320 43370
rect 99320 43200 99380 43310
rect 99200 43190 99380 43200
rect 99200 43030 99320 43090
rect 99320 42910 99380 43030
rect 99460 42900 99470 43490
rect 99510 43430 99590 43440
rect 99590 43370 99600 43430
rect 99490 43310 99610 43370
rect 99510 43290 99590 43300
rect 99590 43210 99600 43290
rect 99610 43190 99670 43310
rect 99510 43150 99590 43160
rect 99590 43090 99600 43150
rect 99490 43030 99610 43090
rect 99510 43010 99590 43020
rect 99590 42930 99600 43010
rect 99610 42910 99670 43030
rect 99725 42900 99735 43540
rect 99740 42900 99750 43580
rect 100265 43540 100315 43550
rect 99790 43310 99910 43370
rect 99910 43200 99970 43310
rect 99790 43190 99970 43200
rect 99790 43030 99910 43090
rect 99910 42910 99970 43030
rect 100050 42900 100060 43490
rect 100100 43430 100180 43440
rect 100180 43370 100190 43430
rect 100080 43310 100200 43370
rect 100100 43290 100180 43300
rect 100180 43210 100190 43290
rect 100200 43190 100260 43310
rect 100100 43150 100180 43160
rect 100180 43090 100190 43150
rect 100080 43030 100200 43090
rect 100100 43010 100180 43020
rect 100180 42930 100190 43010
rect 100200 42910 100260 43030
rect 86830 42860 86970 42870
rect 87360 42860 87440 42870
rect 89060 42860 89140 42870
rect 100245 42860 100250 42870
rect 86745 42730 86850 42790
rect 87440 42780 87450 42860
rect 87740 42800 87820 42810
rect 88060 42800 88140 42810
rect 88480 42800 88560 42810
rect 88800 42800 88880 42810
rect 75560 42720 75640 42730
rect 73940 42640 73950 42720
rect 74080 42640 74160 42650
rect 74400 42640 74480 42650
rect 74820 42640 74900 42650
rect 75140 42640 75220 42650
rect 75640 42640 75650 42720
rect 62060 42580 62140 42590
rect 73860 42580 73940 42590
rect 62140 42500 62150 42580
rect 73245 42560 73380 42570
rect 73940 42500 73950 42580
rect 74160 42560 74170 42640
rect 74480 42560 74490 42640
rect 74900 42560 74910 42640
rect 75220 42560 75230 42640
rect 86850 42610 86910 42730
rect 87360 42720 87440 42730
rect 87820 42720 87830 42800
rect 88140 42720 88150 42800
rect 88560 42720 88570 42800
rect 88880 42720 88890 42800
rect 89140 42780 89150 42860
rect 100315 42790 100325 43540
rect 100330 42870 100340 43580
rect 100860 43560 100940 43570
rect 100940 43480 100950 43560
rect 101160 43520 101170 43600
rect 101480 43520 101490 43600
rect 101900 43520 101910 43600
rect 102220 43520 102230 43600
rect 110450 43580 110510 43700
rect 110710 43580 110770 43700
rect 110970 43580 111030 43700
rect 111230 43580 111290 43700
rect 114440 43620 114450 43700
rect 116140 43620 116150 43700
rect 114580 43600 114660 43610
rect 114900 43600 114980 43610
rect 115320 43600 115400 43610
rect 115640 43600 115720 43610
rect 112860 43580 113250 43590
rect 113450 43580 113840 43590
rect 102560 43560 102640 43570
rect 102640 43480 102650 43560
rect 110340 43550 110700 43560
rect 110340 43470 110350 43550
rect 101240 43440 101320 43450
rect 101560 43440 101640 43450
rect 101980 43440 102060 43450
rect 102300 43440 102380 43450
rect 100400 43430 100480 43440
rect 100480 43370 100490 43430
rect 100860 43420 100940 43430
rect 100380 43310 100500 43370
rect 100940 43340 100950 43420
rect 101320 43360 101330 43440
rect 101640 43360 101650 43440
rect 102060 43360 102070 43440
rect 102380 43360 102390 43440
rect 102560 43420 102640 43430
rect 102640 43340 102650 43420
rect 100500 43190 100560 43310
rect 100860 43280 100940 43290
rect 101080 43280 101160 43290
rect 101400 43280 101480 43290
rect 101820 43280 101900 43290
rect 102140 43280 102220 43290
rect 102560 43280 102640 43290
rect 100940 43200 100950 43280
rect 101160 43200 101170 43280
rect 101480 43200 101490 43280
rect 101900 43200 101910 43280
rect 102220 43200 102230 43280
rect 102640 43200 102650 43280
rect 100400 43150 100480 43160
rect 100480 43090 100490 43150
rect 100860 43140 100940 43150
rect 102560 43140 102640 43150
rect 100380 43030 100500 43090
rect 100940 43060 100950 43140
rect 101240 43120 101320 43130
rect 101560 43120 101640 43130
rect 101980 43120 102060 43130
rect 102300 43120 102380 43130
rect 101320 43040 101330 43120
rect 101640 43040 101650 43120
rect 102060 43040 102070 43120
rect 102380 43040 102390 43120
rect 102640 43060 102650 43140
rect 110320 43030 110380 43390
rect 100500 42910 100560 43030
rect 100860 43000 100940 43010
rect 102560 43000 102640 43010
rect 100940 42920 100950 43000
rect 101080 42960 101160 42970
rect 101400 42960 101480 42970
rect 101820 42960 101900 42970
rect 102140 42960 102220 42970
rect 101160 42880 101170 42960
rect 101480 42880 101490 42960
rect 101900 42880 101910 42960
rect 102220 42880 102230 42960
rect 102640 42920 102650 43000
rect 110415 42910 110425 43550
rect 110430 42950 110440 43470
rect 110580 43030 110640 43390
rect 110675 42910 110685 43550
rect 110690 42950 110700 43550
rect 110860 43550 111220 43560
rect 110860 43470 110870 43550
rect 110840 43030 110900 43390
rect 110935 42910 110945 43550
rect 110950 42950 110960 43470
rect 111100 43030 111160 43390
rect 111195 42910 111205 43550
rect 111210 42950 111220 43550
rect 111705 43540 111755 43550
rect 112585 43540 112635 43550
rect 111360 43030 111420 43390
rect 111490 42960 111500 43490
rect 111540 43430 111620 43440
rect 111620 43370 111630 43430
rect 111520 43310 111640 43370
rect 111540 43290 111620 43300
rect 111620 43210 111630 43290
rect 111640 43190 111700 43310
rect 111540 43150 111620 43160
rect 111620 43090 111630 43150
rect 111520 43030 111640 43090
rect 111540 43010 111620 43020
rect 111620 42930 111630 43010
rect 111640 42910 111700 43030
rect 110365 42900 110415 42910
rect 110625 42900 110675 42910
rect 110885 42900 110935 42910
rect 111145 42900 111195 42910
rect 100330 42860 100470 42870
rect 100860 42860 100940 42870
rect 102560 42860 102640 42870
rect 100245 42730 100350 42790
rect 100940 42780 100950 42860
rect 101240 42800 101320 42810
rect 101560 42800 101640 42810
rect 101980 42800 102060 42810
rect 102300 42800 102380 42810
rect 89060 42720 89140 42730
rect 87440 42640 87450 42720
rect 87580 42640 87660 42650
rect 87900 42640 87980 42650
rect 88320 42640 88400 42650
rect 88640 42640 88720 42650
rect 89140 42640 89150 42720
rect 75560 42580 75640 42590
rect 87360 42580 87440 42590
rect 75640 42500 75650 42580
rect 86745 42560 86880 42570
rect 87440 42500 87450 42580
rect 87660 42560 87670 42640
rect 87980 42560 87990 42640
rect 88400 42560 88410 42640
rect 88720 42560 88730 42640
rect 100350 42610 100410 42730
rect 100860 42720 100940 42730
rect 101320 42720 101330 42800
rect 101640 42720 101650 42800
rect 102060 42720 102070 42800
rect 102380 42720 102390 42800
rect 102640 42780 102650 42860
rect 110540 42850 110680 42892
rect 110740 42850 110880 42892
rect 110940 42850 111080 42892
rect 111480 42860 111690 42870
rect 111755 42850 111765 43540
rect 111770 42870 111780 43500
rect 111840 43430 111920 43440
rect 112420 43430 112500 43440
rect 111920 43370 111930 43430
rect 112500 43370 112510 43430
rect 111820 43310 111940 43370
rect 112400 43310 112520 43370
rect 111940 43190 112000 43310
rect 112420 43290 112500 43300
rect 112500 43210 112510 43290
rect 112520 43190 112580 43310
rect 111840 43150 111920 43160
rect 112420 43150 112500 43160
rect 111920 43090 111930 43150
rect 112500 43090 112510 43150
rect 111820 43030 111940 43090
rect 112400 43030 112520 43090
rect 111940 42910 112000 43030
rect 112420 43010 112500 43020
rect 112500 42930 112510 43010
rect 112520 42910 112580 43030
rect 111770 42860 111910 42870
rect 112430 42860 112570 42870
rect 112635 42850 112645 43540
rect 112650 42870 112660 43580
rect 113175 43540 113225 43550
rect 112700 43310 112820 43370
rect 112820 43200 112880 43310
rect 112700 43190 112880 43200
rect 112700 43030 112820 43090
rect 112820 42910 112880 43030
rect 112960 42870 112970 43490
rect 113010 43430 113090 43440
rect 113090 43370 113100 43430
rect 112990 43310 113110 43370
rect 113010 43290 113090 43300
rect 113090 43210 113100 43290
rect 113110 43190 113170 43310
rect 113010 43150 113090 43160
rect 113090 43090 113100 43150
rect 112990 43030 113110 43090
rect 113010 43010 113090 43020
rect 113090 42930 113100 43010
rect 113110 42910 113170 43030
rect 112650 42860 112860 42870
rect 112950 42860 113160 42870
rect 113225 42850 113235 43540
rect 113240 42870 113250 43580
rect 113765 43540 113815 43550
rect 113290 43310 113410 43370
rect 113410 43200 113470 43310
rect 113290 43190 113470 43200
rect 113290 43030 113410 43090
rect 113410 42910 113470 43030
rect 113550 42870 113560 43490
rect 113600 43430 113680 43440
rect 113680 43370 113690 43430
rect 113580 43310 113700 43370
rect 113600 43290 113680 43300
rect 113680 43210 113690 43290
rect 113700 43190 113760 43310
rect 113600 43150 113680 43160
rect 113680 43090 113690 43150
rect 113580 43030 113700 43090
rect 113600 43010 113680 43020
rect 113680 42930 113690 43010
rect 113700 42910 113760 43030
rect 113240 42860 113450 42870
rect 113540 42860 113750 42870
rect 113815 42790 113825 43540
rect 113830 42870 113840 43580
rect 114360 43560 114440 43570
rect 114440 43480 114450 43560
rect 114660 43520 114670 43600
rect 114980 43520 114990 43600
rect 115400 43520 115410 43600
rect 115720 43520 115730 43600
rect 123950 43580 124010 43700
rect 124210 43580 124270 43700
rect 124470 43580 124530 43700
rect 124730 43580 124790 43700
rect 127940 43620 127950 43700
rect 129640 43620 129650 43700
rect 128080 43600 128160 43610
rect 128400 43600 128480 43610
rect 128820 43600 128900 43610
rect 129140 43600 129220 43610
rect 126360 43580 126750 43590
rect 126950 43580 127340 43590
rect 116060 43560 116140 43570
rect 116140 43480 116150 43560
rect 123840 43550 124200 43560
rect 123840 43470 123850 43550
rect 114740 43440 114820 43450
rect 115060 43440 115140 43450
rect 115480 43440 115560 43450
rect 115800 43440 115880 43450
rect 113900 43430 113980 43440
rect 113980 43370 113990 43430
rect 114360 43420 114440 43430
rect 113880 43310 114000 43370
rect 114440 43340 114450 43420
rect 114820 43360 114830 43440
rect 115140 43360 115150 43440
rect 115560 43360 115570 43440
rect 115880 43360 115890 43440
rect 116060 43420 116140 43430
rect 116140 43340 116150 43420
rect 114000 43190 114060 43310
rect 114360 43280 114440 43290
rect 114580 43280 114660 43290
rect 114900 43280 114980 43290
rect 115320 43280 115400 43290
rect 115640 43280 115720 43290
rect 116060 43280 116140 43290
rect 114440 43200 114450 43280
rect 114660 43200 114670 43280
rect 114980 43200 114990 43280
rect 115400 43200 115410 43280
rect 115720 43200 115730 43280
rect 116140 43200 116150 43280
rect 113900 43150 113980 43160
rect 113980 43090 113990 43150
rect 114360 43140 114440 43150
rect 116060 43140 116140 43150
rect 113880 43030 114000 43090
rect 114440 43060 114450 43140
rect 114740 43120 114820 43130
rect 115060 43120 115140 43130
rect 115480 43120 115560 43130
rect 115800 43120 115880 43130
rect 114820 43040 114830 43120
rect 115140 43040 115150 43120
rect 115560 43040 115570 43120
rect 115880 43040 115890 43120
rect 116140 43060 116150 43140
rect 123820 43030 123880 43390
rect 114000 42910 114060 43030
rect 114360 43000 114440 43010
rect 116060 43000 116140 43010
rect 114440 42920 114450 43000
rect 114580 42960 114660 42970
rect 114900 42960 114980 42970
rect 115320 42960 115400 42970
rect 115640 42960 115720 42970
rect 114660 42880 114670 42960
rect 114980 42880 114990 42960
rect 115400 42880 115410 42960
rect 115720 42880 115730 42960
rect 116140 42920 116150 43000
rect 123915 42910 123925 43550
rect 123930 42950 123940 43470
rect 124080 43030 124140 43390
rect 124175 42910 124185 43550
rect 124190 42950 124200 43550
rect 124360 43550 124720 43560
rect 124360 43470 124370 43550
rect 124340 43030 124400 43390
rect 124435 42910 124445 43550
rect 124450 42950 124460 43470
rect 124600 43030 124660 43390
rect 124695 42910 124705 43550
rect 124710 42950 124720 43550
rect 125205 43540 125255 43550
rect 126085 43540 126135 43550
rect 124860 43030 124920 43390
rect 124990 42960 125000 43490
rect 125040 43430 125120 43440
rect 125120 43370 125130 43430
rect 125020 43310 125140 43370
rect 125040 43290 125120 43300
rect 125120 43210 125130 43290
rect 125140 43190 125200 43310
rect 125040 43150 125120 43160
rect 125120 43090 125130 43150
rect 125020 43030 125140 43090
rect 125040 43010 125120 43020
rect 125120 42930 125130 43010
rect 125140 42910 125200 43030
rect 123865 42900 123915 42910
rect 124125 42900 124175 42910
rect 124385 42900 124435 42910
rect 124645 42900 124695 42910
rect 113830 42860 113970 42870
rect 114360 42860 114440 42870
rect 116060 42860 116140 42870
rect 124040 42860 124180 42892
rect 124240 42860 124380 42892
rect 124440 42860 124580 42892
rect 124980 42860 125190 42870
rect 125255 42860 125265 43540
rect 125270 42870 125280 43500
rect 125340 43430 125420 43440
rect 125920 43430 126000 43440
rect 125420 43370 125430 43430
rect 126000 43370 126010 43430
rect 125320 43310 125440 43370
rect 125900 43310 126020 43370
rect 125440 43190 125500 43310
rect 125920 43290 126000 43300
rect 126000 43210 126010 43290
rect 126020 43190 126080 43310
rect 125340 43150 125420 43160
rect 125920 43150 126000 43160
rect 125420 43090 125430 43150
rect 126000 43090 126010 43150
rect 125320 43030 125440 43090
rect 125900 43030 126020 43090
rect 125440 42910 125500 43030
rect 125920 43010 126000 43020
rect 126000 42930 126010 43010
rect 126020 42910 126080 43030
rect 125270 42860 125410 42870
rect 125930 42860 126070 42870
rect 126135 42860 126145 43540
rect 126150 42870 126160 43580
rect 126675 43540 126725 43550
rect 126200 43310 126320 43370
rect 126320 43200 126380 43310
rect 126200 43190 126380 43200
rect 126200 43030 126320 43090
rect 126320 42910 126380 43030
rect 126460 42870 126470 43490
rect 126510 43430 126590 43440
rect 126590 43370 126600 43430
rect 126490 43310 126610 43370
rect 126510 43290 126590 43300
rect 126590 43210 126600 43290
rect 126610 43190 126670 43310
rect 126510 43150 126590 43160
rect 126590 43090 126600 43150
rect 126490 43030 126610 43090
rect 126510 43010 126590 43020
rect 126590 42930 126600 43010
rect 126610 42910 126670 43030
rect 126150 42860 126360 42870
rect 126450 42860 126660 42870
rect 126725 42860 126735 43540
rect 126740 42870 126750 43580
rect 127265 43540 127315 43550
rect 126790 43310 126910 43370
rect 126910 43200 126970 43310
rect 126790 43190 126970 43200
rect 126790 43030 126910 43090
rect 126910 42910 126970 43030
rect 127050 42870 127060 43490
rect 127100 43430 127180 43440
rect 127180 43370 127190 43430
rect 127080 43310 127200 43370
rect 127100 43290 127180 43300
rect 127180 43210 127190 43290
rect 127200 43190 127260 43310
rect 127100 43150 127180 43160
rect 127180 43090 127190 43150
rect 127080 43030 127200 43090
rect 127100 43010 127180 43020
rect 127180 42930 127190 43010
rect 127200 42910 127260 43030
rect 126740 42860 126950 42870
rect 127040 42860 127250 42870
rect 113745 42730 113850 42790
rect 114440 42780 114450 42860
rect 114740 42800 114820 42810
rect 115060 42800 115140 42810
rect 115480 42800 115560 42810
rect 115800 42800 115880 42810
rect 102560 42720 102640 42730
rect 100940 42640 100950 42720
rect 101080 42640 101160 42650
rect 101400 42640 101480 42650
rect 101820 42640 101900 42650
rect 102140 42640 102220 42650
rect 102640 42640 102650 42720
rect 89060 42580 89140 42590
rect 100860 42580 100940 42590
rect 89140 42500 89150 42580
rect 100245 42560 100380 42570
rect 100940 42500 100950 42580
rect 101160 42560 101170 42640
rect 101480 42560 101490 42640
rect 101900 42560 101910 42640
rect 102220 42560 102230 42640
rect 113850 42610 113910 42730
rect 114360 42720 114440 42730
rect 114820 42720 114830 42800
rect 115140 42720 115150 42800
rect 115560 42720 115570 42800
rect 115880 42720 115890 42800
rect 116140 42780 116150 42860
rect 127315 42790 127325 43540
rect 127330 42870 127340 43580
rect 127860 43560 127940 43570
rect 127940 43480 127950 43560
rect 128160 43520 128170 43600
rect 128480 43520 128490 43600
rect 128900 43520 128910 43600
rect 129220 43520 129230 43600
rect 137450 43580 137510 43700
rect 137710 43580 137770 43700
rect 137970 43580 138030 43700
rect 138230 43580 138290 43700
rect 141440 43620 141450 43700
rect 139860 43580 140250 43590
rect 140450 43580 140840 43590
rect 129560 43560 129640 43570
rect 129640 43480 129650 43560
rect 137340 43550 137700 43560
rect 137340 43470 137350 43550
rect 128240 43440 128320 43450
rect 128560 43440 128640 43450
rect 128980 43440 129060 43450
rect 129300 43440 129380 43450
rect 127400 43430 127480 43440
rect 127480 43370 127490 43430
rect 127860 43420 127940 43430
rect 127380 43310 127500 43370
rect 127940 43340 127950 43420
rect 128320 43360 128330 43440
rect 128640 43360 128650 43440
rect 129060 43360 129070 43440
rect 129380 43360 129390 43440
rect 129560 43420 129640 43430
rect 129640 43340 129650 43420
rect 127500 43190 127560 43310
rect 127860 43280 127940 43290
rect 128080 43280 128160 43290
rect 128400 43280 128480 43290
rect 128820 43280 128900 43290
rect 129140 43280 129220 43290
rect 129560 43280 129640 43290
rect 127940 43200 127950 43280
rect 128160 43200 128170 43280
rect 128480 43200 128490 43280
rect 128900 43200 128910 43280
rect 129220 43200 129230 43280
rect 129640 43200 129650 43280
rect 127400 43150 127480 43160
rect 127480 43090 127490 43150
rect 127860 43140 127940 43150
rect 129560 43140 129640 43150
rect 127380 43030 127500 43090
rect 127940 43060 127950 43140
rect 128240 43120 128320 43130
rect 128560 43120 128640 43130
rect 128980 43120 129060 43130
rect 129300 43120 129380 43130
rect 128320 43040 128330 43120
rect 128640 43040 128650 43120
rect 129060 43040 129070 43120
rect 129380 43040 129390 43120
rect 129640 43060 129650 43140
rect 137320 43030 137380 43390
rect 127500 42910 127560 43030
rect 127860 43000 127940 43010
rect 129560 43000 129640 43010
rect 127940 42920 127950 43000
rect 128080 42960 128160 42970
rect 128400 42960 128480 42970
rect 128820 42960 128900 42970
rect 129140 42960 129220 42970
rect 128160 42880 128170 42960
rect 128480 42880 128490 42960
rect 128900 42880 128910 42960
rect 129220 42880 129230 42960
rect 129640 42920 129650 43000
rect 137415 42910 137425 43550
rect 137430 42950 137440 43470
rect 137580 43030 137640 43390
rect 137675 42910 137685 43550
rect 137690 42950 137700 43550
rect 137860 43550 138220 43560
rect 137860 43470 137870 43550
rect 137840 43030 137900 43390
rect 137935 42910 137945 43550
rect 137950 42950 137960 43470
rect 138100 43030 138160 43390
rect 138195 42910 138205 43550
rect 138210 42950 138220 43550
rect 138705 43540 138755 43550
rect 139585 43540 139635 43550
rect 138360 43030 138420 43390
rect 138490 42960 138500 43490
rect 138540 43430 138620 43440
rect 138620 43370 138630 43430
rect 138520 43310 138640 43370
rect 138540 43290 138620 43300
rect 138620 43210 138630 43290
rect 138640 43190 138700 43310
rect 138540 43150 138620 43160
rect 138620 43090 138630 43150
rect 138520 43030 138640 43090
rect 138540 43010 138620 43020
rect 138620 42930 138630 43010
rect 138640 42910 138700 43030
rect 137365 42900 137415 42910
rect 137625 42900 137675 42910
rect 137885 42900 137935 42910
rect 138145 42900 138195 42910
rect 127330 42860 127470 42870
rect 127860 42860 127940 42870
rect 129560 42860 129640 42870
rect 137540 42860 137680 42892
rect 137740 42860 137880 42892
rect 137940 42860 138080 42892
rect 138480 42860 138690 42870
rect 138755 42860 138765 43540
rect 138770 42870 138780 43500
rect 138840 43430 138920 43440
rect 139420 43430 139500 43440
rect 138920 43370 138930 43430
rect 139500 43370 139510 43430
rect 138820 43310 138940 43370
rect 139400 43310 139520 43370
rect 138940 43190 139000 43310
rect 139420 43290 139500 43300
rect 139500 43210 139510 43290
rect 139520 43190 139580 43310
rect 138840 43150 138920 43160
rect 139420 43150 139500 43160
rect 138920 43090 138930 43150
rect 139500 43090 139510 43150
rect 138820 43030 138940 43090
rect 139400 43030 139520 43090
rect 138940 42910 139000 43030
rect 139420 43010 139500 43020
rect 139500 42930 139510 43010
rect 139520 42910 139580 43030
rect 138770 42860 138910 42870
rect 139430 42860 139570 42870
rect 139635 42860 139645 43540
rect 139650 42870 139660 43580
rect 140175 43540 140225 43550
rect 139700 43310 139820 43370
rect 139820 43200 139880 43310
rect 139700 43190 139880 43200
rect 139700 43030 139820 43090
rect 139820 42910 139880 43030
rect 139960 42870 139970 43490
rect 140010 43430 140090 43440
rect 140090 43370 140100 43430
rect 139990 43310 140110 43370
rect 140010 43290 140090 43300
rect 140090 43210 140100 43290
rect 140110 43190 140170 43310
rect 140010 43150 140090 43160
rect 140090 43090 140100 43150
rect 139990 43030 140110 43090
rect 140010 43010 140090 43020
rect 140090 42930 140100 43010
rect 140110 42910 140170 43030
rect 139650 42860 139860 42870
rect 139950 42860 140160 42870
rect 140225 42860 140235 43540
rect 140240 42870 140250 43580
rect 140765 43540 140815 43550
rect 140290 43310 140410 43370
rect 140410 43200 140470 43310
rect 140290 43190 140470 43200
rect 140290 43030 140410 43090
rect 140410 42910 140470 43030
rect 140550 42870 140560 43490
rect 140600 43430 140680 43440
rect 140680 43370 140690 43430
rect 140580 43310 140700 43370
rect 140600 43290 140680 43300
rect 140680 43210 140690 43290
rect 140700 43190 140760 43310
rect 140600 43150 140680 43160
rect 140680 43090 140690 43150
rect 140580 43030 140700 43090
rect 140600 43010 140680 43020
rect 140680 42930 140690 43010
rect 140700 42910 140760 43030
rect 140240 42860 140450 42870
rect 140540 42860 140750 42870
rect 140815 42860 140825 43540
rect 140830 42870 140840 43580
rect 141360 43560 141440 43570
rect 141440 43480 141450 43560
rect 140900 43430 140980 43440
rect 140980 43370 140990 43430
rect 141360 43420 141440 43430
rect 140880 43310 141000 43370
rect 141440 43340 141450 43420
rect 141000 43190 141060 43310
rect 141360 43280 141440 43290
rect 141440 43200 141450 43280
rect 140900 43150 140980 43160
rect 140980 43090 140990 43150
rect 141360 43140 141440 43150
rect 140880 43030 141000 43090
rect 141440 43060 141450 43140
rect 141000 42910 141060 43030
rect 141360 43000 141440 43010
rect 141440 42920 141450 43000
rect 140830 42860 140970 42870
rect 141360 42860 141440 42870
rect 127245 42730 127350 42790
rect 127940 42780 127950 42860
rect 128240 42800 128320 42810
rect 128560 42800 128640 42810
rect 128980 42800 129060 42810
rect 129300 42800 129380 42810
rect 116060 42720 116140 42730
rect 114440 42640 114450 42720
rect 114580 42640 114660 42650
rect 114900 42640 114980 42650
rect 115320 42640 115400 42650
rect 115640 42640 115720 42650
rect 116140 42640 116150 42720
rect 102560 42580 102640 42590
rect 114360 42580 114440 42590
rect 102640 42500 102650 42580
rect 113745 42560 113880 42570
rect 114440 42500 114450 42580
rect 114660 42560 114670 42640
rect 114980 42560 114990 42640
rect 115400 42560 115410 42640
rect 115720 42560 115730 42640
rect 127350 42610 127410 42730
rect 127860 42720 127940 42730
rect 128320 42720 128330 42800
rect 128640 42720 128650 42800
rect 129060 42720 129070 42800
rect 129380 42720 129390 42800
rect 129640 42780 129650 42860
rect 140830 42730 140850 42790
rect 141440 42780 141450 42860
rect 129560 42720 129640 42730
rect 127940 42640 127950 42720
rect 128080 42640 128160 42650
rect 128400 42640 128480 42650
rect 128820 42640 128900 42650
rect 129140 42640 129220 42650
rect 129640 42640 129650 42720
rect 116060 42580 116140 42590
rect 127860 42580 127940 42590
rect 116140 42500 116150 42580
rect 127245 42560 127380 42570
rect 127940 42500 127950 42580
rect 128160 42560 128170 42640
rect 128480 42560 128490 42640
rect 128900 42560 128910 42640
rect 129220 42560 129230 42640
rect 140850 42610 140910 42730
rect 141360 42720 141440 42730
rect 141440 42640 141450 42720
rect 129560 42580 129640 42590
rect 141360 42580 141440 42590
rect 129640 42500 129650 42580
rect 140830 42560 140880 42570
rect 141440 42500 141450 42580
rect 48500 42440 48640 42450
rect 60360 42440 60440 42450
rect 62060 42440 62140 42450
rect 73860 42440 73940 42450
rect 75560 42440 75640 42450
rect 87360 42440 87440 42450
rect 89060 42440 89140 42450
rect 100860 42440 100940 42450
rect 102560 42440 102640 42450
rect 114360 42440 114440 42450
rect 116060 42440 116140 42450
rect 127860 42440 127940 42450
rect 129560 42440 129640 42450
rect 141360 42440 141440 42450
rect 36180 42340 36260 42350
rect 36500 42340 36580 42350
rect 36820 42340 36900 42350
rect 37140 42340 37220 42350
rect 37460 42340 37540 42350
rect 40340 42340 40420 42350
rect 40660 42340 40740 42350
rect 40980 42340 41060 42350
rect 36260 42260 36270 42340
rect 36580 42260 36590 42340
rect 36900 42260 36910 42340
rect 37220 42260 37230 42340
rect 37540 42260 37550 42340
rect 40420 42260 40430 42340
rect 40740 42260 40750 42340
rect 41060 42260 41070 42340
rect 48500 42300 48605 42440
rect 48640 42360 48650 42440
rect 48870 42360 48900 42420
rect 48990 42360 49020 42420
rect 49110 42360 49140 42420
rect 49230 42360 49260 42420
rect 49350 42360 49380 42420
rect 49470 42360 49500 42420
rect 49590 42360 49620 42420
rect 49710 42360 49740 42420
rect 49830 42360 49860 42420
rect 49950 42360 49980 42420
rect 50070 42360 50100 42420
rect 50190 42360 50220 42420
rect 50310 42360 50340 42420
rect 50430 42360 50460 42420
rect 50550 42360 50580 42420
rect 50670 42360 50700 42420
rect 50790 42360 50820 42420
rect 50910 42360 50940 42420
rect 51030 42360 51060 42420
rect 51150 42360 51180 42420
rect 51270 42360 51300 42420
rect 51390 42360 51420 42420
rect 51510 42360 51540 42420
rect 51630 42360 51660 42420
rect 51750 42360 51780 42420
rect 51870 42360 51900 42420
rect 51990 42360 52020 42420
rect 52110 42360 52140 42420
rect 52230 42360 52260 42420
rect 52350 42360 52380 42420
rect 52470 42360 52500 42420
rect 52590 42360 52620 42420
rect 52710 42360 52740 42420
rect 52830 42360 52860 42420
rect 52950 42360 52980 42420
rect 53070 42360 53100 42420
rect 53190 42360 53220 42420
rect 53310 42360 53340 42420
rect 53430 42360 53460 42420
rect 53550 42360 53580 42420
rect 53670 42360 53700 42420
rect 53790 42360 53820 42420
rect 53910 42360 53940 42420
rect 54030 42360 54060 42420
rect 54150 42360 54180 42420
rect 54270 42360 54300 42420
rect 54390 42360 54420 42420
rect 54510 42360 54540 42420
rect 54630 42360 54660 42420
rect 54750 42360 54780 42420
rect 54870 42360 54900 42420
rect 54990 42360 55020 42420
rect 55110 42360 55140 42420
rect 55230 42360 55260 42420
rect 55350 42360 55380 42420
rect 55470 42360 55500 42420
rect 55590 42360 55620 42420
rect 55710 42360 55740 42420
rect 55830 42360 55860 42420
rect 55950 42360 55980 42420
rect 56070 42360 56100 42420
rect 56190 42360 56220 42420
rect 56310 42360 56340 42420
rect 56430 42360 56460 42420
rect 56550 42360 56580 42420
rect 56670 42360 56700 42420
rect 56790 42360 56820 42420
rect 56910 42360 56940 42420
rect 57030 42360 57060 42420
rect 57150 42360 57180 42420
rect 57270 42360 57300 42420
rect 57390 42360 57420 42420
rect 57510 42360 57540 42420
rect 57630 42360 57660 42420
rect 57750 42360 57780 42420
rect 57870 42360 57900 42420
rect 57990 42360 58020 42420
rect 58110 42360 58140 42420
rect 58230 42360 58260 42420
rect 58350 42360 58380 42420
rect 58470 42360 58500 42420
rect 58590 42360 58620 42420
rect 58710 42360 58740 42420
rect 58830 42360 58860 42420
rect 58950 42360 58980 42420
rect 59070 42360 59100 42420
rect 59190 42360 59220 42420
rect 59310 42360 59340 42420
rect 59430 42360 59460 42420
rect 59550 42360 59580 42420
rect 59670 42360 59700 42420
rect 59790 42360 59820 42420
rect 59910 42360 59940 42420
rect 60030 42360 60060 42420
rect 60150 42360 60180 42420
rect 60440 42360 60450 42440
rect 62140 42360 62150 42440
rect 62370 42360 62400 42420
rect 62490 42360 62520 42420
rect 62610 42360 62640 42420
rect 62730 42360 62760 42420
rect 62850 42360 62880 42420
rect 62970 42360 63000 42420
rect 63090 42360 63120 42420
rect 63210 42360 63240 42420
rect 63330 42360 63360 42420
rect 63450 42360 63480 42420
rect 63570 42360 63600 42420
rect 63690 42360 63720 42420
rect 63810 42360 63840 42420
rect 63930 42360 63960 42420
rect 64050 42360 64080 42420
rect 64170 42360 64200 42420
rect 64290 42360 64320 42420
rect 64410 42360 64440 42420
rect 64530 42360 64560 42420
rect 64650 42360 64680 42420
rect 64770 42360 64800 42420
rect 64890 42360 64920 42420
rect 65010 42360 65040 42420
rect 65130 42360 65160 42420
rect 65250 42360 65280 42420
rect 65370 42360 65400 42420
rect 65490 42360 65520 42420
rect 65610 42360 65640 42420
rect 65730 42360 65760 42420
rect 65850 42360 65880 42420
rect 65970 42360 66000 42420
rect 66090 42360 66120 42420
rect 66210 42360 66240 42420
rect 66330 42360 66360 42420
rect 66450 42360 66480 42420
rect 66570 42360 66600 42420
rect 66690 42360 66720 42420
rect 66810 42360 66840 42420
rect 66930 42360 66960 42420
rect 67050 42360 67080 42420
rect 67170 42360 67200 42420
rect 67290 42360 67320 42420
rect 67410 42360 67440 42420
rect 67530 42360 67560 42420
rect 67650 42360 67680 42420
rect 67770 42360 67800 42420
rect 67890 42360 67920 42420
rect 68010 42360 68040 42420
rect 68130 42360 68160 42420
rect 68250 42360 68280 42420
rect 68370 42360 68400 42420
rect 68490 42360 68520 42420
rect 68610 42360 68640 42420
rect 68730 42360 68760 42420
rect 68850 42360 68880 42420
rect 73290 42360 73320 42420
rect 73410 42360 73440 42420
rect 73530 42360 73560 42420
rect 73650 42360 73680 42420
rect 73940 42360 73950 42440
rect 75640 42360 75650 42440
rect 75870 42360 75900 42420
rect 75990 42360 76020 42420
rect 76110 42360 76140 42420
rect 76230 42360 76255 42420
rect 86790 42360 86820 42420
rect 86910 42360 86940 42420
rect 87030 42360 87060 42420
rect 87150 42360 87180 42420
rect 87440 42360 87450 42440
rect 89140 42360 89150 42440
rect 89370 42360 89400 42420
rect 89490 42360 89520 42420
rect 89610 42360 89640 42420
rect 89730 42360 89755 42420
rect 100290 42360 100320 42420
rect 100410 42360 100440 42420
rect 100530 42360 100560 42420
rect 100650 42360 100680 42420
rect 100940 42360 100950 42440
rect 102640 42360 102650 42440
rect 102870 42360 102900 42420
rect 102990 42360 103020 42420
rect 103110 42360 103140 42420
rect 103230 42360 103255 42420
rect 113790 42360 113820 42420
rect 113910 42360 113940 42420
rect 114030 42360 114060 42420
rect 114150 42360 114180 42420
rect 114440 42360 114450 42440
rect 116140 42360 116150 42440
rect 116370 42360 116400 42420
rect 116490 42360 116520 42420
rect 116610 42360 116640 42420
rect 116730 42360 116755 42420
rect 127290 42360 127320 42420
rect 127410 42360 127440 42420
rect 127530 42360 127560 42420
rect 127650 42360 127680 42420
rect 127940 42360 127950 42440
rect 129640 42360 129650 42440
rect 129870 42360 129900 42420
rect 129990 42360 130020 42420
rect 130110 42360 130140 42420
rect 130230 42360 130255 42420
rect 140910 42360 140940 42420
rect 141030 42360 141060 42420
rect 141150 42360 141180 42420
rect 141440 42360 141450 42440
rect 141565 42300 141620 43960
rect 146480 43895 146490 43975
rect 146800 43895 146810 43975
rect 147120 43895 147130 43975
rect 147440 43895 147450 43975
rect 148860 43895 148870 43975
rect 149180 43895 149190 43975
rect 149500 43895 149510 43975
rect 149820 43895 149830 43975
rect 152280 43895 152290 43975
rect 152600 43895 152610 43975
rect 152920 43895 152930 43975
rect 153240 43895 153250 43975
rect 153560 43895 153570 43975
rect 153880 43895 153890 43975
rect 154200 43895 154210 43975
rect 154520 43895 154530 43975
rect 154840 43895 154850 43975
rect 155160 43895 155170 43975
rect 155480 43895 155490 43975
rect 155800 43895 155810 43975
rect 156120 43895 156130 43975
rect 156440 43895 156450 43975
rect 156760 43895 156770 43975
rect 157080 43895 157090 43975
rect 157400 43895 157410 43975
rect 157720 43895 157730 43975
rect 158040 43895 158050 43975
rect 158360 43895 158370 43975
rect 158680 43895 158690 43975
rect 159000 43895 159010 43975
rect 159320 43895 159330 43975
rect 159640 43895 159650 43975
rect 163670 43935 163680 44015
rect 163990 43935 164000 44015
rect 164310 43935 164320 44015
rect 164630 43935 164640 44015
rect 164950 43935 164960 44015
rect 165270 43935 165280 44015
rect 165590 43935 165600 44015
rect 165910 43935 165920 44015
rect 166230 43935 166240 44015
rect 166550 43935 166560 44015
rect 166870 43935 166880 44015
rect 167190 43935 167200 44015
rect 167510 43935 167520 44015
rect 167830 43935 167840 44015
rect 168150 43935 168160 44015
rect 168470 43935 168480 44015
rect 168790 43935 168800 44015
rect 169110 43935 169120 44015
rect 169430 43935 169440 44015
rect 169750 43935 169760 44015
rect 170070 43935 170080 44015
rect 170390 43935 170400 44015
rect 170710 43935 170720 44015
rect 171030 43935 171040 44015
rect 146220 43780 146300 43790
rect 146540 43780 146620 43790
rect 146860 43780 146940 43790
rect 147180 43780 147260 43790
rect 147500 43780 147580 43790
rect 146300 43700 146310 43780
rect 146620 43700 146630 43780
rect 146940 43700 146950 43780
rect 147260 43700 147270 43780
rect 147580 43700 147590 43780
rect 146380 43620 146460 43630
rect 146700 43620 146780 43630
rect 147020 43620 147100 43630
rect 147340 43620 147420 43630
rect 141665 43600 141745 43610
rect 141985 43600 142065 43610
rect 145200 43600 145265 43610
rect 145505 43600 145585 43610
rect 145825 43600 145905 43610
rect 146145 43600 146225 43610
rect 141745 43520 141755 43600
rect 142065 43520 142075 43600
rect 145265 43520 145275 43600
rect 145585 43520 145595 43600
rect 145905 43520 145915 43600
rect 146225 43550 146235 43600
rect 146145 43520 146235 43550
rect 146460 43540 146470 43620
rect 146780 43540 146790 43620
rect 147100 43540 147110 43620
rect 147420 43540 147430 43620
rect 146220 43460 146300 43470
rect 146540 43460 146620 43470
rect 146860 43460 146940 43470
rect 147180 43460 147260 43470
rect 147500 43460 147580 43470
rect 148780 43460 148860 43470
rect 149100 43460 149180 43470
rect 149420 43460 149500 43470
rect 149740 43460 149820 43470
rect 152300 43460 152380 43470
rect 152620 43460 152700 43470
rect 152940 43460 153020 43470
rect 153260 43460 153340 43470
rect 153580 43460 153660 43470
rect 153900 43460 153980 43470
rect 154220 43460 154300 43470
rect 154540 43460 154620 43470
rect 154860 43460 154940 43470
rect 155180 43460 155260 43470
rect 155500 43460 155580 43470
rect 155820 43460 155900 43470
rect 156140 43460 156220 43470
rect 156460 43460 156540 43470
rect 156780 43460 156860 43470
rect 157100 43460 157180 43470
rect 157420 43460 157500 43470
rect 157740 43460 157820 43470
rect 158060 43460 158140 43470
rect 158380 43460 158460 43470
rect 158700 43460 158780 43470
rect 159020 43460 159100 43470
rect 159340 43460 159420 43470
rect 163500 43460 163580 43470
rect 163820 43460 163900 43470
rect 164140 43460 164220 43470
rect 164460 43460 164540 43470
rect 164780 43460 164860 43470
rect 165100 43460 165180 43470
rect 165420 43460 165500 43470
rect 165740 43460 165820 43470
rect 166060 43460 166140 43470
rect 166380 43460 166460 43470
rect 166700 43460 166780 43470
rect 167020 43460 167100 43470
rect 167340 43460 167420 43470
rect 167660 43460 167740 43470
rect 167980 43460 168060 43470
rect 168300 43460 168380 43470
rect 168620 43460 168700 43470
rect 168940 43460 169020 43470
rect 169260 43460 169340 43470
rect 169580 43460 169660 43470
rect 169900 43460 169980 43470
rect 170220 43460 170300 43470
rect 170540 43460 170620 43470
rect 170860 43460 170940 43470
rect 141825 43440 141905 43450
rect 142145 43440 142200 43450
rect 145345 43440 145425 43450
rect 145665 43440 145745 43450
rect 145985 43440 146065 43450
rect 141905 43360 141915 43440
rect 145425 43360 145435 43440
rect 145745 43360 145755 43440
rect 146065 43360 146075 43440
rect 146300 43380 146310 43460
rect 146620 43380 146630 43460
rect 146940 43380 146950 43460
rect 147260 43380 147270 43460
rect 147580 43380 147590 43460
rect 148860 43380 148870 43460
rect 149180 43380 149190 43460
rect 149500 43380 149510 43460
rect 149820 43380 149830 43460
rect 152380 43380 152390 43460
rect 152700 43380 152710 43460
rect 153020 43380 153030 43460
rect 153340 43380 153350 43460
rect 153660 43380 153670 43460
rect 153980 43380 153990 43460
rect 154300 43380 154310 43460
rect 154620 43380 154630 43460
rect 154940 43380 154950 43460
rect 155260 43380 155270 43460
rect 155580 43380 155590 43460
rect 155900 43380 155910 43460
rect 156220 43380 156230 43460
rect 156540 43380 156550 43460
rect 156860 43380 156870 43460
rect 157180 43380 157190 43460
rect 157500 43380 157510 43460
rect 157820 43380 157830 43460
rect 158140 43380 158150 43460
rect 158460 43380 158470 43460
rect 158780 43380 158790 43460
rect 159100 43380 159110 43460
rect 159420 43380 159430 43460
rect 163580 43380 163590 43460
rect 163900 43380 163910 43460
rect 164220 43380 164230 43460
rect 164540 43380 164550 43460
rect 164860 43380 164870 43460
rect 165180 43380 165190 43460
rect 165500 43380 165510 43460
rect 165820 43380 165830 43460
rect 166140 43380 166150 43460
rect 166460 43380 166470 43460
rect 166780 43380 166790 43460
rect 167100 43380 167110 43460
rect 167420 43380 167430 43460
rect 167740 43380 167750 43460
rect 168060 43380 168070 43460
rect 168380 43380 168390 43460
rect 168700 43380 168710 43460
rect 169020 43380 169030 43460
rect 169340 43380 169350 43460
rect 169660 43380 169670 43460
rect 169980 43380 169990 43460
rect 170300 43380 170310 43460
rect 170620 43380 170630 43460
rect 170940 43380 170950 43460
rect 146380 43300 146460 43310
rect 146700 43300 146780 43310
rect 147020 43300 147100 43310
rect 147340 43300 147420 43310
rect 148940 43300 149020 43310
rect 149260 43300 149340 43310
rect 149580 43300 149660 43310
rect 152460 43300 152540 43310
rect 152780 43300 152860 43310
rect 153100 43300 153180 43310
rect 153420 43300 153500 43310
rect 153740 43300 153820 43310
rect 154060 43300 154140 43310
rect 154380 43300 154460 43310
rect 154700 43300 154780 43310
rect 155020 43300 155100 43310
rect 155340 43300 155420 43310
rect 155660 43300 155740 43310
rect 155980 43300 156060 43310
rect 156300 43300 156380 43310
rect 156620 43300 156700 43310
rect 156940 43300 157020 43310
rect 157260 43300 157340 43310
rect 157580 43300 157660 43310
rect 157900 43300 157980 43310
rect 158220 43300 158300 43310
rect 158540 43300 158620 43310
rect 158860 43300 158940 43310
rect 159180 43300 159260 43310
rect 159500 43300 159580 43310
rect 163660 43300 163740 43310
rect 163980 43300 164060 43310
rect 164300 43300 164380 43310
rect 164620 43300 164700 43310
rect 164940 43300 165020 43310
rect 165260 43300 165340 43310
rect 165580 43300 165660 43310
rect 165900 43300 165980 43310
rect 166220 43300 166300 43310
rect 166540 43300 166620 43310
rect 166860 43300 166940 43310
rect 167180 43300 167260 43310
rect 167500 43300 167580 43310
rect 167820 43300 167900 43310
rect 168140 43300 168220 43310
rect 168460 43300 168540 43310
rect 168780 43300 168860 43310
rect 169100 43300 169180 43310
rect 169420 43300 169500 43310
rect 169740 43300 169820 43310
rect 170060 43300 170140 43310
rect 170380 43300 170460 43310
rect 170700 43300 170780 43310
rect 141665 43280 141745 43290
rect 141985 43280 142065 43290
rect 145200 43280 145265 43290
rect 145505 43280 145585 43290
rect 145825 43280 145905 43290
rect 146145 43280 146225 43290
rect 141745 43200 141755 43280
rect 142065 43200 142075 43280
rect 145265 43200 145275 43280
rect 145585 43200 145595 43280
rect 145905 43200 145915 43280
rect 146225 43230 146235 43280
rect 146145 43200 146235 43230
rect 146460 43220 146470 43300
rect 146780 43220 146790 43300
rect 147100 43220 147110 43300
rect 147420 43220 147430 43300
rect 149020 43220 149030 43300
rect 149340 43220 149350 43300
rect 149660 43220 149670 43300
rect 152540 43220 152550 43300
rect 152860 43220 152870 43300
rect 153180 43220 153190 43300
rect 153500 43220 153510 43300
rect 153820 43220 153830 43300
rect 154140 43220 154150 43300
rect 154460 43220 154470 43300
rect 154780 43220 154790 43300
rect 155100 43220 155110 43300
rect 155420 43220 155430 43300
rect 155740 43220 155750 43300
rect 156060 43220 156070 43300
rect 156380 43220 156390 43300
rect 156700 43220 156710 43300
rect 157020 43220 157030 43300
rect 157340 43220 157350 43300
rect 157660 43220 157670 43300
rect 157980 43220 157990 43300
rect 158300 43220 158310 43300
rect 158620 43220 158630 43300
rect 158940 43220 158950 43300
rect 159260 43220 159270 43300
rect 159580 43220 159590 43300
rect 163740 43220 163750 43300
rect 164060 43220 164070 43300
rect 164380 43220 164390 43300
rect 164700 43220 164710 43300
rect 165020 43220 165030 43300
rect 165340 43220 165350 43300
rect 165660 43220 165670 43300
rect 165980 43220 165990 43300
rect 166300 43220 166310 43300
rect 166620 43220 166630 43300
rect 166940 43220 166950 43300
rect 167260 43220 167270 43300
rect 167580 43220 167590 43300
rect 167900 43220 167910 43300
rect 168220 43220 168230 43300
rect 168540 43220 168550 43300
rect 168860 43220 168870 43300
rect 169180 43220 169190 43300
rect 169500 43220 169510 43300
rect 169820 43220 169830 43300
rect 170140 43220 170150 43300
rect 170460 43220 170470 43300
rect 170780 43220 170790 43300
rect 146220 43140 146300 43150
rect 146540 43140 146620 43150
rect 146860 43140 146940 43150
rect 147180 43140 147260 43150
rect 147500 43140 147580 43150
rect 148780 43140 148860 43150
rect 149100 43140 149180 43150
rect 149420 43140 149500 43150
rect 149740 43140 149820 43150
rect 152300 43140 152380 43150
rect 152620 43140 152700 43150
rect 152940 43140 153020 43150
rect 153260 43140 153340 43150
rect 153580 43140 153660 43150
rect 153900 43140 153980 43150
rect 154220 43140 154300 43150
rect 154540 43140 154620 43150
rect 154860 43140 154940 43150
rect 155180 43140 155260 43150
rect 155500 43140 155580 43150
rect 155820 43140 155900 43150
rect 156140 43140 156220 43150
rect 156460 43140 156540 43150
rect 156780 43140 156860 43150
rect 157100 43140 157180 43150
rect 157420 43140 157500 43150
rect 157740 43140 157820 43150
rect 158060 43140 158140 43150
rect 158380 43140 158460 43150
rect 158700 43140 158780 43150
rect 159020 43140 159100 43150
rect 159340 43140 159420 43150
rect 163500 43140 163580 43150
rect 163820 43140 163900 43150
rect 164140 43140 164220 43150
rect 164460 43140 164540 43150
rect 164780 43140 164860 43150
rect 165100 43140 165180 43150
rect 165420 43140 165500 43150
rect 165740 43140 165820 43150
rect 166060 43140 166140 43150
rect 166380 43140 166460 43150
rect 166700 43140 166780 43150
rect 167020 43140 167100 43150
rect 167340 43140 167420 43150
rect 167660 43140 167740 43150
rect 167980 43140 168060 43150
rect 168300 43140 168380 43150
rect 168620 43140 168700 43150
rect 168940 43140 169020 43150
rect 169260 43140 169340 43150
rect 169580 43140 169660 43150
rect 169900 43140 169980 43150
rect 170220 43140 170300 43150
rect 170540 43140 170620 43150
rect 170860 43140 170940 43150
rect 141825 43120 141905 43130
rect 142145 43120 142200 43130
rect 145345 43120 145425 43130
rect 145665 43120 145745 43130
rect 145985 43120 146065 43130
rect 141905 43040 141915 43120
rect 145425 43040 145435 43120
rect 145745 43040 145755 43120
rect 146065 43040 146075 43120
rect 146300 43060 146310 43140
rect 146620 43060 146630 43140
rect 146940 43060 146950 43140
rect 147260 43060 147270 43140
rect 147580 43060 147590 43140
rect 148860 43060 148870 43140
rect 149180 43060 149190 43140
rect 149500 43060 149510 43140
rect 149820 43060 149830 43140
rect 152380 43060 152390 43140
rect 152700 43060 152710 43140
rect 153020 43060 153030 43140
rect 153340 43060 153350 43140
rect 153660 43060 153670 43140
rect 153980 43060 153990 43140
rect 154300 43060 154310 43140
rect 154620 43060 154630 43140
rect 154940 43060 154950 43140
rect 155260 43060 155270 43140
rect 155580 43060 155590 43140
rect 155900 43060 155910 43140
rect 156220 43060 156230 43140
rect 156540 43060 156550 43140
rect 156860 43060 156870 43140
rect 157180 43060 157190 43140
rect 157500 43060 157510 43140
rect 157820 43060 157830 43140
rect 158140 43060 158150 43140
rect 158460 43060 158470 43140
rect 158780 43060 158790 43140
rect 159100 43060 159110 43140
rect 159420 43060 159430 43140
rect 163580 43060 163590 43140
rect 163900 43060 163910 43140
rect 164220 43060 164230 43140
rect 164540 43060 164550 43140
rect 164860 43060 164870 43140
rect 165180 43060 165190 43140
rect 165500 43060 165510 43140
rect 165820 43060 165830 43140
rect 166140 43060 166150 43140
rect 166460 43060 166470 43140
rect 166780 43060 166790 43140
rect 167100 43060 167110 43140
rect 167420 43060 167430 43140
rect 167740 43060 167750 43140
rect 168060 43060 168070 43140
rect 168380 43060 168390 43140
rect 168700 43060 168710 43140
rect 169020 43060 169030 43140
rect 169340 43060 169350 43140
rect 169660 43060 169670 43140
rect 169980 43060 169990 43140
rect 170300 43060 170310 43140
rect 170620 43060 170630 43140
rect 170940 43060 170950 43140
rect 146380 42980 146460 42990
rect 146700 42980 146780 42990
rect 147020 42980 147100 42990
rect 147340 42980 147420 42990
rect 148940 42980 149020 42990
rect 149260 42980 149340 42990
rect 149580 42980 149660 42990
rect 152460 42980 152540 42990
rect 152780 42980 152860 42990
rect 153100 42980 153180 42990
rect 153420 42980 153500 42990
rect 153740 42980 153820 42990
rect 154060 42980 154140 42990
rect 154380 42980 154460 42990
rect 154700 42980 154780 42990
rect 155020 42980 155100 42990
rect 155340 42980 155420 42990
rect 155660 42980 155740 42990
rect 155980 42980 156000 42990
rect 141665 42960 141745 42970
rect 141985 42960 142065 42970
rect 145200 42960 145265 42970
rect 145505 42960 145585 42970
rect 145825 42960 145905 42970
rect 146145 42960 146225 42970
rect 141745 42880 141755 42960
rect 142065 42880 142075 42960
rect 145265 42880 145275 42960
rect 145585 42880 145595 42960
rect 145905 42880 145915 42960
rect 146225 42910 146235 42960
rect 146145 42880 146235 42910
rect 146460 42900 146470 42980
rect 146780 42900 146790 42980
rect 147100 42900 147110 42980
rect 147420 42900 147430 42980
rect 149020 42900 149030 42980
rect 149340 42900 149350 42980
rect 149660 42900 149670 42980
rect 152540 42900 152550 42980
rect 152860 42900 152870 42980
rect 153180 42900 153190 42980
rect 153500 42900 153510 42980
rect 153820 42900 153830 42980
rect 154140 42900 154150 42980
rect 154460 42900 154470 42980
rect 154780 42900 154790 42980
rect 155100 42900 155110 42980
rect 155420 42900 155430 42980
rect 155740 42900 155750 42980
rect 146220 42820 146300 42830
rect 146540 42820 146620 42830
rect 146860 42820 146940 42830
rect 147180 42820 147260 42830
rect 148780 42820 148860 42830
rect 149100 42820 149180 42830
rect 149420 42820 149500 42830
rect 149740 42820 149820 42830
rect 152300 42820 152380 42830
rect 152620 42820 152700 42830
rect 152940 42820 153020 42830
rect 153260 42820 153340 42830
rect 153580 42820 153660 42830
rect 153900 42820 153980 42830
rect 154220 42820 154300 42830
rect 154540 42820 154620 42830
rect 154860 42820 154940 42830
rect 155180 42820 155260 42830
rect 155500 42820 155580 42830
rect 155820 42820 155900 42830
rect 141825 42800 141905 42810
rect 142145 42800 142200 42810
rect 145345 42800 145425 42810
rect 145665 42800 145745 42810
rect 145985 42800 146065 42810
rect 141905 42720 141915 42800
rect 145425 42720 145435 42800
rect 145745 42720 145755 42800
rect 146065 42720 146075 42800
rect 146300 42740 146310 42820
rect 146620 42740 146630 42820
rect 146940 42740 146950 42820
rect 147260 42740 147270 42820
rect 148860 42740 148870 42820
rect 149180 42740 149190 42820
rect 149500 42740 149510 42820
rect 149820 42740 149830 42820
rect 152380 42740 152390 42820
rect 152700 42740 152710 42820
rect 153020 42740 153030 42820
rect 153340 42740 153350 42820
rect 153660 42740 153670 42820
rect 153980 42740 153990 42820
rect 154300 42740 154310 42820
rect 154620 42740 154630 42820
rect 154940 42740 154950 42820
rect 155260 42740 155270 42820
rect 155580 42740 155590 42820
rect 155900 42740 155910 42820
rect 146380 42660 146460 42670
rect 146700 42660 146780 42670
rect 147020 42660 147100 42670
rect 148940 42660 149020 42670
rect 149260 42660 149340 42670
rect 149580 42660 149660 42670
rect 152460 42660 152540 42670
rect 152780 42660 152860 42670
rect 153100 42660 153180 42670
rect 153420 42660 153500 42670
rect 153740 42660 153820 42670
rect 154060 42660 154140 42670
rect 154380 42660 154460 42670
rect 154700 42660 154780 42670
rect 155020 42660 155100 42670
rect 155340 42660 155420 42670
rect 155660 42660 155740 42670
rect 155980 42660 156000 42670
rect 141665 42640 141745 42650
rect 141985 42640 142065 42650
rect 145200 42640 145265 42650
rect 145505 42640 145585 42650
rect 145825 42640 145905 42650
rect 146145 42640 146225 42650
rect 141745 42560 141755 42640
rect 142065 42560 142075 42640
rect 145265 42560 145275 42640
rect 145585 42560 145595 42640
rect 145905 42560 145915 42640
rect 146225 42590 146235 42640
rect 146145 42560 146235 42590
rect 146460 42580 146470 42660
rect 146780 42580 146790 42660
rect 147100 42580 147110 42660
rect 149020 42580 149030 42660
rect 149340 42580 149350 42660
rect 149660 42580 149670 42660
rect 152540 42580 152550 42660
rect 152860 42580 152870 42660
rect 153180 42580 153190 42660
rect 153500 42580 153510 42660
rect 153820 42580 153830 42660
rect 154140 42580 154150 42660
rect 154460 42580 154470 42660
rect 154780 42580 154790 42660
rect 155100 42580 155110 42660
rect 155420 42580 155430 42660
rect 155740 42580 155750 42660
rect 146220 42500 146300 42510
rect 146540 42500 146620 42510
rect 146860 42500 146940 42510
rect 148780 42500 148860 42510
rect 149100 42500 149180 42510
rect 149420 42500 149500 42510
rect 149740 42500 149820 42510
rect 152300 42500 152380 42510
rect 152620 42500 152700 42510
rect 152940 42500 153020 42510
rect 153260 42500 153340 42510
rect 153580 42500 153660 42510
rect 153900 42500 153980 42510
rect 154220 42500 154300 42510
rect 154540 42500 154620 42510
rect 154860 42500 154940 42510
rect 155180 42500 155260 42510
rect 155500 42500 155580 42510
rect 155820 42500 155900 42510
rect 146300 42420 146310 42500
rect 146620 42420 146630 42500
rect 146940 42420 146950 42500
rect 148860 42420 148870 42500
rect 149180 42420 149190 42500
rect 149500 42420 149510 42500
rect 149820 42420 149830 42500
rect 152380 42420 152390 42500
rect 152700 42420 152710 42500
rect 153020 42420 153030 42500
rect 153340 42420 153350 42500
rect 153660 42420 153670 42500
rect 153980 42420 153990 42500
rect 154300 42420 154310 42500
rect 154620 42420 154630 42500
rect 154940 42420 154950 42500
rect 155260 42420 155270 42500
rect 155580 42420 155590 42500
rect 155900 42420 155910 42500
rect 148940 42340 149020 42350
rect 149260 42340 149340 42350
rect 149580 42340 149660 42350
rect 152460 42340 152540 42350
rect 152780 42340 152860 42350
rect 153100 42340 153180 42350
rect 153420 42340 153500 42350
rect 153740 42340 153820 42350
rect 154060 42340 154140 42350
rect 154380 42340 154460 42350
rect 154700 42340 154780 42350
rect 155020 42340 155100 42350
rect 155340 42340 155420 42350
rect 155660 42340 155740 42350
rect 155980 42340 156000 42350
rect 149020 42260 149030 42340
rect 149340 42260 149350 42340
rect 149660 42260 149670 42340
rect 152540 42260 152550 42340
rect 152860 42260 152870 42340
rect 153180 42260 153190 42340
rect 153500 42260 153510 42340
rect 153820 42260 153830 42340
rect 154140 42260 154150 42340
rect 154460 42260 154470 42340
rect 154780 42260 154790 42340
rect 155100 42260 155110 42340
rect 155420 42260 155430 42340
rect 155740 42260 155750 42340
rect 36020 42180 36100 42190
rect 36340 42180 36420 42190
rect 36660 42180 36740 42190
rect 36980 42180 37060 42190
rect 37300 42180 37380 42190
rect 37620 42180 37700 42190
rect 40180 42180 40260 42190
rect 40500 42180 40580 42190
rect 40820 42180 40900 42190
rect 41140 42180 41220 42190
rect 148780 42180 148860 42190
rect 149100 42180 149180 42190
rect 149420 42180 149500 42190
rect 149740 42180 149820 42190
rect 152300 42180 152380 42190
rect 152620 42180 152700 42190
rect 152940 42180 153020 42190
rect 153260 42180 153340 42190
rect 153580 42180 153660 42190
rect 153900 42180 153980 42190
rect 154220 42180 154300 42190
rect 154540 42180 154620 42190
rect 154860 42180 154940 42190
rect 155180 42180 155260 42190
rect 155500 42180 155580 42190
rect 155820 42180 155900 42190
rect 36100 42100 36110 42180
rect 36420 42100 36430 42180
rect 36740 42100 36750 42180
rect 37060 42100 37070 42180
rect 37380 42100 37390 42180
rect 37700 42100 37710 42180
rect 40260 42100 40270 42180
rect 40580 42100 40590 42180
rect 40900 42100 40910 42180
rect 41220 42100 41230 42180
rect 148860 42100 148870 42180
rect 149180 42100 149190 42180
rect 149500 42100 149510 42180
rect 149820 42100 149830 42180
rect 152380 42100 152390 42180
rect 152700 42100 152710 42180
rect 153020 42100 153030 42180
rect 153340 42100 153350 42180
rect 153660 42100 153670 42180
rect 153980 42100 153990 42180
rect 154300 42100 154310 42180
rect 154620 42100 154630 42180
rect 154940 42100 154950 42180
rect 155260 42100 155270 42180
rect 155580 42100 155590 42180
rect 155900 42100 155910 42180
rect 36180 42020 36260 42030
rect 36500 42020 36580 42030
rect 36820 42020 36900 42030
rect 37140 42020 37220 42030
rect 37460 42020 37540 42030
rect 40340 42020 40420 42030
rect 40660 42020 40740 42030
rect 40980 42020 41060 42030
rect 41300 42020 41380 42030
rect 148620 42020 148700 42030
rect 148940 42020 149020 42030
rect 149260 42020 149340 42030
rect 149580 42020 149660 42030
rect 152460 42020 152540 42030
rect 152780 42020 152860 42030
rect 153100 42020 153180 42030
rect 153420 42020 153500 42030
rect 153740 42020 153820 42030
rect 154060 42020 154140 42030
rect 154380 42020 154460 42030
rect 154700 42020 154780 42030
rect 155020 42020 155100 42030
rect 155340 42020 155420 42030
rect 155660 42020 155740 42030
rect 155980 42020 156000 42030
rect 36260 41940 36270 42020
rect 36580 41940 36590 42020
rect 36900 41940 36910 42020
rect 37220 41940 37230 42020
rect 37540 41940 37550 42020
rect 40420 41940 40430 42020
rect 40740 41940 40750 42020
rect 41060 41940 41070 42020
rect 41380 41940 41390 42020
rect 148700 41940 148710 42020
rect 149020 41940 149030 42020
rect 149340 41940 149350 42020
rect 149660 41940 149670 42020
rect 152540 41940 152550 42020
rect 152860 41940 152870 42020
rect 153180 41940 153190 42020
rect 153500 41940 153510 42020
rect 153820 41940 153830 42020
rect 154140 41940 154150 42020
rect 154460 41940 154470 42020
rect 154780 41940 154790 42020
rect 155100 41940 155110 42020
rect 155420 41940 155430 42020
rect 155740 41940 155750 42020
rect 36020 41860 36100 41870
rect 36340 41860 36420 41870
rect 36660 41860 36740 41870
rect 36980 41860 37060 41870
rect 37300 41860 37380 41870
rect 37620 41860 37700 41870
rect 40180 41860 40260 41870
rect 40500 41860 40580 41870
rect 40820 41860 40900 41870
rect 41140 41860 41220 41870
rect 41460 41860 41540 41870
rect 148460 41860 148540 41870
rect 148780 41860 148860 41870
rect 149100 41860 149180 41870
rect 149420 41860 149500 41870
rect 149740 41860 149820 41870
rect 152300 41860 152380 41870
rect 152620 41860 152700 41870
rect 152940 41860 153020 41870
rect 153260 41860 153340 41870
rect 153580 41860 153660 41870
rect 153900 41860 153980 41870
rect 154220 41860 154300 41870
rect 154540 41860 154620 41870
rect 154860 41860 154940 41870
rect 155180 41860 155260 41870
rect 155500 41860 155580 41870
rect 155820 41860 155900 41870
rect 36100 41780 36110 41860
rect 36420 41780 36430 41860
rect 36740 41780 36750 41860
rect 37060 41780 37070 41860
rect 37380 41780 37390 41860
rect 37700 41780 37710 41860
rect 40260 41780 40270 41860
rect 40580 41780 40590 41860
rect 40900 41780 40910 41860
rect 41220 41780 41230 41860
rect 41540 41780 41550 41860
rect 148540 41780 148550 41860
rect 148860 41780 148870 41860
rect 149180 41780 149190 41860
rect 149500 41780 149510 41860
rect 149820 41780 149830 41860
rect 152380 41780 152390 41860
rect 152700 41780 152710 41860
rect 153020 41780 153030 41860
rect 153340 41780 153350 41860
rect 153660 41780 153670 41860
rect 153980 41780 153990 41860
rect 154300 41780 154310 41860
rect 154620 41780 154630 41860
rect 154940 41780 154950 41860
rect 155260 41780 155270 41860
rect 155580 41780 155590 41860
rect 155900 41780 155910 41860
rect 36180 41700 36260 41710
rect 36500 41700 36580 41710
rect 36820 41700 36900 41710
rect 37140 41700 37220 41710
rect 37460 41700 37540 41710
rect 40340 41700 40420 41710
rect 40660 41700 40740 41710
rect 40980 41700 41060 41710
rect 41300 41700 41380 41710
rect 41620 41700 41700 41710
rect 148300 41700 148380 41710
rect 148620 41700 148700 41710
rect 148940 41700 149020 41710
rect 149260 41700 149340 41710
rect 149580 41700 149660 41710
rect 152460 41700 152540 41710
rect 152780 41700 152860 41710
rect 153100 41700 153180 41710
rect 153420 41700 153500 41710
rect 153740 41700 153820 41710
rect 154060 41700 154140 41710
rect 154380 41700 154460 41710
rect 154700 41700 154780 41710
rect 155020 41700 155100 41710
rect 155340 41700 155420 41710
rect 155660 41700 155740 41710
rect 155980 41700 156000 41710
rect 36260 41620 36270 41700
rect 36580 41620 36590 41700
rect 36900 41620 36910 41700
rect 37220 41620 37230 41700
rect 37540 41620 37550 41700
rect 40420 41620 40430 41700
rect 40740 41620 40750 41700
rect 41060 41620 41070 41700
rect 41380 41620 41390 41700
rect 41700 41620 41710 41700
rect 36020 41540 36100 41550
rect 36340 41540 36420 41550
rect 36660 41540 36740 41550
rect 36980 41540 37060 41550
rect 37300 41540 37380 41550
rect 37620 41540 37700 41550
rect 40180 41540 40260 41550
rect 40500 41540 40580 41550
rect 40820 41540 40900 41550
rect 41140 41540 41220 41550
rect 41460 41540 41540 41550
rect 41780 41540 41860 41550
rect 36100 41460 36110 41540
rect 36420 41460 36430 41540
rect 36740 41460 36750 41540
rect 37060 41460 37070 41540
rect 37380 41460 37390 41540
rect 37700 41460 37710 41540
rect 40260 41460 40270 41540
rect 40580 41460 40590 41540
rect 40900 41460 40910 41540
rect 41220 41460 41230 41540
rect 41540 41460 41550 41540
rect 41860 41460 41870 41540
rect 48500 41410 48605 41660
rect 48870 41540 48900 41600
rect 48990 41540 49020 41600
rect 49110 41540 49140 41600
rect 49230 41540 49260 41600
rect 49350 41540 49380 41600
rect 49470 41540 49500 41600
rect 49590 41540 49620 41600
rect 49710 41540 49740 41600
rect 49830 41540 49860 41600
rect 49950 41540 49980 41600
rect 50070 41540 50100 41600
rect 50190 41540 50220 41600
rect 50310 41540 50340 41600
rect 50430 41540 50460 41600
rect 50550 41540 50580 41600
rect 50670 41540 50700 41600
rect 50790 41540 50820 41600
rect 50910 41540 50940 41600
rect 51030 41540 51060 41600
rect 51150 41540 51180 41600
rect 51270 41540 51300 41600
rect 51390 41540 51420 41600
rect 51510 41540 51540 41600
rect 51630 41540 51660 41600
rect 51750 41540 51780 41600
rect 51870 41540 51900 41600
rect 51990 41540 52020 41600
rect 52110 41540 52140 41600
rect 52230 41540 52260 41600
rect 52350 41540 52380 41600
rect 52470 41540 52500 41600
rect 52590 41540 52620 41600
rect 52710 41540 52740 41600
rect 52830 41540 52860 41600
rect 52950 41540 52980 41600
rect 53070 41540 53100 41600
rect 53190 41540 53220 41600
rect 53310 41540 53340 41600
rect 53430 41540 53460 41600
rect 53550 41540 53580 41600
rect 53670 41540 53700 41600
rect 53790 41540 53820 41600
rect 53910 41540 53940 41600
rect 54030 41540 54060 41600
rect 54150 41540 54180 41600
rect 54270 41540 54300 41600
rect 54390 41540 54420 41600
rect 54510 41540 54540 41600
rect 54630 41540 54660 41600
rect 54750 41540 54780 41600
rect 54870 41540 54900 41600
rect 54990 41540 55020 41600
rect 55110 41540 55140 41600
rect 55230 41540 55260 41600
rect 55350 41540 55380 41600
rect 55470 41540 55500 41600
rect 55590 41540 55620 41600
rect 55710 41540 55740 41600
rect 55830 41540 55860 41600
rect 55950 41540 55980 41600
rect 56070 41540 56100 41600
rect 56190 41540 56220 41600
rect 56310 41540 56340 41600
rect 56430 41540 56460 41600
rect 56550 41540 56580 41600
rect 56670 41540 56700 41600
rect 56790 41540 56820 41600
rect 56910 41540 56940 41600
rect 57030 41540 57060 41600
rect 57150 41540 57180 41600
rect 57270 41540 57300 41600
rect 57390 41540 57420 41600
rect 57510 41540 57540 41600
rect 57630 41540 57660 41600
rect 57750 41540 57780 41600
rect 57870 41540 57900 41600
rect 57990 41540 58020 41600
rect 58110 41540 58140 41600
rect 58230 41540 58260 41600
rect 58350 41540 58380 41600
rect 58470 41540 58500 41600
rect 58590 41540 58620 41600
rect 58710 41540 58740 41600
rect 58830 41540 58860 41600
rect 58950 41540 58980 41600
rect 59070 41540 59100 41600
rect 59190 41540 59220 41600
rect 59310 41540 59340 41600
rect 59430 41540 59460 41600
rect 59550 41540 59580 41600
rect 59670 41540 59700 41600
rect 59790 41540 59820 41600
rect 59910 41540 59940 41600
rect 60030 41540 60060 41600
rect 60150 41540 60180 41600
rect 62370 41540 62400 41600
rect 62490 41540 62520 41600
rect 62610 41540 62640 41600
rect 62730 41540 62760 41600
rect 62850 41540 62880 41600
rect 62970 41540 63000 41600
rect 63090 41540 63120 41600
rect 63210 41540 63240 41600
rect 63330 41540 63360 41600
rect 63450 41540 63480 41600
rect 63570 41540 63600 41600
rect 63690 41540 63720 41600
rect 63810 41540 63840 41600
rect 63930 41540 63960 41600
rect 64050 41540 64080 41600
rect 64170 41540 64200 41600
rect 64290 41540 64320 41600
rect 64410 41540 64440 41600
rect 64530 41540 64560 41600
rect 64650 41540 64680 41600
rect 64770 41540 64800 41600
rect 64890 41540 64920 41600
rect 65010 41540 65040 41600
rect 65130 41540 65160 41600
rect 65250 41540 65280 41600
rect 65370 41540 65400 41600
rect 65490 41540 65520 41600
rect 65610 41540 65640 41600
rect 65730 41540 65760 41600
rect 65850 41540 65880 41600
rect 65970 41540 66000 41600
rect 66090 41540 66120 41600
rect 66210 41540 66240 41600
rect 66330 41540 66360 41600
rect 66450 41540 66480 41600
rect 66570 41540 66600 41600
rect 66690 41540 66720 41600
rect 66810 41540 66840 41600
rect 66930 41540 66960 41600
rect 67050 41540 67080 41600
rect 67170 41540 67200 41600
rect 67290 41540 67320 41600
rect 67410 41540 67440 41600
rect 67530 41540 67560 41600
rect 67650 41540 67680 41600
rect 67770 41540 67800 41600
rect 67890 41540 67920 41600
rect 68010 41540 68040 41600
rect 68130 41540 68160 41600
rect 68250 41540 68280 41600
rect 68370 41540 68400 41600
rect 68490 41540 68520 41600
rect 68610 41540 68640 41600
rect 68730 41540 68760 41600
rect 68850 41540 68880 41600
rect 73290 41540 73320 41600
rect 73410 41540 73440 41600
rect 73530 41540 73560 41600
rect 73650 41540 73680 41600
rect 75870 41540 75900 41600
rect 75990 41540 76020 41600
rect 76110 41540 76140 41600
rect 76230 41540 76255 41600
rect 86790 41540 86820 41600
rect 86910 41540 86940 41600
rect 87030 41540 87060 41600
rect 87150 41540 87180 41600
rect 89370 41540 89400 41600
rect 89490 41540 89520 41600
rect 89610 41540 89640 41600
rect 89730 41540 89755 41600
rect 100290 41540 100320 41600
rect 100410 41540 100440 41600
rect 100530 41540 100560 41600
rect 100650 41540 100680 41600
rect 102870 41540 102900 41600
rect 102990 41540 103020 41600
rect 103110 41540 103140 41600
rect 103230 41540 103255 41600
rect 113790 41540 113820 41600
rect 113910 41540 113940 41600
rect 114030 41540 114060 41600
rect 114150 41540 114180 41600
rect 116370 41540 116400 41600
rect 116490 41540 116520 41600
rect 116610 41540 116640 41600
rect 116730 41540 116755 41600
rect 127290 41540 127320 41600
rect 127410 41540 127440 41600
rect 127530 41540 127560 41600
rect 127650 41540 127680 41600
rect 129870 41540 129900 41600
rect 129990 41540 130020 41600
rect 130110 41540 130140 41600
rect 130230 41540 130255 41600
rect 140910 41540 140940 41600
rect 141030 41540 141060 41600
rect 141150 41540 141180 41600
rect 57110 41480 57910 41490
rect 58130 41480 59990 41490
rect 73245 41480 73490 41490
rect 86745 41480 86990 41490
rect 100245 41480 100490 41490
rect 113745 41480 113990 41490
rect 127245 41480 127490 41490
rect 140830 41480 140990 41490
rect 48500 41400 48640 41410
rect 36180 41380 36260 41390
rect 36500 41380 36580 41390
rect 36820 41380 36900 41390
rect 37140 41380 37220 41390
rect 37460 41380 37540 41390
rect 40340 41380 40420 41390
rect 40660 41380 40740 41390
rect 40980 41380 41060 41390
rect 41300 41380 41380 41390
rect 41620 41380 41700 41390
rect 41940 41380 42020 41390
rect 36260 41300 36270 41380
rect 36580 41300 36590 41380
rect 36900 41300 36910 41380
rect 37220 41300 37230 41380
rect 37540 41300 37550 41380
rect 40420 41300 40430 41380
rect 40740 41300 40750 41380
rect 41060 41300 41070 41380
rect 41380 41300 41390 41380
rect 41700 41300 41710 41380
rect 42020 41300 42030 41380
rect 48500 41270 48605 41400
rect 48640 41320 48650 41400
rect 57370 41350 57490 41410
rect 57670 41350 57790 41410
rect 58250 41350 58370 41410
rect 58550 41350 58670 41410
rect 58850 41350 58970 41410
rect 59150 41350 59270 41410
rect 59450 41350 59570 41410
rect 59750 41350 59870 41410
rect 60360 41400 60440 41410
rect 62060 41400 62140 41410
rect 57260 41340 57340 41350
rect 57490 41340 57620 41350
rect 48500 41260 48640 41270
rect 57340 41260 57350 41340
rect 36020 41220 36100 41230
rect 36340 41220 36420 41230
rect 36660 41220 36740 41230
rect 36980 41220 37060 41230
rect 37300 41220 37380 41230
rect 37620 41220 37700 41230
rect 40500 41220 40580 41230
rect 40820 41220 40900 41230
rect 41140 41220 41220 41230
rect 41460 41220 41540 41230
rect 41780 41220 41860 41230
rect 42100 41220 42180 41230
rect 42420 41220 42500 41230
rect 42740 41220 42820 41230
rect 43060 41220 43140 41230
rect 43380 41220 43460 41230
rect 43785 41220 43865 41230
rect 44105 41220 44185 41230
rect 44425 41220 44505 41230
rect 44745 41220 44825 41230
rect 45065 41220 45145 41230
rect 45385 41220 45465 41230
rect 45705 41220 45785 41230
rect 46025 41220 46105 41230
rect 46345 41220 46425 41230
rect 46665 41220 46745 41230
rect 46985 41220 47065 41230
rect 47305 41220 47385 41230
rect 47625 41220 47705 41230
rect 47945 41220 48025 41230
rect 48265 41220 48345 41230
rect 36100 41140 36110 41220
rect 36420 41140 36430 41220
rect 36740 41140 36750 41220
rect 37060 41140 37070 41220
rect 37380 41140 37390 41220
rect 37700 41140 37710 41220
rect 40580 41140 40590 41220
rect 40900 41140 40910 41220
rect 41220 41140 41230 41220
rect 41540 41140 41550 41220
rect 41860 41140 41870 41220
rect 42180 41140 42190 41220
rect 42500 41140 42510 41220
rect 42820 41140 42830 41220
rect 43140 41140 43150 41220
rect 43460 41140 43470 41220
rect 43865 41140 43875 41220
rect 44185 41140 44195 41220
rect 44505 41140 44515 41220
rect 44825 41140 44835 41220
rect 45145 41140 45155 41220
rect 45465 41140 45475 41220
rect 45785 41140 45795 41220
rect 46105 41140 46115 41220
rect 46425 41140 46435 41220
rect 46745 41140 46755 41220
rect 47065 41140 47075 41220
rect 47385 41140 47395 41220
rect 47705 41140 47715 41220
rect 48025 41140 48035 41220
rect 48345 41140 48355 41220
rect 48500 41130 48605 41260
rect 48640 41180 48650 41260
rect 57490 41230 57550 41340
rect 57620 41260 57630 41340
rect 57790 41230 57850 41350
rect 58370 41340 58500 41350
rect 58670 41340 58800 41350
rect 58970 41340 59100 41350
rect 59270 41340 59400 41350
rect 59570 41340 59710 41350
rect 58370 41230 58430 41340
rect 58500 41260 58510 41340
rect 58670 41230 58730 41340
rect 58800 41260 58810 41340
rect 58970 41230 59030 41340
rect 59100 41260 59110 41340
rect 59270 41230 59330 41340
rect 59400 41260 59410 41340
rect 59570 41230 59630 41340
rect 59710 41260 59720 41340
rect 59870 41230 59930 41350
rect 60440 41320 60450 41400
rect 62140 41320 62150 41400
rect 73250 41350 73370 41410
rect 73860 41400 73940 41410
rect 75560 41400 75640 41410
rect 60360 41260 60440 41270
rect 62060 41260 62140 41270
rect 57455 41180 57465 41210
rect 57755 41180 57765 41210
rect 58335 41180 58345 41210
rect 58635 41180 58645 41210
rect 58935 41180 58945 41210
rect 59235 41180 59245 41210
rect 59535 41180 59545 41210
rect 59835 41180 59845 41210
rect 60440 41180 60450 41260
rect 60580 41220 60660 41230
rect 60900 41220 60980 41230
rect 61320 41220 61400 41230
rect 61640 41220 61720 41230
rect 48500 41120 48640 41130
rect 36180 41060 36260 41070
rect 36500 41060 36580 41070
rect 36820 41060 36900 41070
rect 37140 41060 37220 41070
rect 37460 41060 37540 41070
rect 40660 41060 40740 41070
rect 40980 41060 41060 41070
rect 41300 41060 41380 41070
rect 41620 41060 41700 41070
rect 41940 41060 42020 41070
rect 42260 41060 42340 41070
rect 42580 41060 42660 41070
rect 42900 41060 42980 41070
rect 43220 41060 43300 41070
rect 43945 41060 44025 41070
rect 44265 41060 44345 41070
rect 44585 41060 44665 41070
rect 44905 41060 44985 41070
rect 45225 41060 45305 41070
rect 45545 41060 45625 41070
rect 45865 41060 45945 41070
rect 46185 41060 46265 41070
rect 46505 41060 46585 41070
rect 46825 41060 46905 41070
rect 47145 41060 47225 41070
rect 47465 41060 47545 41070
rect 47785 41060 47865 41070
rect 48105 41060 48185 41070
rect 36260 40980 36270 41060
rect 36580 40980 36590 41060
rect 36900 40980 36910 41060
rect 37220 40980 37230 41060
rect 37540 40980 37550 41060
rect 40740 40980 40750 41060
rect 41060 40980 41070 41060
rect 41380 40980 41390 41060
rect 41700 40980 41710 41060
rect 42020 40980 42030 41060
rect 42340 40980 42350 41060
rect 42660 40980 42670 41060
rect 42980 40980 42990 41060
rect 43300 40980 43310 41060
rect 44025 40980 44035 41060
rect 44345 40980 44355 41060
rect 44665 40980 44675 41060
rect 44985 40980 44995 41060
rect 45305 40980 45315 41060
rect 45625 40980 45635 41060
rect 45945 40980 45955 41060
rect 46265 40980 46275 41060
rect 46585 40980 46595 41060
rect 46905 40980 46915 41060
rect 47225 40980 47235 41060
rect 47545 40980 47555 41060
rect 47865 40980 47875 41060
rect 48185 40980 48195 41060
rect 48500 40990 48605 41120
rect 48640 41040 48650 41120
rect 57100 41090 60140 41180
rect 60660 41140 60670 41220
rect 60980 41140 60990 41220
rect 61400 41140 61410 41220
rect 61720 41140 61730 41220
rect 62140 41180 62150 41260
rect 73370 41230 73430 41350
rect 73940 41320 73950 41400
rect 75640 41320 75650 41400
rect 86750 41350 86870 41410
rect 87360 41400 87440 41410
rect 89060 41400 89140 41410
rect 73860 41260 73940 41270
rect 75560 41260 75640 41270
rect 73335 41180 73345 41210
rect 73940 41180 73950 41260
rect 74080 41220 74160 41230
rect 74400 41220 74480 41230
rect 74820 41220 74900 41230
rect 75140 41220 75220 41230
rect 60360 41120 60440 41130
rect 62060 41120 62140 41130
rect 57220 41050 57340 41090
rect 57375 41050 57405 41090
rect 48500 40980 48640 40990
rect 36020 40900 36100 40910
rect 36340 40900 36420 40910
rect 36660 40900 36740 40910
rect 36980 40900 37060 40910
rect 37300 40900 37380 40910
rect 37620 40900 37700 40910
rect 40820 40900 40900 40910
rect 41140 40900 41220 40910
rect 41460 40900 41540 40910
rect 41780 40900 41860 40910
rect 42100 40900 42180 40910
rect 42420 40900 42500 40910
rect 42740 40900 42820 40910
rect 43060 40900 43140 40910
rect 43380 40900 43460 40910
rect 43785 40900 43865 40910
rect 44105 40900 44185 40910
rect 44425 40900 44505 40910
rect 44745 40900 44825 40910
rect 45065 40900 45145 40910
rect 45385 40900 45465 40910
rect 45705 40900 45785 40910
rect 46025 40900 46105 40910
rect 46345 40900 46425 40910
rect 46665 40900 46745 40910
rect 46985 40900 47065 40910
rect 47305 40900 47385 40910
rect 47625 40900 47705 40910
rect 47945 40900 48025 40910
rect 48265 40900 48345 40910
rect 36100 40820 36110 40900
rect 36420 40820 36430 40900
rect 36740 40820 36750 40900
rect 37060 40820 37070 40900
rect 37380 40820 37390 40900
rect 37700 40820 37710 40900
rect 40900 40820 40910 40900
rect 41220 40820 41230 40900
rect 41540 40820 41550 40900
rect 41860 40820 41870 40900
rect 42180 40820 42190 40900
rect 42500 40820 42510 40900
rect 42820 40820 42830 40900
rect 43140 40820 43150 40900
rect 43460 40820 43470 40900
rect 43865 40820 43875 40900
rect 44185 40820 44195 40900
rect 44505 40820 44515 40900
rect 44825 40820 44835 40900
rect 45145 40820 45155 40900
rect 45465 40820 45475 40900
rect 45785 40820 45795 40900
rect 46105 40820 46115 40900
rect 46425 40820 46435 40900
rect 46745 40820 46755 40900
rect 47065 40820 47075 40900
rect 47385 40820 47395 40900
rect 47705 40820 47715 40900
rect 48025 40820 48035 40900
rect 48345 40820 48355 40900
rect 48500 40850 48605 40980
rect 48640 40900 48650 40980
rect 57340 40940 57405 41050
rect 57220 40930 57405 40940
rect 54260 40895 54380 40925
rect 54996 40918 55076 40928
rect 55156 40918 55236 40928
rect 56601 40918 56681 40928
rect 54260 40865 54290 40895
rect 54350 40865 54380 40895
rect 48500 40840 48640 40850
rect 36180 40740 36260 40750
rect 36500 40740 36580 40750
rect 36820 40740 36900 40750
rect 37140 40740 37220 40750
rect 37460 40740 37540 40750
rect 40980 40740 41060 40750
rect 41300 40740 41380 40750
rect 41620 40740 41700 40750
rect 41940 40740 42020 40750
rect 42260 40740 42340 40750
rect 42580 40740 42660 40750
rect 42900 40740 42980 40750
rect 43220 40740 43300 40750
rect 43945 40740 44025 40750
rect 44265 40740 44345 40750
rect 44585 40740 44665 40750
rect 44905 40740 44985 40750
rect 45225 40740 45305 40750
rect 45545 40740 45625 40750
rect 45865 40740 45945 40750
rect 46185 40740 46265 40750
rect 46505 40740 46585 40750
rect 46825 40740 46905 40750
rect 47145 40740 47225 40750
rect 47465 40740 47545 40750
rect 47785 40740 47865 40750
rect 48105 40740 48185 40750
rect 36260 40660 36270 40740
rect 36580 40660 36590 40740
rect 36900 40660 36910 40740
rect 37220 40660 37230 40740
rect 37540 40660 37550 40740
rect 41060 40660 41070 40740
rect 41380 40660 41390 40740
rect 41700 40660 41710 40740
rect 42020 40660 42030 40740
rect 42340 40660 42350 40740
rect 42660 40660 42670 40740
rect 42980 40660 42990 40740
rect 43300 40660 43310 40740
rect 44025 40660 44035 40740
rect 44345 40660 44355 40740
rect 44665 40660 44675 40740
rect 44985 40660 44995 40740
rect 45305 40660 45315 40740
rect 45625 40660 45635 40740
rect 45945 40660 45955 40740
rect 46265 40660 46275 40740
rect 46585 40660 46595 40740
rect 46905 40660 46915 40740
rect 47225 40660 47235 40740
rect 47545 40660 47555 40740
rect 47865 40660 47875 40740
rect 48185 40660 48195 40740
rect 48500 40710 48605 40840
rect 48640 40760 48650 40840
rect 54260 40775 54380 40865
rect 55076 40848 55086 40918
rect 54996 40838 55086 40848
rect 55156 40848 55166 40918
rect 55236 40848 55246 40918
rect 56681 40848 56691 40918
rect 55156 40838 55246 40848
rect 56601 40838 56691 40848
rect 56720 40895 56840 40925
rect 56871 40918 56951 40928
rect 56720 40865 56750 40895
rect 56810 40865 56840 40895
rect 54260 40715 54290 40775
rect 54350 40715 54380 40775
rect 56720 40775 56840 40865
rect 56951 40848 56961 40918
rect 56871 40838 56961 40848
rect 54996 40758 55076 40768
rect 55156 40758 55236 40768
rect 56601 40758 56681 40768
rect 48500 40700 48640 40710
rect 36020 40580 36100 40590
rect 36340 40580 36420 40590
rect 36660 40580 36740 40590
rect 36980 40580 37060 40590
rect 37300 40580 37380 40590
rect 37620 40580 37700 40590
rect 41140 40580 41220 40590
rect 41460 40580 41540 40590
rect 41780 40580 41860 40590
rect 42100 40580 42180 40590
rect 42420 40580 42500 40590
rect 42740 40580 42820 40590
rect 43060 40580 43140 40590
rect 43380 40580 43460 40590
rect 43785 40580 43865 40590
rect 44105 40580 44185 40590
rect 44425 40580 44505 40590
rect 44745 40580 44825 40590
rect 45065 40580 45145 40590
rect 45385 40580 45465 40590
rect 45705 40580 45785 40590
rect 46025 40580 46105 40590
rect 46345 40580 46425 40590
rect 46665 40580 46745 40590
rect 46985 40580 47065 40590
rect 47305 40580 47385 40590
rect 47625 40580 47705 40590
rect 47945 40580 48025 40590
rect 48265 40580 48345 40590
rect 36100 40500 36110 40580
rect 36420 40500 36430 40580
rect 36740 40500 36750 40580
rect 37060 40500 37070 40580
rect 37380 40500 37390 40580
rect 37700 40500 37710 40580
rect 41220 40500 41230 40580
rect 41540 40500 41550 40580
rect 41860 40500 41870 40580
rect 42180 40500 42190 40580
rect 42500 40500 42510 40580
rect 42820 40500 42830 40580
rect 43140 40500 43150 40580
rect 43460 40500 43470 40580
rect 43865 40500 43875 40580
rect 44185 40500 44195 40580
rect 44505 40500 44515 40580
rect 44825 40500 44835 40580
rect 45145 40500 45155 40580
rect 45465 40500 45475 40580
rect 45785 40500 45795 40580
rect 46105 40500 46115 40580
rect 46425 40500 46435 40580
rect 46745 40500 46755 40580
rect 47065 40500 47075 40580
rect 47385 40500 47395 40580
rect 47705 40500 47715 40580
rect 48025 40500 48035 40580
rect 48345 40500 48355 40580
rect 48500 40570 48605 40700
rect 48640 40620 48650 40700
rect 54260 40685 54380 40715
rect 55076 40678 55086 40758
rect 55156 40678 55166 40758
rect 55236 40678 55246 40758
rect 56681 40678 56691 40758
rect 56720 40715 56750 40775
rect 56810 40715 56840 40775
rect 57220 40770 57340 40830
rect 57375 40770 57405 40930
rect 56871 40758 56951 40768
rect 56720 40685 56840 40715
rect 56951 40678 56961 40758
rect 57340 40660 57405 40770
rect 57220 40650 57405 40660
rect 48500 40560 48640 40570
rect 48500 40430 48605 40560
rect 48640 40480 48650 40560
rect 57375 40470 57405 40650
rect 57455 40470 57485 41090
rect 57520 41050 57640 41090
rect 57675 41050 57705 41090
rect 57540 41030 57620 41040
rect 57620 40950 57630 41030
rect 57640 40930 57705 41050
rect 57540 40890 57620 40900
rect 57620 40830 57630 40890
rect 57520 40770 57640 40830
rect 57675 40770 57705 40930
rect 57540 40750 57620 40760
rect 57620 40670 57630 40750
rect 57640 40650 57705 40770
rect 57540 40610 57620 40620
rect 57620 40530 57630 40610
rect 57675 40470 57705 40650
rect 57755 40470 57785 41090
rect 57820 41050 57940 41090
rect 57970 41050 58090 41090
rect 58100 41050 58220 41090
rect 58255 41050 58285 41090
rect 57940 40930 58090 41050
rect 58220 40940 58285 41050
rect 58100 40930 58285 40940
rect 57840 40890 57920 40900
rect 57920 40830 57930 40890
rect 57820 40770 57940 40830
rect 57970 40770 58090 40930
rect 58100 40770 58220 40830
rect 58255 40770 58285 40930
rect 57940 40650 58090 40770
rect 58220 40660 58285 40770
rect 58100 40650 58285 40660
rect 57840 40610 57920 40620
rect 57920 40530 57930 40610
rect 57970 40470 58090 40650
rect 58255 40470 58285 40650
rect 58335 40470 58365 41090
rect 58400 41050 58520 41090
rect 58555 41050 58585 41090
rect 58420 41030 58500 41040
rect 58500 40950 58510 41030
rect 58520 40930 58585 41050
rect 58420 40890 58500 40900
rect 58500 40830 58510 40890
rect 58400 40770 58520 40830
rect 58555 40770 58585 40930
rect 58420 40750 58500 40760
rect 58500 40670 58510 40750
rect 58520 40650 58585 40770
rect 58420 40610 58500 40620
rect 58500 40530 58510 40610
rect 58555 40470 58585 40650
rect 58635 40470 58665 41090
rect 58700 41050 58820 41090
rect 58855 41050 58885 41090
rect 58820 40940 58885 41050
rect 58700 40930 58885 40940
rect 58700 40770 58820 40830
rect 58855 40770 58885 40930
rect 58820 40660 58885 40770
rect 58700 40650 58885 40660
rect 58855 40470 58885 40650
rect 58935 40470 58965 41090
rect 59000 41050 59120 41090
rect 59155 41050 59185 41090
rect 59020 41030 59100 41040
rect 59100 40950 59110 41030
rect 59120 40930 59185 41050
rect 59020 40890 59100 40900
rect 59100 40830 59110 40890
rect 59000 40770 59120 40830
rect 59155 40770 59185 40930
rect 59020 40750 59100 40760
rect 59100 40670 59110 40750
rect 59120 40650 59185 40770
rect 59020 40610 59100 40620
rect 59100 40530 59110 40610
rect 59155 40470 59185 40650
rect 59235 40470 59265 41090
rect 59300 41050 59420 41090
rect 59455 41050 59485 41090
rect 59420 40940 59485 41050
rect 59300 40930 59485 40940
rect 59300 40770 59420 40830
rect 59455 40770 59485 40930
rect 59420 40660 59485 40770
rect 59300 40650 59485 40660
rect 59455 40470 59485 40650
rect 59535 40470 59565 41090
rect 59600 41050 59720 41090
rect 59755 41050 59785 41090
rect 59620 41030 59700 41040
rect 59700 40950 59710 41030
rect 59720 40930 59785 41050
rect 59620 40890 59700 40900
rect 59700 40830 59710 40890
rect 59600 40770 59720 40830
rect 59755 40770 59785 40930
rect 59620 40750 59700 40760
rect 59700 40670 59710 40750
rect 59720 40650 59785 40770
rect 59620 40610 59700 40620
rect 59700 40530 59710 40610
rect 59755 40470 59785 40650
rect 59835 40470 59865 41090
rect 59900 41050 60020 41090
rect 60050 41050 60140 41090
rect 60020 40930 60140 41050
rect 60440 41040 60450 41120
rect 60740 41060 60820 41070
rect 61060 41060 61140 41070
rect 61480 41060 61560 41070
rect 61800 41060 61880 41070
rect 60360 40980 60440 40990
rect 60820 40980 60830 41060
rect 61140 40980 61150 41060
rect 61560 40980 61570 41060
rect 61880 40980 61890 41060
rect 62140 41040 62150 41120
rect 73245 41090 73640 41180
rect 74160 41140 74170 41220
rect 74480 41140 74490 41220
rect 74900 41140 74910 41220
rect 75220 41140 75230 41220
rect 75640 41180 75650 41260
rect 86870 41230 86930 41350
rect 87440 41320 87450 41400
rect 89140 41320 89150 41400
rect 100250 41350 100370 41410
rect 100860 41400 100940 41410
rect 102560 41400 102640 41410
rect 87360 41260 87440 41270
rect 89060 41260 89140 41270
rect 86835 41180 86845 41210
rect 87440 41180 87450 41260
rect 87580 41220 87660 41230
rect 87900 41220 87980 41230
rect 88320 41220 88400 41230
rect 88640 41220 88720 41230
rect 73860 41120 73940 41130
rect 75560 41120 75640 41130
rect 73255 41050 73285 41090
rect 62060 40980 62140 40990
rect 59920 40890 60000 40900
rect 60000 40830 60010 40890
rect 59900 40770 60020 40830
rect 60050 40770 60140 40930
rect 60440 40900 60450 40980
rect 60580 40900 60660 40910
rect 60900 40900 60980 40910
rect 61320 40900 61400 40910
rect 61640 40900 61720 40910
rect 62140 40900 62150 40980
rect 73245 40930 73285 41050
rect 60360 40840 60440 40850
rect 60020 40650 60140 40770
rect 60440 40760 60450 40840
rect 60660 40820 60670 40900
rect 60980 40820 60990 40900
rect 61400 40820 61410 40900
rect 61720 40820 61730 40900
rect 67760 40895 67880 40925
rect 68496 40918 68576 40928
rect 68656 40918 68736 40928
rect 67760 40865 67790 40895
rect 67850 40865 67880 40895
rect 62060 40840 62140 40850
rect 62140 40760 62150 40840
rect 67760 40775 67880 40865
rect 68576 40848 68586 40918
rect 68496 40838 68586 40848
rect 68656 40848 68666 40918
rect 68736 40848 68746 40918
rect 68656 40838 68746 40848
rect 60740 40740 60820 40750
rect 61060 40740 61140 40750
rect 61480 40740 61560 40750
rect 61800 40740 61880 40750
rect 60360 40700 60440 40710
rect 59920 40610 60000 40620
rect 60000 40530 60010 40610
rect 60050 40470 60140 40650
rect 60440 40620 60450 40700
rect 60820 40660 60830 40740
rect 61140 40660 61150 40740
rect 61560 40660 61570 40740
rect 61880 40660 61890 40740
rect 67760 40715 67790 40775
rect 67850 40715 67880 40775
rect 73255 40770 73285 40930
rect 68496 40758 68576 40768
rect 68656 40758 68736 40768
rect 62060 40700 62140 40710
rect 62140 40620 62150 40700
rect 67760 40685 67880 40715
rect 68576 40678 68586 40758
rect 68656 40678 68666 40758
rect 68736 40678 68746 40758
rect 73245 40650 73285 40770
rect 60580 40580 60660 40590
rect 60900 40580 60980 40590
rect 61320 40580 61400 40590
rect 61640 40580 61720 40590
rect 60360 40560 60440 40570
rect 60440 40480 60450 40560
rect 60660 40500 60670 40580
rect 60980 40500 60990 40580
rect 61400 40500 61410 40580
rect 61720 40500 61730 40580
rect 62060 40560 62140 40570
rect 62140 40480 62150 40560
rect 73255 40470 73285 40650
rect 73335 40470 73365 41090
rect 73400 41050 73520 41090
rect 73550 41050 73640 41090
rect 73520 40930 73640 41050
rect 73940 41040 73950 41120
rect 74240 41060 74320 41070
rect 74560 41060 74640 41070
rect 74980 41060 75060 41070
rect 75300 41060 75380 41070
rect 73860 40980 73940 40990
rect 74320 40980 74330 41060
rect 74640 40980 74650 41060
rect 75060 40980 75070 41060
rect 75380 40980 75390 41060
rect 75640 41040 75650 41120
rect 86745 41090 87140 41180
rect 87660 41140 87670 41220
rect 87980 41140 87990 41220
rect 88400 41140 88410 41220
rect 88720 41140 88730 41220
rect 89140 41180 89150 41260
rect 100370 41230 100430 41350
rect 100940 41320 100950 41400
rect 102640 41320 102650 41400
rect 113750 41350 113870 41410
rect 114360 41400 114440 41410
rect 116060 41400 116140 41410
rect 100860 41260 100940 41270
rect 102560 41260 102640 41270
rect 100335 41180 100345 41210
rect 100940 41180 100950 41260
rect 101080 41220 101160 41230
rect 101400 41220 101480 41230
rect 101820 41220 101900 41230
rect 102140 41220 102220 41230
rect 87360 41120 87440 41130
rect 89060 41120 89140 41130
rect 86755 41050 86785 41090
rect 75560 40980 75640 40990
rect 73420 40890 73500 40900
rect 73500 40830 73510 40890
rect 73400 40770 73520 40830
rect 73550 40770 73640 40930
rect 73940 40900 73950 40980
rect 74080 40900 74160 40910
rect 74400 40900 74480 40910
rect 74820 40900 74900 40910
rect 75140 40900 75220 40910
rect 75640 40900 75650 40980
rect 86745 40930 86785 41050
rect 73860 40840 73940 40850
rect 73520 40650 73640 40770
rect 73940 40760 73950 40840
rect 74160 40820 74170 40900
rect 74480 40820 74490 40900
rect 74900 40820 74910 40900
rect 75220 40820 75230 40900
rect 75560 40840 75640 40850
rect 75640 40760 75650 40840
rect 86755 40770 86785 40930
rect 74240 40740 74320 40750
rect 74560 40740 74640 40750
rect 74980 40740 75060 40750
rect 75300 40740 75380 40750
rect 73860 40700 73940 40710
rect 73420 40610 73500 40620
rect 73500 40530 73510 40610
rect 73550 40470 73640 40650
rect 73940 40620 73950 40700
rect 74320 40660 74330 40740
rect 74640 40660 74650 40740
rect 75060 40660 75070 40740
rect 75380 40660 75390 40740
rect 75560 40700 75640 40710
rect 75640 40620 75650 40700
rect 86745 40650 86785 40770
rect 74080 40580 74160 40590
rect 74400 40580 74480 40590
rect 74820 40580 74900 40590
rect 75140 40580 75220 40590
rect 73860 40560 73940 40570
rect 73940 40480 73950 40560
rect 74160 40500 74170 40580
rect 74480 40500 74490 40580
rect 74900 40500 74910 40580
rect 75220 40500 75230 40580
rect 75560 40560 75640 40570
rect 75640 40480 75650 40560
rect 86755 40470 86785 40650
rect 86835 40470 86865 41090
rect 86900 41050 87020 41090
rect 87050 41050 87140 41090
rect 87020 40930 87140 41050
rect 87440 41040 87450 41120
rect 87740 41060 87820 41070
rect 88060 41060 88140 41070
rect 88480 41060 88560 41070
rect 88800 41060 88880 41070
rect 87360 40980 87440 40990
rect 87820 40980 87830 41060
rect 88140 40980 88150 41060
rect 88560 40980 88570 41060
rect 88880 40980 88890 41060
rect 89140 41040 89150 41120
rect 100245 41090 100640 41180
rect 101160 41140 101170 41220
rect 101480 41140 101490 41220
rect 101900 41140 101910 41220
rect 102220 41140 102230 41220
rect 102640 41180 102650 41260
rect 113870 41230 113930 41350
rect 114440 41320 114450 41400
rect 116140 41320 116150 41400
rect 127250 41350 127370 41410
rect 127860 41400 127940 41410
rect 129560 41400 129640 41410
rect 114360 41260 114440 41270
rect 116060 41260 116140 41270
rect 113835 41180 113845 41210
rect 114440 41180 114450 41260
rect 114580 41220 114660 41230
rect 114900 41220 114980 41230
rect 115320 41220 115400 41230
rect 115640 41220 115720 41230
rect 100860 41120 100940 41130
rect 102560 41120 102640 41130
rect 100255 41050 100285 41090
rect 89060 40980 89140 40990
rect 86920 40890 87000 40900
rect 87000 40830 87010 40890
rect 86900 40770 87020 40830
rect 87050 40770 87140 40930
rect 87440 40900 87450 40980
rect 87580 40900 87660 40910
rect 87900 40900 87980 40910
rect 88320 40900 88400 40910
rect 88640 40900 88720 40910
rect 89140 40900 89150 40980
rect 100245 40930 100285 41050
rect 87360 40840 87440 40850
rect 87020 40650 87140 40770
rect 87440 40760 87450 40840
rect 87660 40820 87670 40900
rect 87980 40820 87990 40900
rect 88400 40820 88410 40900
rect 88720 40820 88730 40900
rect 89060 40840 89140 40850
rect 89140 40760 89150 40840
rect 100255 40770 100285 40930
rect 87740 40740 87820 40750
rect 88060 40740 88140 40750
rect 88480 40740 88560 40750
rect 88800 40740 88880 40750
rect 87360 40700 87440 40710
rect 86920 40610 87000 40620
rect 87000 40530 87010 40610
rect 87050 40470 87140 40650
rect 87440 40620 87450 40700
rect 87820 40660 87830 40740
rect 88140 40660 88150 40740
rect 88560 40660 88570 40740
rect 88880 40660 88890 40740
rect 89060 40700 89140 40710
rect 89140 40620 89150 40700
rect 100245 40650 100285 40770
rect 87580 40580 87660 40590
rect 87900 40580 87980 40590
rect 88320 40580 88400 40590
rect 88640 40580 88720 40590
rect 87360 40560 87440 40570
rect 87440 40480 87450 40560
rect 87660 40500 87670 40580
rect 87980 40500 87990 40580
rect 88400 40500 88410 40580
rect 88720 40500 88730 40580
rect 89060 40560 89140 40570
rect 89140 40480 89150 40560
rect 100255 40470 100285 40650
rect 100335 40470 100365 41090
rect 100400 41050 100520 41090
rect 100550 41050 100640 41090
rect 100520 40930 100640 41050
rect 100940 41040 100950 41120
rect 101240 41060 101320 41070
rect 101560 41060 101640 41070
rect 101980 41060 102060 41070
rect 102300 41060 102380 41070
rect 100860 40980 100940 40990
rect 101320 40980 101330 41060
rect 101640 40980 101650 41060
rect 102060 40980 102070 41060
rect 102380 40980 102390 41060
rect 102640 41040 102650 41120
rect 113745 41090 114140 41180
rect 114660 41140 114670 41220
rect 114980 41140 114990 41220
rect 115400 41140 115410 41220
rect 115720 41140 115730 41220
rect 116140 41180 116150 41260
rect 127370 41230 127430 41350
rect 127940 41320 127950 41400
rect 129640 41320 129650 41400
rect 140830 41350 140870 41410
rect 141360 41400 141440 41410
rect 127860 41260 127940 41270
rect 129560 41260 129640 41270
rect 127335 41180 127345 41210
rect 127940 41180 127950 41260
rect 128080 41220 128160 41230
rect 128400 41220 128480 41230
rect 128820 41220 128900 41230
rect 129140 41220 129220 41230
rect 114360 41120 114440 41130
rect 116060 41120 116140 41130
rect 113755 41050 113785 41090
rect 102560 40980 102640 40990
rect 100420 40890 100500 40900
rect 100500 40830 100510 40890
rect 100400 40770 100520 40830
rect 100550 40770 100640 40930
rect 100940 40900 100950 40980
rect 101080 40900 101160 40910
rect 101400 40900 101480 40910
rect 101820 40900 101900 40910
rect 102140 40900 102220 40910
rect 102640 40900 102650 40980
rect 113745 40930 113785 41050
rect 100860 40840 100940 40850
rect 100520 40650 100640 40770
rect 100940 40760 100950 40840
rect 101160 40820 101170 40900
rect 101480 40820 101490 40900
rect 101900 40820 101910 40900
rect 102220 40820 102230 40900
rect 102560 40840 102640 40850
rect 102640 40760 102650 40840
rect 113755 40770 113785 40930
rect 101240 40740 101320 40750
rect 101560 40740 101640 40750
rect 101980 40740 102060 40750
rect 102300 40740 102380 40750
rect 100860 40700 100940 40710
rect 100420 40610 100500 40620
rect 100500 40530 100510 40610
rect 100550 40470 100640 40650
rect 100940 40620 100950 40700
rect 101320 40660 101330 40740
rect 101640 40660 101650 40740
rect 102060 40660 102070 40740
rect 102380 40660 102390 40740
rect 102560 40700 102640 40710
rect 102640 40620 102650 40700
rect 113745 40650 113785 40770
rect 101080 40580 101160 40590
rect 101400 40580 101480 40590
rect 101820 40580 101900 40590
rect 102140 40580 102220 40590
rect 100860 40560 100940 40570
rect 100940 40480 100950 40560
rect 101160 40500 101170 40580
rect 101480 40500 101490 40580
rect 101900 40500 101910 40580
rect 102220 40500 102230 40580
rect 102560 40560 102640 40570
rect 102640 40480 102650 40560
rect 113755 40470 113785 40650
rect 113835 40470 113865 41090
rect 113900 41050 114020 41090
rect 114050 41050 114140 41090
rect 114020 40930 114140 41050
rect 114440 41040 114450 41120
rect 114740 41060 114820 41070
rect 115060 41060 115140 41070
rect 115480 41060 115560 41070
rect 115800 41060 115880 41070
rect 114360 40980 114440 40990
rect 114820 40980 114830 41060
rect 115140 40980 115150 41060
rect 115560 40980 115570 41060
rect 115880 40980 115890 41060
rect 116140 41040 116150 41120
rect 127245 41090 127640 41180
rect 128160 41140 128170 41220
rect 128480 41140 128490 41220
rect 128900 41140 128910 41220
rect 129220 41140 129230 41220
rect 129640 41180 129650 41260
rect 140870 41230 140930 41350
rect 141440 41320 141450 41400
rect 141360 41260 141440 41270
rect 140835 41180 140845 41210
rect 141440 41180 141450 41260
rect 127860 41120 127940 41130
rect 129560 41120 129640 41130
rect 127255 41050 127285 41090
rect 116060 40980 116140 40990
rect 113920 40890 114000 40900
rect 114000 40830 114010 40890
rect 113900 40770 114020 40830
rect 114050 40770 114140 40930
rect 114440 40900 114450 40980
rect 114580 40900 114660 40910
rect 114900 40900 114980 40910
rect 115320 40900 115400 40910
rect 115640 40900 115720 40910
rect 116140 40900 116150 40980
rect 127245 40930 127285 41050
rect 114360 40840 114440 40850
rect 114020 40650 114140 40770
rect 114440 40760 114450 40840
rect 114660 40820 114670 40900
rect 114980 40820 114990 40900
rect 115400 40820 115410 40900
rect 115720 40820 115730 40900
rect 116060 40840 116140 40850
rect 116140 40760 116150 40840
rect 127255 40770 127285 40930
rect 114740 40740 114820 40750
rect 115060 40740 115140 40750
rect 115480 40740 115560 40750
rect 115800 40740 115880 40750
rect 114360 40700 114440 40710
rect 113920 40610 114000 40620
rect 114000 40530 114010 40610
rect 114050 40470 114140 40650
rect 114440 40620 114450 40700
rect 114820 40660 114830 40740
rect 115140 40660 115150 40740
rect 115560 40660 115570 40740
rect 115880 40660 115890 40740
rect 116060 40700 116140 40710
rect 116140 40620 116150 40700
rect 127245 40650 127285 40770
rect 114580 40580 114660 40590
rect 114900 40580 114980 40590
rect 115320 40580 115400 40590
rect 115640 40580 115720 40590
rect 114360 40560 114440 40570
rect 114440 40480 114450 40560
rect 114660 40500 114670 40580
rect 114980 40500 114990 40580
rect 115400 40500 115410 40580
rect 115720 40500 115730 40580
rect 116060 40560 116140 40570
rect 116140 40480 116150 40560
rect 127255 40470 127285 40650
rect 127335 40470 127365 41090
rect 127400 41050 127520 41090
rect 127550 41050 127640 41090
rect 127520 40930 127640 41050
rect 127940 41040 127950 41120
rect 128240 41060 128320 41070
rect 128560 41060 128640 41070
rect 128980 41060 129060 41070
rect 129300 41060 129380 41070
rect 127860 40980 127940 40990
rect 128320 40980 128330 41060
rect 128640 40980 128650 41060
rect 129060 40980 129070 41060
rect 129380 40980 129390 41060
rect 129640 41040 129650 41120
rect 140830 41090 141140 41180
rect 141360 41120 141440 41130
rect 129560 40980 129640 40990
rect 127420 40890 127500 40900
rect 127500 40830 127510 40890
rect 127400 40770 127520 40830
rect 127550 40770 127640 40930
rect 127940 40900 127950 40980
rect 128080 40900 128160 40910
rect 128400 40900 128480 40910
rect 128820 40900 128900 40910
rect 129140 40900 129220 40910
rect 129640 40900 129650 40980
rect 127860 40840 127940 40850
rect 127520 40650 127640 40770
rect 127940 40760 127950 40840
rect 128160 40820 128170 40900
rect 128480 40820 128490 40900
rect 128900 40820 128910 40900
rect 129220 40820 129230 40900
rect 129560 40840 129640 40850
rect 129640 40760 129650 40840
rect 128240 40740 128320 40750
rect 128560 40740 128640 40750
rect 128980 40740 129060 40750
rect 129300 40740 129380 40750
rect 127860 40700 127940 40710
rect 127420 40610 127500 40620
rect 127500 40530 127510 40610
rect 127550 40470 127640 40650
rect 127940 40620 127950 40700
rect 128320 40660 128330 40740
rect 128640 40660 128650 40740
rect 129060 40660 129070 40740
rect 129380 40660 129390 40740
rect 129560 40700 129640 40710
rect 129640 40620 129650 40700
rect 128080 40580 128160 40590
rect 128400 40580 128480 40590
rect 128820 40580 128900 40590
rect 129140 40580 129220 40590
rect 127860 40560 127940 40570
rect 127940 40480 127950 40560
rect 128160 40500 128170 40580
rect 128480 40500 128490 40580
rect 128900 40500 128910 40580
rect 129220 40500 129230 40580
rect 129560 40560 129640 40570
rect 129640 40480 129650 40560
rect 140835 40470 140865 41090
rect 140900 41050 141020 41090
rect 141050 41050 141140 41090
rect 141020 40930 141140 41050
rect 141440 41040 141450 41120
rect 141360 40980 141440 40990
rect 140920 40890 141000 40900
rect 141000 40830 141010 40890
rect 140900 40770 141020 40830
rect 141050 40770 141140 40930
rect 141440 40900 141450 40980
rect 141360 40840 141440 40850
rect 141020 40650 141140 40770
rect 141440 40760 141450 40840
rect 141360 40700 141440 40710
rect 140920 40610 141000 40620
rect 141000 40530 141010 40610
rect 141050 40470 141140 40650
rect 141440 40620 141450 40700
rect 141360 40560 141440 40570
rect 141440 40480 141450 40560
rect 36180 40420 36260 40430
rect 36500 40420 36580 40430
rect 36820 40420 36900 40430
rect 37140 40420 37220 40430
rect 37460 40420 37540 40430
rect 41300 40420 41380 40430
rect 41620 40420 41700 40430
rect 41940 40420 42020 40430
rect 42260 40420 42340 40430
rect 42580 40420 42660 40430
rect 42900 40420 42980 40430
rect 43220 40420 43300 40430
rect 43945 40420 44025 40430
rect 44265 40420 44345 40430
rect 44585 40420 44665 40430
rect 44905 40420 44985 40430
rect 45225 40420 45305 40430
rect 45545 40420 45625 40430
rect 45865 40420 45945 40430
rect 46185 40420 46265 40430
rect 46505 40420 46585 40430
rect 46825 40420 46905 40430
rect 47145 40420 47225 40430
rect 47465 40420 47545 40430
rect 47785 40420 47865 40430
rect 48105 40420 48185 40430
rect 48500 40420 48640 40430
rect 57455 40420 57465 40470
rect 57470 40460 57690 40470
rect 57755 40420 57765 40470
rect 57770 40460 57780 40470
rect 36260 40340 36270 40420
rect 36580 40340 36590 40420
rect 36900 40340 36910 40420
rect 37220 40340 37230 40420
rect 37540 40340 37550 40420
rect 41380 40340 41390 40420
rect 41700 40340 41710 40420
rect 42020 40340 42030 40420
rect 42340 40340 42350 40420
rect 42660 40340 42670 40420
rect 42980 40340 42990 40420
rect 43300 40340 43310 40420
rect 44025 40340 44035 40420
rect 44345 40340 44355 40420
rect 44665 40340 44675 40420
rect 44985 40340 44995 40420
rect 45305 40340 45315 40420
rect 45625 40340 45635 40420
rect 45945 40340 45955 40420
rect 46265 40340 46275 40420
rect 46585 40340 46595 40420
rect 46905 40340 46915 40420
rect 47225 40340 47235 40420
rect 47545 40340 47555 40420
rect 47865 40340 47875 40420
rect 48185 40340 48195 40420
rect 48500 40290 48605 40420
rect 48640 40340 48650 40420
rect 48500 40280 48640 40290
rect 36020 40260 36100 40270
rect 36340 40260 36420 40270
rect 36660 40260 36740 40270
rect 36980 40260 37060 40270
rect 37300 40260 37380 40270
rect 37620 40260 37700 40270
rect 41460 40260 41540 40270
rect 41780 40260 41860 40270
rect 42100 40260 42180 40270
rect 42420 40260 42500 40270
rect 42740 40260 42820 40270
rect 43060 40260 43140 40270
rect 43380 40260 43460 40270
rect 43785 40260 43865 40270
rect 44105 40260 44185 40270
rect 44425 40260 44505 40270
rect 44745 40260 44825 40270
rect 45065 40260 45145 40270
rect 45385 40260 45465 40270
rect 45705 40260 45785 40270
rect 46025 40260 46105 40270
rect 46345 40260 46425 40270
rect 46665 40260 46745 40270
rect 46985 40260 47065 40270
rect 47305 40260 47385 40270
rect 47625 40260 47705 40270
rect 47945 40260 48025 40270
rect 48265 40260 48345 40270
rect 36100 40180 36110 40260
rect 36420 40180 36430 40260
rect 36740 40180 36750 40260
rect 37060 40180 37070 40260
rect 37380 40180 37390 40260
rect 37700 40180 37710 40260
rect 41540 40180 41550 40260
rect 41860 40180 41870 40260
rect 42180 40180 42190 40260
rect 42500 40180 42510 40260
rect 42820 40180 42830 40260
rect 43140 40180 43150 40260
rect 43460 40180 43470 40260
rect 43865 40180 43875 40260
rect 44185 40180 44195 40260
rect 44505 40180 44515 40260
rect 44825 40180 44835 40260
rect 45145 40180 45155 40260
rect 45465 40180 45475 40260
rect 45785 40180 45795 40260
rect 46105 40180 46115 40260
rect 46425 40180 46435 40260
rect 46745 40180 46755 40260
rect 47065 40180 47075 40260
rect 47385 40180 47395 40260
rect 47705 40180 47715 40260
rect 48025 40180 48035 40260
rect 48345 40180 48355 40260
rect 48500 40150 48605 40280
rect 48640 40200 48650 40280
rect 58060 40270 58070 40470
rect 58335 40420 58345 40470
rect 58350 40460 58570 40470
rect 58635 40420 58645 40470
rect 58650 40460 58660 40470
rect 58935 40420 58945 40470
rect 58950 40460 59170 40470
rect 59235 40420 59245 40470
rect 59250 40460 59260 40470
rect 59535 40420 59545 40470
rect 59550 40460 59770 40470
rect 59835 40420 59845 40470
rect 59850 40460 59860 40470
rect 73245 40460 73270 40470
rect 60360 40420 60440 40430
rect 60740 40420 60820 40430
rect 61060 40420 61140 40430
rect 61480 40420 61560 40430
rect 61800 40420 61880 40430
rect 62060 40420 62140 40430
rect 73335 40420 73345 40470
rect 73350 40460 73360 40470
rect 86745 40460 86770 40470
rect 73860 40420 73940 40430
rect 74240 40420 74320 40430
rect 74560 40420 74640 40430
rect 74980 40420 75060 40430
rect 75300 40420 75380 40430
rect 75560 40420 75640 40430
rect 86835 40420 86845 40470
rect 86850 40460 86860 40470
rect 100245 40460 100270 40470
rect 87360 40420 87440 40430
rect 87740 40420 87820 40430
rect 88060 40420 88140 40430
rect 88480 40420 88560 40430
rect 88800 40420 88880 40430
rect 89060 40420 89140 40430
rect 100335 40420 100345 40470
rect 100350 40460 100360 40470
rect 113745 40460 113770 40470
rect 100860 40420 100940 40430
rect 101240 40420 101320 40430
rect 101560 40420 101640 40430
rect 101980 40420 102060 40430
rect 102300 40420 102380 40430
rect 102560 40420 102640 40430
rect 113835 40420 113845 40470
rect 113850 40460 113860 40470
rect 127245 40460 127270 40470
rect 114360 40420 114440 40430
rect 114740 40420 114820 40430
rect 115060 40420 115140 40430
rect 115480 40420 115560 40430
rect 115800 40420 115880 40430
rect 116060 40420 116140 40430
rect 127335 40420 127345 40470
rect 127350 40460 127360 40470
rect 127860 40420 127940 40430
rect 128240 40420 128320 40430
rect 128560 40420 128640 40430
rect 128980 40420 129060 40430
rect 129300 40420 129380 40430
rect 129560 40420 129640 40430
rect 140835 40420 140845 40470
rect 140850 40460 140860 40470
rect 141360 40420 141440 40430
rect 60440 40340 60450 40420
rect 60820 40340 60830 40420
rect 61140 40340 61150 40420
rect 61560 40340 61570 40420
rect 61880 40340 61890 40420
rect 62140 40340 62150 40420
rect 73940 40340 73950 40420
rect 74320 40340 74330 40420
rect 74640 40340 74650 40420
rect 75060 40340 75070 40420
rect 75380 40340 75390 40420
rect 75640 40340 75650 40420
rect 87440 40340 87450 40420
rect 87820 40340 87830 40420
rect 88140 40340 88150 40420
rect 88560 40340 88570 40420
rect 88880 40340 88890 40420
rect 89140 40340 89150 40420
rect 100940 40340 100950 40420
rect 101320 40340 101330 40420
rect 101640 40340 101650 40420
rect 102060 40340 102070 40420
rect 102380 40340 102390 40420
rect 102640 40340 102650 40420
rect 114440 40340 114450 40420
rect 114820 40340 114830 40420
rect 115140 40340 115150 40420
rect 115560 40340 115570 40420
rect 115880 40340 115890 40420
rect 116140 40340 116150 40420
rect 127940 40340 127950 40420
rect 128320 40340 128330 40420
rect 128640 40340 128650 40420
rect 129060 40340 129070 40420
rect 129380 40340 129390 40420
rect 129640 40340 129650 40420
rect 141440 40340 141450 40420
rect 60360 40280 60440 40290
rect 62060 40280 62140 40290
rect 73860 40280 73940 40290
rect 75560 40280 75640 40290
rect 87360 40280 87440 40290
rect 89060 40280 89140 40290
rect 100860 40280 100940 40290
rect 102560 40280 102640 40290
rect 114360 40280 114440 40290
rect 116060 40280 116140 40290
rect 127860 40280 127940 40290
rect 129560 40280 129640 40290
rect 141360 40280 141440 40290
rect 57180 40260 57980 40270
rect 58060 40260 60060 40270
rect 60440 40200 60450 40280
rect 60580 40260 60660 40270
rect 60900 40260 60980 40270
rect 61320 40260 61400 40270
rect 61640 40260 61720 40270
rect 60660 40180 60670 40260
rect 60980 40180 60990 40260
rect 61400 40180 61410 40260
rect 61720 40180 61730 40260
rect 62140 40200 62150 40280
rect 73245 40260 73560 40270
rect 73940 40200 73950 40280
rect 74080 40260 74160 40270
rect 74400 40260 74480 40270
rect 74820 40260 74900 40270
rect 75140 40260 75220 40270
rect 74160 40180 74170 40260
rect 74480 40180 74490 40260
rect 74900 40180 74910 40260
rect 75220 40180 75230 40260
rect 75640 40200 75650 40280
rect 86745 40260 87060 40270
rect 87440 40200 87450 40280
rect 87580 40260 87660 40270
rect 87900 40260 87980 40270
rect 88320 40260 88400 40270
rect 88640 40260 88720 40270
rect 87660 40180 87670 40260
rect 87980 40180 87990 40260
rect 88400 40180 88410 40260
rect 88720 40180 88730 40260
rect 89140 40200 89150 40280
rect 100245 40260 100560 40270
rect 100940 40200 100950 40280
rect 101080 40260 101160 40270
rect 101400 40260 101480 40270
rect 101820 40260 101900 40270
rect 102140 40260 102220 40270
rect 101160 40180 101170 40260
rect 101480 40180 101490 40260
rect 101900 40180 101910 40260
rect 102220 40180 102230 40260
rect 102640 40200 102650 40280
rect 113745 40260 114060 40270
rect 114440 40200 114450 40280
rect 114580 40260 114660 40270
rect 114900 40260 114980 40270
rect 115320 40260 115400 40270
rect 115640 40260 115720 40270
rect 114660 40180 114670 40260
rect 114980 40180 114990 40260
rect 115400 40180 115410 40260
rect 115720 40180 115730 40260
rect 116140 40200 116150 40280
rect 127245 40260 127560 40270
rect 127940 40200 127950 40280
rect 128080 40260 128160 40270
rect 128400 40260 128480 40270
rect 128820 40260 128900 40270
rect 129140 40260 129220 40270
rect 128160 40180 128170 40260
rect 128480 40180 128490 40260
rect 128900 40180 128910 40260
rect 129220 40180 129230 40260
rect 129640 40200 129650 40280
rect 140830 40260 141060 40270
rect 141440 40200 141450 40280
rect 48500 40140 48640 40150
rect 60360 40140 60440 40150
rect 62060 40140 62140 40150
rect 73860 40140 73940 40150
rect 75560 40140 75640 40150
rect 87360 40140 87440 40150
rect 89060 40140 89140 40150
rect 100860 40140 100940 40150
rect 102560 40140 102640 40150
rect 114360 40140 114440 40150
rect 116060 40140 116140 40150
rect 127860 40140 127940 40150
rect 129560 40140 129640 40150
rect 141360 40140 141440 40150
rect 36180 40100 36260 40110
rect 36500 40100 36580 40110
rect 36820 40100 36900 40110
rect 37140 40100 37220 40110
rect 37460 40100 37540 40110
rect 36260 40020 36270 40100
rect 36580 40020 36590 40100
rect 36900 40020 36910 40100
rect 37220 40020 37230 40100
rect 37540 40020 37550 40100
rect 48500 40000 48605 40140
rect 48640 40060 48650 40140
rect 48870 40060 48900 40120
rect 48990 40060 49020 40120
rect 49110 40060 49140 40120
rect 49230 40060 49260 40120
rect 49350 40060 49380 40120
rect 49470 40060 49500 40120
rect 49590 40060 49620 40120
rect 49710 40060 49740 40120
rect 49830 40060 49860 40120
rect 49950 40060 49980 40120
rect 50070 40060 50100 40120
rect 50190 40060 50220 40120
rect 50310 40060 50340 40120
rect 50430 40060 50460 40120
rect 50550 40060 50580 40120
rect 50670 40060 50700 40120
rect 50790 40060 50820 40120
rect 50910 40060 50940 40120
rect 51030 40060 51060 40120
rect 51150 40060 51180 40120
rect 51270 40060 51300 40120
rect 51390 40060 51420 40120
rect 51510 40060 51540 40120
rect 51630 40060 51660 40120
rect 51750 40060 51780 40120
rect 51870 40060 51900 40120
rect 51990 40060 52020 40120
rect 52110 40060 52140 40120
rect 52230 40060 52260 40120
rect 52350 40060 52380 40120
rect 52470 40060 52500 40120
rect 52590 40060 52620 40120
rect 52710 40060 52740 40120
rect 52830 40060 52860 40120
rect 52950 40060 52980 40120
rect 53070 40060 53100 40120
rect 53190 40060 53220 40120
rect 53310 40060 53340 40120
rect 53430 40060 53460 40120
rect 53550 40060 53580 40120
rect 53670 40060 53700 40120
rect 53790 40060 53820 40120
rect 53910 40060 53940 40120
rect 54030 40060 54060 40120
rect 54150 40060 54180 40120
rect 54270 40060 54300 40120
rect 54390 40060 54420 40120
rect 54510 40060 54540 40120
rect 54630 40060 54660 40120
rect 54750 40060 54780 40120
rect 54870 40060 54900 40120
rect 54990 40060 55020 40120
rect 55110 40060 55140 40120
rect 55230 40060 55260 40120
rect 55350 40060 55380 40120
rect 55470 40060 55500 40120
rect 55590 40060 55620 40120
rect 55710 40060 55740 40120
rect 55830 40060 55860 40120
rect 55950 40060 55980 40120
rect 56070 40060 56100 40120
rect 56190 40060 56220 40120
rect 56310 40060 56340 40120
rect 56430 40060 56460 40120
rect 56550 40060 56580 40120
rect 56670 40060 56700 40120
rect 56790 40060 56820 40120
rect 56910 40060 56940 40120
rect 57030 40060 57060 40120
rect 57150 40060 57180 40120
rect 57270 40060 57300 40120
rect 57390 40060 57420 40120
rect 57510 40060 57540 40120
rect 57630 40060 57660 40120
rect 57750 40060 57780 40120
rect 57870 40060 57900 40120
rect 57990 40060 58020 40120
rect 58110 40060 58140 40120
rect 58230 40060 58260 40120
rect 58350 40060 58380 40120
rect 58470 40060 58500 40120
rect 58590 40060 58620 40120
rect 58710 40060 58740 40120
rect 58830 40060 58860 40120
rect 58950 40060 58980 40120
rect 59070 40060 59100 40120
rect 59190 40060 59220 40120
rect 59310 40060 59340 40120
rect 59430 40060 59460 40120
rect 59550 40060 59580 40120
rect 59670 40060 59700 40120
rect 59790 40060 59820 40120
rect 59910 40060 59940 40120
rect 60030 40060 60060 40120
rect 60150 40060 60180 40120
rect 60440 40060 60450 40140
rect 62140 40060 62150 40140
rect 62370 40060 62400 40120
rect 62490 40060 62520 40120
rect 62610 40060 62640 40120
rect 62730 40060 62760 40120
rect 62850 40060 62880 40120
rect 62970 40060 63000 40120
rect 63090 40060 63120 40120
rect 63210 40060 63240 40120
rect 63330 40060 63360 40120
rect 63450 40060 63480 40120
rect 63570 40060 63600 40120
rect 63690 40060 63720 40120
rect 63810 40060 63840 40120
rect 63930 40060 63960 40120
rect 64050 40060 64080 40120
rect 64170 40060 64200 40120
rect 64290 40060 64320 40120
rect 64410 40060 64440 40120
rect 64530 40060 64560 40120
rect 64650 40060 64680 40120
rect 64770 40060 64800 40120
rect 64890 40060 64920 40120
rect 65010 40060 65040 40120
rect 65130 40060 65160 40120
rect 65250 40060 65280 40120
rect 65370 40060 65400 40120
rect 65490 40060 65520 40120
rect 65610 40060 65640 40120
rect 65730 40060 65760 40120
rect 65850 40060 65880 40120
rect 65970 40060 66000 40120
rect 66090 40060 66120 40120
rect 66210 40060 66240 40120
rect 66330 40060 66360 40120
rect 66450 40060 66480 40120
rect 66570 40060 66600 40120
rect 66690 40060 66720 40120
rect 66810 40060 66840 40120
rect 66930 40060 66960 40120
rect 67050 40060 67080 40120
rect 67170 40060 67200 40120
rect 67290 40060 67320 40120
rect 67410 40060 67440 40120
rect 67530 40060 67560 40120
rect 67650 40060 67680 40120
rect 67770 40060 67800 40120
rect 67890 40060 67920 40120
rect 68010 40060 68040 40120
rect 68130 40060 68160 40120
rect 68250 40060 68280 40120
rect 68370 40060 68400 40120
rect 68490 40060 68520 40120
rect 68610 40060 68640 40120
rect 68730 40060 68760 40120
rect 68850 40060 68880 40120
rect 73290 40060 73320 40120
rect 73410 40060 73440 40120
rect 73530 40060 73560 40120
rect 73650 40060 73680 40120
rect 73940 40060 73950 40140
rect 75640 40060 75650 40140
rect 75870 40060 75900 40120
rect 75990 40060 76020 40120
rect 76110 40060 76140 40120
rect 76230 40060 76255 40120
rect 86790 40060 86820 40120
rect 86910 40060 86940 40120
rect 87030 40060 87060 40120
rect 87150 40060 87180 40120
rect 87440 40060 87450 40140
rect 89140 40060 89150 40140
rect 89370 40060 89400 40120
rect 89490 40060 89520 40120
rect 89610 40060 89640 40120
rect 89730 40060 89755 40120
rect 100290 40060 100320 40120
rect 100410 40060 100440 40120
rect 100530 40060 100560 40120
rect 100650 40060 100680 40120
rect 100940 40060 100950 40140
rect 102640 40060 102650 40140
rect 102870 40060 102900 40120
rect 102990 40060 103020 40120
rect 103110 40060 103140 40120
rect 103230 40060 103255 40120
rect 113790 40060 113820 40120
rect 113910 40060 113940 40120
rect 114030 40060 114060 40120
rect 114150 40060 114180 40120
rect 114440 40060 114450 40140
rect 116140 40060 116150 40140
rect 116370 40060 116400 40120
rect 116490 40060 116520 40120
rect 116610 40060 116640 40120
rect 116730 40060 116755 40120
rect 127290 40060 127320 40120
rect 127410 40060 127440 40120
rect 127530 40060 127560 40120
rect 127650 40060 127680 40120
rect 127940 40060 127950 40140
rect 129640 40060 129650 40140
rect 129870 40060 129900 40120
rect 129990 40060 130020 40120
rect 130110 40060 130140 40120
rect 130230 40060 130255 40120
rect 140910 40060 140940 40120
rect 141030 40060 141060 40120
rect 141150 40060 141180 40120
rect 141440 40060 141450 40140
rect 141565 40000 141620 41660
rect 148380 41620 148390 41700
rect 148700 41620 148710 41700
rect 149020 41620 149030 41700
rect 149340 41620 149350 41700
rect 149660 41620 149670 41700
rect 152540 41620 152550 41700
rect 152860 41620 152870 41700
rect 153180 41620 153190 41700
rect 153500 41620 153510 41700
rect 153820 41620 153830 41700
rect 154140 41620 154150 41700
rect 154460 41620 154470 41700
rect 154780 41620 154790 41700
rect 155100 41620 155110 41700
rect 155420 41620 155430 41700
rect 155740 41620 155750 41700
rect 148140 41540 148220 41550
rect 148460 41540 148540 41550
rect 148780 41540 148860 41550
rect 149100 41540 149180 41550
rect 149420 41540 149500 41550
rect 149740 41540 149820 41550
rect 152300 41540 152380 41550
rect 152620 41540 152700 41550
rect 152940 41540 153020 41550
rect 153260 41540 153340 41550
rect 153580 41540 153660 41550
rect 153900 41540 153980 41550
rect 154220 41540 154300 41550
rect 154540 41540 154620 41550
rect 154860 41540 154940 41550
rect 155180 41540 155260 41550
rect 155500 41540 155580 41550
rect 155820 41540 155900 41550
rect 148220 41460 148230 41540
rect 148540 41460 148550 41540
rect 148860 41460 148870 41540
rect 149180 41460 149190 41540
rect 149500 41460 149510 41540
rect 149820 41460 149830 41540
rect 152380 41460 152390 41540
rect 152700 41460 152710 41540
rect 153020 41460 153030 41540
rect 153340 41460 153350 41540
rect 153660 41460 153670 41540
rect 153980 41460 153990 41540
rect 154300 41460 154310 41540
rect 154620 41460 154630 41540
rect 154940 41460 154950 41540
rect 155260 41460 155270 41540
rect 155580 41460 155590 41540
rect 155900 41460 155910 41540
rect 147980 41380 148060 41390
rect 148300 41380 148380 41390
rect 148620 41380 148700 41390
rect 148940 41380 149020 41390
rect 149260 41380 149340 41390
rect 149580 41380 149660 41390
rect 152460 41380 152540 41390
rect 152780 41380 152860 41390
rect 153100 41380 153180 41390
rect 153420 41380 153500 41390
rect 153740 41380 153820 41390
rect 154060 41380 154140 41390
rect 154380 41380 154460 41390
rect 154700 41380 154780 41390
rect 155020 41380 155100 41390
rect 155340 41380 155420 41390
rect 155660 41380 155740 41390
rect 155980 41380 156000 41390
rect 148060 41300 148070 41380
rect 148380 41300 148390 41380
rect 148700 41300 148710 41380
rect 149020 41300 149030 41380
rect 149340 41300 149350 41380
rect 149660 41300 149670 41380
rect 152540 41300 152550 41380
rect 152860 41300 152870 41380
rect 153180 41300 153190 41380
rect 153500 41300 153510 41380
rect 153820 41300 153830 41380
rect 154140 41300 154150 41380
rect 154460 41300 154470 41380
rect 154780 41300 154790 41380
rect 155100 41300 155110 41380
rect 155420 41300 155430 41380
rect 155740 41300 155750 41380
rect 141665 41220 141745 41230
rect 141985 41220 142065 41230
rect 145200 41220 145265 41230
rect 145505 41220 145585 41230
rect 145825 41220 145905 41230
rect 146145 41220 146225 41230
rect 146540 41220 146620 41230
rect 146860 41220 146940 41230
rect 147180 41220 147260 41230
rect 147500 41220 147580 41230
rect 147820 41220 147900 41230
rect 148140 41220 148220 41230
rect 148460 41220 148540 41230
rect 148780 41220 148860 41230
rect 149100 41220 149180 41230
rect 149420 41220 149500 41230
rect 152300 41220 152380 41230
rect 152620 41220 152700 41230
rect 152940 41220 153020 41230
rect 153260 41220 153340 41230
rect 153580 41220 153660 41230
rect 153900 41220 153980 41230
rect 154220 41220 154300 41230
rect 154540 41220 154620 41230
rect 154860 41220 154940 41230
rect 155180 41220 155260 41230
rect 155500 41220 155580 41230
rect 155820 41220 155900 41230
rect 141745 41140 141755 41220
rect 142065 41140 142075 41220
rect 145265 41140 145275 41220
rect 145585 41140 145595 41220
rect 145905 41140 145915 41220
rect 146225 41140 146235 41220
rect 146620 41140 146630 41220
rect 146940 41140 146950 41220
rect 147260 41140 147270 41220
rect 147580 41140 147590 41220
rect 147900 41140 147910 41220
rect 148220 41140 148230 41220
rect 148540 41140 148550 41220
rect 148860 41140 148870 41220
rect 149180 41140 149190 41220
rect 149500 41140 149510 41220
rect 152380 41140 152390 41220
rect 152700 41140 152710 41220
rect 153020 41140 153030 41220
rect 153340 41140 153350 41220
rect 153660 41140 153670 41220
rect 153980 41140 153990 41220
rect 154300 41140 154310 41220
rect 154620 41140 154630 41220
rect 154940 41140 154950 41220
rect 155260 41140 155270 41220
rect 155580 41140 155590 41220
rect 155900 41140 155910 41220
rect 141825 41060 141905 41070
rect 142145 41060 142200 41070
rect 145345 41060 145425 41070
rect 145665 41060 145745 41070
rect 145985 41060 146065 41070
rect 146700 41060 146780 41070
rect 147020 41060 147100 41070
rect 147340 41060 147420 41070
rect 147660 41060 147740 41070
rect 147980 41060 148060 41070
rect 148300 41060 148380 41070
rect 148620 41060 148700 41070
rect 148940 41060 149020 41070
rect 149260 41060 149340 41070
rect 152460 41060 152540 41070
rect 152780 41060 152860 41070
rect 153100 41060 153180 41070
rect 153420 41060 153500 41070
rect 153740 41060 153820 41070
rect 154060 41060 154140 41070
rect 154380 41060 154460 41070
rect 154700 41060 154780 41070
rect 155020 41060 155100 41070
rect 155340 41060 155420 41070
rect 155660 41060 155740 41070
rect 155980 41060 156000 41070
rect 141905 40980 141915 41060
rect 145425 40980 145435 41060
rect 145745 40980 145755 41060
rect 146065 40980 146075 41060
rect 146780 40980 146790 41060
rect 147100 40980 147110 41060
rect 147420 40980 147430 41060
rect 147740 40980 147750 41060
rect 148060 40980 148070 41060
rect 148380 40980 148390 41060
rect 148700 40980 148710 41060
rect 149020 40980 149030 41060
rect 149340 40980 149350 41060
rect 152540 40980 152550 41060
rect 152860 40980 152870 41060
rect 153180 40980 153190 41060
rect 153500 40980 153510 41060
rect 153820 40980 153830 41060
rect 154140 40980 154150 41060
rect 154460 40980 154470 41060
rect 154780 40980 154790 41060
rect 155100 40980 155110 41060
rect 155420 40980 155430 41060
rect 155740 40980 155750 41060
rect 141665 40900 141745 40910
rect 141985 40900 142065 40910
rect 145200 40900 145265 40910
rect 145505 40900 145585 40910
rect 145825 40900 145905 40910
rect 146145 40900 146225 40910
rect 146540 40900 146620 40910
rect 146860 40900 146940 40910
rect 147180 40900 147260 40910
rect 147500 40900 147580 40910
rect 147820 40900 147900 40910
rect 148140 40900 148220 40910
rect 148460 40900 148540 40910
rect 148780 40900 148860 40910
rect 149100 40900 149180 40910
rect 152300 40900 152380 40910
rect 152620 40900 152700 40910
rect 152940 40900 153020 40910
rect 153260 40900 153340 40910
rect 153580 40900 153660 40910
rect 153900 40900 153980 40910
rect 154220 40900 154300 40910
rect 154540 40900 154620 40910
rect 154860 40900 154940 40910
rect 155180 40900 155260 40910
rect 155500 40900 155580 40910
rect 155820 40900 155900 40910
rect 141745 40820 141755 40900
rect 142065 40820 142075 40900
rect 145265 40820 145275 40900
rect 145585 40820 145595 40900
rect 145905 40820 145915 40900
rect 146225 40820 146235 40900
rect 146620 40820 146630 40900
rect 146940 40820 146950 40900
rect 147260 40820 147270 40900
rect 147580 40820 147590 40900
rect 147900 40820 147910 40900
rect 148220 40820 148230 40900
rect 148540 40820 148550 40900
rect 148860 40820 148870 40900
rect 149180 40820 149190 40900
rect 152380 40820 152390 40900
rect 152700 40820 152710 40900
rect 153020 40820 153030 40900
rect 153340 40820 153350 40900
rect 153660 40820 153670 40900
rect 153980 40820 153990 40900
rect 154300 40820 154310 40900
rect 154620 40820 154630 40900
rect 154940 40820 154950 40900
rect 155260 40820 155270 40900
rect 155580 40820 155590 40900
rect 155900 40820 155910 40900
rect 141825 40740 141905 40750
rect 142145 40740 142200 40750
rect 145345 40740 145425 40750
rect 145665 40740 145745 40750
rect 145985 40740 146065 40750
rect 146700 40740 146780 40750
rect 147020 40740 147100 40750
rect 147340 40740 147420 40750
rect 147660 40740 147740 40750
rect 147980 40740 148060 40750
rect 148300 40740 148380 40750
rect 148620 40740 148700 40750
rect 148940 40740 149020 40750
rect 152460 40740 152540 40750
rect 152780 40740 152860 40750
rect 153100 40740 153180 40750
rect 153420 40740 153500 40750
rect 153740 40740 153820 40750
rect 154060 40740 154140 40750
rect 154380 40740 154460 40750
rect 154700 40740 154780 40750
rect 155020 40740 155100 40750
rect 155340 40740 155420 40750
rect 155660 40740 155740 40750
rect 155980 40740 156000 40750
rect 141905 40660 141915 40740
rect 145425 40660 145435 40740
rect 145745 40660 145755 40740
rect 146065 40660 146075 40740
rect 146780 40660 146790 40740
rect 147100 40660 147110 40740
rect 147420 40660 147430 40740
rect 147740 40660 147750 40740
rect 148060 40660 148070 40740
rect 148380 40660 148390 40740
rect 148700 40660 148710 40740
rect 149020 40660 149030 40740
rect 152540 40660 152550 40740
rect 152860 40660 152870 40740
rect 153180 40660 153190 40740
rect 153500 40660 153510 40740
rect 153820 40660 153830 40740
rect 154140 40660 154150 40740
rect 154460 40660 154470 40740
rect 154780 40660 154790 40740
rect 155100 40660 155110 40740
rect 155420 40660 155430 40740
rect 155740 40660 155750 40740
rect 141665 40580 141745 40590
rect 141985 40580 142065 40590
rect 145200 40580 145265 40590
rect 145505 40580 145585 40590
rect 145825 40580 145905 40590
rect 146145 40580 146225 40590
rect 146540 40580 146620 40590
rect 146860 40580 146940 40590
rect 147180 40580 147260 40590
rect 147500 40580 147580 40590
rect 147820 40580 147900 40590
rect 148140 40580 148220 40590
rect 148460 40580 148540 40590
rect 148780 40580 148860 40590
rect 152300 40580 152380 40590
rect 152620 40580 152700 40590
rect 152940 40580 153020 40590
rect 153260 40580 153340 40590
rect 153580 40580 153660 40590
rect 153900 40580 153980 40590
rect 154220 40580 154300 40590
rect 154540 40580 154620 40590
rect 154860 40580 154940 40590
rect 155180 40580 155260 40590
rect 155500 40580 155580 40590
rect 155820 40580 155900 40590
rect 141745 40500 141755 40580
rect 142065 40500 142075 40580
rect 145265 40500 145275 40580
rect 145585 40500 145595 40580
rect 145905 40500 145915 40580
rect 146225 40500 146235 40580
rect 146620 40500 146630 40580
rect 146940 40500 146950 40580
rect 147260 40500 147270 40580
rect 147580 40500 147590 40580
rect 147900 40500 147910 40580
rect 148220 40500 148230 40580
rect 148540 40500 148550 40580
rect 148860 40500 148870 40580
rect 152380 40500 152390 40580
rect 152700 40500 152710 40580
rect 153020 40500 153030 40580
rect 153340 40500 153350 40580
rect 153660 40500 153670 40580
rect 153980 40500 153990 40580
rect 154300 40500 154310 40580
rect 154620 40500 154630 40580
rect 154940 40500 154950 40580
rect 155260 40500 155270 40580
rect 155580 40500 155590 40580
rect 155900 40500 155910 40580
rect 141825 40420 141905 40430
rect 142145 40420 142200 40430
rect 145345 40420 145425 40430
rect 145665 40420 145745 40430
rect 145985 40420 146065 40430
rect 146700 40420 146780 40430
rect 147020 40420 147100 40430
rect 147340 40420 147420 40430
rect 147660 40420 147740 40430
rect 147980 40420 148060 40430
rect 148300 40420 148380 40430
rect 148620 40420 148700 40430
rect 152460 40420 152540 40430
rect 152780 40420 152860 40430
rect 153100 40420 153180 40430
rect 153420 40420 153500 40430
rect 153740 40420 153820 40430
rect 154060 40420 154140 40430
rect 154380 40420 154460 40430
rect 154700 40420 154780 40430
rect 155020 40420 155100 40430
rect 155340 40420 155420 40430
rect 155660 40420 155740 40430
rect 155980 40420 156000 40430
rect 141905 40340 141915 40420
rect 145425 40340 145435 40420
rect 145745 40340 145755 40420
rect 146065 40340 146075 40420
rect 146780 40340 146790 40420
rect 147100 40340 147110 40420
rect 147420 40340 147430 40420
rect 147740 40340 147750 40420
rect 148060 40340 148070 40420
rect 148380 40340 148390 40420
rect 148700 40340 148710 40420
rect 152540 40340 152550 40420
rect 152860 40340 152870 40420
rect 153180 40340 153190 40420
rect 153500 40340 153510 40420
rect 153820 40340 153830 40420
rect 154140 40340 154150 40420
rect 154460 40340 154470 40420
rect 154780 40340 154790 40420
rect 155100 40340 155110 40420
rect 155420 40340 155430 40420
rect 155740 40340 155750 40420
rect 141665 40260 141745 40270
rect 141985 40260 142065 40270
rect 145200 40260 145265 40270
rect 145505 40260 145585 40270
rect 145825 40260 145905 40270
rect 146145 40260 146225 40270
rect 146540 40260 146620 40270
rect 146860 40260 146940 40270
rect 147180 40260 147260 40270
rect 147500 40260 147580 40270
rect 147820 40260 147900 40270
rect 148140 40260 148220 40270
rect 148460 40260 148540 40270
rect 152300 40260 152380 40270
rect 152620 40260 152700 40270
rect 152940 40260 153020 40270
rect 153260 40260 153340 40270
rect 153580 40260 153660 40270
rect 153900 40260 153980 40270
rect 154220 40260 154300 40270
rect 154540 40260 154620 40270
rect 154860 40260 154940 40270
rect 155180 40260 155260 40270
rect 155500 40260 155580 40270
rect 155820 40260 155900 40270
rect 141745 40180 141755 40260
rect 142065 40180 142075 40260
rect 145265 40180 145275 40260
rect 145585 40180 145595 40260
rect 145905 40180 145915 40260
rect 146225 40180 146235 40260
rect 146620 40180 146630 40260
rect 146940 40180 146950 40260
rect 147260 40180 147270 40260
rect 147580 40180 147590 40260
rect 147900 40180 147910 40260
rect 148220 40180 148230 40260
rect 148540 40180 148550 40260
rect 152380 40180 152390 40260
rect 152700 40180 152710 40260
rect 153020 40180 153030 40260
rect 153340 40180 153350 40260
rect 153660 40180 153670 40260
rect 153980 40180 153990 40260
rect 154300 40180 154310 40260
rect 154620 40180 154630 40260
rect 154940 40180 154950 40260
rect 155260 40180 155270 40260
rect 155580 40180 155590 40260
rect 155900 40180 155910 40260
rect 152460 40100 152540 40110
rect 152780 40100 152860 40110
rect 153100 40100 153180 40110
rect 153420 40100 153500 40110
rect 153740 40100 153820 40110
rect 154060 40100 154140 40110
rect 154380 40100 154460 40110
rect 154700 40100 154780 40110
rect 155020 40100 155100 40110
rect 155340 40100 155420 40110
rect 155660 40100 155740 40110
rect 155980 40100 156000 40110
rect 152540 40020 152550 40100
rect 152860 40020 152870 40100
rect 153180 40020 153190 40100
rect 153500 40020 153510 40100
rect 153820 40020 153830 40100
rect 154140 40020 154150 40100
rect 154460 40020 154470 40100
rect 154780 40020 154790 40100
rect 155100 40020 155110 40100
rect 155420 40020 155430 40100
rect 155740 40020 155750 40100
rect 36020 39940 36100 39950
rect 36340 39940 36420 39950
rect 36660 39940 36740 39950
rect 36980 39940 37060 39950
rect 37300 39940 37380 39950
rect 37620 39940 37700 39950
rect 152300 39940 152380 39950
rect 152620 39940 152700 39950
rect 152940 39940 153020 39950
rect 153260 39940 153340 39950
rect 153580 39940 153660 39950
rect 153900 39940 153980 39950
rect 154220 39940 154300 39950
rect 154540 39940 154620 39950
rect 154860 39940 154940 39950
rect 155180 39940 155260 39950
rect 155500 39940 155580 39950
rect 155820 39940 155900 39950
rect 36100 39860 36110 39940
rect 36420 39860 36430 39940
rect 36740 39860 36750 39940
rect 37060 39860 37070 39940
rect 37380 39860 37390 39940
rect 37700 39860 37710 39940
rect 152380 39860 152390 39940
rect 152700 39860 152710 39940
rect 153020 39860 153030 39940
rect 153340 39860 153350 39940
rect 153660 39860 153670 39940
rect 153980 39860 153990 39940
rect 154300 39860 154310 39940
rect 154620 39860 154630 39940
rect 154940 39860 154950 39940
rect 155260 39860 155270 39940
rect 155580 39860 155590 39940
rect 155900 39860 155910 39940
rect 36180 39780 36260 39790
rect 36500 39780 36580 39790
rect 36820 39780 36900 39790
rect 37140 39780 37220 39790
rect 37460 39780 37540 39790
rect 37780 39780 37860 39790
rect 152140 39780 152220 39790
rect 152460 39780 152540 39790
rect 152780 39780 152860 39790
rect 153100 39780 153180 39790
rect 153420 39780 153500 39790
rect 153740 39780 153820 39790
rect 154060 39780 154140 39790
rect 154380 39780 154460 39790
rect 154700 39780 154780 39790
rect 155020 39780 155100 39790
rect 155340 39780 155420 39790
rect 155660 39780 155740 39790
rect 155980 39780 156000 39790
rect 36260 39700 36270 39780
rect 36580 39700 36590 39780
rect 36900 39700 36910 39780
rect 37220 39700 37230 39780
rect 37540 39700 37550 39780
rect 37860 39700 37870 39780
rect 152220 39700 152230 39780
rect 152540 39700 152550 39780
rect 152860 39700 152870 39780
rect 153180 39700 153190 39780
rect 153500 39700 153510 39780
rect 153820 39700 153830 39780
rect 154140 39700 154150 39780
rect 154460 39700 154470 39780
rect 154780 39700 154790 39780
rect 155100 39700 155110 39780
rect 155420 39700 155430 39780
rect 155740 39700 155750 39780
rect 36020 39620 36100 39630
rect 36340 39620 36420 39630
rect 36660 39620 36740 39630
rect 36980 39620 37060 39630
rect 37300 39620 37380 39630
rect 37620 39620 37700 39630
rect 37940 39620 38020 39630
rect 151980 39620 152060 39630
rect 152300 39620 152380 39630
rect 152620 39620 152700 39630
rect 152940 39620 153020 39630
rect 153260 39620 153340 39630
rect 153580 39620 153660 39630
rect 153900 39620 153980 39630
rect 154220 39620 154300 39630
rect 154540 39620 154620 39630
rect 154860 39620 154940 39630
rect 155180 39620 155260 39630
rect 155500 39620 155580 39630
rect 155820 39620 155900 39630
rect 36100 39540 36110 39620
rect 36420 39540 36430 39620
rect 36740 39540 36750 39620
rect 37060 39540 37070 39620
rect 37380 39540 37390 39620
rect 37700 39540 37710 39620
rect 38020 39540 38030 39620
rect 152060 39540 152070 39620
rect 152380 39540 152390 39620
rect 152700 39540 152710 39620
rect 153020 39540 153030 39620
rect 153340 39540 153350 39620
rect 153660 39540 153670 39620
rect 153980 39540 153990 39620
rect 154300 39540 154310 39620
rect 154620 39540 154630 39620
rect 154940 39540 154950 39620
rect 155260 39540 155270 39620
rect 155580 39540 155590 39620
rect 155900 39540 155910 39620
rect 36180 39460 36260 39470
rect 36500 39460 36580 39470
rect 36820 39460 36900 39470
rect 37140 39460 37220 39470
rect 37460 39460 37540 39470
rect 37780 39460 37860 39470
rect 38100 39460 38180 39470
rect 151820 39460 151900 39470
rect 152140 39460 152220 39470
rect 152460 39460 152540 39470
rect 152780 39460 152860 39470
rect 153100 39460 153180 39470
rect 153420 39460 153500 39470
rect 153740 39460 153820 39470
rect 154060 39460 154140 39470
rect 154380 39460 154460 39470
rect 154700 39460 154780 39470
rect 155020 39460 155100 39470
rect 155340 39460 155420 39470
rect 155660 39460 155740 39470
rect 155980 39460 156000 39470
rect 36260 39380 36270 39460
rect 36580 39380 36590 39460
rect 36900 39380 36910 39460
rect 37220 39380 37230 39460
rect 37540 39380 37550 39460
rect 37860 39380 37870 39460
rect 38180 39380 38190 39460
rect 56285 39395 56365 39405
rect 56465 39395 56545 39405
rect 56645 39395 56725 39405
rect 56825 39395 56905 39405
rect 57005 39395 57085 39405
rect 56365 39315 56375 39395
rect 56545 39315 56555 39395
rect 56725 39315 56735 39395
rect 56905 39315 56915 39395
rect 57085 39315 57095 39395
rect 151900 39380 151910 39460
rect 152220 39380 152230 39460
rect 152540 39380 152550 39460
rect 152860 39380 152870 39460
rect 153180 39380 153190 39460
rect 153500 39380 153510 39460
rect 153820 39380 153830 39460
rect 154140 39380 154150 39460
rect 154460 39380 154470 39460
rect 154780 39380 154790 39460
rect 155100 39380 155110 39460
rect 155420 39380 155430 39460
rect 155740 39380 155750 39460
rect 36020 39300 36100 39310
rect 36340 39300 36420 39310
rect 36660 39300 36740 39310
rect 36980 39300 37060 39310
rect 37300 39300 37380 39310
rect 37620 39300 37700 39310
rect 37940 39300 38020 39310
rect 38260 39300 38340 39310
rect 151660 39300 151740 39310
rect 151980 39300 152060 39310
rect 152300 39300 152380 39310
rect 152620 39300 152700 39310
rect 152940 39300 153020 39310
rect 153260 39300 153340 39310
rect 153580 39300 153660 39310
rect 153900 39300 153980 39310
rect 154220 39300 154300 39310
rect 154540 39300 154620 39310
rect 154860 39300 154940 39310
rect 155180 39300 155260 39310
rect 155500 39300 155580 39310
rect 155820 39300 155900 39310
rect 36100 39220 36110 39300
rect 36420 39220 36430 39300
rect 36740 39220 36750 39300
rect 37060 39220 37070 39300
rect 37380 39220 37390 39300
rect 37700 39220 37710 39300
rect 38020 39220 38030 39300
rect 38340 39220 38350 39300
rect 56285 39215 56365 39225
rect 56465 39215 56545 39225
rect 56645 39215 56725 39225
rect 56825 39215 56905 39225
rect 57005 39215 57085 39225
rect 151740 39220 151750 39300
rect 152060 39220 152070 39300
rect 152380 39220 152390 39300
rect 152700 39220 152710 39300
rect 153020 39220 153030 39300
rect 153340 39220 153350 39300
rect 153660 39220 153670 39300
rect 153980 39220 153990 39300
rect 154300 39220 154310 39300
rect 154620 39220 154630 39300
rect 154940 39220 154950 39300
rect 155260 39220 155270 39300
rect 155580 39220 155590 39300
rect 155900 39220 155910 39300
rect 36180 39140 36260 39150
rect 36500 39140 36580 39150
rect 36820 39140 36900 39150
rect 37140 39140 37220 39150
rect 37460 39140 37540 39150
rect 37780 39140 37860 39150
rect 38100 39140 38180 39150
rect 38420 39140 38500 39150
rect 36260 39060 36270 39140
rect 36580 39060 36590 39140
rect 36900 39060 36910 39140
rect 37220 39060 37230 39140
rect 37540 39060 37550 39140
rect 37860 39060 37870 39140
rect 38180 39060 38190 39140
rect 38500 39060 38510 39140
rect 56365 39135 56375 39215
rect 56545 39135 56555 39215
rect 56725 39135 56735 39215
rect 56905 39135 56915 39215
rect 57085 39135 57095 39215
rect 151500 39140 151580 39150
rect 151820 39140 151900 39150
rect 152140 39140 152220 39150
rect 152460 39140 152540 39150
rect 152780 39140 152860 39150
rect 153100 39140 153180 39150
rect 153420 39140 153500 39150
rect 153740 39140 153820 39150
rect 154060 39140 154140 39150
rect 154380 39140 154460 39150
rect 154700 39140 154780 39150
rect 155020 39140 155100 39150
rect 155340 39140 155420 39150
rect 155660 39140 155740 39150
rect 155980 39140 156000 39150
rect 151580 39060 151590 39140
rect 151900 39060 151910 39140
rect 152220 39060 152230 39140
rect 152540 39060 152550 39140
rect 152860 39060 152870 39140
rect 153180 39060 153190 39140
rect 153500 39060 153510 39140
rect 153820 39060 153830 39140
rect 154140 39060 154150 39140
rect 154460 39060 154470 39140
rect 154780 39060 154790 39140
rect 155100 39060 155110 39140
rect 155420 39060 155430 39140
rect 155740 39060 155750 39140
rect 56285 39035 56365 39045
rect 56465 39035 56545 39045
rect 56645 39035 56725 39045
rect 56825 39035 56905 39045
rect 57005 39035 57085 39045
rect 36020 38980 36100 38990
rect 36340 38980 36420 38990
rect 36660 38980 36740 38990
rect 36980 38980 37060 38990
rect 37300 38980 37380 38990
rect 37620 38980 37700 38990
rect 37940 38980 38020 38990
rect 38260 38980 38340 38990
rect 38580 38980 38660 38990
rect 36100 38900 36110 38980
rect 36420 38900 36430 38980
rect 36740 38900 36750 38980
rect 37060 38900 37070 38980
rect 37380 38900 37390 38980
rect 37700 38900 37710 38980
rect 38020 38900 38030 38980
rect 38340 38900 38350 38980
rect 38660 38900 38670 38980
rect 56365 38955 56375 39035
rect 56545 38955 56555 39035
rect 56725 38955 56735 39035
rect 56905 38955 56915 39035
rect 57085 38955 57095 39035
rect 151340 38980 151420 38990
rect 151660 38980 151740 38990
rect 151980 38980 152060 38990
rect 152300 38980 152380 38990
rect 152620 38980 152700 38990
rect 152940 38980 153020 38990
rect 153260 38980 153340 38990
rect 153580 38980 153660 38990
rect 153900 38980 153980 38990
rect 154220 38980 154300 38990
rect 154540 38980 154620 38990
rect 154860 38980 154940 38990
rect 155180 38980 155260 38990
rect 155500 38980 155580 38990
rect 155820 38980 155900 38990
rect 151420 38900 151430 38980
rect 151740 38900 151750 38980
rect 152060 38900 152070 38980
rect 152380 38900 152390 38980
rect 152700 38900 152710 38980
rect 153020 38900 153030 38980
rect 153340 38900 153350 38980
rect 153660 38900 153670 38980
rect 153980 38900 153990 38980
rect 154300 38900 154310 38980
rect 154620 38900 154630 38980
rect 154940 38900 154950 38980
rect 155260 38900 155270 38980
rect 155580 38900 155590 38980
rect 155900 38900 155910 38980
rect 56285 38855 56365 38865
rect 56465 38855 56545 38865
rect 56645 38855 56725 38865
rect 56825 38855 56905 38865
rect 57005 38855 57085 38865
rect 36180 38820 36260 38830
rect 36500 38820 36580 38830
rect 36820 38820 36900 38830
rect 37140 38820 37220 38830
rect 37460 38820 37540 38830
rect 37780 38820 37860 38830
rect 38100 38820 38180 38830
rect 38420 38820 38500 38830
rect 38740 38820 38820 38830
rect 36260 38740 36270 38820
rect 36580 38740 36590 38820
rect 36900 38740 36910 38820
rect 37220 38740 37230 38820
rect 37540 38740 37550 38820
rect 37860 38740 37870 38820
rect 38180 38740 38190 38820
rect 38500 38740 38510 38820
rect 38820 38740 38830 38820
rect 56365 38775 56375 38855
rect 56545 38775 56555 38855
rect 56725 38775 56735 38855
rect 56905 38775 56915 38855
rect 57085 38775 57095 38855
rect 151180 38820 151260 38830
rect 151500 38820 151580 38830
rect 151820 38820 151900 38830
rect 152140 38820 152220 38830
rect 152460 38820 152540 38830
rect 152780 38820 152860 38830
rect 153100 38820 153180 38830
rect 153420 38820 153500 38830
rect 153740 38820 153820 38830
rect 154060 38820 154140 38830
rect 154380 38820 154460 38830
rect 154700 38820 154780 38830
rect 155020 38820 155100 38830
rect 155340 38820 155420 38830
rect 155660 38820 155740 38830
rect 155980 38820 156000 38830
rect 151260 38740 151270 38820
rect 151580 38740 151590 38820
rect 151900 38740 151910 38820
rect 152220 38740 152230 38820
rect 152540 38740 152550 38820
rect 152860 38740 152870 38820
rect 153180 38740 153190 38820
rect 153500 38740 153510 38820
rect 153820 38740 153830 38820
rect 154140 38740 154150 38820
rect 154460 38740 154470 38820
rect 154780 38740 154790 38820
rect 155100 38740 155110 38820
rect 155420 38740 155430 38820
rect 155740 38740 155750 38820
rect 56285 38675 56365 38685
rect 56465 38675 56545 38685
rect 56645 38675 56725 38685
rect 56825 38675 56905 38685
rect 57005 38675 57085 38685
rect 36020 38660 36100 38670
rect 36340 38660 36420 38670
rect 36660 38660 36740 38670
rect 36980 38660 37060 38670
rect 37300 38660 37380 38670
rect 37620 38660 37700 38670
rect 37940 38660 38020 38670
rect 38260 38660 38340 38670
rect 38580 38660 38660 38670
rect 38900 38660 38980 38670
rect 36100 38580 36110 38660
rect 36420 38580 36430 38660
rect 36740 38580 36750 38660
rect 37060 38580 37070 38660
rect 37380 38580 37390 38660
rect 37700 38580 37710 38660
rect 38020 38580 38030 38660
rect 38340 38580 38350 38660
rect 38660 38580 38670 38660
rect 38980 38580 38990 38660
rect 56365 38595 56375 38675
rect 56545 38595 56555 38675
rect 56725 38595 56735 38675
rect 56905 38595 56915 38675
rect 57085 38595 57095 38675
rect 151020 38660 151100 38670
rect 151340 38660 151420 38670
rect 151660 38660 151740 38670
rect 151980 38660 152060 38670
rect 152300 38660 152380 38670
rect 152620 38660 152700 38670
rect 152940 38660 153020 38670
rect 153260 38660 153340 38670
rect 153580 38660 153660 38670
rect 153900 38660 153980 38670
rect 154220 38660 154300 38670
rect 154540 38660 154620 38670
rect 154860 38660 154940 38670
rect 155180 38660 155260 38670
rect 155500 38660 155580 38670
rect 155820 38660 155900 38670
rect 151100 38580 151110 38660
rect 151420 38580 151430 38660
rect 151740 38580 151750 38660
rect 152060 38580 152070 38660
rect 152380 38580 152390 38660
rect 152700 38580 152710 38660
rect 153020 38580 153030 38660
rect 153340 38580 153350 38660
rect 153660 38580 153670 38660
rect 153980 38580 153990 38660
rect 154300 38580 154310 38660
rect 154620 38580 154630 38660
rect 154940 38580 154950 38660
rect 155260 38580 155270 38660
rect 155580 38580 155590 38660
rect 155900 38580 155910 38660
rect 36180 38500 36260 38510
rect 36500 38500 36580 38510
rect 36820 38500 36900 38510
rect 37140 38500 37220 38510
rect 37460 38500 37540 38510
rect 37780 38500 37860 38510
rect 38100 38500 38180 38510
rect 38420 38500 38500 38510
rect 38740 38500 38820 38510
rect 39060 38500 39140 38510
rect 150860 38500 150940 38510
rect 151180 38500 151260 38510
rect 151500 38500 151580 38510
rect 151820 38500 151900 38510
rect 152140 38500 152220 38510
rect 152460 38500 152540 38510
rect 152780 38500 152860 38510
rect 153100 38500 153180 38510
rect 153420 38500 153500 38510
rect 153740 38500 153820 38510
rect 154060 38500 154140 38510
rect 154380 38500 154460 38510
rect 154700 38500 154780 38510
rect 155020 38500 155100 38510
rect 155340 38500 155420 38510
rect 155660 38500 155740 38510
rect 155980 38500 156000 38510
rect 36260 38420 36270 38500
rect 36580 38420 36590 38500
rect 36900 38420 36910 38500
rect 37220 38420 37230 38500
rect 37540 38420 37550 38500
rect 37860 38420 37870 38500
rect 38180 38420 38190 38500
rect 38500 38420 38510 38500
rect 38820 38420 38830 38500
rect 39140 38420 39150 38500
rect 150940 38420 150950 38500
rect 151260 38420 151270 38500
rect 151580 38420 151590 38500
rect 151900 38420 151910 38500
rect 152220 38420 152230 38500
rect 152540 38420 152550 38500
rect 152860 38420 152870 38500
rect 153180 38420 153190 38500
rect 153500 38420 153510 38500
rect 153820 38420 153830 38500
rect 154140 38420 154150 38500
rect 154460 38420 154470 38500
rect 154780 38420 154790 38500
rect 155100 38420 155110 38500
rect 155420 38420 155430 38500
rect 155740 38420 155750 38500
rect 36020 38340 36100 38350
rect 36340 38340 36420 38350
rect 36660 38340 36740 38350
rect 36980 38340 37060 38350
rect 37300 38340 37380 38350
rect 37620 38340 37700 38350
rect 37940 38340 38020 38350
rect 38260 38340 38340 38350
rect 38580 38340 38660 38350
rect 38900 38340 38980 38350
rect 39220 38340 39300 38350
rect 150700 38340 150780 38350
rect 151020 38340 151100 38350
rect 151340 38340 151420 38350
rect 151660 38340 151740 38350
rect 151980 38340 152060 38350
rect 152300 38340 152380 38350
rect 152620 38340 152700 38350
rect 152940 38340 153020 38350
rect 153260 38340 153340 38350
rect 153580 38340 153660 38350
rect 153900 38340 153980 38350
rect 154220 38340 154300 38350
rect 154540 38340 154620 38350
rect 154860 38340 154940 38350
rect 155180 38340 155260 38350
rect 155500 38340 155580 38350
rect 155820 38340 155900 38350
rect 36100 38260 36110 38340
rect 36420 38260 36430 38340
rect 36740 38260 36750 38340
rect 37060 38260 37070 38340
rect 37380 38260 37390 38340
rect 37700 38260 37710 38340
rect 38020 38260 38030 38340
rect 38340 38260 38350 38340
rect 38660 38260 38670 38340
rect 38980 38260 38990 38340
rect 39300 38260 39310 38340
rect 150780 38260 150790 38340
rect 151100 38260 151110 38340
rect 151420 38260 151430 38340
rect 151740 38260 151750 38340
rect 152060 38260 152070 38340
rect 152380 38260 152390 38340
rect 152700 38260 152710 38340
rect 153020 38260 153030 38340
rect 153340 38260 153350 38340
rect 153660 38260 153670 38340
rect 153980 38260 153990 38340
rect 154300 38260 154310 38340
rect 154620 38260 154630 38340
rect 154940 38260 154950 38340
rect 155260 38260 155270 38340
rect 155580 38260 155590 38340
rect 155900 38260 155910 38340
rect 36180 38180 36260 38190
rect 36500 38180 36580 38190
rect 36820 38180 36900 38190
rect 37140 38180 37220 38190
rect 37460 38180 37540 38190
rect 37780 38180 37860 38190
rect 38100 38180 38180 38190
rect 38420 38180 38500 38190
rect 38740 38180 38820 38190
rect 39060 38180 39140 38190
rect 39380 38180 39460 38190
rect 150540 38180 150620 38190
rect 150860 38180 150940 38190
rect 151180 38180 151260 38190
rect 151500 38180 151580 38190
rect 151820 38180 151900 38190
rect 152140 38180 152220 38190
rect 152460 38180 152540 38190
rect 152780 38180 152860 38190
rect 153100 38180 153180 38190
rect 153420 38180 153500 38190
rect 153740 38180 153820 38190
rect 154060 38180 154140 38190
rect 154380 38180 154460 38190
rect 154700 38180 154780 38190
rect 155020 38180 155100 38190
rect 155340 38180 155420 38190
rect 155660 38180 155740 38190
rect 155980 38180 156000 38190
rect 36260 38100 36270 38180
rect 36580 38100 36590 38180
rect 36900 38100 36910 38180
rect 37220 38100 37230 38180
rect 37540 38100 37550 38180
rect 37860 38100 37870 38180
rect 38180 38100 38190 38180
rect 38500 38100 38510 38180
rect 38820 38100 38830 38180
rect 39140 38100 39150 38180
rect 39460 38100 39470 38180
rect 150620 38100 150630 38180
rect 150940 38100 150950 38180
rect 151260 38100 151270 38180
rect 151580 38100 151590 38180
rect 151900 38100 151910 38180
rect 152220 38100 152230 38180
rect 152540 38100 152550 38180
rect 152860 38100 152870 38180
rect 153180 38100 153190 38180
rect 153500 38100 153510 38180
rect 153820 38100 153830 38180
rect 154140 38100 154150 38180
rect 154460 38100 154470 38180
rect 154780 38100 154790 38180
rect 155100 38100 155110 38180
rect 155420 38100 155430 38180
rect 155740 38100 155750 38180
rect 36020 38020 36100 38030
rect 36340 38020 36420 38030
rect 36660 38020 36740 38030
rect 36980 38020 37060 38030
rect 37300 38020 37380 38030
rect 37620 38020 37700 38030
rect 37940 38020 38020 38030
rect 38260 38020 38340 38030
rect 38580 38020 38660 38030
rect 38900 38020 38980 38030
rect 39220 38020 39300 38030
rect 39540 38020 39620 38030
rect 150380 38020 150460 38030
rect 150700 38020 150780 38030
rect 151020 38020 151100 38030
rect 151340 38020 151420 38030
rect 151660 38020 151740 38030
rect 151980 38020 152060 38030
rect 152300 38020 152380 38030
rect 152620 38020 152700 38030
rect 152940 38020 153020 38030
rect 153260 38020 153340 38030
rect 153580 38020 153660 38030
rect 153900 38020 153980 38030
rect 154220 38020 154300 38030
rect 154540 38020 154620 38030
rect 154860 38020 154940 38030
rect 155180 38020 155260 38030
rect 155500 38020 155580 38030
rect 155820 38020 155900 38030
rect 36100 37940 36110 38020
rect 36420 37940 36430 38020
rect 36740 37940 36750 38020
rect 37060 37940 37070 38020
rect 37380 37940 37390 38020
rect 37700 37940 37710 38020
rect 38020 37940 38030 38020
rect 38340 37940 38350 38020
rect 38660 37940 38670 38020
rect 38980 37940 38990 38020
rect 39300 37940 39310 38020
rect 39620 37940 39630 38020
rect 48500 37930 48605 38000
rect 48500 37920 48640 37930
rect 48710 37920 48790 37930
rect 60060 37920 60140 37930
rect 60210 37920 60290 37930
rect 60360 37920 60440 37930
rect 62060 37920 62140 37930
rect 62210 37920 62290 37930
rect 73560 37920 73640 37930
rect 73710 37920 73790 37930
rect 73860 37920 73940 37930
rect 75560 37920 75640 37930
rect 75710 37920 75790 37930
rect 87060 37920 87140 37930
rect 87210 37920 87290 37930
rect 87360 37920 87440 37930
rect 89060 37920 89140 37930
rect 89210 37920 89290 37930
rect 100560 37920 100640 37930
rect 100710 37920 100790 37930
rect 100860 37920 100940 37930
rect 102560 37920 102640 37930
rect 102710 37920 102790 37930
rect 114060 37920 114140 37930
rect 114210 37920 114290 37930
rect 114360 37920 114440 37930
rect 116060 37920 116140 37930
rect 116210 37920 116290 37930
rect 127560 37920 127640 37930
rect 127710 37920 127790 37930
rect 127860 37920 127940 37930
rect 129560 37920 129640 37930
rect 129710 37920 129790 37930
rect 141060 37920 141140 37930
rect 141210 37920 141290 37930
rect 141360 37920 141440 37930
rect 36180 37860 36260 37870
rect 36500 37860 36580 37870
rect 36820 37860 36900 37870
rect 37140 37860 37220 37870
rect 37460 37860 37540 37870
rect 37780 37860 37860 37870
rect 38100 37860 38180 37870
rect 38420 37860 38500 37870
rect 38740 37860 38820 37870
rect 39060 37860 39140 37870
rect 39380 37860 39460 37870
rect 39700 37860 39780 37870
rect 36260 37780 36270 37860
rect 36580 37780 36590 37860
rect 36900 37780 36910 37860
rect 37220 37780 37230 37860
rect 37540 37780 37550 37860
rect 37860 37780 37870 37860
rect 38180 37780 38190 37860
rect 38500 37780 38510 37860
rect 38820 37780 38830 37860
rect 39140 37780 39150 37860
rect 39460 37780 39470 37860
rect 39780 37780 39790 37860
rect 43785 37800 43865 37810
rect 44105 37800 44185 37810
rect 44425 37800 44505 37810
rect 44745 37800 44825 37810
rect 45065 37800 45145 37810
rect 45385 37800 45465 37810
rect 45705 37800 45785 37810
rect 46025 37800 46105 37810
rect 46345 37800 46425 37810
rect 46665 37800 46745 37810
rect 46985 37800 47065 37810
rect 47305 37800 47385 37810
rect 47625 37800 47705 37810
rect 47945 37800 48025 37810
rect 48265 37800 48345 37810
rect 43865 37720 43875 37800
rect 44185 37720 44195 37800
rect 44505 37720 44515 37800
rect 44825 37720 44835 37800
rect 45145 37720 45155 37800
rect 45465 37720 45475 37800
rect 45785 37720 45795 37800
rect 46105 37720 46115 37800
rect 46425 37720 46435 37800
rect 46745 37720 46755 37800
rect 47065 37720 47075 37800
rect 47385 37720 47395 37800
rect 47705 37720 47715 37800
rect 48025 37720 48035 37800
rect 48345 37720 48355 37800
rect 48500 37750 48605 37920
rect 48640 37840 48650 37920
rect 48790 37840 48800 37920
rect 49180 37870 49210 37900
rect 49300 37870 49330 37900
rect 49420 37870 49450 37900
rect 49540 37870 49570 37900
rect 49660 37870 49690 37900
rect 49780 37870 49810 37900
rect 49900 37870 49930 37900
rect 50020 37870 50050 37900
rect 50140 37870 50170 37900
rect 50260 37870 50290 37900
rect 50380 37870 50410 37900
rect 50500 37870 50530 37900
rect 50620 37870 50650 37900
rect 50740 37870 50770 37900
rect 50860 37870 50890 37900
rect 50980 37870 51010 37900
rect 51100 37870 51130 37900
rect 51220 37870 51250 37900
rect 51340 37870 51370 37900
rect 51460 37870 51490 37900
rect 51580 37870 51610 37900
rect 51700 37870 51730 37900
rect 51820 37870 51850 37900
rect 51940 37870 51970 37900
rect 52060 37870 52090 37900
rect 52180 37870 52210 37900
rect 52300 37870 52330 37900
rect 52420 37870 52450 37900
rect 52540 37870 52570 37900
rect 52660 37870 52690 37900
rect 52780 37870 52810 37900
rect 52900 37870 52930 37900
rect 53020 37870 53050 37900
rect 53140 37870 53170 37900
rect 53260 37870 53290 37900
rect 53380 37870 53410 37900
rect 53500 37870 53530 37900
rect 53620 37870 53650 37900
rect 53740 37870 53770 37900
rect 53860 37870 53890 37900
rect 53980 37870 54010 37900
rect 54100 37870 54130 37900
rect 54220 37870 54250 37900
rect 54340 37870 54370 37900
rect 54460 37870 54490 37900
rect 54580 37870 54610 37900
rect 54700 37870 54730 37900
rect 54820 37870 54850 37900
rect 54940 37870 54970 37900
rect 55060 37870 55090 37900
rect 55180 37870 55210 37900
rect 55300 37870 55330 37900
rect 55420 37870 55450 37900
rect 55540 37870 55570 37900
rect 55660 37870 55690 37900
rect 55780 37870 55810 37900
rect 55900 37870 55930 37900
rect 56020 37870 56050 37900
rect 56140 37870 56170 37900
rect 56260 37870 56290 37900
rect 56380 37870 56410 37900
rect 56500 37870 56530 37900
rect 56620 37870 56650 37900
rect 56740 37870 56770 37900
rect 56860 37870 56890 37900
rect 56980 37870 57010 37900
rect 57100 37870 57130 37900
rect 57220 37870 57250 37900
rect 57340 37870 57370 37900
rect 57460 37870 57490 37900
rect 57580 37870 57610 37900
rect 57700 37870 57730 37900
rect 57820 37870 57850 37900
rect 57940 37870 57970 37900
rect 58060 37870 58090 37900
rect 58180 37870 58210 37900
rect 58300 37870 58330 37900
rect 58420 37870 58450 37900
rect 58540 37870 58570 37900
rect 58660 37870 58690 37900
rect 58780 37870 58810 37900
rect 58900 37870 58930 37900
rect 59020 37870 59050 37900
rect 59140 37870 59170 37900
rect 59260 37870 59290 37900
rect 59380 37870 59410 37900
rect 59500 37870 59530 37900
rect 59620 37870 59650 37900
rect 59740 37870 59770 37900
rect 59860 37870 59890 37900
rect 49060 37840 49120 37870
rect 49180 37840 49240 37870
rect 49300 37840 49360 37870
rect 49420 37840 49480 37870
rect 49540 37840 49600 37870
rect 49660 37840 49720 37870
rect 49780 37840 49840 37870
rect 49900 37840 49960 37870
rect 50020 37840 50080 37870
rect 50140 37840 50200 37870
rect 50260 37840 50320 37870
rect 50380 37840 50440 37870
rect 50500 37840 50560 37870
rect 50620 37840 50680 37870
rect 50740 37840 50800 37870
rect 50860 37840 50920 37870
rect 50980 37840 51040 37870
rect 51100 37840 51160 37870
rect 51220 37840 51280 37870
rect 51340 37840 51400 37870
rect 51460 37840 51520 37870
rect 51580 37840 51640 37870
rect 51700 37840 51760 37870
rect 51820 37840 51880 37870
rect 51940 37840 52000 37870
rect 52060 37840 52120 37870
rect 52180 37840 52240 37870
rect 52300 37840 52360 37870
rect 52420 37840 52480 37870
rect 52540 37840 52600 37870
rect 52660 37840 52720 37870
rect 52780 37840 52840 37870
rect 52900 37840 52960 37870
rect 53020 37840 53080 37870
rect 53140 37840 53200 37870
rect 53260 37840 53320 37870
rect 53380 37840 53440 37870
rect 53500 37840 53560 37870
rect 53620 37840 53680 37870
rect 53740 37840 53800 37870
rect 53860 37840 53920 37870
rect 53980 37840 54040 37870
rect 54100 37840 54160 37870
rect 54220 37840 54280 37870
rect 54340 37840 54400 37870
rect 54460 37840 54520 37870
rect 54580 37840 54640 37870
rect 54700 37840 54760 37870
rect 54820 37840 54880 37870
rect 54940 37840 55000 37870
rect 55060 37840 55120 37870
rect 55180 37840 55240 37870
rect 55300 37840 55360 37870
rect 55420 37840 55480 37870
rect 55540 37840 55600 37870
rect 55660 37840 55720 37870
rect 55780 37840 55840 37870
rect 55900 37840 55960 37870
rect 56020 37840 56080 37870
rect 56140 37840 56200 37870
rect 56260 37840 56320 37870
rect 56380 37840 56440 37870
rect 56500 37840 56560 37870
rect 56620 37840 56680 37870
rect 56740 37840 56800 37870
rect 56860 37840 56920 37870
rect 56980 37840 57040 37870
rect 57100 37840 57160 37870
rect 57220 37840 57280 37870
rect 57340 37840 57400 37870
rect 57460 37840 57520 37870
rect 57580 37840 57640 37870
rect 57700 37840 57760 37870
rect 57820 37840 57880 37870
rect 57940 37840 58000 37870
rect 58060 37840 58120 37870
rect 58180 37840 58240 37870
rect 58300 37840 58360 37870
rect 58420 37840 58480 37870
rect 58540 37840 58600 37870
rect 58660 37840 58720 37870
rect 58780 37840 58840 37870
rect 58900 37840 58960 37870
rect 59020 37840 59080 37870
rect 59140 37840 59200 37870
rect 59260 37840 59320 37870
rect 59380 37840 59440 37870
rect 59500 37840 59560 37870
rect 59620 37840 59680 37870
rect 59740 37840 59800 37870
rect 59860 37840 59920 37870
rect 60140 37840 60150 37920
rect 60290 37840 60300 37920
rect 60440 37840 60450 37920
rect 62140 37840 62150 37920
rect 62290 37840 62300 37920
rect 62680 37870 62710 37900
rect 62800 37870 62830 37900
rect 62920 37870 62950 37900
rect 63040 37870 63070 37900
rect 63160 37870 63190 37900
rect 63280 37870 63310 37900
rect 63400 37870 63430 37900
rect 63520 37870 63550 37900
rect 63640 37870 63670 37900
rect 63760 37870 63790 37900
rect 63880 37870 63910 37900
rect 64000 37870 64030 37900
rect 64120 37870 64150 37900
rect 64240 37870 64270 37900
rect 64360 37870 64390 37900
rect 64480 37870 64510 37900
rect 64600 37870 64630 37900
rect 64720 37870 64750 37900
rect 64840 37870 64870 37900
rect 64960 37870 64990 37900
rect 65080 37870 65110 37900
rect 65200 37870 65230 37900
rect 65320 37870 65350 37900
rect 65440 37870 65470 37900
rect 65560 37870 65590 37900
rect 65680 37870 65710 37900
rect 65800 37870 65830 37900
rect 65920 37870 65950 37900
rect 66040 37870 66070 37900
rect 66160 37870 66190 37900
rect 66280 37870 66310 37900
rect 66400 37870 66430 37900
rect 66520 37870 66550 37900
rect 66640 37870 66670 37900
rect 66760 37870 66790 37900
rect 66880 37870 66910 37900
rect 67000 37870 67030 37900
rect 67120 37870 67150 37900
rect 67240 37870 67270 37900
rect 67360 37870 67390 37900
rect 67480 37870 67510 37900
rect 67600 37870 67630 37900
rect 67720 37870 67750 37900
rect 67840 37870 67870 37900
rect 67960 37870 67990 37900
rect 68080 37870 68110 37900
rect 68200 37870 68230 37900
rect 68320 37870 68350 37900
rect 68440 37870 68470 37900
rect 68560 37870 68590 37900
rect 68680 37870 68710 37900
rect 68800 37870 68830 37900
rect 62560 37840 62620 37870
rect 62680 37840 62740 37870
rect 62800 37840 62860 37870
rect 62920 37840 62980 37870
rect 63040 37840 63100 37870
rect 63160 37840 63220 37870
rect 63280 37840 63340 37870
rect 63400 37840 63460 37870
rect 63520 37840 63580 37870
rect 63640 37840 63700 37870
rect 63760 37840 63820 37870
rect 63880 37840 63940 37870
rect 64000 37840 64060 37870
rect 64120 37840 64180 37870
rect 64240 37840 64300 37870
rect 64360 37840 64420 37870
rect 64480 37840 64540 37870
rect 64600 37840 64660 37870
rect 64720 37840 64780 37870
rect 64840 37840 64900 37870
rect 64960 37840 65020 37870
rect 65080 37840 65140 37870
rect 65200 37840 65260 37870
rect 65320 37840 65380 37870
rect 65440 37840 65500 37870
rect 65560 37840 65620 37870
rect 65680 37840 65740 37870
rect 65800 37840 65860 37870
rect 65920 37840 65980 37870
rect 66040 37840 66100 37870
rect 66160 37840 66220 37870
rect 66280 37840 66340 37870
rect 66400 37840 66460 37870
rect 66520 37840 66580 37870
rect 66640 37840 66700 37870
rect 66760 37840 66820 37870
rect 66880 37840 66940 37870
rect 67000 37840 67060 37870
rect 67120 37840 67180 37870
rect 67240 37840 67300 37870
rect 67360 37840 67420 37870
rect 67480 37840 67540 37870
rect 67600 37840 67660 37870
rect 67720 37840 67780 37870
rect 67840 37840 67900 37870
rect 67960 37840 68020 37870
rect 68080 37840 68140 37870
rect 68200 37840 68260 37870
rect 68320 37840 68380 37870
rect 68440 37840 68500 37870
rect 68560 37840 68620 37870
rect 68680 37840 68740 37870
rect 68800 37840 68860 37870
rect 68920 37840 68950 37900
rect 73245 37870 73270 37900
rect 73360 37870 73390 37900
rect 73245 37840 73300 37870
rect 73360 37840 73420 37870
rect 73640 37840 73650 37920
rect 73790 37840 73800 37920
rect 73940 37840 73950 37920
rect 75640 37840 75650 37920
rect 75790 37840 75800 37920
rect 76180 37870 76210 37900
rect 86745 37870 86770 37900
rect 86860 37870 86890 37900
rect 76060 37840 76120 37870
rect 76180 37840 76240 37870
rect 86745 37840 86800 37870
rect 86860 37840 86920 37870
rect 87140 37840 87150 37920
rect 87290 37840 87300 37920
rect 87440 37840 87450 37920
rect 89140 37840 89150 37920
rect 89290 37840 89300 37920
rect 89680 37870 89710 37900
rect 100245 37870 100270 37900
rect 100360 37870 100390 37900
rect 89560 37840 89620 37870
rect 89680 37840 89740 37870
rect 100245 37840 100300 37870
rect 100360 37840 100420 37870
rect 100640 37840 100650 37920
rect 100790 37840 100800 37920
rect 100940 37840 100950 37920
rect 102640 37840 102650 37920
rect 102790 37840 102800 37920
rect 103180 37870 103210 37900
rect 113745 37870 113770 37900
rect 113860 37870 113890 37900
rect 103060 37840 103120 37870
rect 103180 37840 103240 37870
rect 113745 37840 113800 37870
rect 113860 37840 113920 37870
rect 114140 37840 114150 37920
rect 114290 37840 114300 37920
rect 114440 37840 114450 37920
rect 116140 37840 116150 37920
rect 116290 37840 116300 37920
rect 116680 37870 116710 37900
rect 127245 37870 127270 37900
rect 127360 37870 127390 37900
rect 116560 37840 116620 37870
rect 116680 37840 116740 37870
rect 127245 37840 127300 37870
rect 127360 37840 127420 37870
rect 127640 37840 127650 37920
rect 127790 37840 127800 37920
rect 127940 37840 127950 37920
rect 129640 37840 129650 37920
rect 129790 37840 129800 37920
rect 130180 37870 130210 37900
rect 140860 37870 140890 37900
rect 130060 37840 130120 37870
rect 130180 37840 130240 37870
rect 140860 37840 140920 37870
rect 141140 37840 141150 37920
rect 141290 37840 141300 37920
rect 141440 37840 141450 37920
rect 60580 37800 60660 37810
rect 60900 37800 60980 37810
rect 61320 37800 61400 37810
rect 61640 37800 61720 37810
rect 74080 37800 74160 37810
rect 74400 37800 74480 37810
rect 74820 37800 74900 37810
rect 75140 37800 75220 37810
rect 87580 37800 87660 37810
rect 87900 37800 87980 37810
rect 88320 37800 88400 37810
rect 88640 37800 88720 37810
rect 101080 37800 101160 37810
rect 101400 37800 101480 37810
rect 101820 37800 101900 37810
rect 102140 37800 102220 37810
rect 114580 37800 114660 37810
rect 114900 37800 114980 37810
rect 115320 37800 115400 37810
rect 115640 37800 115720 37810
rect 128080 37800 128160 37810
rect 128400 37800 128480 37810
rect 128820 37800 128900 37810
rect 129140 37800 129220 37810
rect 49180 37750 49210 37780
rect 49300 37750 49330 37780
rect 49420 37750 49450 37780
rect 49540 37750 49570 37780
rect 49660 37750 49690 37780
rect 49780 37750 49810 37780
rect 49900 37750 49930 37780
rect 50020 37750 50050 37780
rect 50140 37750 50170 37780
rect 50260 37750 50290 37780
rect 50380 37750 50410 37780
rect 50500 37750 50530 37780
rect 50620 37750 50650 37780
rect 50740 37750 50770 37780
rect 50860 37750 50890 37780
rect 50980 37750 51010 37780
rect 51100 37750 51130 37780
rect 51220 37750 51250 37780
rect 51340 37750 51370 37780
rect 51460 37750 51490 37780
rect 51580 37750 51610 37780
rect 51700 37750 51730 37780
rect 51820 37750 51850 37780
rect 51940 37750 51970 37780
rect 52060 37750 52090 37780
rect 52180 37750 52210 37780
rect 52300 37750 52330 37780
rect 52420 37750 52450 37780
rect 52540 37750 52570 37780
rect 52660 37750 52690 37780
rect 52780 37750 52810 37780
rect 52900 37750 52930 37780
rect 53020 37750 53050 37780
rect 53140 37750 53170 37780
rect 53260 37750 53290 37780
rect 53380 37750 53410 37780
rect 53500 37750 53530 37780
rect 53620 37750 53650 37780
rect 53740 37750 53770 37780
rect 53860 37750 53890 37780
rect 53980 37750 54010 37780
rect 54100 37750 54130 37780
rect 54220 37750 54250 37780
rect 54340 37750 54370 37780
rect 54460 37750 54490 37780
rect 54580 37750 54610 37780
rect 54700 37750 54730 37780
rect 54820 37750 54850 37780
rect 54940 37750 54970 37780
rect 55060 37750 55090 37780
rect 55180 37750 55210 37780
rect 55300 37750 55330 37780
rect 55420 37750 55450 37780
rect 55540 37750 55570 37780
rect 55660 37750 55690 37780
rect 55780 37750 55810 37780
rect 55900 37750 55930 37780
rect 56020 37750 56050 37780
rect 56140 37750 56170 37780
rect 56260 37750 56290 37780
rect 56380 37750 56410 37780
rect 56500 37750 56530 37780
rect 56620 37750 56650 37780
rect 56740 37750 56770 37780
rect 56860 37750 56890 37780
rect 56980 37750 57010 37780
rect 57100 37750 57130 37780
rect 57220 37750 57250 37780
rect 57340 37750 57370 37780
rect 57460 37750 57490 37780
rect 57580 37750 57610 37780
rect 57700 37750 57730 37780
rect 57820 37750 57850 37780
rect 57940 37750 57970 37780
rect 58060 37750 58090 37780
rect 58180 37750 58210 37780
rect 58300 37750 58330 37780
rect 58420 37750 58450 37780
rect 58540 37750 58570 37780
rect 58660 37750 58690 37780
rect 58780 37750 58810 37780
rect 58900 37750 58930 37780
rect 59020 37750 59050 37780
rect 59140 37750 59170 37780
rect 59260 37750 59290 37780
rect 59380 37750 59410 37780
rect 59500 37750 59530 37780
rect 59620 37750 59650 37780
rect 59740 37750 59770 37780
rect 59860 37750 59890 37780
rect 48500 37740 48640 37750
rect 48710 37740 48790 37750
rect 36020 37700 36100 37710
rect 36340 37700 36420 37710
rect 36660 37700 36740 37710
rect 36980 37700 37060 37710
rect 37300 37700 37380 37710
rect 37620 37700 37700 37710
rect 37940 37700 38020 37710
rect 38260 37700 38340 37710
rect 38580 37700 38660 37710
rect 38900 37700 38980 37710
rect 39220 37700 39300 37710
rect 39540 37700 39620 37710
rect 39860 37700 39940 37710
rect 40180 37700 40260 37710
rect 40500 37700 40580 37710
rect 40820 37700 40900 37710
rect 41140 37700 41220 37710
rect 41460 37700 41540 37710
rect 41780 37700 41860 37710
rect 42100 37700 42180 37710
rect 42420 37700 42500 37710
rect 42740 37700 42820 37710
rect 43060 37700 43140 37710
rect 43380 37700 43460 37710
rect 36100 37620 36110 37700
rect 36420 37620 36430 37700
rect 36740 37620 36750 37700
rect 37060 37620 37070 37700
rect 37380 37620 37390 37700
rect 37700 37620 37710 37700
rect 38020 37620 38030 37700
rect 38340 37620 38350 37700
rect 38660 37620 38670 37700
rect 38980 37620 38990 37700
rect 39300 37620 39310 37700
rect 39620 37620 39630 37700
rect 39940 37620 39950 37700
rect 40260 37620 40270 37700
rect 40580 37620 40590 37700
rect 40900 37620 40910 37700
rect 41220 37620 41230 37700
rect 41540 37620 41550 37700
rect 41860 37620 41870 37700
rect 42180 37620 42190 37700
rect 42500 37620 42510 37700
rect 42820 37620 42830 37700
rect 43140 37620 43150 37700
rect 43460 37620 43470 37700
rect 43945 37640 44025 37650
rect 44265 37640 44345 37650
rect 44585 37640 44665 37650
rect 44905 37640 44985 37650
rect 45225 37640 45305 37650
rect 45545 37640 45625 37650
rect 45865 37640 45945 37650
rect 46185 37640 46265 37650
rect 46505 37640 46585 37650
rect 46825 37640 46905 37650
rect 47145 37640 47225 37650
rect 47465 37640 47545 37650
rect 47785 37640 47865 37650
rect 48105 37640 48185 37650
rect 44025 37560 44035 37640
rect 44345 37560 44355 37640
rect 44665 37560 44675 37640
rect 44985 37560 44995 37640
rect 45305 37560 45315 37640
rect 45625 37560 45635 37640
rect 45945 37560 45955 37640
rect 46265 37560 46275 37640
rect 46585 37560 46595 37640
rect 46905 37560 46915 37640
rect 47225 37560 47235 37640
rect 47545 37560 47555 37640
rect 47865 37560 47875 37640
rect 48185 37560 48195 37640
rect 48500 37570 48605 37740
rect 48640 37660 48650 37740
rect 48790 37660 48800 37740
rect 49060 37720 49120 37750
rect 49180 37720 49240 37750
rect 49300 37720 49360 37750
rect 49420 37720 49480 37750
rect 49540 37720 49600 37750
rect 49660 37720 49720 37750
rect 49780 37720 49840 37750
rect 49900 37720 49960 37750
rect 50020 37720 50080 37750
rect 50140 37720 50200 37750
rect 50260 37720 50320 37750
rect 50380 37720 50440 37750
rect 50500 37720 50560 37750
rect 50620 37720 50680 37750
rect 50740 37720 50800 37750
rect 50860 37720 50920 37750
rect 50980 37720 51040 37750
rect 51100 37720 51160 37750
rect 51220 37720 51280 37750
rect 51340 37720 51400 37750
rect 51460 37720 51520 37750
rect 51580 37720 51640 37750
rect 51700 37720 51760 37750
rect 51820 37720 51880 37750
rect 51940 37720 52000 37750
rect 52060 37720 52120 37750
rect 52180 37720 52240 37750
rect 52300 37720 52360 37750
rect 52420 37720 52480 37750
rect 52540 37720 52600 37750
rect 52660 37720 52720 37750
rect 52780 37720 52840 37750
rect 52900 37720 52960 37750
rect 53020 37720 53080 37750
rect 53140 37720 53200 37750
rect 53260 37720 53320 37750
rect 53380 37720 53440 37750
rect 53500 37720 53560 37750
rect 53620 37720 53680 37750
rect 53740 37720 53800 37750
rect 53860 37720 53920 37750
rect 53980 37720 54040 37750
rect 54100 37720 54160 37750
rect 54220 37720 54280 37750
rect 54340 37720 54400 37750
rect 54460 37720 54520 37750
rect 54580 37720 54640 37750
rect 54700 37720 54760 37750
rect 54820 37720 54880 37750
rect 54940 37720 55000 37750
rect 55060 37720 55120 37750
rect 55180 37720 55240 37750
rect 55300 37720 55360 37750
rect 55420 37720 55480 37750
rect 55540 37720 55600 37750
rect 55660 37720 55720 37750
rect 55780 37720 55840 37750
rect 55900 37720 55960 37750
rect 56020 37720 56080 37750
rect 56140 37720 56200 37750
rect 56260 37720 56320 37750
rect 56380 37720 56440 37750
rect 56500 37720 56560 37750
rect 56620 37720 56680 37750
rect 56740 37720 56800 37750
rect 56860 37720 56920 37750
rect 56980 37720 57040 37750
rect 57100 37720 57160 37750
rect 57220 37720 57280 37750
rect 57340 37720 57400 37750
rect 57460 37720 57520 37750
rect 57580 37720 57640 37750
rect 57700 37720 57760 37750
rect 57820 37720 57880 37750
rect 57940 37720 58000 37750
rect 58060 37720 58120 37750
rect 58180 37720 58240 37750
rect 58300 37720 58360 37750
rect 58420 37720 58480 37750
rect 58540 37720 58600 37750
rect 58660 37720 58720 37750
rect 58780 37720 58840 37750
rect 58900 37720 58960 37750
rect 59020 37720 59080 37750
rect 59140 37720 59200 37750
rect 59260 37720 59320 37750
rect 59380 37720 59440 37750
rect 59500 37720 59560 37750
rect 59620 37720 59680 37750
rect 59740 37720 59800 37750
rect 59860 37720 59920 37750
rect 60060 37740 60140 37750
rect 60210 37740 60290 37750
rect 60360 37740 60440 37750
rect 60140 37660 60150 37740
rect 60290 37660 60300 37740
rect 60440 37660 60450 37740
rect 60660 37720 60670 37800
rect 60980 37720 60990 37800
rect 61400 37720 61410 37800
rect 61720 37720 61730 37800
rect 62680 37750 62710 37780
rect 62800 37750 62830 37780
rect 62920 37750 62950 37780
rect 63040 37750 63070 37780
rect 63160 37750 63190 37780
rect 63280 37750 63310 37780
rect 63400 37750 63430 37780
rect 63520 37750 63550 37780
rect 63640 37750 63670 37780
rect 63760 37750 63790 37780
rect 63880 37750 63910 37780
rect 64000 37750 64030 37780
rect 64120 37750 64150 37780
rect 64240 37750 64270 37780
rect 64360 37750 64390 37780
rect 64480 37750 64510 37780
rect 64600 37750 64630 37780
rect 64720 37750 64750 37780
rect 64840 37750 64870 37780
rect 64960 37750 64990 37780
rect 65080 37750 65110 37780
rect 65200 37750 65230 37780
rect 65320 37750 65350 37780
rect 65440 37750 65470 37780
rect 65560 37750 65590 37780
rect 65680 37750 65710 37780
rect 65800 37750 65830 37780
rect 65920 37750 65950 37780
rect 66040 37750 66070 37780
rect 66160 37750 66190 37780
rect 66280 37750 66310 37780
rect 66400 37750 66430 37780
rect 66520 37750 66550 37780
rect 66640 37750 66670 37780
rect 66760 37750 66790 37780
rect 66880 37750 66910 37780
rect 67000 37750 67030 37780
rect 67120 37750 67150 37780
rect 67240 37750 67270 37780
rect 67360 37750 67390 37780
rect 67480 37750 67510 37780
rect 67600 37750 67630 37780
rect 67720 37750 67750 37780
rect 67840 37750 67870 37780
rect 67960 37750 67990 37780
rect 68080 37750 68110 37780
rect 68200 37750 68230 37780
rect 68320 37750 68350 37780
rect 68440 37750 68470 37780
rect 68560 37750 68590 37780
rect 68680 37750 68710 37780
rect 68800 37750 68830 37780
rect 62060 37740 62140 37750
rect 62210 37740 62290 37750
rect 62140 37660 62150 37740
rect 62290 37660 62300 37740
rect 62560 37720 62620 37750
rect 62680 37720 62740 37750
rect 62800 37720 62860 37750
rect 62920 37720 62980 37750
rect 63040 37720 63100 37750
rect 63160 37720 63220 37750
rect 63280 37720 63340 37750
rect 63400 37720 63460 37750
rect 63520 37720 63580 37750
rect 63640 37720 63700 37750
rect 63760 37720 63820 37750
rect 63880 37720 63940 37750
rect 64000 37720 64060 37750
rect 64120 37720 64180 37750
rect 64240 37720 64300 37750
rect 64360 37720 64420 37750
rect 64480 37720 64540 37750
rect 64600 37720 64660 37750
rect 64720 37720 64780 37750
rect 64840 37720 64900 37750
rect 64960 37720 65020 37750
rect 65080 37720 65140 37750
rect 65200 37720 65260 37750
rect 65320 37720 65380 37750
rect 65440 37720 65500 37750
rect 65560 37720 65620 37750
rect 65680 37720 65740 37750
rect 65800 37720 65860 37750
rect 65920 37720 65980 37750
rect 66040 37720 66100 37750
rect 66160 37720 66220 37750
rect 66280 37720 66340 37750
rect 66400 37720 66460 37750
rect 66520 37720 66580 37750
rect 66640 37720 66700 37750
rect 66760 37720 66820 37750
rect 66880 37720 66940 37750
rect 67000 37720 67060 37750
rect 67120 37720 67180 37750
rect 67240 37720 67300 37750
rect 67360 37720 67420 37750
rect 67480 37720 67540 37750
rect 67600 37720 67660 37750
rect 67720 37720 67780 37750
rect 67840 37720 67900 37750
rect 67960 37720 68020 37750
rect 68080 37720 68140 37750
rect 68200 37720 68260 37750
rect 68320 37720 68380 37750
rect 68440 37720 68500 37750
rect 68560 37720 68620 37750
rect 68680 37720 68740 37750
rect 68800 37720 68860 37750
rect 68920 37720 68950 37780
rect 73245 37750 73270 37780
rect 73360 37750 73390 37780
rect 73245 37720 73300 37750
rect 73360 37720 73420 37750
rect 73560 37740 73640 37750
rect 73710 37740 73790 37750
rect 73860 37740 73940 37750
rect 73640 37660 73650 37740
rect 73790 37660 73800 37740
rect 73940 37660 73950 37740
rect 74160 37720 74170 37800
rect 74480 37720 74490 37800
rect 74900 37720 74910 37800
rect 75220 37720 75230 37800
rect 76180 37750 76210 37780
rect 86745 37750 86770 37780
rect 86860 37750 86890 37780
rect 75560 37740 75640 37750
rect 75710 37740 75790 37750
rect 75640 37660 75650 37740
rect 75790 37660 75800 37740
rect 76060 37720 76120 37750
rect 76180 37720 76240 37750
rect 86745 37720 86800 37750
rect 86860 37720 86920 37750
rect 87060 37740 87140 37750
rect 87210 37740 87290 37750
rect 87360 37740 87440 37750
rect 87140 37660 87150 37740
rect 87290 37660 87300 37740
rect 87440 37660 87450 37740
rect 87660 37720 87670 37800
rect 87980 37720 87990 37800
rect 88400 37720 88410 37800
rect 88720 37720 88730 37800
rect 89680 37750 89710 37780
rect 100245 37750 100270 37780
rect 100360 37750 100390 37780
rect 89060 37740 89140 37750
rect 89210 37740 89290 37750
rect 89140 37660 89150 37740
rect 89290 37660 89300 37740
rect 89560 37720 89620 37750
rect 89680 37720 89740 37750
rect 100245 37720 100300 37750
rect 100360 37720 100420 37750
rect 100560 37740 100640 37750
rect 100710 37740 100790 37750
rect 100860 37740 100940 37750
rect 100640 37660 100650 37740
rect 100790 37660 100800 37740
rect 100940 37660 100950 37740
rect 101160 37720 101170 37800
rect 101480 37720 101490 37800
rect 101900 37720 101910 37800
rect 102220 37720 102230 37800
rect 103180 37750 103210 37780
rect 113745 37750 113770 37780
rect 113860 37750 113890 37780
rect 102560 37740 102640 37750
rect 102710 37740 102790 37750
rect 102640 37660 102650 37740
rect 102790 37660 102800 37740
rect 103060 37720 103120 37750
rect 103180 37720 103240 37750
rect 113745 37720 113800 37750
rect 113860 37720 113920 37750
rect 114060 37740 114140 37750
rect 114210 37740 114290 37750
rect 114360 37740 114440 37750
rect 114140 37660 114150 37740
rect 114290 37660 114300 37740
rect 114440 37660 114450 37740
rect 114660 37720 114670 37800
rect 114980 37720 114990 37800
rect 115400 37720 115410 37800
rect 115720 37720 115730 37800
rect 116680 37750 116710 37780
rect 127245 37750 127270 37780
rect 127360 37750 127390 37780
rect 116060 37740 116140 37750
rect 116210 37740 116290 37750
rect 116140 37660 116150 37740
rect 116290 37660 116300 37740
rect 116560 37720 116620 37750
rect 116680 37720 116740 37750
rect 127245 37720 127300 37750
rect 127360 37720 127420 37750
rect 127560 37740 127640 37750
rect 127710 37740 127790 37750
rect 127860 37740 127940 37750
rect 127640 37660 127650 37740
rect 127790 37660 127800 37740
rect 127940 37660 127950 37740
rect 128160 37720 128170 37800
rect 128480 37720 128490 37800
rect 128900 37720 128910 37800
rect 129220 37720 129230 37800
rect 130180 37750 130210 37780
rect 140860 37750 140890 37780
rect 129560 37740 129640 37750
rect 129710 37740 129790 37750
rect 129640 37660 129650 37740
rect 129790 37660 129800 37740
rect 130060 37720 130120 37750
rect 130180 37720 130240 37750
rect 140860 37720 140920 37750
rect 141060 37740 141140 37750
rect 141210 37740 141290 37750
rect 141360 37740 141440 37750
rect 141140 37660 141150 37740
rect 141290 37660 141300 37740
rect 141440 37660 141450 37740
rect 49180 37600 49210 37660
rect 49300 37600 49330 37660
rect 49420 37600 49450 37660
rect 49540 37600 49570 37660
rect 49660 37600 49690 37660
rect 49780 37600 49810 37660
rect 49900 37600 49930 37660
rect 50020 37600 50050 37660
rect 50140 37600 50170 37660
rect 50260 37600 50290 37660
rect 50380 37600 50410 37660
rect 50500 37600 50530 37660
rect 50620 37600 50650 37660
rect 50740 37600 50770 37660
rect 50860 37600 50890 37660
rect 50980 37600 51010 37660
rect 51100 37600 51130 37660
rect 51220 37600 51250 37660
rect 51340 37600 51370 37660
rect 51460 37600 51490 37660
rect 51580 37600 51610 37660
rect 51700 37600 51730 37660
rect 51820 37600 51850 37660
rect 51940 37600 51970 37660
rect 52060 37600 52090 37660
rect 52180 37600 52210 37660
rect 52300 37600 52330 37660
rect 52420 37600 52450 37660
rect 52540 37600 52570 37660
rect 52660 37600 52690 37660
rect 52780 37600 52810 37660
rect 52900 37600 52930 37660
rect 53020 37600 53050 37660
rect 53140 37600 53170 37660
rect 53260 37600 53290 37660
rect 53380 37600 53410 37660
rect 53500 37600 53530 37660
rect 53620 37600 53650 37660
rect 53740 37600 53770 37660
rect 53860 37600 53890 37660
rect 53980 37600 54010 37660
rect 54100 37600 54130 37660
rect 54220 37600 54250 37660
rect 54340 37600 54370 37660
rect 54460 37600 54490 37660
rect 54580 37600 54610 37660
rect 54700 37600 54730 37660
rect 54820 37600 54850 37660
rect 54940 37600 54970 37660
rect 55060 37600 55090 37660
rect 55180 37600 55210 37660
rect 55300 37600 55330 37660
rect 55420 37600 55450 37660
rect 55540 37600 55570 37660
rect 55660 37600 55690 37660
rect 55780 37600 55810 37660
rect 55900 37600 55930 37660
rect 56020 37600 56050 37660
rect 56140 37600 56170 37660
rect 56260 37600 56290 37660
rect 56380 37600 56410 37660
rect 56500 37600 56530 37660
rect 56620 37600 56650 37660
rect 56740 37600 56770 37660
rect 56860 37600 56890 37660
rect 56980 37600 57010 37660
rect 57100 37600 57130 37660
rect 57220 37600 57250 37660
rect 57340 37600 57370 37660
rect 57460 37600 57490 37660
rect 57580 37600 57610 37660
rect 57700 37600 57730 37660
rect 57820 37600 57850 37660
rect 57940 37600 57970 37660
rect 58060 37600 58090 37660
rect 58180 37600 58210 37660
rect 58300 37600 58330 37660
rect 58420 37600 58450 37660
rect 58540 37600 58570 37660
rect 58660 37600 58690 37660
rect 58780 37600 58810 37660
rect 58900 37600 58930 37660
rect 59020 37600 59050 37660
rect 59140 37600 59170 37660
rect 59260 37600 59290 37660
rect 59380 37600 59410 37660
rect 59500 37600 59530 37660
rect 59620 37600 59650 37660
rect 59740 37600 59770 37660
rect 59860 37600 59890 37660
rect 60740 37640 60820 37650
rect 61060 37640 61140 37650
rect 61480 37640 61560 37650
rect 61800 37640 61880 37650
rect 48500 37560 48640 37570
rect 48710 37560 48790 37570
rect 60060 37560 60140 37570
rect 60210 37560 60290 37570
rect 60360 37560 60440 37570
rect 60820 37560 60830 37640
rect 61140 37560 61150 37640
rect 61560 37560 61570 37640
rect 61880 37560 61890 37640
rect 62680 37600 62710 37660
rect 62800 37600 62830 37660
rect 62920 37600 62950 37660
rect 63040 37600 63070 37660
rect 63160 37600 63190 37660
rect 63280 37600 63310 37660
rect 63400 37600 63430 37660
rect 63520 37600 63550 37660
rect 63640 37600 63670 37660
rect 63760 37600 63790 37660
rect 63880 37600 63910 37660
rect 64000 37600 64030 37660
rect 64120 37600 64150 37660
rect 64240 37600 64270 37660
rect 64360 37600 64390 37660
rect 64480 37600 64510 37660
rect 64600 37600 64630 37660
rect 64720 37600 64750 37660
rect 64840 37600 64870 37660
rect 64960 37600 64990 37660
rect 65080 37600 65110 37660
rect 65200 37600 65230 37660
rect 65320 37600 65350 37660
rect 65440 37600 65470 37660
rect 65560 37600 65590 37660
rect 65680 37600 65710 37660
rect 65800 37600 65830 37660
rect 65920 37600 65950 37660
rect 66040 37600 66070 37660
rect 66160 37600 66190 37660
rect 66280 37600 66310 37660
rect 66400 37600 66430 37660
rect 66520 37600 66550 37660
rect 66640 37600 66670 37660
rect 66760 37600 66790 37660
rect 66880 37600 66910 37660
rect 67000 37600 67030 37660
rect 67120 37600 67150 37660
rect 67240 37600 67270 37660
rect 67360 37600 67390 37660
rect 67480 37600 67510 37660
rect 67600 37600 67630 37660
rect 67720 37600 67750 37660
rect 67840 37600 67870 37660
rect 67960 37600 67990 37660
rect 68080 37600 68110 37660
rect 68200 37600 68230 37660
rect 68320 37600 68350 37660
rect 68440 37600 68470 37660
rect 68560 37600 68590 37660
rect 68680 37600 68710 37660
rect 68800 37600 68830 37660
rect 68920 37600 68950 37660
rect 73245 37600 73270 37660
rect 73360 37600 73390 37660
rect 74240 37640 74320 37650
rect 74560 37640 74640 37650
rect 74980 37640 75060 37650
rect 75300 37640 75380 37650
rect 62060 37560 62140 37570
rect 62210 37560 62290 37570
rect 73560 37560 73640 37570
rect 73710 37560 73790 37570
rect 73860 37560 73940 37570
rect 74320 37560 74330 37640
rect 74640 37560 74650 37640
rect 75060 37560 75070 37640
rect 75380 37560 75390 37640
rect 76180 37600 76210 37660
rect 86745 37600 86770 37660
rect 86860 37600 86890 37660
rect 87740 37640 87820 37650
rect 88060 37640 88140 37650
rect 88480 37640 88560 37650
rect 88800 37640 88880 37650
rect 75560 37560 75640 37570
rect 75710 37560 75790 37570
rect 87060 37560 87140 37570
rect 87210 37560 87290 37570
rect 87360 37560 87440 37570
rect 87820 37560 87830 37640
rect 88140 37560 88150 37640
rect 88560 37560 88570 37640
rect 88880 37560 88890 37640
rect 89680 37600 89710 37660
rect 100245 37600 100270 37660
rect 100360 37600 100390 37660
rect 101240 37640 101320 37650
rect 101560 37640 101640 37650
rect 101980 37640 102060 37650
rect 102300 37640 102380 37650
rect 89060 37560 89140 37570
rect 89210 37560 89290 37570
rect 100560 37560 100640 37570
rect 100710 37560 100790 37570
rect 100860 37560 100940 37570
rect 101320 37560 101330 37640
rect 101640 37560 101650 37640
rect 102060 37560 102070 37640
rect 102380 37560 102390 37640
rect 103180 37600 103210 37660
rect 113745 37600 113770 37660
rect 113860 37600 113890 37660
rect 114740 37640 114820 37650
rect 115060 37640 115140 37650
rect 115480 37640 115560 37650
rect 115800 37640 115880 37650
rect 102560 37560 102640 37570
rect 102710 37560 102790 37570
rect 114060 37560 114140 37570
rect 114210 37560 114290 37570
rect 114360 37560 114440 37570
rect 114820 37560 114830 37640
rect 115140 37560 115150 37640
rect 115560 37560 115570 37640
rect 115880 37560 115890 37640
rect 116680 37600 116710 37660
rect 127245 37600 127270 37660
rect 127360 37600 127390 37660
rect 128240 37640 128320 37650
rect 128560 37640 128640 37650
rect 128980 37640 129060 37650
rect 129300 37640 129380 37650
rect 116060 37560 116140 37570
rect 116210 37560 116290 37570
rect 127560 37560 127640 37570
rect 127710 37560 127790 37570
rect 127860 37560 127940 37570
rect 128320 37560 128330 37640
rect 128640 37560 128650 37640
rect 129060 37560 129070 37640
rect 129380 37560 129390 37640
rect 130180 37600 130210 37660
rect 140860 37600 140890 37660
rect 129560 37560 129640 37570
rect 129710 37560 129790 37570
rect 141060 37560 141140 37570
rect 141210 37560 141290 37570
rect 141360 37560 141440 37570
rect 36180 37540 36260 37550
rect 36500 37540 36580 37550
rect 36820 37540 36900 37550
rect 37140 37540 37220 37550
rect 37460 37540 37540 37550
rect 37780 37540 37860 37550
rect 38100 37540 38180 37550
rect 38420 37540 38500 37550
rect 38740 37540 38820 37550
rect 39060 37540 39140 37550
rect 39380 37540 39460 37550
rect 39700 37540 39780 37550
rect 40020 37540 40100 37550
rect 40340 37540 40420 37550
rect 40660 37540 40740 37550
rect 40980 37540 41060 37550
rect 41300 37540 41380 37550
rect 41620 37540 41700 37550
rect 41940 37540 42020 37550
rect 42260 37540 42340 37550
rect 42580 37540 42660 37550
rect 42900 37540 42980 37550
rect 43220 37540 43300 37550
rect 36260 37460 36270 37540
rect 36580 37460 36590 37540
rect 36900 37460 36910 37540
rect 37220 37460 37230 37540
rect 37540 37460 37550 37540
rect 37860 37460 37870 37540
rect 38180 37460 38190 37540
rect 38500 37460 38510 37540
rect 38820 37460 38830 37540
rect 39140 37460 39150 37540
rect 39460 37460 39470 37540
rect 39780 37460 39790 37540
rect 40100 37460 40110 37540
rect 40420 37460 40430 37540
rect 40740 37460 40750 37540
rect 41060 37460 41070 37540
rect 41380 37460 41390 37540
rect 41700 37460 41710 37540
rect 42020 37460 42030 37540
rect 42340 37460 42350 37540
rect 42660 37460 42670 37540
rect 42980 37460 42990 37540
rect 43300 37460 43310 37540
rect 43785 37480 43865 37490
rect 44105 37480 44185 37490
rect 44425 37480 44505 37490
rect 44745 37480 44825 37490
rect 45065 37480 45145 37490
rect 45385 37480 45465 37490
rect 45705 37480 45785 37490
rect 46025 37480 46105 37490
rect 46345 37480 46425 37490
rect 46665 37480 46745 37490
rect 46985 37480 47065 37490
rect 47305 37480 47385 37490
rect 47625 37480 47705 37490
rect 47945 37480 48025 37490
rect 48265 37480 48345 37490
rect 43865 37400 43875 37480
rect 44185 37400 44195 37480
rect 44505 37400 44515 37480
rect 44825 37400 44835 37480
rect 45145 37400 45155 37480
rect 45465 37400 45475 37480
rect 45785 37400 45795 37480
rect 46105 37400 46115 37480
rect 46425 37400 46435 37480
rect 46745 37400 46755 37480
rect 47065 37400 47075 37480
rect 47385 37400 47395 37480
rect 47705 37400 47715 37480
rect 48025 37400 48035 37480
rect 48345 37400 48355 37480
rect 48500 37390 48605 37560
rect 48640 37480 48650 37560
rect 48790 37480 48800 37560
rect 60140 37480 60150 37560
rect 60290 37480 60300 37560
rect 60440 37480 60450 37560
rect 60580 37480 60660 37490
rect 60900 37480 60980 37490
rect 61320 37480 61400 37490
rect 61640 37480 61720 37490
rect 62140 37480 62150 37560
rect 62290 37480 62300 37560
rect 73640 37480 73650 37560
rect 73790 37480 73800 37560
rect 73940 37480 73950 37560
rect 74080 37480 74160 37490
rect 74400 37480 74480 37490
rect 74820 37480 74900 37490
rect 75140 37480 75220 37490
rect 75640 37480 75650 37560
rect 75790 37480 75800 37560
rect 87140 37480 87150 37560
rect 87290 37480 87300 37560
rect 87440 37480 87450 37560
rect 87580 37480 87660 37490
rect 87900 37480 87980 37490
rect 88320 37480 88400 37490
rect 88640 37480 88720 37490
rect 89140 37480 89150 37560
rect 89290 37480 89300 37560
rect 100640 37480 100650 37560
rect 100790 37480 100800 37560
rect 100940 37480 100950 37560
rect 101080 37480 101160 37490
rect 101400 37480 101480 37490
rect 101820 37480 101900 37490
rect 102140 37480 102220 37490
rect 102640 37480 102650 37560
rect 102790 37480 102800 37560
rect 114140 37480 114150 37560
rect 114290 37480 114300 37560
rect 114440 37480 114450 37560
rect 114580 37480 114660 37490
rect 114900 37480 114980 37490
rect 115320 37480 115400 37490
rect 115640 37480 115720 37490
rect 116140 37480 116150 37560
rect 116290 37480 116300 37560
rect 127640 37480 127650 37560
rect 127790 37480 127800 37560
rect 127940 37480 127950 37560
rect 128080 37480 128160 37490
rect 128400 37480 128480 37490
rect 128820 37480 128900 37490
rect 129140 37480 129220 37490
rect 129640 37480 129650 37560
rect 129790 37480 129800 37560
rect 141140 37480 141150 37560
rect 141290 37480 141300 37560
rect 141440 37480 141450 37560
rect 60660 37400 60670 37480
rect 60980 37400 60990 37480
rect 61400 37400 61410 37480
rect 61720 37400 61730 37480
rect 74160 37400 74170 37480
rect 74480 37400 74490 37480
rect 74900 37400 74910 37480
rect 75220 37400 75230 37480
rect 87660 37400 87670 37480
rect 87980 37400 87990 37480
rect 88400 37400 88410 37480
rect 88720 37400 88730 37480
rect 101160 37400 101170 37480
rect 101480 37400 101490 37480
rect 101900 37400 101910 37480
rect 102220 37400 102230 37480
rect 114660 37400 114670 37480
rect 114980 37400 114990 37480
rect 115400 37400 115410 37480
rect 115720 37400 115730 37480
rect 128160 37400 128170 37480
rect 128480 37400 128490 37480
rect 128900 37400 128910 37480
rect 129220 37400 129230 37480
rect 36020 37380 36100 37390
rect 36340 37380 36420 37390
rect 36660 37380 36740 37390
rect 36980 37380 37060 37390
rect 37300 37380 37380 37390
rect 37620 37380 37700 37390
rect 37940 37380 38020 37390
rect 38260 37380 38340 37390
rect 38580 37380 38660 37390
rect 38900 37380 38980 37390
rect 39220 37380 39300 37390
rect 39540 37380 39620 37390
rect 39860 37380 39940 37390
rect 40180 37380 40260 37390
rect 40500 37380 40580 37390
rect 40820 37380 40900 37390
rect 41140 37380 41220 37390
rect 41460 37380 41540 37390
rect 41780 37380 41860 37390
rect 42100 37380 42180 37390
rect 42420 37380 42500 37390
rect 42740 37380 42820 37390
rect 43060 37380 43140 37390
rect 43380 37380 43460 37390
rect 48500 37380 48640 37390
rect 48710 37380 48790 37390
rect 60060 37380 60140 37390
rect 60210 37380 60290 37390
rect 60360 37380 60440 37390
rect 62060 37380 62140 37390
rect 62210 37380 62290 37390
rect 73560 37380 73640 37390
rect 73710 37380 73790 37390
rect 73860 37380 73940 37390
rect 75560 37380 75640 37390
rect 75710 37380 75790 37390
rect 87060 37380 87140 37390
rect 87210 37380 87290 37390
rect 87360 37380 87440 37390
rect 89060 37380 89140 37390
rect 89210 37380 89290 37390
rect 100560 37380 100640 37390
rect 100710 37380 100790 37390
rect 100860 37380 100940 37390
rect 102560 37380 102640 37390
rect 102710 37380 102790 37390
rect 114060 37380 114140 37390
rect 114210 37380 114290 37390
rect 114360 37380 114440 37390
rect 116060 37380 116140 37390
rect 116210 37380 116290 37390
rect 127560 37380 127640 37390
rect 127710 37380 127790 37390
rect 127860 37380 127940 37390
rect 129560 37380 129640 37390
rect 129710 37380 129790 37390
rect 141060 37380 141140 37390
rect 141210 37380 141290 37390
rect 141360 37380 141440 37390
rect 36100 37300 36110 37380
rect 36420 37300 36430 37380
rect 36740 37300 36750 37380
rect 37060 37300 37070 37380
rect 37380 37300 37390 37380
rect 37700 37300 37710 37380
rect 38020 37300 38030 37380
rect 38340 37300 38350 37380
rect 38660 37300 38670 37380
rect 38980 37300 38990 37380
rect 39300 37300 39310 37380
rect 39620 37300 39630 37380
rect 39940 37300 39950 37380
rect 40260 37300 40270 37380
rect 40580 37300 40590 37380
rect 40900 37300 40910 37380
rect 41220 37300 41230 37380
rect 41540 37300 41550 37380
rect 41860 37300 41870 37380
rect 42180 37300 42190 37380
rect 42500 37300 42510 37380
rect 42820 37300 42830 37380
rect 43140 37300 43150 37380
rect 43460 37300 43470 37380
rect 43945 37320 44025 37330
rect 44265 37320 44345 37330
rect 44585 37320 44665 37330
rect 44905 37320 44985 37330
rect 45225 37320 45305 37330
rect 45545 37320 45625 37330
rect 45865 37320 45945 37330
rect 46185 37320 46265 37330
rect 46505 37320 46585 37330
rect 46825 37320 46905 37330
rect 47145 37320 47225 37330
rect 47465 37320 47545 37330
rect 47785 37320 47865 37330
rect 48105 37320 48185 37330
rect 44025 37240 44035 37320
rect 44345 37240 44355 37320
rect 44665 37240 44675 37320
rect 44985 37240 44995 37320
rect 45305 37240 45315 37320
rect 45625 37240 45635 37320
rect 45945 37240 45955 37320
rect 46265 37240 46275 37320
rect 46585 37240 46595 37320
rect 46905 37240 46915 37320
rect 47225 37240 47235 37320
rect 47545 37240 47555 37320
rect 47865 37240 47875 37320
rect 48185 37240 48195 37320
rect 36180 37220 36260 37230
rect 36500 37220 36580 37230
rect 36820 37220 36900 37230
rect 37140 37220 37220 37230
rect 37460 37220 37540 37230
rect 37780 37220 37860 37230
rect 38100 37220 38180 37230
rect 38420 37220 38500 37230
rect 38740 37220 38820 37230
rect 39060 37220 39140 37230
rect 39380 37220 39460 37230
rect 39700 37220 39780 37230
rect 40020 37220 40100 37230
rect 40340 37220 40420 37230
rect 40660 37220 40740 37230
rect 40980 37220 41060 37230
rect 41300 37220 41380 37230
rect 41620 37220 41700 37230
rect 41940 37220 42020 37230
rect 42260 37220 42340 37230
rect 42580 37220 42660 37230
rect 42900 37220 42980 37230
rect 43220 37220 43300 37230
rect 36260 37140 36270 37220
rect 36580 37140 36590 37220
rect 36900 37140 36910 37220
rect 37220 37140 37230 37220
rect 37540 37140 37550 37220
rect 37860 37140 37870 37220
rect 38180 37140 38190 37220
rect 38500 37140 38510 37220
rect 38820 37140 38830 37220
rect 39140 37140 39150 37220
rect 39460 37140 39470 37220
rect 39780 37140 39790 37220
rect 40100 37140 40110 37220
rect 40420 37140 40430 37220
rect 40740 37140 40750 37220
rect 41060 37140 41070 37220
rect 41380 37140 41390 37220
rect 41700 37140 41710 37220
rect 42020 37140 42030 37220
rect 42340 37140 42350 37220
rect 42660 37140 42670 37220
rect 42980 37140 42990 37220
rect 43300 37140 43310 37220
rect 48500 37210 48605 37380
rect 48640 37300 48650 37380
rect 48790 37300 48800 37380
rect 60140 37300 60150 37380
rect 60290 37300 60300 37380
rect 60440 37300 60450 37380
rect 60740 37320 60820 37330
rect 61060 37320 61140 37330
rect 61480 37320 61560 37330
rect 61800 37320 61880 37330
rect 60820 37240 60830 37320
rect 61140 37240 61150 37320
rect 61560 37240 61570 37320
rect 61880 37240 61890 37320
rect 62140 37300 62150 37380
rect 62290 37300 62300 37380
rect 73640 37300 73650 37380
rect 73790 37300 73800 37380
rect 73940 37300 73950 37380
rect 74240 37320 74320 37330
rect 74560 37320 74640 37330
rect 74980 37320 75060 37330
rect 75300 37320 75380 37330
rect 74320 37240 74330 37320
rect 74640 37240 74650 37320
rect 75060 37240 75070 37320
rect 75380 37240 75390 37320
rect 75640 37300 75650 37380
rect 75790 37300 75800 37380
rect 87140 37300 87150 37380
rect 87290 37300 87300 37380
rect 87440 37300 87450 37380
rect 87740 37320 87820 37330
rect 88060 37320 88140 37330
rect 88480 37320 88560 37330
rect 88800 37320 88880 37330
rect 87820 37240 87830 37320
rect 88140 37240 88150 37320
rect 88560 37240 88570 37320
rect 88880 37240 88890 37320
rect 89140 37300 89150 37380
rect 89290 37300 89300 37380
rect 100640 37300 100650 37380
rect 100790 37300 100800 37380
rect 100940 37300 100950 37380
rect 101240 37320 101320 37330
rect 101560 37320 101640 37330
rect 101980 37320 102060 37330
rect 102300 37320 102380 37330
rect 101320 37240 101330 37320
rect 101640 37240 101650 37320
rect 102060 37240 102070 37320
rect 102380 37240 102390 37320
rect 102640 37300 102650 37380
rect 102790 37300 102800 37380
rect 114140 37300 114150 37380
rect 114290 37300 114300 37380
rect 114440 37300 114450 37380
rect 114740 37320 114820 37330
rect 115060 37320 115140 37330
rect 115480 37320 115560 37330
rect 115800 37320 115880 37330
rect 114820 37240 114830 37320
rect 115140 37240 115150 37320
rect 115560 37240 115570 37320
rect 115880 37240 115890 37320
rect 116140 37300 116150 37380
rect 116290 37300 116300 37380
rect 127640 37300 127650 37380
rect 127790 37300 127800 37380
rect 127940 37300 127950 37380
rect 128240 37320 128320 37330
rect 128560 37320 128640 37330
rect 128980 37320 129060 37330
rect 129300 37320 129380 37330
rect 128320 37240 128330 37320
rect 128640 37240 128650 37320
rect 129060 37240 129070 37320
rect 129380 37240 129390 37320
rect 129640 37300 129650 37380
rect 129790 37300 129800 37380
rect 141140 37300 141150 37380
rect 141290 37300 141300 37380
rect 141440 37300 141450 37380
rect 48500 37200 48640 37210
rect 48710 37200 48790 37210
rect 60060 37200 60140 37210
rect 60210 37200 60290 37210
rect 60360 37200 60440 37210
rect 62060 37200 62140 37210
rect 62210 37200 62290 37210
rect 73560 37200 73640 37210
rect 73710 37200 73790 37210
rect 73860 37200 73940 37210
rect 75560 37200 75640 37210
rect 75710 37200 75790 37210
rect 87060 37200 87140 37210
rect 87210 37200 87290 37210
rect 87360 37200 87440 37210
rect 89060 37200 89140 37210
rect 89210 37200 89290 37210
rect 100560 37200 100640 37210
rect 100710 37200 100790 37210
rect 100860 37200 100940 37210
rect 102560 37200 102640 37210
rect 102710 37200 102790 37210
rect 114060 37200 114140 37210
rect 114210 37200 114290 37210
rect 114360 37200 114440 37210
rect 116060 37200 116140 37210
rect 116210 37200 116290 37210
rect 127560 37200 127640 37210
rect 127710 37200 127790 37210
rect 127860 37200 127940 37210
rect 129560 37200 129640 37210
rect 129710 37200 129790 37210
rect 141060 37200 141140 37210
rect 141210 37200 141290 37210
rect 141360 37200 141440 37210
rect 43785 37160 43865 37170
rect 44105 37160 44185 37170
rect 44425 37160 44505 37170
rect 44745 37160 44825 37170
rect 45065 37160 45145 37170
rect 45385 37160 45465 37170
rect 45705 37160 45785 37170
rect 46025 37160 46105 37170
rect 46345 37160 46425 37170
rect 46665 37160 46745 37170
rect 46985 37160 47065 37170
rect 47305 37160 47385 37170
rect 47625 37160 47705 37170
rect 47945 37160 48025 37170
rect 48265 37160 48345 37170
rect 43865 37080 43875 37160
rect 44185 37080 44195 37160
rect 44505 37080 44515 37160
rect 44825 37080 44835 37160
rect 45145 37080 45155 37160
rect 45465 37080 45475 37160
rect 45785 37080 45795 37160
rect 46105 37080 46115 37160
rect 46425 37080 46435 37160
rect 46745 37080 46755 37160
rect 47065 37080 47075 37160
rect 47385 37080 47395 37160
rect 47705 37080 47715 37160
rect 48025 37080 48035 37160
rect 48345 37080 48355 37160
rect 36020 37060 36100 37070
rect 36340 37060 36420 37070
rect 36660 37060 36740 37070
rect 36980 37060 37060 37070
rect 37300 37060 37380 37070
rect 37620 37060 37700 37070
rect 37940 37060 38020 37070
rect 38260 37060 38340 37070
rect 38580 37060 38660 37070
rect 38900 37060 38980 37070
rect 39220 37060 39300 37070
rect 39540 37060 39620 37070
rect 39860 37060 39940 37070
rect 40180 37060 40260 37070
rect 40500 37060 40580 37070
rect 40820 37060 40900 37070
rect 41140 37060 41220 37070
rect 41460 37060 41540 37070
rect 41780 37060 41860 37070
rect 42100 37060 42180 37070
rect 42420 37060 42500 37070
rect 42740 37060 42820 37070
rect 43060 37060 43140 37070
rect 43380 37060 43460 37070
rect 36100 36980 36110 37060
rect 36420 36980 36430 37060
rect 36740 36980 36750 37060
rect 37060 36980 37070 37060
rect 37380 36980 37390 37060
rect 37700 36980 37710 37060
rect 38020 36980 38030 37060
rect 38340 36980 38350 37060
rect 38660 36980 38670 37060
rect 38980 36980 38990 37060
rect 39300 36980 39310 37060
rect 39620 36980 39630 37060
rect 39940 36980 39950 37060
rect 40260 36980 40270 37060
rect 40580 36980 40590 37060
rect 40900 36980 40910 37060
rect 41220 36980 41230 37060
rect 41540 36980 41550 37060
rect 41860 36980 41870 37060
rect 42180 36980 42190 37060
rect 42500 36980 42510 37060
rect 42820 36980 42830 37060
rect 43140 36980 43150 37060
rect 43460 36980 43470 37060
rect 48500 37030 48605 37200
rect 48640 37120 48650 37200
rect 48790 37120 48800 37200
rect 49240 37100 59760 37190
rect 60140 37120 60150 37200
rect 60290 37120 60300 37200
rect 60440 37120 60450 37200
rect 60580 37160 60660 37170
rect 60900 37160 60980 37170
rect 61320 37160 61400 37170
rect 61640 37160 61720 37170
rect 49560 37030 49590 37100
rect 48500 37020 48640 37030
rect 48710 37020 48790 37030
rect 49270 37020 49350 37030
rect 49420 37020 49500 37030
rect 49560 37020 49650 37030
rect 49660 37020 49690 37100
rect 43945 37000 44025 37010
rect 44265 37000 44345 37010
rect 44585 37000 44665 37010
rect 44905 37000 44985 37010
rect 45225 37000 45305 37010
rect 45545 37000 45625 37010
rect 45865 37000 45945 37010
rect 46185 37000 46265 37010
rect 46505 37000 46585 37010
rect 46825 37000 46905 37010
rect 47145 37000 47225 37010
rect 47465 37000 47545 37010
rect 47785 37000 47865 37010
rect 48105 37000 48185 37010
rect 44025 36920 44035 37000
rect 44345 36920 44355 37000
rect 44665 36920 44675 37000
rect 44985 36920 44995 37000
rect 45305 36920 45315 37000
rect 45625 36920 45635 37000
rect 45945 36920 45955 37000
rect 46265 36920 46275 37000
rect 46585 36920 46595 37000
rect 46905 36920 46915 37000
rect 47225 36920 47235 37000
rect 47545 36920 47555 37000
rect 47865 36920 47875 37000
rect 48185 36920 48195 37000
rect 36180 36900 36260 36910
rect 36500 36900 36580 36910
rect 36820 36900 36900 36910
rect 37140 36900 37220 36910
rect 37460 36900 37540 36910
rect 37780 36900 37860 36910
rect 38100 36900 38180 36910
rect 38420 36900 38500 36910
rect 38740 36900 38820 36910
rect 39060 36900 39140 36910
rect 39380 36900 39460 36910
rect 39700 36900 39780 36910
rect 40020 36900 40100 36910
rect 40340 36900 40420 36910
rect 40660 36900 40740 36910
rect 40980 36900 41060 36910
rect 41300 36900 41380 36910
rect 41620 36900 41700 36910
rect 41940 36900 42020 36910
rect 42260 36900 42340 36910
rect 42580 36900 42660 36910
rect 42900 36900 42980 36910
rect 43220 36900 43300 36910
rect 36260 36820 36270 36900
rect 36580 36820 36590 36900
rect 36900 36820 36910 36900
rect 37220 36820 37230 36900
rect 37540 36820 37550 36900
rect 37860 36820 37870 36900
rect 38180 36820 38190 36900
rect 38500 36820 38510 36900
rect 38820 36820 38830 36900
rect 39140 36820 39150 36900
rect 39460 36820 39470 36900
rect 39780 36820 39790 36900
rect 40100 36820 40110 36900
rect 40420 36820 40430 36900
rect 40740 36820 40750 36900
rect 41060 36820 41070 36900
rect 41380 36820 41390 36900
rect 41700 36820 41710 36900
rect 42020 36820 42030 36900
rect 42340 36820 42350 36900
rect 42660 36820 42670 36900
rect 42980 36820 42990 36900
rect 43300 36820 43310 36900
rect 48500 36850 48605 37020
rect 48640 36940 48650 37020
rect 48790 36940 48800 37020
rect 49350 36940 49360 37020
rect 49500 36940 49510 37020
rect 49560 36850 49590 37020
rect 49650 36940 49690 37020
rect 43785 36840 43865 36850
rect 44105 36840 44185 36850
rect 44425 36840 44505 36850
rect 44745 36840 44825 36850
rect 45065 36840 45145 36850
rect 45385 36840 45465 36850
rect 45705 36840 45785 36850
rect 46025 36840 46105 36850
rect 46345 36840 46425 36850
rect 46665 36840 46745 36850
rect 46985 36840 47065 36850
rect 47305 36840 47385 36850
rect 47625 36840 47705 36850
rect 47945 36840 48025 36850
rect 48265 36840 48345 36850
rect 48500 36840 48640 36850
rect 48710 36840 48790 36850
rect 49270 36840 49350 36850
rect 49420 36840 49500 36850
rect 49560 36840 49650 36850
rect 49660 36840 49690 36940
rect 43865 36760 43875 36840
rect 44185 36760 44195 36840
rect 44505 36760 44515 36840
rect 44825 36760 44835 36840
rect 45145 36760 45155 36840
rect 45465 36760 45475 36840
rect 45785 36760 45795 36840
rect 46105 36760 46115 36840
rect 46425 36760 46435 36840
rect 46745 36760 46755 36840
rect 47065 36760 47075 36840
rect 47385 36760 47395 36840
rect 47705 36760 47715 36840
rect 48025 36760 48035 36840
rect 48345 36760 48355 36840
rect 36020 36740 36100 36750
rect 36340 36740 36420 36750
rect 36660 36740 36740 36750
rect 36980 36740 37060 36750
rect 37300 36740 37380 36750
rect 37620 36740 37700 36750
rect 37940 36740 38020 36750
rect 38260 36740 38340 36750
rect 38580 36740 38660 36750
rect 38900 36740 38980 36750
rect 39220 36740 39300 36750
rect 39540 36740 39620 36750
rect 39860 36740 39940 36750
rect 40180 36740 40260 36750
rect 40500 36740 40580 36750
rect 40820 36740 40900 36750
rect 41140 36740 41220 36750
rect 41460 36740 41540 36750
rect 41780 36740 41860 36750
rect 42100 36740 42180 36750
rect 42420 36740 42500 36750
rect 42740 36740 42820 36750
rect 43060 36740 43140 36750
rect 43380 36740 43460 36750
rect 36100 36660 36110 36740
rect 36420 36660 36430 36740
rect 36740 36660 36750 36740
rect 37060 36660 37070 36740
rect 37380 36660 37390 36740
rect 37700 36660 37710 36740
rect 38020 36660 38030 36740
rect 38340 36660 38350 36740
rect 38660 36660 38670 36740
rect 38980 36660 38990 36740
rect 39300 36660 39310 36740
rect 39620 36660 39630 36740
rect 39940 36660 39950 36740
rect 40260 36660 40270 36740
rect 40580 36660 40590 36740
rect 40900 36660 40910 36740
rect 41220 36660 41230 36740
rect 41540 36660 41550 36740
rect 41860 36660 41870 36740
rect 42180 36660 42190 36740
rect 42500 36660 42510 36740
rect 42820 36660 42830 36740
rect 43140 36660 43150 36740
rect 43460 36660 43470 36740
rect 43945 36680 44025 36690
rect 44265 36680 44345 36690
rect 44585 36680 44665 36690
rect 44905 36680 44985 36690
rect 45225 36680 45305 36690
rect 45545 36680 45625 36690
rect 45865 36680 45945 36690
rect 46185 36680 46265 36690
rect 46505 36680 46585 36690
rect 46825 36680 46905 36690
rect 47145 36680 47225 36690
rect 47465 36680 47545 36690
rect 47785 36680 47865 36690
rect 48105 36680 48185 36690
rect 44025 36600 44035 36680
rect 44345 36600 44355 36680
rect 44665 36600 44675 36680
rect 44985 36600 44995 36680
rect 45305 36600 45315 36680
rect 45625 36600 45635 36680
rect 45945 36600 45955 36680
rect 46265 36600 46275 36680
rect 46585 36600 46595 36680
rect 46905 36600 46915 36680
rect 47225 36600 47235 36680
rect 47545 36600 47555 36680
rect 47865 36600 47875 36680
rect 48185 36600 48195 36680
rect 48500 36670 48605 36840
rect 48640 36760 48650 36840
rect 48790 36760 48800 36840
rect 49350 36760 49360 36840
rect 49500 36760 49510 36840
rect 49560 36670 49590 36840
rect 49650 36760 49690 36840
rect 48500 36660 48640 36670
rect 48710 36660 48790 36670
rect 49270 36660 49350 36670
rect 49420 36660 49500 36670
rect 49560 36660 49650 36670
rect 49660 36660 49690 36760
rect 36180 36580 36260 36590
rect 36500 36580 36580 36590
rect 36820 36580 36900 36590
rect 37140 36580 37220 36590
rect 37460 36580 37540 36590
rect 37780 36580 37860 36590
rect 38100 36580 38180 36590
rect 38420 36580 38500 36590
rect 38740 36580 38820 36590
rect 39060 36580 39140 36590
rect 39380 36580 39460 36590
rect 39700 36580 39780 36590
rect 40020 36580 40100 36590
rect 40340 36580 40420 36590
rect 40660 36580 40740 36590
rect 40980 36580 41060 36590
rect 41300 36580 41380 36590
rect 41620 36580 41700 36590
rect 41940 36580 42020 36590
rect 42260 36580 42340 36590
rect 42580 36580 42660 36590
rect 42900 36580 42980 36590
rect 43220 36580 43300 36590
rect 36260 36500 36270 36580
rect 36580 36500 36590 36580
rect 36900 36500 36910 36580
rect 37220 36500 37230 36580
rect 37540 36500 37550 36580
rect 37860 36500 37870 36580
rect 38180 36500 38190 36580
rect 38500 36500 38510 36580
rect 38820 36500 38830 36580
rect 39140 36500 39150 36580
rect 39460 36500 39470 36580
rect 39780 36500 39790 36580
rect 40100 36500 40110 36580
rect 40420 36500 40430 36580
rect 40740 36500 40750 36580
rect 41060 36500 41070 36580
rect 41380 36500 41390 36580
rect 41700 36500 41710 36580
rect 42020 36500 42030 36580
rect 42340 36500 42350 36580
rect 42660 36500 42670 36580
rect 42980 36500 42990 36580
rect 43300 36500 43310 36580
rect 43785 36520 43865 36530
rect 44105 36520 44185 36530
rect 44425 36520 44505 36530
rect 44745 36520 44825 36530
rect 45065 36520 45145 36530
rect 45385 36520 45465 36530
rect 45705 36520 45785 36530
rect 46025 36520 46105 36530
rect 46345 36520 46425 36530
rect 46665 36520 46745 36530
rect 46985 36520 47065 36530
rect 47305 36520 47385 36530
rect 47625 36520 47705 36530
rect 47945 36520 48025 36530
rect 48265 36520 48345 36530
rect 43865 36440 43875 36520
rect 44185 36440 44195 36520
rect 44505 36440 44515 36520
rect 44825 36440 44835 36520
rect 45145 36440 45155 36520
rect 45465 36440 45475 36520
rect 45785 36440 45795 36520
rect 46105 36440 46115 36520
rect 46425 36440 46435 36520
rect 46745 36440 46755 36520
rect 47065 36440 47075 36520
rect 47385 36440 47395 36520
rect 47705 36440 47715 36520
rect 48025 36440 48035 36520
rect 48345 36440 48355 36520
rect 48500 36490 48605 36660
rect 48640 36580 48650 36660
rect 48790 36580 48800 36660
rect 49350 36580 49360 36660
rect 49500 36580 49510 36660
rect 49560 36490 49590 36660
rect 49650 36580 49690 36660
rect 48500 36480 48640 36490
rect 48710 36480 48790 36490
rect 49270 36480 49350 36490
rect 49420 36480 49500 36490
rect 49560 36480 49650 36490
rect 49660 36480 49690 36580
rect 36020 36420 36100 36430
rect 36340 36420 36420 36430
rect 36660 36420 36740 36430
rect 36980 36420 37060 36430
rect 37300 36420 37380 36430
rect 37620 36420 37700 36430
rect 37940 36420 38020 36430
rect 38260 36420 38340 36430
rect 38580 36420 38660 36430
rect 38900 36420 38980 36430
rect 39220 36420 39300 36430
rect 39540 36420 39620 36430
rect 39860 36420 39940 36430
rect 40180 36420 40260 36430
rect 40500 36420 40580 36430
rect 40820 36420 40900 36430
rect 41140 36420 41220 36430
rect 41460 36420 41540 36430
rect 41780 36420 41860 36430
rect 42100 36420 42180 36430
rect 42420 36420 42500 36430
rect 42740 36420 42820 36430
rect 43060 36420 43140 36430
rect 43380 36420 43460 36430
rect 36100 36340 36110 36420
rect 36420 36340 36430 36420
rect 36740 36340 36750 36420
rect 37060 36340 37070 36420
rect 37380 36340 37390 36420
rect 37700 36340 37710 36420
rect 38020 36340 38030 36420
rect 38340 36340 38350 36420
rect 38660 36340 38670 36420
rect 38980 36340 38990 36420
rect 39300 36340 39310 36420
rect 39620 36340 39630 36420
rect 39940 36340 39950 36420
rect 40260 36340 40270 36420
rect 40580 36340 40590 36420
rect 40900 36340 40910 36420
rect 41220 36340 41230 36420
rect 41540 36340 41550 36420
rect 41860 36340 41870 36420
rect 42180 36340 42190 36420
rect 42500 36340 42510 36420
rect 42820 36340 42830 36420
rect 43140 36340 43150 36420
rect 43460 36340 43470 36420
rect 43945 36360 44025 36370
rect 44265 36360 44345 36370
rect 44585 36360 44665 36370
rect 44905 36360 44985 36370
rect 45225 36360 45305 36370
rect 45545 36360 45625 36370
rect 45865 36360 45945 36370
rect 46185 36360 46265 36370
rect 46505 36360 46585 36370
rect 46825 36360 46905 36370
rect 47145 36360 47225 36370
rect 47465 36360 47545 36370
rect 47785 36360 47865 36370
rect 48105 36360 48185 36370
rect 44025 36280 44035 36360
rect 44345 36280 44355 36360
rect 44665 36280 44675 36360
rect 44985 36280 44995 36360
rect 45305 36280 45315 36360
rect 45625 36280 45635 36360
rect 45945 36280 45955 36360
rect 46265 36280 46275 36360
rect 46585 36280 46595 36360
rect 46905 36280 46915 36360
rect 47225 36280 47235 36360
rect 47545 36280 47555 36360
rect 47865 36280 47875 36360
rect 48185 36280 48195 36360
rect 48500 36310 48605 36480
rect 48640 36400 48650 36480
rect 48790 36400 48800 36480
rect 49350 36400 49360 36480
rect 49500 36400 49510 36480
rect 49560 36310 49590 36480
rect 49650 36400 49690 36480
rect 48500 36300 48640 36310
rect 48710 36300 48790 36310
rect 49270 36300 49350 36310
rect 49420 36300 49500 36310
rect 49560 36300 49650 36310
rect 49660 36300 49690 36400
rect 36180 36260 36260 36270
rect 36500 36260 36580 36270
rect 36820 36260 36900 36270
rect 37140 36260 37220 36270
rect 37460 36260 37540 36270
rect 37780 36260 37860 36270
rect 38100 36260 38180 36270
rect 38420 36260 38500 36270
rect 38740 36260 38820 36270
rect 39060 36260 39140 36270
rect 39380 36260 39460 36270
rect 39700 36260 39780 36270
rect 40020 36260 40100 36270
rect 40340 36260 40420 36270
rect 40660 36260 40740 36270
rect 40980 36260 41060 36270
rect 41300 36260 41380 36270
rect 41620 36260 41700 36270
rect 41940 36260 42020 36270
rect 42260 36260 42340 36270
rect 42580 36260 42660 36270
rect 42900 36260 42980 36270
rect 43220 36260 43300 36270
rect 36260 36180 36270 36260
rect 36580 36180 36590 36260
rect 36900 36180 36910 36260
rect 37220 36180 37230 36260
rect 37540 36180 37550 36260
rect 37860 36180 37870 36260
rect 38180 36180 38190 36260
rect 38500 36180 38510 36260
rect 38820 36180 38830 36260
rect 39140 36180 39150 36260
rect 39460 36180 39470 36260
rect 39780 36180 39790 36260
rect 40100 36180 40110 36260
rect 40420 36180 40430 36260
rect 40740 36180 40750 36260
rect 41060 36180 41070 36260
rect 41380 36180 41390 36260
rect 41700 36180 41710 36260
rect 42020 36180 42030 36260
rect 42340 36180 42350 36260
rect 42660 36180 42670 36260
rect 42980 36180 42990 36260
rect 43300 36180 43310 36260
rect 43785 36200 43865 36210
rect 44105 36200 44185 36210
rect 44425 36200 44505 36210
rect 44745 36200 44825 36210
rect 45065 36200 45145 36210
rect 45385 36200 45465 36210
rect 45705 36200 45785 36210
rect 46025 36200 46105 36210
rect 46345 36200 46425 36210
rect 46665 36200 46745 36210
rect 46985 36200 47065 36210
rect 47305 36200 47385 36210
rect 47625 36200 47705 36210
rect 47945 36200 48025 36210
rect 48265 36200 48345 36210
rect 43865 36120 43875 36200
rect 44185 36120 44195 36200
rect 44505 36120 44515 36200
rect 44825 36120 44835 36200
rect 45145 36120 45155 36200
rect 45465 36120 45475 36200
rect 45785 36120 45795 36200
rect 46105 36120 46115 36200
rect 46425 36120 46435 36200
rect 46745 36120 46755 36200
rect 47065 36120 47075 36200
rect 47385 36120 47395 36200
rect 47705 36120 47715 36200
rect 48025 36120 48035 36200
rect 48345 36120 48355 36200
rect 48500 36130 48605 36300
rect 48640 36220 48650 36300
rect 48790 36220 48800 36300
rect 49350 36220 49360 36300
rect 49500 36220 49510 36300
rect 49560 36130 49590 36300
rect 49650 36220 49690 36300
rect 48500 36120 48640 36130
rect 48710 36120 48790 36130
rect 49270 36120 49350 36130
rect 49420 36120 49500 36130
rect 49560 36120 49650 36130
rect 49660 36120 49690 36220
rect 36020 36100 36100 36110
rect 36340 36100 36420 36110
rect 36660 36100 36740 36110
rect 36980 36100 37060 36110
rect 37300 36100 37380 36110
rect 37620 36100 37700 36110
rect 37940 36100 38020 36110
rect 38260 36100 38340 36110
rect 38580 36100 38660 36110
rect 38900 36100 38980 36110
rect 39220 36100 39300 36110
rect 39540 36100 39620 36110
rect 39860 36100 39940 36110
rect 40180 36100 40260 36110
rect 40500 36100 40580 36110
rect 40820 36100 40900 36110
rect 41140 36100 41220 36110
rect 41460 36100 41540 36110
rect 41780 36100 41860 36110
rect 42100 36100 42180 36110
rect 42420 36100 42500 36110
rect 42740 36100 42820 36110
rect 43060 36100 43140 36110
rect 43380 36100 43460 36110
rect 36100 36020 36110 36100
rect 36420 36020 36430 36100
rect 36740 36020 36750 36100
rect 37060 36020 37070 36100
rect 37380 36020 37390 36100
rect 37700 36020 37710 36100
rect 38020 36020 38030 36100
rect 38340 36020 38350 36100
rect 38660 36020 38670 36100
rect 38980 36020 38990 36100
rect 39300 36020 39310 36100
rect 39620 36020 39630 36100
rect 39940 36020 39950 36100
rect 40260 36020 40270 36100
rect 40580 36020 40590 36100
rect 40900 36020 40910 36100
rect 41220 36020 41230 36100
rect 41540 36020 41550 36100
rect 41860 36020 41870 36100
rect 42180 36020 42190 36100
rect 42500 36020 42510 36100
rect 42820 36020 42830 36100
rect 43140 36020 43150 36100
rect 43460 36020 43470 36100
rect 43945 36040 44025 36050
rect 44265 36040 44345 36050
rect 44585 36040 44665 36050
rect 44905 36040 44985 36050
rect 45225 36040 45305 36050
rect 45545 36040 45625 36050
rect 45865 36040 45945 36050
rect 46185 36040 46265 36050
rect 46505 36040 46585 36050
rect 46825 36040 46905 36050
rect 47145 36040 47225 36050
rect 47465 36040 47545 36050
rect 47785 36040 47865 36050
rect 48105 36040 48185 36050
rect 44025 35960 44035 36040
rect 44345 35960 44355 36040
rect 44665 35960 44675 36040
rect 44985 35960 44995 36040
rect 45305 35960 45315 36040
rect 45625 35960 45635 36040
rect 45945 35960 45955 36040
rect 46265 35960 46275 36040
rect 46585 35960 46595 36040
rect 46905 35960 46915 36040
rect 47225 35960 47235 36040
rect 47545 35960 47555 36040
rect 47865 35960 47875 36040
rect 48185 35960 48195 36040
rect 48500 35950 48605 36120
rect 48640 36040 48650 36120
rect 48790 36040 48800 36120
rect 49350 36040 49360 36120
rect 49500 36040 49510 36120
rect 49560 35950 49590 36120
rect 49650 36040 49690 36120
rect 42950 35940 42980 35950
rect 43220 35940 43300 35950
rect 48500 35940 48640 35950
rect 48710 35940 48790 35950
rect 49270 35940 49350 35950
rect 49420 35940 49500 35950
rect 49560 35940 49650 35950
rect 49660 35940 49690 36040
rect 42980 35860 42990 35940
rect 43300 35860 43310 35940
rect 43785 35880 43865 35890
rect 44105 35880 44185 35890
rect 44425 35880 44505 35890
rect 44745 35880 44825 35890
rect 45065 35880 45145 35890
rect 45385 35880 45465 35890
rect 45705 35880 45785 35890
rect 46025 35880 46105 35890
rect 46345 35880 46425 35890
rect 46665 35880 46745 35890
rect 46985 35880 47065 35890
rect 47305 35880 47385 35890
rect 47625 35880 47705 35890
rect 47945 35880 48025 35890
rect 48265 35880 48345 35890
rect 43865 35800 43875 35880
rect 44185 35800 44195 35880
rect 44505 35800 44515 35880
rect 44825 35800 44835 35880
rect 45145 35800 45155 35880
rect 45465 35800 45475 35880
rect 45785 35800 45795 35880
rect 46105 35800 46115 35880
rect 46425 35800 46435 35880
rect 46745 35800 46755 35880
rect 47065 35800 47075 35880
rect 47385 35800 47395 35880
rect 47705 35800 47715 35880
rect 48025 35800 48035 35880
rect 48345 35800 48355 35880
rect 43060 35780 43140 35790
rect 43380 35780 43460 35790
rect 43140 35700 43150 35780
rect 43460 35700 43470 35780
rect 48500 35770 48605 35940
rect 48640 35860 48650 35940
rect 48790 35860 48800 35940
rect 49350 35860 49360 35940
rect 49500 35860 49510 35940
rect 49560 35770 49590 35940
rect 49650 35860 49690 35940
rect 48500 35760 48640 35770
rect 48710 35760 48790 35770
rect 49270 35760 49350 35770
rect 49420 35760 49500 35770
rect 49560 35760 49650 35770
rect 49660 35760 49690 35860
rect 43945 35720 44025 35730
rect 44265 35720 44345 35730
rect 44585 35720 44665 35730
rect 44905 35720 44985 35730
rect 45225 35720 45305 35730
rect 45545 35720 45625 35730
rect 45865 35720 45945 35730
rect 46185 35720 46265 35730
rect 46505 35720 46585 35730
rect 46825 35720 46905 35730
rect 47145 35720 47225 35730
rect 47465 35720 47545 35730
rect 47785 35720 47865 35730
rect 48105 35720 48185 35730
rect 44025 35640 44035 35720
rect 44345 35640 44355 35720
rect 44665 35640 44675 35720
rect 44985 35640 44995 35720
rect 45305 35640 45315 35720
rect 45625 35640 45635 35720
rect 45945 35640 45955 35720
rect 46265 35640 46275 35720
rect 46585 35640 46595 35720
rect 46905 35640 46915 35720
rect 47225 35640 47235 35720
rect 47545 35640 47555 35720
rect 47865 35640 47875 35720
rect 48185 35640 48195 35720
rect 42950 35620 42980 35630
rect 43220 35620 43300 35630
rect 42980 35540 42990 35620
rect 43300 35540 43310 35620
rect 48500 35590 48605 35760
rect 48640 35680 48650 35760
rect 48790 35680 48800 35760
rect 49350 35680 49360 35760
rect 49500 35680 49510 35760
rect 49560 35590 49590 35760
rect 49650 35680 49690 35760
rect 48500 35580 48640 35590
rect 48710 35580 48790 35590
rect 49270 35580 49350 35590
rect 49420 35580 49500 35590
rect 49560 35580 49650 35590
rect 49660 35580 49690 35680
rect 43785 35560 43865 35570
rect 44105 35560 44185 35570
rect 44425 35560 44505 35570
rect 44745 35560 44825 35570
rect 45065 35560 45145 35570
rect 45385 35560 45465 35570
rect 45705 35560 45785 35570
rect 46025 35560 46105 35570
rect 46345 35560 46425 35570
rect 46665 35560 46745 35570
rect 46985 35560 47065 35570
rect 47305 35560 47385 35570
rect 47625 35560 47705 35570
rect 47945 35560 48025 35570
rect 48265 35560 48345 35570
rect 43865 35480 43875 35560
rect 44185 35480 44195 35560
rect 44505 35480 44515 35560
rect 44825 35480 44835 35560
rect 45145 35480 45155 35560
rect 45465 35480 45475 35560
rect 45785 35480 45795 35560
rect 46105 35480 46115 35560
rect 46425 35480 46435 35560
rect 46745 35480 46755 35560
rect 47065 35480 47075 35560
rect 47385 35480 47395 35560
rect 47705 35480 47715 35560
rect 48025 35480 48035 35560
rect 48345 35480 48355 35560
rect 43060 35460 43140 35470
rect 43380 35460 43460 35470
rect 43140 35380 43150 35460
rect 43460 35380 43470 35460
rect 48500 35410 48605 35580
rect 48640 35500 48650 35580
rect 48790 35500 48800 35580
rect 49350 35500 49360 35580
rect 49500 35500 49510 35580
rect 49560 35410 49590 35580
rect 49650 35500 49690 35580
rect 43945 35400 44025 35410
rect 44265 35400 44345 35410
rect 44585 35400 44665 35410
rect 44905 35400 44985 35410
rect 45225 35400 45305 35410
rect 45545 35400 45625 35410
rect 45865 35400 45945 35410
rect 46185 35400 46265 35410
rect 46505 35400 46585 35410
rect 46825 35400 46905 35410
rect 47145 35400 47225 35410
rect 47465 35400 47545 35410
rect 47785 35400 47865 35410
rect 48105 35400 48185 35410
rect 48500 35400 48640 35410
rect 48710 35400 48790 35410
rect 49270 35400 49350 35410
rect 49420 35400 49500 35410
rect 49560 35400 49650 35410
rect 49660 35400 49690 35500
rect 44025 35320 44035 35400
rect 44345 35320 44355 35400
rect 44665 35320 44675 35400
rect 44985 35320 44995 35400
rect 45305 35320 45315 35400
rect 45625 35320 45635 35400
rect 45945 35320 45955 35400
rect 46265 35320 46275 35400
rect 46585 35320 46595 35400
rect 46905 35320 46915 35400
rect 47225 35320 47235 35400
rect 47545 35320 47555 35400
rect 47865 35320 47875 35400
rect 48185 35320 48195 35400
rect 42950 35300 42980 35310
rect 43220 35300 43300 35310
rect 42980 35220 42990 35300
rect 43300 35220 43310 35300
rect 43785 35240 43865 35250
rect 44105 35240 44185 35250
rect 44425 35240 44505 35250
rect 44745 35240 44825 35250
rect 45065 35240 45145 35250
rect 45385 35240 45465 35250
rect 45705 35240 45785 35250
rect 46025 35240 46105 35250
rect 46345 35240 46425 35250
rect 46665 35240 46745 35250
rect 46985 35240 47065 35250
rect 47305 35240 47385 35250
rect 47625 35240 47705 35250
rect 47945 35240 48025 35250
rect 48265 35240 48345 35250
rect 43865 35160 43875 35240
rect 44185 35160 44195 35240
rect 44505 35160 44515 35240
rect 44825 35160 44835 35240
rect 45145 35160 45155 35240
rect 45465 35160 45475 35240
rect 45785 35160 45795 35240
rect 46105 35160 46115 35240
rect 46425 35160 46435 35240
rect 46745 35160 46755 35240
rect 47065 35160 47075 35240
rect 47385 35160 47395 35240
rect 47705 35160 47715 35240
rect 48025 35160 48035 35240
rect 48345 35160 48355 35240
rect 48500 35230 48605 35400
rect 48640 35320 48650 35400
rect 48790 35320 48800 35400
rect 49350 35320 49360 35400
rect 49500 35320 49510 35400
rect 49560 35230 49590 35400
rect 49650 35320 49690 35400
rect 48500 35220 48640 35230
rect 48710 35220 48790 35230
rect 49270 35220 49350 35230
rect 49420 35220 49500 35230
rect 49560 35220 49650 35230
rect 49660 35220 49690 35320
rect 43060 35140 43140 35150
rect 43380 35140 43460 35150
rect 43140 35060 43150 35140
rect 43460 35060 43470 35140
rect 43945 35080 44025 35090
rect 44265 35080 44345 35090
rect 44585 35080 44665 35090
rect 44905 35080 44985 35090
rect 45225 35080 45305 35090
rect 45545 35080 45625 35090
rect 45865 35080 45945 35090
rect 46185 35080 46265 35090
rect 46505 35080 46585 35090
rect 46825 35080 46905 35090
rect 47145 35080 47225 35090
rect 47465 35080 47545 35090
rect 47785 35080 47865 35090
rect 48105 35080 48185 35090
rect 44025 35000 44035 35080
rect 44345 35000 44355 35080
rect 44665 35000 44675 35080
rect 44985 35000 44995 35080
rect 45305 35000 45315 35080
rect 45625 35000 45635 35080
rect 45945 35000 45955 35080
rect 46265 35000 46275 35080
rect 46585 35000 46595 35080
rect 46905 35000 46915 35080
rect 47225 35000 47235 35080
rect 47545 35000 47555 35080
rect 47865 35000 47875 35080
rect 48185 35000 48195 35080
rect 48500 35050 48605 35220
rect 48640 35140 48650 35220
rect 48790 35140 48800 35220
rect 49350 35140 49360 35220
rect 49500 35140 49510 35220
rect 49560 35050 49590 35220
rect 49650 35140 49690 35220
rect 48500 35040 48640 35050
rect 48710 35040 48790 35050
rect 49270 35040 49350 35050
rect 49420 35040 49500 35050
rect 49560 35040 49650 35050
rect 49660 35040 49690 35140
rect 42950 34980 42980 34990
rect 43220 34980 43300 34990
rect 42980 34900 42990 34980
rect 43300 34900 43310 34980
rect 43785 34920 43865 34930
rect 44105 34920 44185 34930
rect 44425 34920 44505 34930
rect 44745 34920 44825 34930
rect 45065 34920 45145 34930
rect 45385 34920 45465 34930
rect 45705 34920 45785 34930
rect 46025 34920 46105 34930
rect 46345 34920 46425 34930
rect 46665 34920 46745 34930
rect 46985 34920 47065 34930
rect 47305 34920 47385 34930
rect 47625 34920 47705 34930
rect 47945 34920 48025 34930
rect 48265 34920 48345 34930
rect 43865 34840 43875 34920
rect 44185 34840 44195 34920
rect 44505 34840 44515 34920
rect 44825 34840 44835 34920
rect 45145 34840 45155 34920
rect 45465 34840 45475 34920
rect 45785 34840 45795 34920
rect 46105 34840 46115 34920
rect 46425 34840 46435 34920
rect 46745 34840 46755 34920
rect 47065 34840 47075 34920
rect 47385 34840 47395 34920
rect 47705 34840 47715 34920
rect 48025 34840 48035 34920
rect 48345 34840 48355 34920
rect 48500 34870 48605 35040
rect 48640 34960 48650 35040
rect 48790 34960 48800 35040
rect 49350 34960 49360 35040
rect 49500 34960 49510 35040
rect 49560 34870 49590 35040
rect 49650 34960 49690 35040
rect 48500 34860 48640 34870
rect 48710 34860 48790 34870
rect 49270 34860 49350 34870
rect 49420 34860 49500 34870
rect 49560 34860 49650 34870
rect 49660 34860 49690 34960
rect 43060 34820 43140 34830
rect 43380 34820 43460 34830
rect 43140 34740 43150 34820
rect 43460 34740 43470 34820
rect 43945 34760 44025 34770
rect 44265 34760 44345 34770
rect 44585 34760 44665 34770
rect 44905 34760 44985 34770
rect 45225 34760 45305 34770
rect 45545 34760 45625 34770
rect 45865 34760 45945 34770
rect 46185 34760 46265 34770
rect 46505 34760 46585 34770
rect 46825 34760 46905 34770
rect 47145 34760 47225 34770
rect 47465 34760 47545 34770
rect 47785 34760 47865 34770
rect 48105 34760 48185 34770
rect 44025 34680 44035 34760
rect 44345 34680 44355 34760
rect 44665 34680 44675 34760
rect 44985 34680 44995 34760
rect 45305 34680 45315 34760
rect 45625 34680 45635 34760
rect 45945 34680 45955 34760
rect 46265 34680 46275 34760
rect 46585 34680 46595 34760
rect 46905 34680 46915 34760
rect 47225 34680 47235 34760
rect 47545 34680 47555 34760
rect 47865 34680 47875 34760
rect 48185 34680 48195 34760
rect 48500 34690 48605 34860
rect 48640 34780 48650 34860
rect 48790 34780 48800 34860
rect 49350 34780 49360 34860
rect 49500 34780 49510 34860
rect 49560 34690 49590 34860
rect 49650 34780 49690 34860
rect 48500 34680 48640 34690
rect 48710 34680 48790 34690
rect 49270 34680 49350 34690
rect 49420 34680 49500 34690
rect 49560 34680 49650 34690
rect 49660 34680 49690 34780
rect 42950 34660 42980 34670
rect 43220 34660 43300 34670
rect 42980 34580 42990 34660
rect 43300 34580 43310 34660
rect 43785 34600 43865 34610
rect 44105 34600 44185 34610
rect 44425 34600 44505 34610
rect 44745 34600 44825 34610
rect 45065 34600 45145 34610
rect 45385 34600 45465 34610
rect 45705 34600 45785 34610
rect 46025 34600 46105 34610
rect 46345 34600 46425 34610
rect 46665 34600 46745 34610
rect 46985 34600 47065 34610
rect 47305 34600 47385 34610
rect 47625 34600 47705 34610
rect 47945 34600 48025 34610
rect 48265 34600 48345 34610
rect 43865 34520 43875 34600
rect 44185 34520 44195 34600
rect 44505 34520 44515 34600
rect 44825 34520 44835 34600
rect 45145 34520 45155 34600
rect 45465 34520 45475 34600
rect 45785 34520 45795 34600
rect 46105 34520 46115 34600
rect 46425 34520 46435 34600
rect 46745 34520 46755 34600
rect 47065 34520 47075 34600
rect 47385 34520 47395 34600
rect 47705 34520 47715 34600
rect 48025 34520 48035 34600
rect 48345 34520 48355 34600
rect 48500 34510 48605 34680
rect 48640 34600 48650 34680
rect 48790 34600 48800 34680
rect 49350 34600 49360 34680
rect 49500 34600 49510 34680
rect 49560 34510 49590 34680
rect 49650 34600 49690 34680
rect 43060 34500 43140 34510
rect 43380 34500 43460 34510
rect 48500 34500 48640 34510
rect 48710 34500 48790 34510
rect 49270 34500 49350 34510
rect 49420 34500 49500 34510
rect 49560 34500 49650 34510
rect 49660 34500 49690 34600
rect 43140 34420 43150 34500
rect 43460 34420 43470 34500
rect 43945 34440 44025 34450
rect 44265 34440 44345 34450
rect 44585 34440 44665 34450
rect 44905 34440 44985 34450
rect 45225 34440 45305 34450
rect 45545 34440 45625 34450
rect 45865 34440 45945 34450
rect 46185 34440 46265 34450
rect 46505 34440 46585 34450
rect 46825 34440 46905 34450
rect 47145 34440 47225 34450
rect 47465 34440 47545 34450
rect 47785 34440 47865 34450
rect 48105 34440 48185 34450
rect 44025 34360 44035 34440
rect 44345 34360 44355 34440
rect 44665 34360 44675 34440
rect 44985 34360 44995 34440
rect 45305 34360 45315 34440
rect 45625 34360 45635 34440
rect 45945 34360 45955 34440
rect 46265 34360 46275 34440
rect 46585 34360 46595 34440
rect 46905 34360 46915 34440
rect 47225 34360 47235 34440
rect 47545 34360 47555 34440
rect 47865 34360 47875 34440
rect 48185 34360 48195 34440
rect 42950 34340 42980 34350
rect 43220 34340 43300 34350
rect 42980 34260 42990 34340
rect 43300 34260 43310 34340
rect 48500 34330 48605 34500
rect 48640 34420 48650 34500
rect 48790 34420 48800 34500
rect 49350 34420 49360 34500
rect 49500 34420 49510 34500
rect 49560 34330 49590 34500
rect 49650 34420 49690 34500
rect 48500 34320 48640 34330
rect 48710 34320 48790 34330
rect 49270 34320 49350 34330
rect 49420 34320 49500 34330
rect 49560 34320 49650 34330
rect 49660 34320 49690 34420
rect 43785 34280 43865 34290
rect 44105 34280 44185 34290
rect 44425 34280 44505 34290
rect 44745 34280 44825 34290
rect 45065 34280 45145 34290
rect 45385 34280 45465 34290
rect 45705 34280 45785 34290
rect 46025 34280 46105 34290
rect 46345 34280 46425 34290
rect 46665 34280 46745 34290
rect 46985 34280 47065 34290
rect 47305 34280 47385 34290
rect 47625 34280 47705 34290
rect 47945 34280 48025 34290
rect 48265 34280 48345 34290
rect 43865 34200 43875 34280
rect 44185 34200 44195 34280
rect 44505 34200 44515 34280
rect 44825 34200 44835 34280
rect 45145 34200 45155 34280
rect 45465 34200 45475 34280
rect 45785 34200 45795 34280
rect 46105 34200 46115 34280
rect 46425 34200 46435 34280
rect 46745 34200 46755 34280
rect 47065 34200 47075 34280
rect 47385 34200 47395 34280
rect 47705 34200 47715 34280
rect 48025 34200 48035 34280
rect 48345 34200 48355 34280
rect 43060 34180 43140 34190
rect 43380 34180 43460 34190
rect 43140 34100 43150 34180
rect 43460 34100 43470 34180
rect 48500 34150 48605 34320
rect 48640 34240 48650 34320
rect 48790 34240 48800 34320
rect 49350 34240 49360 34320
rect 49500 34240 49510 34320
rect 49560 34150 49590 34320
rect 49650 34240 49690 34320
rect 48500 34140 48640 34150
rect 48710 34140 48790 34150
rect 49270 34140 49350 34150
rect 49420 34140 49500 34150
rect 49560 34140 49650 34150
rect 49660 34140 49690 34240
rect 43945 34120 44025 34130
rect 44265 34120 44345 34130
rect 44585 34120 44665 34130
rect 44905 34120 44985 34130
rect 45225 34120 45305 34130
rect 45545 34120 45625 34130
rect 45865 34120 45945 34130
rect 46185 34120 46265 34130
rect 46505 34120 46585 34130
rect 46825 34120 46905 34130
rect 47145 34120 47225 34130
rect 47465 34120 47545 34130
rect 47785 34120 47865 34130
rect 48105 34120 48185 34130
rect 44025 34040 44035 34120
rect 44345 34040 44355 34120
rect 44665 34040 44675 34120
rect 44985 34040 44995 34120
rect 45305 34040 45315 34120
rect 45625 34040 45635 34120
rect 45945 34040 45955 34120
rect 46265 34040 46275 34120
rect 46585 34040 46595 34120
rect 46905 34040 46915 34120
rect 47225 34040 47235 34120
rect 47545 34040 47555 34120
rect 47865 34040 47875 34120
rect 48185 34040 48195 34120
rect 42950 34020 42980 34030
rect 43220 34020 43300 34030
rect 42980 33940 42990 34020
rect 43300 33940 43310 34020
rect 48500 33970 48605 34140
rect 48640 34060 48650 34140
rect 48790 34060 48800 34140
rect 49350 34060 49360 34140
rect 49500 34060 49510 34140
rect 49560 33970 49590 34140
rect 49650 34060 49690 34140
rect 43785 33960 43865 33970
rect 44105 33960 44185 33970
rect 44425 33960 44505 33970
rect 44745 33960 44825 33970
rect 45065 33960 45145 33970
rect 45385 33960 45465 33970
rect 45705 33960 45785 33970
rect 46025 33960 46105 33970
rect 46345 33960 46425 33970
rect 46665 33960 46745 33970
rect 46985 33960 47065 33970
rect 47305 33960 47385 33970
rect 47625 33960 47705 33970
rect 47945 33960 48025 33970
rect 48265 33960 48345 33970
rect 48500 33960 48640 33970
rect 48710 33960 48790 33970
rect 49270 33960 49350 33970
rect 49420 33960 49500 33970
rect 49560 33960 49650 33970
rect 49660 33960 49690 34060
rect 43865 33880 43875 33960
rect 44185 33880 44195 33960
rect 44505 33880 44515 33960
rect 44825 33880 44835 33960
rect 45145 33880 45155 33960
rect 45465 33880 45475 33960
rect 45785 33880 45795 33960
rect 46105 33880 46115 33960
rect 46425 33880 46435 33960
rect 46745 33880 46755 33960
rect 47065 33880 47075 33960
rect 47385 33880 47395 33960
rect 47705 33880 47715 33960
rect 48025 33880 48035 33960
rect 48345 33880 48355 33960
rect 43060 33860 43140 33870
rect 43380 33860 43460 33870
rect 43140 33780 43150 33860
rect 43460 33780 43470 33860
rect 43945 33800 44025 33810
rect 44265 33800 44345 33810
rect 44585 33800 44665 33810
rect 44905 33800 44985 33810
rect 45225 33800 45305 33810
rect 45545 33800 45625 33810
rect 45865 33800 45945 33810
rect 46185 33800 46265 33810
rect 46505 33800 46585 33810
rect 46825 33800 46905 33810
rect 47145 33800 47225 33810
rect 47465 33800 47545 33810
rect 47785 33800 47865 33810
rect 48105 33800 48185 33810
rect 44025 33720 44035 33800
rect 44345 33720 44355 33800
rect 44665 33720 44675 33800
rect 44985 33720 44995 33800
rect 45305 33720 45315 33800
rect 45625 33720 45635 33800
rect 45945 33720 45955 33800
rect 46265 33720 46275 33800
rect 46585 33720 46595 33800
rect 46905 33720 46915 33800
rect 47225 33720 47235 33800
rect 47545 33720 47555 33800
rect 47865 33720 47875 33800
rect 48185 33720 48195 33800
rect 48500 33790 48605 33960
rect 48640 33880 48650 33960
rect 48790 33880 48800 33960
rect 49350 33880 49360 33960
rect 49500 33880 49510 33960
rect 49560 33790 49590 33960
rect 49650 33880 49690 33960
rect 48500 33780 48640 33790
rect 48710 33780 48790 33790
rect 49270 33780 49350 33790
rect 49420 33780 49500 33790
rect 49560 33780 49650 33790
rect 49660 33780 49690 33880
rect 42950 33700 42980 33710
rect 43220 33700 43300 33710
rect 42980 33620 42990 33700
rect 43300 33620 43310 33700
rect 43785 33640 43865 33650
rect 44105 33640 44185 33650
rect 44425 33640 44505 33650
rect 44745 33640 44825 33650
rect 45065 33640 45145 33650
rect 45385 33640 45465 33650
rect 45705 33640 45785 33650
rect 46025 33640 46105 33650
rect 46345 33640 46425 33650
rect 46665 33640 46745 33650
rect 46985 33640 47065 33650
rect 47305 33640 47385 33650
rect 47625 33640 47705 33650
rect 47945 33640 48025 33650
rect 48265 33640 48345 33650
rect 43865 33560 43875 33640
rect 44185 33560 44195 33640
rect 44505 33560 44515 33640
rect 44825 33560 44835 33640
rect 45145 33560 45155 33640
rect 45465 33560 45475 33640
rect 45785 33560 45795 33640
rect 46105 33560 46115 33640
rect 46425 33560 46435 33640
rect 46745 33560 46755 33640
rect 47065 33560 47075 33640
rect 47385 33560 47395 33640
rect 47705 33560 47715 33640
rect 48025 33560 48035 33640
rect 48345 33560 48355 33640
rect 48500 33610 48605 33780
rect 48640 33700 48650 33780
rect 48790 33700 48800 33780
rect 49350 33700 49360 33780
rect 49500 33700 49510 33780
rect 49560 33610 49590 33780
rect 49650 33700 49690 33780
rect 48500 33600 48640 33610
rect 48710 33600 48790 33610
rect 49270 33600 49350 33610
rect 49420 33600 49500 33610
rect 49560 33600 49650 33610
rect 49660 33600 49690 33700
rect 43060 33540 43140 33550
rect 43380 33540 43460 33550
rect 43140 33460 43150 33540
rect 43460 33460 43470 33540
rect 43945 33480 44025 33490
rect 44265 33480 44345 33490
rect 44585 33480 44665 33490
rect 44905 33480 44985 33490
rect 45225 33480 45305 33490
rect 45545 33480 45625 33490
rect 45865 33480 45945 33490
rect 46185 33480 46265 33490
rect 46505 33480 46585 33490
rect 46825 33480 46905 33490
rect 47145 33480 47225 33490
rect 47465 33480 47545 33490
rect 47785 33480 47865 33490
rect 48105 33480 48185 33490
rect 44025 33400 44035 33480
rect 44345 33400 44355 33480
rect 44665 33400 44675 33480
rect 44985 33400 44995 33480
rect 45305 33400 45315 33480
rect 45625 33400 45635 33480
rect 45945 33400 45955 33480
rect 46265 33400 46275 33480
rect 46585 33400 46595 33480
rect 46905 33400 46915 33480
rect 47225 33400 47235 33480
rect 47545 33400 47555 33480
rect 47865 33400 47875 33480
rect 48185 33400 48195 33480
rect 48500 33430 48605 33600
rect 48640 33520 48650 33600
rect 48790 33520 48800 33600
rect 49350 33520 49360 33600
rect 49500 33520 49510 33600
rect 49560 33430 49590 33600
rect 49650 33520 49690 33600
rect 48500 33420 48640 33430
rect 48710 33420 48790 33430
rect 49270 33420 49350 33430
rect 49420 33420 49500 33430
rect 49560 33420 49650 33430
rect 49660 33420 49690 33520
rect 42950 33380 42980 33390
rect 43220 33380 43300 33390
rect 42980 33300 42990 33380
rect 43300 33300 43310 33380
rect 43785 33320 43865 33330
rect 44105 33320 44185 33330
rect 44425 33320 44505 33330
rect 44745 33320 44825 33330
rect 45065 33320 45145 33330
rect 45385 33320 45465 33330
rect 45705 33320 45785 33330
rect 46025 33320 46105 33330
rect 46345 33320 46425 33330
rect 46665 33320 46745 33330
rect 46985 33320 47065 33330
rect 47305 33320 47385 33330
rect 47625 33320 47705 33330
rect 47945 33320 48025 33330
rect 48265 33320 48345 33330
rect 43865 33240 43875 33320
rect 44185 33240 44195 33320
rect 44505 33240 44515 33320
rect 44825 33240 44835 33320
rect 45145 33240 45155 33320
rect 45465 33240 45475 33320
rect 45785 33240 45795 33320
rect 46105 33240 46115 33320
rect 46425 33240 46435 33320
rect 46745 33240 46755 33320
rect 47065 33240 47075 33320
rect 47385 33240 47395 33320
rect 47705 33240 47715 33320
rect 48025 33240 48035 33320
rect 48345 33240 48355 33320
rect 48500 33250 48605 33420
rect 48640 33340 48650 33420
rect 48790 33340 48800 33420
rect 49350 33340 49360 33420
rect 49500 33340 49510 33420
rect 49560 33250 49590 33420
rect 49650 33340 49690 33420
rect 48500 33240 48640 33250
rect 48710 33240 48790 33250
rect 49270 33240 49350 33250
rect 49420 33240 49500 33250
rect 49560 33240 49650 33250
rect 49660 33240 49690 33340
rect 43060 33220 43140 33230
rect 43380 33220 43460 33230
rect 43140 33140 43150 33220
rect 43460 33140 43470 33220
rect 43945 33160 44025 33170
rect 44265 33160 44345 33170
rect 44585 33160 44665 33170
rect 44905 33160 44985 33170
rect 45225 33160 45305 33170
rect 45545 33160 45625 33170
rect 45865 33160 45945 33170
rect 46185 33160 46265 33170
rect 46505 33160 46585 33170
rect 46825 33160 46905 33170
rect 47145 33160 47225 33170
rect 47465 33160 47545 33170
rect 47785 33160 47865 33170
rect 48105 33160 48185 33170
rect 44025 33080 44035 33160
rect 44345 33080 44355 33160
rect 44665 33080 44675 33160
rect 44985 33080 44995 33160
rect 45305 33080 45315 33160
rect 45625 33080 45635 33160
rect 45945 33080 45955 33160
rect 46265 33080 46275 33160
rect 46585 33080 46595 33160
rect 46905 33080 46915 33160
rect 47225 33080 47235 33160
rect 47545 33080 47555 33160
rect 47865 33080 47875 33160
rect 48185 33080 48195 33160
rect 48500 33070 48605 33240
rect 48640 33160 48650 33240
rect 48790 33160 48800 33240
rect 49350 33160 49360 33240
rect 49500 33160 49510 33240
rect 49560 33070 49590 33240
rect 49650 33160 49690 33240
rect 42950 33060 42980 33070
rect 43220 33060 43300 33070
rect 48500 33060 48640 33070
rect 48710 33060 48790 33070
rect 49270 33060 49350 33070
rect 49420 33060 49500 33070
rect 49560 33060 49650 33070
rect 49660 33060 49690 33160
rect 42980 32980 42990 33060
rect 43300 32980 43310 33060
rect 43785 33000 43865 33010
rect 44105 33000 44185 33010
rect 44425 33000 44505 33010
rect 44745 33000 44825 33010
rect 45065 33000 45145 33010
rect 45385 33000 45465 33010
rect 45705 33000 45785 33010
rect 46025 33000 46105 33010
rect 46345 33000 46425 33010
rect 46665 33000 46745 33010
rect 46985 33000 47065 33010
rect 47305 33000 47385 33010
rect 47625 33000 47705 33010
rect 47945 33000 48025 33010
rect 48265 33000 48345 33010
rect 43865 32920 43875 33000
rect 44185 32920 44195 33000
rect 44505 32920 44515 33000
rect 44825 32920 44835 33000
rect 45145 32920 45155 33000
rect 45465 32920 45475 33000
rect 45785 32920 45795 33000
rect 46105 32920 46115 33000
rect 46425 32920 46435 33000
rect 46745 32920 46755 33000
rect 47065 32920 47075 33000
rect 47385 32920 47395 33000
rect 47705 32920 47715 33000
rect 48025 32920 48035 33000
rect 48345 32920 48355 33000
rect 43060 32900 43140 32910
rect 43380 32900 43460 32910
rect 43140 32820 43150 32900
rect 43460 32820 43470 32900
rect 48500 32890 48605 33060
rect 48640 32980 48650 33060
rect 48790 32980 48800 33060
rect 49350 32980 49360 33060
rect 49500 32980 49510 33060
rect 49560 32890 49590 33060
rect 49650 32980 49690 33060
rect 48500 32880 48640 32890
rect 48710 32880 48790 32890
rect 49270 32880 49350 32890
rect 49420 32880 49500 32890
rect 49560 32880 49650 32890
rect 49660 32880 49690 32980
rect 43945 32840 44025 32850
rect 44265 32840 44345 32850
rect 44585 32840 44665 32850
rect 44905 32840 44985 32850
rect 45225 32840 45305 32850
rect 45545 32840 45625 32850
rect 45865 32840 45945 32850
rect 46185 32840 46265 32850
rect 46505 32840 46585 32850
rect 46825 32840 46905 32850
rect 47145 32840 47225 32850
rect 47465 32840 47545 32850
rect 47785 32840 47865 32850
rect 48105 32840 48185 32850
rect 44025 32760 44035 32840
rect 44345 32760 44355 32840
rect 44665 32760 44675 32840
rect 44985 32760 44995 32840
rect 45305 32760 45315 32840
rect 45625 32760 45635 32840
rect 45945 32760 45955 32840
rect 46265 32760 46275 32840
rect 46585 32760 46595 32840
rect 46905 32760 46915 32840
rect 47225 32760 47235 32840
rect 47545 32760 47555 32840
rect 47865 32760 47875 32840
rect 48185 32760 48195 32840
rect 42950 32740 42980 32750
rect 43220 32740 43300 32750
rect 42980 32660 42990 32740
rect 43300 32660 43310 32740
rect 48500 32710 48605 32880
rect 48640 32800 48650 32880
rect 48790 32800 48800 32880
rect 49350 32800 49360 32880
rect 49500 32800 49510 32880
rect 49560 32710 49590 32880
rect 49650 32800 49690 32880
rect 48500 32700 48640 32710
rect 48710 32700 48790 32710
rect 49270 32700 49350 32710
rect 49420 32700 49500 32710
rect 49560 32700 49650 32710
rect 49660 32700 49690 32800
rect 43785 32680 43865 32690
rect 44105 32680 44185 32690
rect 44425 32680 44505 32690
rect 44745 32680 44825 32690
rect 45065 32680 45145 32690
rect 45385 32680 45465 32690
rect 45705 32680 45785 32690
rect 46025 32680 46105 32690
rect 46345 32680 46425 32690
rect 46665 32680 46745 32690
rect 46985 32680 47065 32690
rect 47305 32680 47385 32690
rect 47625 32680 47705 32690
rect 47945 32680 48025 32690
rect 48265 32680 48345 32690
rect 43865 32600 43875 32680
rect 44185 32600 44195 32680
rect 44505 32600 44515 32680
rect 44825 32600 44835 32680
rect 45145 32600 45155 32680
rect 45465 32600 45475 32680
rect 45785 32600 45795 32680
rect 46105 32600 46115 32680
rect 46425 32600 46435 32680
rect 46745 32600 46755 32680
rect 47065 32600 47075 32680
rect 47385 32600 47395 32680
rect 47705 32600 47715 32680
rect 48025 32600 48035 32680
rect 48345 32600 48355 32680
rect 43060 32580 43140 32590
rect 43380 32580 43460 32590
rect 43140 32500 43150 32580
rect 43460 32500 43470 32580
rect 48500 32530 48605 32700
rect 48640 32620 48650 32700
rect 48790 32620 48800 32700
rect 49350 32620 49360 32700
rect 49500 32620 49510 32700
rect 49560 32530 49590 32700
rect 49650 32620 49690 32700
rect 43945 32520 44025 32530
rect 44265 32520 44345 32530
rect 44585 32520 44665 32530
rect 44905 32520 44985 32530
rect 45225 32520 45305 32530
rect 45545 32520 45625 32530
rect 45865 32520 45945 32530
rect 46185 32520 46265 32530
rect 46505 32520 46585 32530
rect 46825 32520 46905 32530
rect 47145 32520 47225 32530
rect 47465 32520 47545 32530
rect 47785 32520 47865 32530
rect 48105 32520 48185 32530
rect 48500 32520 48640 32530
rect 48710 32520 48790 32530
rect 49270 32520 49350 32530
rect 49420 32520 49500 32530
rect 49560 32520 49650 32530
rect 49660 32520 49690 32620
rect 44025 32440 44035 32520
rect 44345 32440 44355 32520
rect 44665 32440 44675 32520
rect 44985 32440 44995 32520
rect 45305 32440 45315 32520
rect 45625 32440 45635 32520
rect 45945 32440 45955 32520
rect 46265 32440 46275 32520
rect 46585 32440 46595 32520
rect 46905 32440 46915 32520
rect 47225 32440 47235 32520
rect 47545 32440 47555 32520
rect 47865 32440 47875 32520
rect 48185 32440 48195 32520
rect 42950 32420 42980 32430
rect 43220 32420 43300 32430
rect 42980 32340 42990 32420
rect 43300 32340 43310 32420
rect 43785 32360 43865 32370
rect 44105 32360 44185 32370
rect 44425 32360 44505 32370
rect 44745 32360 44825 32370
rect 45065 32360 45145 32370
rect 45385 32360 45465 32370
rect 45705 32360 45785 32370
rect 46025 32360 46105 32370
rect 46345 32360 46425 32370
rect 46665 32360 46745 32370
rect 46985 32360 47065 32370
rect 47305 32360 47385 32370
rect 47625 32360 47705 32370
rect 47945 32360 48025 32370
rect 48265 32360 48345 32370
rect 43865 32280 43875 32360
rect 44185 32280 44195 32360
rect 44505 32280 44515 32360
rect 44825 32280 44835 32360
rect 45145 32280 45155 32360
rect 45465 32280 45475 32360
rect 45785 32280 45795 32360
rect 46105 32280 46115 32360
rect 46425 32280 46435 32360
rect 46745 32280 46755 32360
rect 47065 32280 47075 32360
rect 47385 32280 47395 32360
rect 47705 32280 47715 32360
rect 48025 32280 48035 32360
rect 48345 32280 48355 32360
rect 48500 32350 48605 32520
rect 48640 32440 48650 32520
rect 48790 32440 48800 32520
rect 49350 32440 49360 32520
rect 49500 32440 49510 32520
rect 49560 32350 49590 32520
rect 49650 32440 49690 32520
rect 48500 32340 48640 32350
rect 48710 32340 48790 32350
rect 49270 32340 49350 32350
rect 49420 32340 49500 32350
rect 49560 32340 49650 32350
rect 49660 32340 49690 32440
rect 43060 32260 43140 32270
rect 43380 32260 43460 32270
rect 43140 32180 43150 32260
rect 43460 32180 43470 32260
rect 43945 32200 44025 32210
rect 44265 32200 44345 32210
rect 44585 32200 44665 32210
rect 44905 32200 44985 32210
rect 45225 32200 45305 32210
rect 45545 32200 45625 32210
rect 45865 32200 45945 32210
rect 46185 32200 46265 32210
rect 46505 32200 46585 32210
rect 46825 32200 46905 32210
rect 47145 32200 47225 32210
rect 47465 32200 47545 32210
rect 47785 32200 47865 32210
rect 48105 32200 48185 32210
rect 44025 32120 44035 32200
rect 44345 32120 44355 32200
rect 44665 32120 44675 32200
rect 44985 32120 44995 32200
rect 45305 32120 45315 32200
rect 45625 32120 45635 32200
rect 45945 32120 45955 32200
rect 46265 32120 46275 32200
rect 46585 32120 46595 32200
rect 46905 32120 46915 32200
rect 47225 32120 47235 32200
rect 47545 32120 47555 32200
rect 47865 32120 47875 32200
rect 48185 32120 48195 32200
rect 48500 32170 48605 32340
rect 48640 32260 48650 32340
rect 48790 32260 48800 32340
rect 49350 32260 49360 32340
rect 49500 32260 49510 32340
rect 49560 32170 49590 32340
rect 49650 32260 49690 32340
rect 48500 32160 48640 32170
rect 48710 32160 48790 32170
rect 49270 32160 49350 32170
rect 49420 32160 49500 32170
rect 49560 32160 49650 32170
rect 49660 32160 49690 32260
rect 42950 32100 42980 32110
rect 43220 32100 43300 32110
rect 42980 32020 42990 32100
rect 43300 32020 43310 32100
rect 43785 32040 43865 32050
rect 44105 32040 44185 32050
rect 44425 32040 44505 32050
rect 44745 32040 44825 32050
rect 45065 32040 45145 32050
rect 45385 32040 45465 32050
rect 45705 32040 45785 32050
rect 46025 32040 46105 32050
rect 46345 32040 46425 32050
rect 46665 32040 46745 32050
rect 46985 32040 47065 32050
rect 47305 32040 47385 32050
rect 47625 32040 47705 32050
rect 47945 32040 48025 32050
rect 48265 32040 48345 32050
rect 43865 31960 43875 32040
rect 44185 31960 44195 32040
rect 44505 31960 44515 32040
rect 44825 31960 44835 32040
rect 45145 31960 45155 32040
rect 45465 31960 45475 32040
rect 45785 31960 45795 32040
rect 46105 31960 46115 32040
rect 46425 31960 46435 32040
rect 46745 31960 46755 32040
rect 47065 31960 47075 32040
rect 47385 31960 47395 32040
rect 47705 31960 47715 32040
rect 48025 31960 48035 32040
rect 48345 31960 48355 32040
rect 48500 31990 48605 32160
rect 48640 32080 48650 32160
rect 48790 32080 48800 32160
rect 49350 32080 49360 32160
rect 49500 32080 49510 32160
rect 49560 31990 49590 32160
rect 49650 32080 49690 32160
rect 48500 31980 48640 31990
rect 48710 31980 48790 31990
rect 49270 31980 49350 31990
rect 49420 31980 49500 31990
rect 49560 31980 49650 31990
rect 49660 31980 49690 32080
rect 43060 31940 43140 31950
rect 43380 31940 43460 31950
rect 43140 31860 43150 31940
rect 43460 31860 43470 31940
rect 43945 31880 44025 31890
rect 44265 31880 44345 31890
rect 44585 31880 44665 31890
rect 44905 31880 44985 31890
rect 45225 31880 45305 31890
rect 45545 31880 45625 31890
rect 45865 31880 45945 31890
rect 46185 31880 46265 31890
rect 46505 31880 46585 31890
rect 46825 31880 46905 31890
rect 47145 31880 47225 31890
rect 47465 31880 47545 31890
rect 47785 31880 47865 31890
rect 48105 31880 48185 31890
rect 44025 31800 44035 31880
rect 44345 31800 44355 31880
rect 44665 31800 44675 31880
rect 44985 31800 44995 31880
rect 45305 31800 45315 31880
rect 45625 31800 45635 31880
rect 45945 31800 45955 31880
rect 46265 31800 46275 31880
rect 46585 31800 46595 31880
rect 46905 31800 46915 31880
rect 47225 31800 47235 31880
rect 47545 31800 47555 31880
rect 47865 31800 47875 31880
rect 48185 31800 48195 31880
rect 48500 31810 48605 31980
rect 48640 31900 48650 31980
rect 48790 31900 48800 31980
rect 49350 31900 49360 31980
rect 49500 31900 49510 31980
rect 49560 31810 49590 31980
rect 49650 31900 49690 31980
rect 48500 31800 48640 31810
rect 48710 31800 48790 31810
rect 49270 31800 49350 31810
rect 49420 31800 49500 31810
rect 49560 31800 49650 31810
rect 49660 31800 49690 31900
rect 42950 31780 42980 31790
rect 43220 31780 43300 31790
rect 42980 31700 42990 31780
rect 43300 31700 43310 31780
rect 43785 31720 43865 31730
rect 44105 31720 44185 31730
rect 44425 31720 44505 31730
rect 44745 31720 44825 31730
rect 45065 31720 45145 31730
rect 45385 31720 45465 31730
rect 45705 31720 45785 31730
rect 46025 31720 46105 31730
rect 46345 31720 46425 31730
rect 46665 31720 46745 31730
rect 46985 31720 47065 31730
rect 47305 31720 47385 31730
rect 47625 31720 47705 31730
rect 47945 31720 48025 31730
rect 48265 31720 48345 31730
rect 43865 31640 43875 31720
rect 44185 31640 44195 31720
rect 44505 31640 44515 31720
rect 44825 31640 44835 31720
rect 45145 31640 45155 31720
rect 45465 31640 45475 31720
rect 45785 31640 45795 31720
rect 46105 31640 46115 31720
rect 46425 31640 46435 31720
rect 46745 31640 46755 31720
rect 47065 31640 47075 31720
rect 47385 31640 47395 31720
rect 47705 31640 47715 31720
rect 48025 31640 48035 31720
rect 48345 31640 48355 31720
rect 48500 31630 48605 31800
rect 48640 31720 48650 31800
rect 48790 31720 48800 31800
rect 49350 31720 49360 31800
rect 49500 31720 49510 31800
rect 49560 31630 49590 31800
rect 49650 31720 49690 31800
rect 43060 31620 43140 31630
rect 43380 31620 43460 31630
rect 48500 31620 48640 31630
rect 48710 31620 48790 31630
rect 49270 31620 49350 31630
rect 49420 31620 49500 31630
rect 49560 31620 49650 31630
rect 49660 31620 49690 31720
rect 43140 31540 43150 31620
rect 43460 31540 43470 31620
rect 43945 31560 44025 31570
rect 44265 31560 44345 31570
rect 44585 31560 44665 31570
rect 44905 31560 44985 31570
rect 45225 31560 45305 31570
rect 45545 31560 45625 31570
rect 45865 31560 45945 31570
rect 46185 31560 46265 31570
rect 46505 31560 46585 31570
rect 46825 31560 46905 31570
rect 47145 31560 47225 31570
rect 47465 31560 47545 31570
rect 47785 31560 47865 31570
rect 48105 31560 48185 31570
rect 44025 31480 44035 31560
rect 44345 31480 44355 31560
rect 44665 31480 44675 31560
rect 44985 31480 44995 31560
rect 45305 31480 45315 31560
rect 45625 31480 45635 31560
rect 45945 31480 45955 31560
rect 46265 31480 46275 31560
rect 46585 31480 46595 31560
rect 46905 31480 46915 31560
rect 47225 31480 47235 31560
rect 47545 31480 47555 31560
rect 47865 31480 47875 31560
rect 48185 31480 48195 31560
rect 42950 31460 42980 31470
rect 43220 31460 43300 31470
rect 42980 31380 42990 31460
rect 43300 31380 43310 31460
rect 48500 31450 48605 31620
rect 48640 31540 48650 31620
rect 48790 31540 48800 31620
rect 49350 31540 49360 31620
rect 49500 31540 49510 31620
rect 49560 31450 49590 31620
rect 49650 31540 49690 31620
rect 48500 31440 48640 31450
rect 48710 31440 48790 31450
rect 49270 31440 49350 31450
rect 49420 31440 49500 31450
rect 49560 31440 49650 31450
rect 49660 31440 49690 31540
rect 43785 31400 43865 31410
rect 44105 31400 44185 31410
rect 44425 31400 44505 31410
rect 44745 31400 44825 31410
rect 45065 31400 45145 31410
rect 45385 31400 45465 31410
rect 45705 31400 45785 31410
rect 46025 31400 46105 31410
rect 46345 31400 46425 31410
rect 46665 31400 46745 31410
rect 46985 31400 47065 31410
rect 47305 31400 47385 31410
rect 47625 31400 47705 31410
rect 47945 31400 48025 31410
rect 48265 31400 48345 31410
rect 43865 31320 43875 31400
rect 44185 31320 44195 31400
rect 44505 31320 44515 31400
rect 44825 31320 44835 31400
rect 45145 31320 45155 31400
rect 45465 31320 45475 31400
rect 45785 31320 45795 31400
rect 46105 31320 46115 31400
rect 46425 31320 46435 31400
rect 46745 31320 46755 31400
rect 47065 31320 47075 31400
rect 47385 31320 47395 31400
rect 47705 31320 47715 31400
rect 48025 31320 48035 31400
rect 48345 31320 48355 31400
rect 43060 31300 43140 31310
rect 43380 31300 43460 31310
rect 43140 31220 43150 31300
rect 43460 31220 43470 31300
rect 48500 31270 48605 31440
rect 48640 31360 48650 31440
rect 48790 31360 48800 31440
rect 49350 31360 49360 31440
rect 49500 31360 49510 31440
rect 49560 31270 49590 31440
rect 49650 31360 49690 31440
rect 48500 31260 48640 31270
rect 48710 31260 48790 31270
rect 49270 31260 49350 31270
rect 49420 31260 49500 31270
rect 49560 31260 49650 31270
rect 49660 31260 49690 31360
rect 43945 31240 44025 31250
rect 44265 31240 44345 31250
rect 44585 31240 44665 31250
rect 44905 31240 44985 31250
rect 45225 31240 45305 31250
rect 45545 31240 45625 31250
rect 45865 31240 45945 31250
rect 46185 31240 46265 31250
rect 46505 31240 46585 31250
rect 46825 31240 46905 31250
rect 47145 31240 47225 31250
rect 47465 31240 47545 31250
rect 47785 31240 47865 31250
rect 48105 31240 48185 31250
rect 44025 31160 44035 31240
rect 44345 31160 44355 31240
rect 44665 31160 44675 31240
rect 44985 31160 44995 31240
rect 45305 31160 45315 31240
rect 45625 31160 45635 31240
rect 45945 31160 45955 31240
rect 46265 31160 46275 31240
rect 46585 31160 46595 31240
rect 46905 31160 46915 31240
rect 47225 31160 47235 31240
rect 47545 31160 47555 31240
rect 47865 31160 47875 31240
rect 48185 31160 48195 31240
rect 42950 31140 42980 31150
rect 43220 31140 43300 31150
rect 42980 31060 42990 31140
rect 43300 31060 43310 31140
rect 48500 31090 48605 31260
rect 48640 31180 48650 31260
rect 48790 31180 48800 31260
rect 49350 31180 49360 31260
rect 49500 31180 49510 31260
rect 49560 31100 49590 31260
rect 49650 31180 49690 31260
rect 49660 31100 49690 31180
rect 49790 31100 49800 37100
rect 49890 37020 49970 37030
rect 50210 37020 50290 37030
rect 49970 36940 49980 37020
rect 50290 36940 50300 37020
rect 49890 36840 49970 36850
rect 50210 36840 50290 36850
rect 49970 36760 49980 36840
rect 50290 36760 50300 36840
rect 49890 36660 49970 36670
rect 50210 36660 50290 36670
rect 49970 36580 49980 36660
rect 50290 36580 50300 36660
rect 49890 36480 49970 36490
rect 50210 36480 50290 36490
rect 49970 36400 49980 36480
rect 50290 36400 50300 36480
rect 49890 36300 49970 36310
rect 50210 36300 50290 36310
rect 49970 36220 49980 36300
rect 50290 36220 50300 36300
rect 49890 36120 49970 36130
rect 50210 36120 50290 36130
rect 49970 36040 49980 36120
rect 50290 36040 50300 36120
rect 49890 35940 49970 35950
rect 50210 35940 50290 35950
rect 49970 35860 49980 35940
rect 50290 35860 50300 35940
rect 49890 35760 49970 35770
rect 50210 35760 50290 35770
rect 49970 35680 49980 35760
rect 50290 35680 50300 35760
rect 49890 35580 49970 35590
rect 50210 35580 50290 35590
rect 49970 35500 49980 35580
rect 50290 35500 50300 35580
rect 49890 35400 49970 35410
rect 50210 35400 50290 35410
rect 49970 35320 49980 35400
rect 50290 35320 50300 35400
rect 49890 35220 49970 35230
rect 50210 35220 50290 35230
rect 49970 35140 49980 35220
rect 50290 35140 50300 35220
rect 49890 35040 49970 35050
rect 50210 35040 50290 35050
rect 49970 34960 49980 35040
rect 50290 34960 50300 35040
rect 49890 34860 49970 34870
rect 50210 34860 50290 34870
rect 49970 34780 49980 34860
rect 50290 34780 50300 34860
rect 49890 34680 49970 34690
rect 50210 34680 50290 34690
rect 49970 34600 49980 34680
rect 50290 34600 50300 34680
rect 49890 34500 49970 34510
rect 50210 34500 50290 34510
rect 49970 34420 49980 34500
rect 50290 34420 50300 34500
rect 49890 34320 49970 34330
rect 50210 34320 50290 34330
rect 49970 34240 49980 34320
rect 50290 34240 50300 34320
rect 49890 34140 49970 34150
rect 50210 34140 50290 34150
rect 49970 34060 49980 34140
rect 50290 34060 50300 34140
rect 49890 33960 49970 33970
rect 50210 33960 50290 33970
rect 49970 33880 49980 33960
rect 50290 33880 50300 33960
rect 49890 33780 49970 33790
rect 50210 33780 50290 33790
rect 49970 33700 49980 33780
rect 50290 33700 50300 33780
rect 49890 33600 49970 33610
rect 50210 33600 50290 33610
rect 49970 33520 49980 33600
rect 50290 33520 50300 33600
rect 49890 33420 49970 33430
rect 50210 33420 50290 33430
rect 49970 33340 49980 33420
rect 50290 33340 50300 33420
rect 49890 33240 49970 33250
rect 50210 33240 50290 33250
rect 49970 33160 49980 33240
rect 50290 33160 50300 33240
rect 49890 33060 49970 33070
rect 50210 33060 50290 33070
rect 49970 32980 49980 33060
rect 50290 32980 50300 33060
rect 49890 32880 49970 32890
rect 50210 32880 50290 32890
rect 49970 32800 49980 32880
rect 50290 32800 50300 32880
rect 49890 32700 49970 32710
rect 50210 32700 50290 32710
rect 49970 32620 49980 32700
rect 50290 32620 50300 32700
rect 49890 32520 49970 32530
rect 50210 32520 50290 32530
rect 49970 32440 49980 32520
rect 50290 32440 50300 32520
rect 49890 32340 49970 32350
rect 50210 32340 50290 32350
rect 49970 32260 49980 32340
rect 50290 32260 50300 32340
rect 49890 32160 49970 32170
rect 50210 32160 50290 32170
rect 49970 32080 49980 32160
rect 50290 32080 50300 32160
rect 49890 31980 49970 31990
rect 50210 31980 50290 31990
rect 49970 31900 49980 31980
rect 50290 31900 50300 31980
rect 49890 31800 49970 31810
rect 50210 31800 50290 31810
rect 49970 31720 49980 31800
rect 50290 31720 50300 31800
rect 49890 31620 49970 31630
rect 50210 31620 50290 31630
rect 49970 31540 49980 31620
rect 50290 31540 50300 31620
rect 49890 31440 49970 31450
rect 50210 31440 50290 31450
rect 49970 31360 49980 31440
rect 50290 31360 50300 31440
rect 49890 31260 49970 31270
rect 50210 31260 50290 31270
rect 49970 31180 49980 31260
rect 50290 31180 50300 31260
rect 50470 31100 50480 37100
rect 50490 31100 50520 37100
rect 50590 37030 50620 37100
rect 50820 37030 50850 37100
rect 50530 37020 50620 37030
rect 50680 37020 50760 37030
rect 50820 37020 50910 37030
rect 50920 37020 50950 37100
rect 50590 36850 50620 37020
rect 50760 36940 50770 37020
rect 50820 36850 50850 37020
rect 50910 36940 50950 37020
rect 50530 36840 50620 36850
rect 50680 36840 50760 36850
rect 50820 36840 50910 36850
rect 50920 36840 50950 36940
rect 50590 36670 50620 36840
rect 50760 36760 50770 36840
rect 50820 36670 50850 36840
rect 50910 36760 50950 36840
rect 50530 36660 50620 36670
rect 50680 36660 50760 36670
rect 50820 36660 50910 36670
rect 50920 36660 50950 36760
rect 50590 36490 50620 36660
rect 50760 36580 50770 36660
rect 50820 36490 50850 36660
rect 50910 36580 50950 36660
rect 50530 36480 50620 36490
rect 50680 36480 50760 36490
rect 50820 36480 50910 36490
rect 50920 36480 50950 36580
rect 50590 36310 50620 36480
rect 50760 36400 50770 36480
rect 50820 36310 50850 36480
rect 50910 36400 50950 36480
rect 50530 36300 50620 36310
rect 50680 36300 50760 36310
rect 50820 36300 50910 36310
rect 50920 36300 50950 36400
rect 50590 36130 50620 36300
rect 50760 36220 50770 36300
rect 50820 36130 50850 36300
rect 50910 36220 50950 36300
rect 50530 36120 50620 36130
rect 50680 36120 50760 36130
rect 50820 36120 50910 36130
rect 50920 36120 50950 36220
rect 50590 35950 50620 36120
rect 50760 36040 50770 36120
rect 50820 35950 50850 36120
rect 50910 36040 50950 36120
rect 50530 35940 50620 35950
rect 50680 35940 50760 35950
rect 50820 35940 50910 35950
rect 50920 35940 50950 36040
rect 50590 35770 50620 35940
rect 50760 35860 50770 35940
rect 50820 35770 50850 35940
rect 50910 35860 50950 35940
rect 50530 35760 50620 35770
rect 50680 35760 50760 35770
rect 50820 35760 50910 35770
rect 50920 35760 50950 35860
rect 50590 35590 50620 35760
rect 50760 35680 50770 35760
rect 50820 35590 50850 35760
rect 50910 35680 50950 35760
rect 50530 35580 50620 35590
rect 50680 35580 50760 35590
rect 50820 35580 50910 35590
rect 50920 35580 50950 35680
rect 50590 35410 50620 35580
rect 50760 35500 50770 35580
rect 50820 35410 50850 35580
rect 50910 35500 50950 35580
rect 50530 35400 50620 35410
rect 50680 35400 50760 35410
rect 50820 35400 50910 35410
rect 50920 35400 50950 35500
rect 50590 35230 50620 35400
rect 50760 35320 50770 35400
rect 50820 35230 50850 35400
rect 50910 35320 50950 35400
rect 50530 35220 50620 35230
rect 50680 35220 50760 35230
rect 50820 35220 50910 35230
rect 50920 35220 50950 35320
rect 50590 35050 50620 35220
rect 50760 35140 50770 35220
rect 50820 35050 50850 35220
rect 50910 35140 50950 35220
rect 50530 35040 50620 35050
rect 50680 35040 50760 35050
rect 50820 35040 50910 35050
rect 50920 35040 50950 35140
rect 50590 34870 50620 35040
rect 50760 34960 50770 35040
rect 50820 34870 50850 35040
rect 50910 34960 50950 35040
rect 50530 34860 50620 34870
rect 50680 34860 50760 34870
rect 50820 34860 50910 34870
rect 50920 34860 50950 34960
rect 50590 34690 50620 34860
rect 50760 34780 50770 34860
rect 50820 34690 50850 34860
rect 50910 34780 50950 34860
rect 50530 34680 50620 34690
rect 50680 34680 50760 34690
rect 50820 34680 50910 34690
rect 50920 34680 50950 34780
rect 50590 34510 50620 34680
rect 50760 34600 50770 34680
rect 50820 34510 50850 34680
rect 50910 34600 50950 34680
rect 50530 34500 50620 34510
rect 50680 34500 50760 34510
rect 50820 34500 50910 34510
rect 50920 34500 50950 34600
rect 50590 34330 50620 34500
rect 50760 34420 50770 34500
rect 50820 34330 50850 34500
rect 50910 34420 50950 34500
rect 50530 34320 50620 34330
rect 50680 34320 50760 34330
rect 50820 34320 50910 34330
rect 50920 34320 50950 34420
rect 50590 34150 50620 34320
rect 50760 34240 50770 34320
rect 50820 34150 50850 34320
rect 50910 34240 50950 34320
rect 50530 34140 50620 34150
rect 50680 34140 50760 34150
rect 50820 34140 50910 34150
rect 50920 34140 50950 34240
rect 50590 33970 50620 34140
rect 50760 34060 50770 34140
rect 50820 33970 50850 34140
rect 50910 34060 50950 34140
rect 50530 33960 50620 33970
rect 50680 33960 50760 33970
rect 50820 33960 50910 33970
rect 50920 33960 50950 34060
rect 50590 33790 50620 33960
rect 50760 33880 50770 33960
rect 50820 33790 50850 33960
rect 50910 33880 50950 33960
rect 50530 33780 50620 33790
rect 50680 33780 50760 33790
rect 50820 33780 50910 33790
rect 50920 33780 50950 33880
rect 50590 33610 50620 33780
rect 50760 33700 50770 33780
rect 50820 33610 50850 33780
rect 50910 33700 50950 33780
rect 50530 33600 50620 33610
rect 50680 33600 50760 33610
rect 50820 33600 50910 33610
rect 50920 33600 50950 33700
rect 50590 33430 50620 33600
rect 50760 33520 50770 33600
rect 50820 33430 50850 33600
rect 50910 33520 50950 33600
rect 50530 33420 50620 33430
rect 50680 33420 50760 33430
rect 50820 33420 50910 33430
rect 50920 33420 50950 33520
rect 50590 33250 50620 33420
rect 50760 33340 50770 33420
rect 50820 33250 50850 33420
rect 50910 33340 50950 33420
rect 50530 33240 50620 33250
rect 50680 33240 50760 33250
rect 50820 33240 50910 33250
rect 50920 33240 50950 33340
rect 50590 33070 50620 33240
rect 50760 33160 50770 33240
rect 50820 33070 50850 33240
rect 50910 33160 50950 33240
rect 50530 33060 50620 33070
rect 50680 33060 50760 33070
rect 50820 33060 50910 33070
rect 50920 33060 50950 33160
rect 50590 32890 50620 33060
rect 50760 32980 50770 33060
rect 50820 32890 50850 33060
rect 50910 32980 50950 33060
rect 50530 32880 50620 32890
rect 50680 32880 50760 32890
rect 50820 32880 50910 32890
rect 50920 32880 50950 32980
rect 50590 32710 50620 32880
rect 50760 32800 50770 32880
rect 50820 32710 50850 32880
rect 50910 32800 50950 32880
rect 50530 32700 50620 32710
rect 50680 32700 50760 32710
rect 50820 32700 50910 32710
rect 50920 32700 50950 32800
rect 50590 32530 50620 32700
rect 50760 32620 50770 32700
rect 50820 32530 50850 32700
rect 50910 32620 50950 32700
rect 50530 32520 50620 32530
rect 50680 32520 50760 32530
rect 50820 32520 50910 32530
rect 50920 32520 50950 32620
rect 50590 32350 50620 32520
rect 50760 32440 50770 32520
rect 50820 32350 50850 32520
rect 50910 32440 50950 32520
rect 50530 32340 50620 32350
rect 50680 32340 50760 32350
rect 50820 32340 50910 32350
rect 50920 32340 50950 32440
rect 50590 32170 50620 32340
rect 50760 32260 50770 32340
rect 50820 32170 50850 32340
rect 50910 32260 50950 32340
rect 50530 32160 50620 32170
rect 50680 32160 50760 32170
rect 50820 32160 50910 32170
rect 50920 32160 50950 32260
rect 50590 31990 50620 32160
rect 50760 32080 50770 32160
rect 50820 31990 50850 32160
rect 50910 32080 50950 32160
rect 50530 31980 50620 31990
rect 50680 31980 50760 31990
rect 50820 31980 50910 31990
rect 50920 31980 50950 32080
rect 50590 31810 50620 31980
rect 50760 31900 50770 31980
rect 50820 31810 50850 31980
rect 50910 31900 50950 31980
rect 50530 31800 50620 31810
rect 50680 31800 50760 31810
rect 50820 31800 50910 31810
rect 50920 31800 50950 31900
rect 50590 31630 50620 31800
rect 50760 31720 50770 31800
rect 50820 31630 50850 31800
rect 50910 31720 50950 31800
rect 50530 31620 50620 31630
rect 50680 31620 50760 31630
rect 50820 31620 50910 31630
rect 50920 31620 50950 31720
rect 50590 31450 50620 31620
rect 50760 31540 50770 31620
rect 50820 31450 50850 31620
rect 50910 31540 50950 31620
rect 50530 31440 50620 31450
rect 50680 31440 50760 31450
rect 50820 31440 50910 31450
rect 50920 31440 50950 31540
rect 50590 31270 50620 31440
rect 50760 31360 50770 31440
rect 50820 31270 50850 31440
rect 50910 31360 50950 31440
rect 50530 31260 50620 31270
rect 50680 31260 50760 31270
rect 50820 31260 50910 31270
rect 50920 31260 50950 31360
rect 50590 31100 50620 31260
rect 50760 31180 50770 31260
rect 50820 31100 50850 31260
rect 50910 31180 50950 31260
rect 50920 31100 50950 31180
rect 51050 31100 51060 37100
rect 51150 37020 51230 37030
rect 51470 37020 51550 37030
rect 51230 36940 51240 37020
rect 51550 36940 51560 37020
rect 51150 36840 51230 36850
rect 51470 36840 51550 36850
rect 51230 36760 51240 36840
rect 51550 36760 51560 36840
rect 51150 36660 51230 36670
rect 51470 36660 51550 36670
rect 51230 36580 51240 36660
rect 51550 36580 51560 36660
rect 51150 36480 51230 36490
rect 51470 36480 51550 36490
rect 51230 36400 51240 36480
rect 51550 36400 51560 36480
rect 51150 36300 51230 36310
rect 51470 36300 51550 36310
rect 51230 36220 51240 36300
rect 51550 36220 51560 36300
rect 51150 36120 51230 36130
rect 51470 36120 51550 36130
rect 51230 36040 51240 36120
rect 51550 36040 51560 36120
rect 51150 35940 51230 35950
rect 51470 35940 51550 35950
rect 51230 35860 51240 35940
rect 51550 35860 51560 35940
rect 51150 35760 51230 35770
rect 51470 35760 51550 35770
rect 51230 35680 51240 35760
rect 51550 35680 51560 35760
rect 51150 35580 51230 35590
rect 51470 35580 51550 35590
rect 51230 35500 51240 35580
rect 51550 35500 51560 35580
rect 51150 35400 51230 35410
rect 51470 35400 51550 35410
rect 51230 35320 51240 35400
rect 51550 35320 51560 35400
rect 51150 35220 51230 35230
rect 51470 35220 51550 35230
rect 51230 35140 51240 35220
rect 51550 35140 51560 35220
rect 51150 35040 51230 35050
rect 51470 35040 51550 35050
rect 51230 34960 51240 35040
rect 51550 34960 51560 35040
rect 51150 34860 51230 34870
rect 51470 34860 51550 34870
rect 51230 34780 51240 34860
rect 51550 34780 51560 34860
rect 51150 34680 51230 34690
rect 51470 34680 51550 34690
rect 51230 34600 51240 34680
rect 51550 34600 51560 34680
rect 51150 34500 51230 34510
rect 51470 34500 51550 34510
rect 51230 34420 51240 34500
rect 51550 34420 51560 34500
rect 51150 34320 51230 34330
rect 51470 34320 51550 34330
rect 51230 34240 51240 34320
rect 51550 34240 51560 34320
rect 51150 34140 51230 34150
rect 51470 34140 51550 34150
rect 51230 34060 51240 34140
rect 51550 34060 51560 34140
rect 51150 33960 51230 33970
rect 51470 33960 51550 33970
rect 51230 33880 51240 33960
rect 51550 33880 51560 33960
rect 51150 33780 51230 33790
rect 51470 33780 51550 33790
rect 51230 33700 51240 33780
rect 51550 33700 51560 33780
rect 51150 33600 51230 33610
rect 51470 33600 51550 33610
rect 51230 33520 51240 33600
rect 51550 33520 51560 33600
rect 51150 33420 51230 33430
rect 51470 33420 51550 33430
rect 51230 33340 51240 33420
rect 51550 33340 51560 33420
rect 51150 33240 51230 33250
rect 51470 33240 51550 33250
rect 51230 33160 51240 33240
rect 51550 33160 51560 33240
rect 51150 33060 51230 33070
rect 51470 33060 51550 33070
rect 51230 32980 51240 33060
rect 51550 32980 51560 33060
rect 51150 32880 51230 32890
rect 51470 32880 51550 32890
rect 51230 32800 51240 32880
rect 51550 32800 51560 32880
rect 51150 32700 51230 32710
rect 51470 32700 51550 32710
rect 51230 32620 51240 32700
rect 51550 32620 51560 32700
rect 51150 32520 51230 32530
rect 51470 32520 51550 32530
rect 51230 32440 51240 32520
rect 51550 32440 51560 32520
rect 51150 32340 51230 32350
rect 51470 32340 51550 32350
rect 51230 32260 51240 32340
rect 51550 32260 51560 32340
rect 51150 32160 51230 32170
rect 51470 32160 51550 32170
rect 51230 32080 51240 32160
rect 51550 32080 51560 32160
rect 51150 31980 51230 31990
rect 51470 31980 51550 31990
rect 51230 31900 51240 31980
rect 51550 31900 51560 31980
rect 51150 31800 51230 31810
rect 51470 31800 51550 31810
rect 51230 31720 51240 31800
rect 51550 31720 51560 31800
rect 51150 31620 51230 31630
rect 51470 31620 51550 31630
rect 51230 31540 51240 31620
rect 51550 31540 51560 31620
rect 51150 31440 51230 31450
rect 51470 31440 51550 31450
rect 51230 31360 51240 31440
rect 51550 31360 51560 31440
rect 51150 31260 51230 31270
rect 51470 31260 51550 31270
rect 51230 31180 51240 31260
rect 51550 31180 51560 31260
rect 51730 31100 51740 37100
rect 51750 31100 51780 37100
rect 51850 37030 51880 37100
rect 52080 37030 52110 37100
rect 51790 37020 51880 37030
rect 51940 37020 52020 37030
rect 52080 37020 52170 37030
rect 52180 37020 52210 37100
rect 51850 36850 51880 37020
rect 52020 36940 52030 37020
rect 52080 36850 52110 37020
rect 52170 36940 52210 37020
rect 51790 36840 51880 36850
rect 51940 36840 52020 36850
rect 52080 36840 52170 36850
rect 52180 36840 52210 36940
rect 51850 36670 51880 36840
rect 52020 36760 52030 36840
rect 52080 36670 52110 36840
rect 52170 36760 52210 36840
rect 51790 36660 51880 36670
rect 51940 36660 52020 36670
rect 52080 36660 52170 36670
rect 52180 36660 52210 36760
rect 51850 36490 51880 36660
rect 52020 36580 52030 36660
rect 52080 36490 52110 36660
rect 52170 36580 52210 36660
rect 51790 36480 51880 36490
rect 51940 36480 52020 36490
rect 52080 36480 52170 36490
rect 52180 36480 52210 36580
rect 51850 36310 51880 36480
rect 52020 36400 52030 36480
rect 52080 36310 52110 36480
rect 52170 36400 52210 36480
rect 51790 36300 51880 36310
rect 51940 36300 52020 36310
rect 52080 36300 52170 36310
rect 52180 36300 52210 36400
rect 51850 36130 51880 36300
rect 52020 36220 52030 36300
rect 52080 36130 52110 36300
rect 52170 36220 52210 36300
rect 51790 36120 51880 36130
rect 51940 36120 52020 36130
rect 52080 36120 52170 36130
rect 52180 36120 52210 36220
rect 51850 35950 51880 36120
rect 52020 36040 52030 36120
rect 52080 35950 52110 36120
rect 52170 36040 52210 36120
rect 51790 35940 51880 35950
rect 51940 35940 52020 35950
rect 52080 35940 52170 35950
rect 52180 35940 52210 36040
rect 51850 35770 51880 35940
rect 52020 35860 52030 35940
rect 52080 35770 52110 35940
rect 52170 35860 52210 35940
rect 51790 35760 51880 35770
rect 51940 35760 52020 35770
rect 52080 35760 52170 35770
rect 52180 35760 52210 35860
rect 51850 35590 51880 35760
rect 52020 35680 52030 35760
rect 52080 35590 52110 35760
rect 52170 35680 52210 35760
rect 51790 35580 51880 35590
rect 51940 35580 52020 35590
rect 52080 35580 52170 35590
rect 52180 35580 52210 35680
rect 51850 35410 51880 35580
rect 52020 35500 52030 35580
rect 52080 35410 52110 35580
rect 52170 35500 52210 35580
rect 51790 35400 51880 35410
rect 51940 35400 52020 35410
rect 52080 35400 52170 35410
rect 52180 35400 52210 35500
rect 51850 35230 51880 35400
rect 52020 35320 52030 35400
rect 52080 35230 52110 35400
rect 52170 35320 52210 35400
rect 51790 35220 51880 35230
rect 51940 35220 52020 35230
rect 52080 35220 52170 35230
rect 52180 35220 52210 35320
rect 51850 35050 51880 35220
rect 52020 35140 52030 35220
rect 52080 35050 52110 35220
rect 52170 35140 52210 35220
rect 51790 35040 51880 35050
rect 51940 35040 52020 35050
rect 52080 35040 52170 35050
rect 52180 35040 52210 35140
rect 51850 34870 51880 35040
rect 52020 34960 52030 35040
rect 52080 34870 52110 35040
rect 52170 34960 52210 35040
rect 51790 34860 51880 34870
rect 51940 34860 52020 34870
rect 52080 34860 52170 34870
rect 52180 34860 52210 34960
rect 51850 34690 51880 34860
rect 52020 34780 52030 34860
rect 52080 34690 52110 34860
rect 52170 34780 52210 34860
rect 51790 34680 51880 34690
rect 51940 34680 52020 34690
rect 52080 34680 52170 34690
rect 52180 34680 52210 34780
rect 51850 34510 51880 34680
rect 52020 34600 52030 34680
rect 52080 34510 52110 34680
rect 52170 34600 52210 34680
rect 51790 34500 51880 34510
rect 51940 34500 52020 34510
rect 52080 34500 52170 34510
rect 52180 34500 52210 34600
rect 51850 34330 51880 34500
rect 52020 34420 52030 34500
rect 52080 34330 52110 34500
rect 52170 34420 52210 34500
rect 51790 34320 51880 34330
rect 51940 34320 52020 34330
rect 52080 34320 52170 34330
rect 52180 34320 52210 34420
rect 51850 34150 51880 34320
rect 52020 34240 52030 34320
rect 52080 34150 52110 34320
rect 52170 34240 52210 34320
rect 51790 34140 51880 34150
rect 51940 34140 52020 34150
rect 52080 34140 52170 34150
rect 52180 34140 52210 34240
rect 51850 33970 51880 34140
rect 52020 34060 52030 34140
rect 52080 33970 52110 34140
rect 52170 34060 52210 34140
rect 51790 33960 51880 33970
rect 51940 33960 52020 33970
rect 52080 33960 52170 33970
rect 52180 33960 52210 34060
rect 51850 33790 51880 33960
rect 52020 33880 52030 33960
rect 52080 33790 52110 33960
rect 52170 33880 52210 33960
rect 51790 33780 51880 33790
rect 51940 33780 52020 33790
rect 52080 33780 52170 33790
rect 52180 33780 52210 33880
rect 51850 33610 51880 33780
rect 52020 33700 52030 33780
rect 52080 33610 52110 33780
rect 52170 33700 52210 33780
rect 51790 33600 51880 33610
rect 51940 33600 52020 33610
rect 52080 33600 52170 33610
rect 52180 33600 52210 33700
rect 51850 33430 51880 33600
rect 52020 33520 52030 33600
rect 52080 33430 52110 33600
rect 52170 33520 52210 33600
rect 51790 33420 51880 33430
rect 51940 33420 52020 33430
rect 52080 33420 52170 33430
rect 52180 33420 52210 33520
rect 51850 33250 51880 33420
rect 52020 33340 52030 33420
rect 52080 33250 52110 33420
rect 52170 33340 52210 33420
rect 51790 33240 51880 33250
rect 51940 33240 52020 33250
rect 52080 33240 52170 33250
rect 52180 33240 52210 33340
rect 51850 33070 51880 33240
rect 52020 33160 52030 33240
rect 52080 33070 52110 33240
rect 52170 33160 52210 33240
rect 51790 33060 51880 33070
rect 51940 33060 52020 33070
rect 52080 33060 52170 33070
rect 52180 33060 52210 33160
rect 51850 32890 51880 33060
rect 52020 32980 52030 33060
rect 52080 32890 52110 33060
rect 52170 32980 52210 33060
rect 51790 32880 51880 32890
rect 51940 32880 52020 32890
rect 52080 32880 52170 32890
rect 52180 32880 52210 32980
rect 51850 32710 51880 32880
rect 52020 32800 52030 32880
rect 52080 32710 52110 32880
rect 52170 32800 52210 32880
rect 51790 32700 51880 32710
rect 51940 32700 52020 32710
rect 52080 32700 52170 32710
rect 52180 32700 52210 32800
rect 51850 32530 51880 32700
rect 52020 32620 52030 32700
rect 52080 32530 52110 32700
rect 52170 32620 52210 32700
rect 51790 32520 51880 32530
rect 51940 32520 52020 32530
rect 52080 32520 52170 32530
rect 52180 32520 52210 32620
rect 51850 32350 51880 32520
rect 52020 32440 52030 32520
rect 52080 32350 52110 32520
rect 52170 32440 52210 32520
rect 51790 32340 51880 32350
rect 51940 32340 52020 32350
rect 52080 32340 52170 32350
rect 52180 32340 52210 32440
rect 51850 32170 51880 32340
rect 52020 32260 52030 32340
rect 52080 32170 52110 32340
rect 52170 32260 52210 32340
rect 51790 32160 51880 32170
rect 51940 32160 52020 32170
rect 52080 32160 52170 32170
rect 52180 32160 52210 32260
rect 51850 31990 51880 32160
rect 52020 32080 52030 32160
rect 52080 31990 52110 32160
rect 52170 32080 52210 32160
rect 51790 31980 51880 31990
rect 51940 31980 52020 31990
rect 52080 31980 52170 31990
rect 52180 31980 52210 32080
rect 51850 31810 51880 31980
rect 52020 31900 52030 31980
rect 52080 31810 52110 31980
rect 52170 31900 52210 31980
rect 51790 31800 51880 31810
rect 51940 31800 52020 31810
rect 52080 31800 52170 31810
rect 52180 31800 52210 31900
rect 51850 31630 51880 31800
rect 52020 31720 52030 31800
rect 52080 31630 52110 31800
rect 52170 31720 52210 31800
rect 51790 31620 51880 31630
rect 51940 31620 52020 31630
rect 52080 31620 52170 31630
rect 52180 31620 52210 31720
rect 51850 31450 51880 31620
rect 52020 31540 52030 31620
rect 52080 31450 52110 31620
rect 52170 31540 52210 31620
rect 51790 31440 51880 31450
rect 51940 31440 52020 31450
rect 52080 31440 52170 31450
rect 52180 31440 52210 31540
rect 51850 31270 51880 31440
rect 52020 31360 52030 31440
rect 52080 31270 52110 31440
rect 52170 31360 52210 31440
rect 51790 31260 51880 31270
rect 51940 31260 52020 31270
rect 52080 31260 52170 31270
rect 52180 31260 52210 31360
rect 51850 31100 51880 31260
rect 52020 31180 52030 31260
rect 52080 31100 52110 31260
rect 52170 31180 52210 31260
rect 52180 31100 52210 31180
rect 52310 31100 52320 37100
rect 52410 37020 52490 37030
rect 52730 37020 52810 37030
rect 52490 36940 52500 37020
rect 52810 36940 52820 37020
rect 52410 36840 52490 36850
rect 52730 36840 52810 36850
rect 52490 36760 52500 36840
rect 52810 36760 52820 36840
rect 52410 36660 52490 36670
rect 52730 36660 52810 36670
rect 52490 36580 52500 36660
rect 52810 36580 52820 36660
rect 52410 36480 52490 36490
rect 52730 36480 52810 36490
rect 52490 36400 52500 36480
rect 52810 36400 52820 36480
rect 52410 36300 52490 36310
rect 52730 36300 52810 36310
rect 52490 36220 52500 36300
rect 52810 36220 52820 36300
rect 52410 36120 52490 36130
rect 52730 36120 52810 36130
rect 52490 36040 52500 36120
rect 52810 36040 52820 36120
rect 52410 35940 52490 35950
rect 52730 35940 52810 35950
rect 52490 35860 52500 35940
rect 52810 35860 52820 35940
rect 52410 35760 52490 35770
rect 52730 35760 52810 35770
rect 52490 35680 52500 35760
rect 52810 35680 52820 35760
rect 52410 35580 52490 35590
rect 52730 35580 52810 35590
rect 52490 35500 52500 35580
rect 52810 35500 52820 35580
rect 52410 35400 52490 35410
rect 52730 35400 52810 35410
rect 52490 35320 52500 35400
rect 52810 35320 52820 35400
rect 52410 35220 52490 35230
rect 52730 35220 52810 35230
rect 52490 35140 52500 35220
rect 52810 35140 52820 35220
rect 52410 35040 52490 35050
rect 52730 35040 52810 35050
rect 52490 34960 52500 35040
rect 52810 34960 52820 35040
rect 52410 34860 52490 34870
rect 52730 34860 52810 34870
rect 52490 34780 52500 34860
rect 52810 34780 52820 34860
rect 52410 34680 52490 34690
rect 52730 34680 52810 34690
rect 52490 34600 52500 34680
rect 52810 34600 52820 34680
rect 52410 34500 52490 34510
rect 52730 34500 52810 34510
rect 52490 34420 52500 34500
rect 52810 34420 52820 34500
rect 52410 34320 52490 34330
rect 52730 34320 52810 34330
rect 52490 34240 52500 34320
rect 52810 34240 52820 34320
rect 52410 34140 52490 34150
rect 52730 34140 52810 34150
rect 52490 34060 52500 34140
rect 52810 34060 52820 34140
rect 52410 33960 52490 33970
rect 52730 33960 52810 33970
rect 52490 33880 52500 33960
rect 52810 33880 52820 33960
rect 52410 33780 52490 33790
rect 52730 33780 52810 33790
rect 52490 33700 52500 33780
rect 52810 33700 52820 33780
rect 52410 33600 52490 33610
rect 52730 33600 52810 33610
rect 52490 33520 52500 33600
rect 52810 33520 52820 33600
rect 52410 33420 52490 33430
rect 52730 33420 52810 33430
rect 52490 33340 52500 33420
rect 52810 33340 52820 33420
rect 52410 33240 52490 33250
rect 52730 33240 52810 33250
rect 52490 33160 52500 33240
rect 52810 33160 52820 33240
rect 52410 33060 52490 33070
rect 52730 33060 52810 33070
rect 52490 32980 52500 33060
rect 52810 32980 52820 33060
rect 52410 32880 52490 32890
rect 52730 32880 52810 32890
rect 52490 32800 52500 32880
rect 52810 32800 52820 32880
rect 52410 32700 52490 32710
rect 52730 32700 52810 32710
rect 52490 32620 52500 32700
rect 52810 32620 52820 32700
rect 52410 32520 52490 32530
rect 52730 32520 52810 32530
rect 52490 32440 52500 32520
rect 52810 32440 52820 32520
rect 52410 32340 52490 32350
rect 52730 32340 52810 32350
rect 52490 32260 52500 32340
rect 52810 32260 52820 32340
rect 52410 32160 52490 32170
rect 52730 32160 52810 32170
rect 52490 32080 52500 32160
rect 52810 32080 52820 32160
rect 52410 31980 52490 31990
rect 52730 31980 52810 31990
rect 52490 31900 52500 31980
rect 52810 31900 52820 31980
rect 52410 31800 52490 31810
rect 52730 31800 52810 31810
rect 52490 31720 52500 31800
rect 52810 31720 52820 31800
rect 52410 31620 52490 31630
rect 52730 31620 52810 31630
rect 52490 31540 52500 31620
rect 52810 31540 52820 31620
rect 52410 31440 52490 31450
rect 52730 31440 52810 31450
rect 52490 31360 52500 31440
rect 52810 31360 52820 31440
rect 52410 31260 52490 31270
rect 52730 31260 52810 31270
rect 52490 31180 52500 31260
rect 52810 31180 52820 31260
rect 52990 31100 53000 37100
rect 53010 31100 53040 37100
rect 53110 37030 53140 37100
rect 53340 37030 53370 37100
rect 53050 37020 53140 37030
rect 53200 37020 53280 37030
rect 53340 37020 53430 37030
rect 53440 37020 53470 37100
rect 53110 36850 53140 37020
rect 53280 36940 53290 37020
rect 53340 36850 53370 37020
rect 53430 36940 53470 37020
rect 53050 36840 53140 36850
rect 53200 36840 53280 36850
rect 53340 36840 53430 36850
rect 53440 36840 53470 36940
rect 53110 36670 53140 36840
rect 53280 36760 53290 36840
rect 53340 36670 53370 36840
rect 53430 36760 53470 36840
rect 53050 36660 53140 36670
rect 53200 36660 53280 36670
rect 53340 36660 53430 36670
rect 53440 36660 53470 36760
rect 53110 36490 53140 36660
rect 53280 36580 53290 36660
rect 53340 36490 53370 36660
rect 53430 36580 53470 36660
rect 53050 36480 53140 36490
rect 53200 36480 53280 36490
rect 53340 36480 53430 36490
rect 53440 36480 53470 36580
rect 53110 36310 53140 36480
rect 53280 36400 53290 36480
rect 53340 36310 53370 36480
rect 53430 36400 53470 36480
rect 53050 36300 53140 36310
rect 53200 36300 53280 36310
rect 53340 36300 53430 36310
rect 53440 36300 53470 36400
rect 53110 36130 53140 36300
rect 53280 36220 53290 36300
rect 53340 36130 53370 36300
rect 53430 36220 53470 36300
rect 53050 36120 53140 36130
rect 53200 36120 53280 36130
rect 53340 36120 53430 36130
rect 53440 36120 53470 36220
rect 53110 35950 53140 36120
rect 53280 36040 53290 36120
rect 53340 35950 53370 36120
rect 53430 36040 53470 36120
rect 53050 35940 53140 35950
rect 53200 35940 53280 35950
rect 53340 35940 53430 35950
rect 53440 35940 53470 36040
rect 53110 35770 53140 35940
rect 53280 35860 53290 35940
rect 53340 35770 53370 35940
rect 53430 35860 53470 35940
rect 53050 35760 53140 35770
rect 53200 35760 53280 35770
rect 53340 35760 53430 35770
rect 53440 35760 53470 35860
rect 53110 35590 53140 35760
rect 53280 35680 53290 35760
rect 53340 35590 53370 35760
rect 53430 35680 53470 35760
rect 53050 35580 53140 35590
rect 53200 35580 53280 35590
rect 53340 35580 53430 35590
rect 53440 35580 53470 35680
rect 53110 35410 53140 35580
rect 53280 35500 53290 35580
rect 53340 35410 53370 35580
rect 53430 35500 53470 35580
rect 53050 35400 53140 35410
rect 53200 35400 53280 35410
rect 53340 35400 53430 35410
rect 53440 35400 53470 35500
rect 53110 35230 53140 35400
rect 53280 35320 53290 35400
rect 53340 35230 53370 35400
rect 53430 35320 53470 35400
rect 53050 35220 53140 35230
rect 53200 35220 53280 35230
rect 53340 35220 53430 35230
rect 53440 35220 53470 35320
rect 53110 35050 53140 35220
rect 53280 35140 53290 35220
rect 53340 35050 53370 35220
rect 53430 35140 53470 35220
rect 53050 35040 53140 35050
rect 53200 35040 53280 35050
rect 53340 35040 53430 35050
rect 53440 35040 53470 35140
rect 53110 34870 53140 35040
rect 53280 34960 53290 35040
rect 53340 34870 53370 35040
rect 53430 34960 53470 35040
rect 53050 34860 53140 34870
rect 53200 34860 53280 34870
rect 53340 34860 53430 34870
rect 53440 34860 53470 34960
rect 53110 34690 53140 34860
rect 53280 34780 53290 34860
rect 53340 34690 53370 34860
rect 53430 34780 53470 34860
rect 53050 34680 53140 34690
rect 53200 34680 53280 34690
rect 53340 34680 53430 34690
rect 53440 34680 53470 34780
rect 53110 34510 53140 34680
rect 53280 34600 53290 34680
rect 53340 34510 53370 34680
rect 53430 34600 53470 34680
rect 53050 34500 53140 34510
rect 53200 34500 53280 34510
rect 53340 34500 53430 34510
rect 53440 34500 53470 34600
rect 53110 34330 53140 34500
rect 53280 34420 53290 34500
rect 53340 34330 53370 34500
rect 53430 34420 53470 34500
rect 53050 34320 53140 34330
rect 53200 34320 53280 34330
rect 53340 34320 53430 34330
rect 53440 34320 53470 34420
rect 53110 34150 53140 34320
rect 53280 34240 53290 34320
rect 53340 34150 53370 34320
rect 53430 34240 53470 34320
rect 53050 34140 53140 34150
rect 53200 34140 53280 34150
rect 53340 34140 53430 34150
rect 53440 34140 53470 34240
rect 53110 33970 53140 34140
rect 53280 34060 53290 34140
rect 53340 33970 53370 34140
rect 53430 34060 53470 34140
rect 53050 33960 53140 33970
rect 53200 33960 53280 33970
rect 53340 33960 53430 33970
rect 53440 33960 53470 34060
rect 53110 33790 53140 33960
rect 53280 33880 53290 33960
rect 53340 33790 53370 33960
rect 53430 33880 53470 33960
rect 53050 33780 53140 33790
rect 53200 33780 53280 33790
rect 53340 33780 53430 33790
rect 53440 33780 53470 33880
rect 53110 33610 53140 33780
rect 53280 33700 53290 33780
rect 53340 33610 53370 33780
rect 53430 33700 53470 33780
rect 53050 33600 53140 33610
rect 53200 33600 53280 33610
rect 53340 33600 53430 33610
rect 53440 33600 53470 33700
rect 53110 33430 53140 33600
rect 53280 33520 53290 33600
rect 53340 33430 53370 33600
rect 53430 33520 53470 33600
rect 53050 33420 53140 33430
rect 53200 33420 53280 33430
rect 53340 33420 53430 33430
rect 53440 33420 53470 33520
rect 53110 33250 53140 33420
rect 53280 33340 53290 33420
rect 53340 33250 53370 33420
rect 53430 33340 53470 33420
rect 53050 33240 53140 33250
rect 53200 33240 53280 33250
rect 53340 33240 53430 33250
rect 53440 33240 53470 33340
rect 53110 33070 53140 33240
rect 53280 33160 53290 33240
rect 53340 33070 53370 33240
rect 53430 33160 53470 33240
rect 53050 33060 53140 33070
rect 53200 33060 53280 33070
rect 53340 33060 53430 33070
rect 53440 33060 53470 33160
rect 53110 32890 53140 33060
rect 53280 32980 53290 33060
rect 53340 32890 53370 33060
rect 53430 32980 53470 33060
rect 53050 32880 53140 32890
rect 53200 32880 53280 32890
rect 53340 32880 53430 32890
rect 53440 32880 53470 32980
rect 53110 32710 53140 32880
rect 53280 32800 53290 32880
rect 53340 32710 53370 32880
rect 53430 32800 53470 32880
rect 53050 32700 53140 32710
rect 53200 32700 53280 32710
rect 53340 32700 53430 32710
rect 53440 32700 53470 32800
rect 53110 32530 53140 32700
rect 53280 32620 53290 32700
rect 53340 32530 53370 32700
rect 53430 32620 53470 32700
rect 53050 32520 53140 32530
rect 53200 32520 53280 32530
rect 53340 32520 53430 32530
rect 53440 32520 53470 32620
rect 53110 32350 53140 32520
rect 53280 32440 53290 32520
rect 53340 32350 53370 32520
rect 53430 32440 53470 32520
rect 53050 32340 53140 32350
rect 53200 32340 53280 32350
rect 53340 32340 53430 32350
rect 53440 32340 53470 32440
rect 53110 32170 53140 32340
rect 53280 32260 53290 32340
rect 53340 32170 53370 32340
rect 53430 32260 53470 32340
rect 53050 32160 53140 32170
rect 53200 32160 53280 32170
rect 53340 32160 53430 32170
rect 53440 32160 53470 32260
rect 53110 31990 53140 32160
rect 53280 32080 53290 32160
rect 53340 31990 53370 32160
rect 53430 32080 53470 32160
rect 53050 31980 53140 31990
rect 53200 31980 53280 31990
rect 53340 31980 53430 31990
rect 53440 31980 53470 32080
rect 53110 31810 53140 31980
rect 53280 31900 53290 31980
rect 53340 31810 53370 31980
rect 53430 31900 53470 31980
rect 53050 31800 53140 31810
rect 53200 31800 53280 31810
rect 53340 31800 53430 31810
rect 53440 31800 53470 31900
rect 53110 31630 53140 31800
rect 53280 31720 53290 31800
rect 53340 31630 53370 31800
rect 53430 31720 53470 31800
rect 53050 31620 53140 31630
rect 53200 31620 53280 31630
rect 53340 31620 53430 31630
rect 53440 31620 53470 31720
rect 53110 31450 53140 31620
rect 53280 31540 53290 31620
rect 53340 31450 53370 31620
rect 53430 31540 53470 31620
rect 53050 31440 53140 31450
rect 53200 31440 53280 31450
rect 53340 31440 53430 31450
rect 53440 31440 53470 31540
rect 53110 31270 53140 31440
rect 53280 31360 53290 31440
rect 53340 31270 53370 31440
rect 53430 31360 53470 31440
rect 53050 31260 53140 31270
rect 53200 31260 53280 31270
rect 53340 31260 53430 31270
rect 53440 31260 53470 31360
rect 53110 31100 53140 31260
rect 53280 31180 53290 31260
rect 53340 31100 53370 31260
rect 53430 31180 53470 31260
rect 53440 31100 53470 31180
rect 53570 31100 53580 37100
rect 53670 37020 53750 37030
rect 53990 37020 54070 37030
rect 53750 36940 53760 37020
rect 54070 36940 54080 37020
rect 53670 36840 53750 36850
rect 53990 36840 54070 36850
rect 53750 36760 53760 36840
rect 54070 36760 54080 36840
rect 53670 36660 53750 36670
rect 53990 36660 54070 36670
rect 53750 36580 53760 36660
rect 54070 36580 54080 36660
rect 53670 36480 53750 36490
rect 53990 36480 54070 36490
rect 53750 36400 53760 36480
rect 54070 36400 54080 36480
rect 53670 36300 53750 36310
rect 53990 36300 54070 36310
rect 53750 36220 53760 36300
rect 54070 36220 54080 36300
rect 53670 36120 53750 36130
rect 53990 36120 54070 36130
rect 53750 36040 53760 36120
rect 54070 36040 54080 36120
rect 53670 35940 53750 35950
rect 53990 35940 54070 35950
rect 53750 35860 53760 35940
rect 54070 35860 54080 35940
rect 53670 35760 53750 35770
rect 53990 35760 54070 35770
rect 53750 35680 53760 35760
rect 54070 35680 54080 35760
rect 53670 35580 53750 35590
rect 53990 35580 54070 35590
rect 53750 35500 53760 35580
rect 54070 35500 54080 35580
rect 53670 35400 53750 35410
rect 53990 35400 54070 35410
rect 53750 35320 53760 35400
rect 54070 35320 54080 35400
rect 53670 35220 53750 35230
rect 53990 35220 54070 35230
rect 53750 35140 53760 35220
rect 54070 35140 54080 35220
rect 53670 35040 53750 35050
rect 53990 35040 54070 35050
rect 53750 34960 53760 35040
rect 54070 34960 54080 35040
rect 53670 34860 53750 34870
rect 53990 34860 54070 34870
rect 53750 34780 53760 34860
rect 54070 34780 54080 34860
rect 53670 34680 53750 34690
rect 53990 34680 54070 34690
rect 53750 34600 53760 34680
rect 54070 34600 54080 34680
rect 53670 34500 53750 34510
rect 53990 34500 54070 34510
rect 53750 34420 53760 34500
rect 54070 34420 54080 34500
rect 53670 34320 53750 34330
rect 53990 34320 54070 34330
rect 53750 34240 53760 34320
rect 54070 34240 54080 34320
rect 53670 34140 53750 34150
rect 53990 34140 54070 34150
rect 53750 34060 53760 34140
rect 54070 34060 54080 34140
rect 53670 33960 53750 33970
rect 53990 33960 54070 33970
rect 53750 33880 53760 33960
rect 54070 33880 54080 33960
rect 53670 33780 53750 33790
rect 53990 33780 54070 33790
rect 53750 33700 53760 33780
rect 54070 33700 54080 33780
rect 53670 33600 53750 33610
rect 53990 33600 54070 33610
rect 53750 33520 53760 33600
rect 54070 33520 54080 33600
rect 53670 33420 53750 33430
rect 53990 33420 54070 33430
rect 53750 33340 53760 33420
rect 54070 33340 54080 33420
rect 53670 33240 53750 33250
rect 53990 33240 54070 33250
rect 53750 33160 53760 33240
rect 54070 33160 54080 33240
rect 53670 33060 53750 33070
rect 53990 33060 54070 33070
rect 53750 32980 53760 33060
rect 54070 32980 54080 33060
rect 53670 32880 53750 32890
rect 53990 32880 54070 32890
rect 53750 32800 53760 32880
rect 54070 32800 54080 32880
rect 53670 32700 53750 32710
rect 53990 32700 54070 32710
rect 53750 32620 53760 32700
rect 54070 32620 54080 32700
rect 53670 32520 53750 32530
rect 53990 32520 54070 32530
rect 53750 32440 53760 32520
rect 54070 32440 54080 32520
rect 53670 32340 53750 32350
rect 53990 32340 54070 32350
rect 53750 32260 53760 32340
rect 54070 32260 54080 32340
rect 53670 32160 53750 32170
rect 53990 32160 54070 32170
rect 53750 32080 53760 32160
rect 54070 32080 54080 32160
rect 53670 31980 53750 31990
rect 53990 31980 54070 31990
rect 53750 31900 53760 31980
rect 54070 31900 54080 31980
rect 53670 31800 53750 31810
rect 53990 31800 54070 31810
rect 53750 31720 53760 31800
rect 54070 31720 54080 31800
rect 53670 31620 53750 31630
rect 53990 31620 54070 31630
rect 53750 31540 53760 31620
rect 54070 31540 54080 31620
rect 53670 31440 53750 31450
rect 53990 31440 54070 31450
rect 53750 31360 53760 31440
rect 54070 31360 54080 31440
rect 53670 31260 53750 31270
rect 53990 31260 54070 31270
rect 53750 31180 53760 31260
rect 54070 31180 54080 31260
rect 54250 31100 54260 37100
rect 54270 31100 54300 37100
rect 54370 37030 54400 37100
rect 54600 37030 54630 37100
rect 54310 37020 54400 37030
rect 54460 37020 54540 37030
rect 54600 37020 54690 37030
rect 54700 37020 54730 37100
rect 54370 36850 54400 37020
rect 54540 36940 54550 37020
rect 54600 36850 54630 37020
rect 54690 36940 54730 37020
rect 54310 36840 54400 36850
rect 54460 36840 54540 36850
rect 54600 36840 54690 36850
rect 54700 36840 54730 36940
rect 54370 36670 54400 36840
rect 54540 36760 54550 36840
rect 54600 36670 54630 36840
rect 54690 36760 54730 36840
rect 54310 36660 54400 36670
rect 54460 36660 54540 36670
rect 54600 36660 54690 36670
rect 54700 36660 54730 36760
rect 54370 36490 54400 36660
rect 54540 36580 54550 36660
rect 54600 36490 54630 36660
rect 54690 36580 54730 36660
rect 54310 36480 54400 36490
rect 54460 36480 54540 36490
rect 54600 36480 54690 36490
rect 54700 36480 54730 36580
rect 54370 36310 54400 36480
rect 54540 36400 54550 36480
rect 54600 36310 54630 36480
rect 54690 36400 54730 36480
rect 54310 36300 54400 36310
rect 54460 36300 54540 36310
rect 54600 36300 54690 36310
rect 54700 36300 54730 36400
rect 54370 36130 54400 36300
rect 54540 36220 54550 36300
rect 54600 36130 54630 36300
rect 54690 36220 54730 36300
rect 54310 36120 54400 36130
rect 54460 36120 54540 36130
rect 54600 36120 54690 36130
rect 54700 36120 54730 36220
rect 54370 35950 54400 36120
rect 54540 36040 54550 36120
rect 54600 35950 54630 36120
rect 54690 36040 54730 36120
rect 54310 35940 54400 35950
rect 54460 35940 54540 35950
rect 54600 35940 54690 35950
rect 54700 35940 54730 36040
rect 54370 35770 54400 35940
rect 54540 35860 54550 35940
rect 54600 35770 54630 35940
rect 54690 35860 54730 35940
rect 54310 35760 54400 35770
rect 54460 35760 54540 35770
rect 54600 35760 54690 35770
rect 54700 35760 54730 35860
rect 54370 35590 54400 35760
rect 54540 35680 54550 35760
rect 54600 35590 54630 35760
rect 54690 35680 54730 35760
rect 54310 35580 54400 35590
rect 54460 35580 54540 35590
rect 54600 35580 54690 35590
rect 54700 35580 54730 35680
rect 54370 35410 54400 35580
rect 54540 35500 54550 35580
rect 54600 35410 54630 35580
rect 54690 35500 54730 35580
rect 54310 35400 54400 35410
rect 54460 35400 54540 35410
rect 54600 35400 54690 35410
rect 54700 35400 54730 35500
rect 54370 35230 54400 35400
rect 54540 35320 54550 35400
rect 54600 35230 54630 35400
rect 54690 35320 54730 35400
rect 54310 35220 54400 35230
rect 54460 35220 54540 35230
rect 54600 35220 54690 35230
rect 54700 35220 54730 35320
rect 54370 35050 54400 35220
rect 54540 35140 54550 35220
rect 54600 35050 54630 35220
rect 54690 35140 54730 35220
rect 54310 35040 54400 35050
rect 54460 35040 54540 35050
rect 54600 35040 54690 35050
rect 54700 35040 54730 35140
rect 54370 34870 54400 35040
rect 54540 34960 54550 35040
rect 54600 34870 54630 35040
rect 54690 34960 54730 35040
rect 54310 34860 54400 34870
rect 54460 34860 54540 34870
rect 54600 34860 54690 34870
rect 54700 34860 54730 34960
rect 54370 34690 54400 34860
rect 54540 34780 54550 34860
rect 54600 34690 54630 34860
rect 54690 34780 54730 34860
rect 54310 34680 54400 34690
rect 54460 34680 54540 34690
rect 54600 34680 54690 34690
rect 54700 34680 54730 34780
rect 54370 34510 54400 34680
rect 54540 34600 54550 34680
rect 54600 34510 54630 34680
rect 54690 34600 54730 34680
rect 54310 34500 54400 34510
rect 54460 34500 54540 34510
rect 54600 34500 54690 34510
rect 54700 34500 54730 34600
rect 54370 34330 54400 34500
rect 54540 34420 54550 34500
rect 54600 34330 54630 34500
rect 54690 34420 54730 34500
rect 54310 34320 54400 34330
rect 54460 34320 54540 34330
rect 54600 34320 54690 34330
rect 54700 34320 54730 34420
rect 54370 34150 54400 34320
rect 54540 34240 54550 34320
rect 54600 34150 54630 34320
rect 54690 34240 54730 34320
rect 54310 34140 54400 34150
rect 54460 34140 54540 34150
rect 54600 34140 54690 34150
rect 54700 34140 54730 34240
rect 54370 33970 54400 34140
rect 54540 34060 54550 34140
rect 54600 33970 54630 34140
rect 54690 34060 54730 34140
rect 54310 33960 54400 33970
rect 54460 33960 54540 33970
rect 54600 33960 54690 33970
rect 54700 33960 54730 34060
rect 54370 33790 54400 33960
rect 54540 33880 54550 33960
rect 54600 33790 54630 33960
rect 54690 33880 54730 33960
rect 54310 33780 54400 33790
rect 54460 33780 54540 33790
rect 54600 33780 54690 33790
rect 54700 33780 54730 33880
rect 54370 33610 54400 33780
rect 54540 33700 54550 33780
rect 54600 33610 54630 33780
rect 54690 33700 54730 33780
rect 54310 33600 54400 33610
rect 54460 33600 54540 33610
rect 54600 33600 54690 33610
rect 54700 33600 54730 33700
rect 54370 33430 54400 33600
rect 54540 33520 54550 33600
rect 54600 33430 54630 33600
rect 54690 33520 54730 33600
rect 54310 33420 54400 33430
rect 54460 33420 54540 33430
rect 54600 33420 54690 33430
rect 54700 33420 54730 33520
rect 54370 33250 54400 33420
rect 54540 33340 54550 33420
rect 54600 33250 54630 33420
rect 54690 33340 54730 33420
rect 54310 33240 54400 33250
rect 54460 33240 54540 33250
rect 54600 33240 54690 33250
rect 54700 33240 54730 33340
rect 54370 33070 54400 33240
rect 54540 33160 54550 33240
rect 54600 33070 54630 33240
rect 54690 33160 54730 33240
rect 54310 33060 54400 33070
rect 54460 33060 54540 33070
rect 54600 33060 54690 33070
rect 54700 33060 54730 33160
rect 54370 32890 54400 33060
rect 54540 32980 54550 33060
rect 54600 32890 54630 33060
rect 54690 32980 54730 33060
rect 54310 32880 54400 32890
rect 54460 32880 54540 32890
rect 54600 32880 54690 32890
rect 54700 32880 54730 32980
rect 54370 32710 54400 32880
rect 54540 32800 54550 32880
rect 54600 32710 54630 32880
rect 54690 32800 54730 32880
rect 54310 32700 54400 32710
rect 54460 32700 54540 32710
rect 54600 32700 54690 32710
rect 54700 32700 54730 32800
rect 54370 32530 54400 32700
rect 54540 32620 54550 32700
rect 54600 32530 54630 32700
rect 54690 32620 54730 32700
rect 54310 32520 54400 32530
rect 54460 32520 54540 32530
rect 54600 32520 54690 32530
rect 54700 32520 54730 32620
rect 54370 32350 54400 32520
rect 54540 32440 54550 32520
rect 54600 32350 54630 32520
rect 54690 32440 54730 32520
rect 54310 32340 54400 32350
rect 54460 32340 54540 32350
rect 54600 32340 54690 32350
rect 54700 32340 54730 32440
rect 54370 32170 54400 32340
rect 54540 32260 54550 32340
rect 54600 32170 54630 32340
rect 54690 32260 54730 32340
rect 54310 32160 54400 32170
rect 54460 32160 54540 32170
rect 54600 32160 54690 32170
rect 54700 32160 54730 32260
rect 54370 31990 54400 32160
rect 54540 32080 54550 32160
rect 54600 31990 54630 32160
rect 54690 32080 54730 32160
rect 54310 31980 54400 31990
rect 54460 31980 54540 31990
rect 54600 31980 54690 31990
rect 54700 31980 54730 32080
rect 54370 31810 54400 31980
rect 54540 31900 54550 31980
rect 54600 31810 54630 31980
rect 54690 31900 54730 31980
rect 54310 31800 54400 31810
rect 54460 31800 54540 31810
rect 54600 31800 54690 31810
rect 54700 31800 54730 31900
rect 54370 31630 54400 31800
rect 54540 31720 54550 31800
rect 54600 31630 54630 31800
rect 54690 31720 54730 31800
rect 54310 31620 54400 31630
rect 54460 31620 54540 31630
rect 54600 31620 54690 31630
rect 54700 31620 54730 31720
rect 54370 31450 54400 31620
rect 54540 31540 54550 31620
rect 54600 31450 54630 31620
rect 54690 31540 54730 31620
rect 54310 31440 54400 31450
rect 54460 31440 54540 31450
rect 54600 31440 54690 31450
rect 54700 31440 54730 31540
rect 54370 31270 54400 31440
rect 54540 31360 54550 31440
rect 54600 31270 54630 31440
rect 54690 31360 54730 31440
rect 54310 31260 54400 31270
rect 54460 31260 54540 31270
rect 54600 31260 54690 31270
rect 54700 31260 54730 31360
rect 54370 31100 54400 31260
rect 54540 31180 54550 31260
rect 54600 31100 54630 31260
rect 54690 31180 54730 31260
rect 54700 31100 54730 31180
rect 54830 31100 54840 37100
rect 54930 37020 55010 37030
rect 55250 37020 55330 37030
rect 55010 36940 55020 37020
rect 55330 36940 55340 37020
rect 54930 36840 55010 36850
rect 55250 36840 55330 36850
rect 55010 36760 55020 36840
rect 55330 36760 55340 36840
rect 54930 36660 55010 36670
rect 55250 36660 55330 36670
rect 55010 36580 55020 36660
rect 55330 36580 55340 36660
rect 54930 36480 55010 36490
rect 55250 36480 55330 36490
rect 55010 36400 55020 36480
rect 55330 36400 55340 36480
rect 54930 36300 55010 36310
rect 55250 36300 55330 36310
rect 55010 36220 55020 36300
rect 55330 36220 55340 36300
rect 54930 36120 55010 36130
rect 55250 36120 55330 36130
rect 55010 36040 55020 36120
rect 55330 36040 55340 36120
rect 54930 35940 55010 35950
rect 55250 35940 55330 35950
rect 55010 35860 55020 35940
rect 55330 35860 55340 35940
rect 54930 35760 55010 35770
rect 55250 35760 55330 35770
rect 55010 35680 55020 35760
rect 55330 35680 55340 35760
rect 54930 35580 55010 35590
rect 55250 35580 55330 35590
rect 55010 35500 55020 35580
rect 55330 35500 55340 35580
rect 54930 35400 55010 35410
rect 55250 35400 55330 35410
rect 55010 35320 55020 35400
rect 55330 35320 55340 35400
rect 54930 35220 55010 35230
rect 55250 35220 55330 35230
rect 55010 35140 55020 35220
rect 55330 35140 55340 35220
rect 54930 35040 55010 35050
rect 55250 35040 55330 35050
rect 55010 34960 55020 35040
rect 55330 34960 55340 35040
rect 54930 34860 55010 34870
rect 55250 34860 55330 34870
rect 55010 34780 55020 34860
rect 55330 34780 55340 34860
rect 54930 34680 55010 34690
rect 55250 34680 55330 34690
rect 55010 34600 55020 34680
rect 55330 34600 55340 34680
rect 54930 34500 55010 34510
rect 55250 34500 55330 34510
rect 55010 34420 55020 34500
rect 55330 34420 55340 34500
rect 54930 34320 55010 34330
rect 55250 34320 55330 34330
rect 55010 34240 55020 34320
rect 55330 34240 55340 34320
rect 54930 34140 55010 34150
rect 55250 34140 55330 34150
rect 55010 34060 55020 34140
rect 55330 34060 55340 34140
rect 54930 33960 55010 33970
rect 55250 33960 55330 33970
rect 55010 33880 55020 33960
rect 55330 33880 55340 33960
rect 54930 33780 55010 33790
rect 55250 33780 55330 33790
rect 55010 33700 55020 33780
rect 55330 33700 55340 33780
rect 54930 33600 55010 33610
rect 55250 33600 55330 33610
rect 55010 33520 55020 33600
rect 55330 33520 55340 33600
rect 54930 33420 55010 33430
rect 55250 33420 55330 33430
rect 55010 33340 55020 33420
rect 55330 33340 55340 33420
rect 54930 33240 55010 33250
rect 55250 33240 55330 33250
rect 55010 33160 55020 33240
rect 55330 33160 55340 33240
rect 54930 33060 55010 33070
rect 55250 33060 55330 33070
rect 55010 32980 55020 33060
rect 55330 32980 55340 33060
rect 54930 32880 55010 32890
rect 55250 32880 55330 32890
rect 55010 32800 55020 32880
rect 55330 32800 55340 32880
rect 54930 32700 55010 32710
rect 55250 32700 55330 32710
rect 55010 32620 55020 32700
rect 55330 32620 55340 32700
rect 54930 32520 55010 32530
rect 55250 32520 55330 32530
rect 55010 32440 55020 32520
rect 55330 32440 55340 32520
rect 54930 32340 55010 32350
rect 55250 32340 55330 32350
rect 55010 32260 55020 32340
rect 55330 32260 55340 32340
rect 54930 32160 55010 32170
rect 55250 32160 55330 32170
rect 55010 32080 55020 32160
rect 55330 32080 55340 32160
rect 54930 31980 55010 31990
rect 55250 31980 55330 31990
rect 55010 31900 55020 31980
rect 55330 31900 55340 31980
rect 54930 31800 55010 31810
rect 55250 31800 55330 31810
rect 55010 31720 55020 31800
rect 55330 31720 55340 31800
rect 54930 31620 55010 31630
rect 55250 31620 55330 31630
rect 55010 31540 55020 31620
rect 55330 31540 55340 31620
rect 54930 31440 55010 31450
rect 55250 31440 55330 31450
rect 55010 31360 55020 31440
rect 55330 31360 55340 31440
rect 54930 31260 55010 31270
rect 55250 31260 55330 31270
rect 55010 31180 55020 31260
rect 55330 31180 55340 31260
rect 55510 31100 55520 37100
rect 55530 31100 55560 37100
rect 55630 37030 55660 37100
rect 55860 37030 55890 37100
rect 55570 37020 55660 37030
rect 55720 37020 55800 37030
rect 55860 37020 55950 37030
rect 55960 37020 55990 37100
rect 55630 36850 55660 37020
rect 55800 36940 55810 37020
rect 55860 36850 55890 37020
rect 55950 36940 55990 37020
rect 55570 36840 55660 36850
rect 55720 36840 55800 36850
rect 55860 36840 55950 36850
rect 55960 36840 55990 36940
rect 55630 36670 55660 36840
rect 55800 36760 55810 36840
rect 55860 36670 55890 36840
rect 55950 36760 55990 36840
rect 55570 36660 55660 36670
rect 55720 36660 55800 36670
rect 55860 36660 55950 36670
rect 55960 36660 55990 36760
rect 55630 36490 55660 36660
rect 55800 36580 55810 36660
rect 55860 36490 55890 36660
rect 55950 36580 55990 36660
rect 55570 36480 55660 36490
rect 55720 36480 55800 36490
rect 55860 36480 55950 36490
rect 55960 36480 55990 36580
rect 55630 36310 55660 36480
rect 55800 36400 55810 36480
rect 55860 36310 55890 36480
rect 55950 36400 55990 36480
rect 55570 36300 55660 36310
rect 55720 36300 55800 36310
rect 55860 36300 55950 36310
rect 55960 36300 55990 36400
rect 55630 36130 55660 36300
rect 55800 36220 55810 36300
rect 55860 36130 55890 36300
rect 55950 36220 55990 36300
rect 55570 36120 55660 36130
rect 55720 36120 55800 36130
rect 55860 36120 55950 36130
rect 55960 36120 55990 36220
rect 55630 35950 55660 36120
rect 55800 36040 55810 36120
rect 55860 35950 55890 36120
rect 55950 36040 55990 36120
rect 55570 35940 55660 35950
rect 55720 35940 55800 35950
rect 55860 35940 55950 35950
rect 55960 35940 55990 36040
rect 55630 35770 55660 35940
rect 55800 35860 55810 35940
rect 55860 35770 55890 35940
rect 55950 35860 55990 35940
rect 55570 35760 55660 35770
rect 55720 35760 55800 35770
rect 55860 35760 55950 35770
rect 55960 35760 55990 35860
rect 55630 35590 55660 35760
rect 55800 35680 55810 35760
rect 55860 35590 55890 35760
rect 55950 35680 55990 35760
rect 55570 35580 55660 35590
rect 55720 35580 55800 35590
rect 55860 35580 55950 35590
rect 55960 35580 55990 35680
rect 55630 35410 55660 35580
rect 55800 35500 55810 35580
rect 55860 35410 55890 35580
rect 55950 35500 55990 35580
rect 55570 35400 55660 35410
rect 55720 35400 55800 35410
rect 55860 35400 55950 35410
rect 55960 35400 55990 35500
rect 55630 35230 55660 35400
rect 55800 35320 55810 35400
rect 55860 35230 55890 35400
rect 55950 35320 55990 35400
rect 55570 35220 55660 35230
rect 55720 35220 55800 35230
rect 55860 35220 55950 35230
rect 55960 35220 55990 35320
rect 55630 35050 55660 35220
rect 55800 35140 55810 35220
rect 55860 35050 55890 35220
rect 55950 35140 55990 35220
rect 55570 35040 55660 35050
rect 55720 35040 55800 35050
rect 55860 35040 55950 35050
rect 55960 35040 55990 35140
rect 55630 34870 55660 35040
rect 55800 34960 55810 35040
rect 55860 34870 55890 35040
rect 55950 34960 55990 35040
rect 55570 34860 55660 34870
rect 55720 34860 55800 34870
rect 55860 34860 55950 34870
rect 55960 34860 55990 34960
rect 55630 34690 55660 34860
rect 55800 34780 55810 34860
rect 55860 34690 55890 34860
rect 55950 34780 55990 34860
rect 55570 34680 55660 34690
rect 55720 34680 55800 34690
rect 55860 34680 55950 34690
rect 55960 34680 55990 34780
rect 55630 34510 55660 34680
rect 55800 34600 55810 34680
rect 55860 34510 55890 34680
rect 55950 34600 55990 34680
rect 55570 34500 55660 34510
rect 55720 34500 55800 34510
rect 55860 34500 55950 34510
rect 55960 34500 55990 34600
rect 55630 34330 55660 34500
rect 55800 34420 55810 34500
rect 55860 34330 55890 34500
rect 55950 34420 55990 34500
rect 55570 34320 55660 34330
rect 55720 34320 55800 34330
rect 55860 34320 55950 34330
rect 55960 34320 55990 34420
rect 55630 34150 55660 34320
rect 55800 34240 55810 34320
rect 55860 34150 55890 34320
rect 55950 34240 55990 34320
rect 55570 34140 55660 34150
rect 55720 34140 55800 34150
rect 55860 34140 55950 34150
rect 55960 34140 55990 34240
rect 55630 33970 55660 34140
rect 55800 34060 55810 34140
rect 55860 33970 55890 34140
rect 55950 34060 55990 34140
rect 55570 33960 55660 33970
rect 55720 33960 55800 33970
rect 55860 33960 55950 33970
rect 55960 33960 55990 34060
rect 55630 33790 55660 33960
rect 55800 33880 55810 33960
rect 55860 33790 55890 33960
rect 55950 33880 55990 33960
rect 55570 33780 55660 33790
rect 55720 33780 55800 33790
rect 55860 33780 55950 33790
rect 55960 33780 55990 33880
rect 55630 33610 55660 33780
rect 55800 33700 55810 33780
rect 55860 33610 55890 33780
rect 55950 33700 55990 33780
rect 55570 33600 55660 33610
rect 55720 33600 55800 33610
rect 55860 33600 55950 33610
rect 55960 33600 55990 33700
rect 55630 33430 55660 33600
rect 55800 33520 55810 33600
rect 55860 33430 55890 33600
rect 55950 33520 55990 33600
rect 55570 33420 55660 33430
rect 55720 33420 55800 33430
rect 55860 33420 55950 33430
rect 55960 33420 55990 33520
rect 55630 33250 55660 33420
rect 55800 33340 55810 33420
rect 55860 33250 55890 33420
rect 55950 33340 55990 33420
rect 55570 33240 55660 33250
rect 55720 33240 55800 33250
rect 55860 33240 55950 33250
rect 55960 33240 55990 33340
rect 55630 33070 55660 33240
rect 55800 33160 55810 33240
rect 55860 33070 55890 33240
rect 55950 33160 55990 33240
rect 55570 33060 55660 33070
rect 55720 33060 55800 33070
rect 55860 33060 55950 33070
rect 55960 33060 55990 33160
rect 55630 32890 55660 33060
rect 55800 32980 55810 33060
rect 55860 32890 55890 33060
rect 55950 32980 55990 33060
rect 55570 32880 55660 32890
rect 55720 32880 55800 32890
rect 55860 32880 55950 32890
rect 55960 32880 55990 32980
rect 55630 32710 55660 32880
rect 55800 32800 55810 32880
rect 55860 32710 55890 32880
rect 55950 32800 55990 32880
rect 55570 32700 55660 32710
rect 55720 32700 55800 32710
rect 55860 32700 55950 32710
rect 55960 32700 55990 32800
rect 55630 32530 55660 32700
rect 55800 32620 55810 32700
rect 55860 32530 55890 32700
rect 55950 32620 55990 32700
rect 55570 32520 55660 32530
rect 55720 32520 55800 32530
rect 55860 32520 55950 32530
rect 55960 32520 55990 32620
rect 55630 32350 55660 32520
rect 55800 32440 55810 32520
rect 55860 32350 55890 32520
rect 55950 32440 55990 32520
rect 55570 32340 55660 32350
rect 55720 32340 55800 32350
rect 55860 32340 55950 32350
rect 55960 32340 55990 32440
rect 55630 32170 55660 32340
rect 55800 32260 55810 32340
rect 55860 32170 55890 32340
rect 55950 32260 55990 32340
rect 55570 32160 55660 32170
rect 55720 32160 55800 32170
rect 55860 32160 55950 32170
rect 55960 32160 55990 32260
rect 55630 31990 55660 32160
rect 55800 32080 55810 32160
rect 55860 31990 55890 32160
rect 55950 32080 55990 32160
rect 55570 31980 55660 31990
rect 55720 31980 55800 31990
rect 55860 31980 55950 31990
rect 55960 31980 55990 32080
rect 55630 31810 55660 31980
rect 55800 31900 55810 31980
rect 55860 31810 55890 31980
rect 55950 31900 55990 31980
rect 55570 31800 55660 31810
rect 55720 31800 55800 31810
rect 55860 31800 55950 31810
rect 55960 31800 55990 31900
rect 55630 31630 55660 31800
rect 55800 31720 55810 31800
rect 55860 31630 55890 31800
rect 55950 31720 55990 31800
rect 55570 31620 55660 31630
rect 55720 31620 55800 31630
rect 55860 31620 55950 31630
rect 55960 31620 55990 31720
rect 55630 31450 55660 31620
rect 55800 31540 55810 31620
rect 55860 31450 55890 31620
rect 55950 31540 55990 31620
rect 55570 31440 55660 31450
rect 55720 31440 55800 31450
rect 55860 31440 55950 31450
rect 55960 31440 55990 31540
rect 55630 31270 55660 31440
rect 55800 31360 55810 31440
rect 55860 31270 55890 31440
rect 55950 31360 55990 31440
rect 55570 31260 55660 31270
rect 55720 31260 55800 31270
rect 55860 31260 55950 31270
rect 55960 31260 55990 31360
rect 55630 31100 55660 31260
rect 55800 31180 55810 31260
rect 55860 31100 55890 31260
rect 55950 31180 55990 31260
rect 55960 31100 55990 31180
rect 56090 31100 56100 37100
rect 56190 37020 56270 37030
rect 56510 37020 56590 37030
rect 56270 36940 56280 37020
rect 56590 36940 56600 37020
rect 56190 36840 56270 36850
rect 56510 36840 56590 36850
rect 56270 36760 56280 36840
rect 56590 36760 56600 36840
rect 56190 36660 56270 36670
rect 56510 36660 56590 36670
rect 56270 36580 56280 36660
rect 56590 36580 56600 36660
rect 56190 36480 56270 36490
rect 56510 36480 56590 36490
rect 56270 36400 56280 36480
rect 56590 36400 56600 36480
rect 56190 36300 56270 36310
rect 56510 36300 56590 36310
rect 56270 36220 56280 36300
rect 56590 36220 56600 36300
rect 56190 36120 56270 36130
rect 56510 36120 56590 36130
rect 56270 36040 56280 36120
rect 56590 36040 56600 36120
rect 56190 35940 56270 35950
rect 56510 35940 56590 35950
rect 56270 35860 56280 35940
rect 56590 35860 56600 35940
rect 56190 35760 56270 35770
rect 56510 35760 56590 35770
rect 56270 35680 56280 35760
rect 56590 35680 56600 35760
rect 56190 35580 56270 35590
rect 56510 35580 56590 35590
rect 56270 35500 56280 35580
rect 56590 35500 56600 35580
rect 56190 35400 56270 35410
rect 56510 35400 56590 35410
rect 56270 35320 56280 35400
rect 56590 35320 56600 35400
rect 56190 35220 56270 35230
rect 56510 35220 56590 35230
rect 56270 35140 56280 35220
rect 56590 35140 56600 35220
rect 56190 35040 56270 35050
rect 56510 35040 56590 35050
rect 56270 34960 56280 35040
rect 56590 34960 56600 35040
rect 56190 34860 56270 34870
rect 56510 34860 56590 34870
rect 56270 34780 56280 34860
rect 56590 34780 56600 34860
rect 56190 34680 56270 34690
rect 56510 34680 56590 34690
rect 56270 34600 56280 34680
rect 56590 34600 56600 34680
rect 56190 34500 56270 34510
rect 56510 34500 56590 34510
rect 56270 34420 56280 34500
rect 56590 34420 56600 34500
rect 56190 34320 56270 34330
rect 56510 34320 56590 34330
rect 56270 34240 56280 34320
rect 56590 34240 56600 34320
rect 56190 34140 56270 34150
rect 56510 34140 56590 34150
rect 56270 34060 56280 34140
rect 56590 34060 56600 34140
rect 56190 33960 56270 33970
rect 56510 33960 56590 33970
rect 56270 33880 56280 33960
rect 56590 33880 56600 33960
rect 56190 33780 56270 33790
rect 56510 33780 56590 33790
rect 56270 33700 56280 33780
rect 56590 33700 56600 33780
rect 56190 33600 56270 33610
rect 56510 33600 56590 33610
rect 56270 33520 56280 33600
rect 56590 33520 56600 33600
rect 56190 33420 56270 33430
rect 56510 33420 56590 33430
rect 56270 33340 56280 33420
rect 56590 33340 56600 33420
rect 56190 33240 56270 33250
rect 56510 33240 56590 33250
rect 56270 33160 56280 33240
rect 56590 33160 56600 33240
rect 56190 33060 56270 33070
rect 56510 33060 56590 33070
rect 56270 32980 56280 33060
rect 56590 32980 56600 33060
rect 56190 32880 56270 32890
rect 56510 32880 56590 32890
rect 56270 32800 56280 32880
rect 56590 32800 56600 32880
rect 56190 32700 56270 32710
rect 56510 32700 56590 32710
rect 56270 32620 56280 32700
rect 56590 32620 56600 32700
rect 56190 32520 56270 32530
rect 56510 32520 56590 32530
rect 56270 32440 56280 32520
rect 56590 32440 56600 32520
rect 56190 32340 56270 32350
rect 56510 32340 56590 32350
rect 56270 32260 56280 32340
rect 56590 32260 56600 32340
rect 56190 32160 56270 32170
rect 56510 32160 56590 32170
rect 56270 32080 56280 32160
rect 56590 32080 56600 32160
rect 56190 31980 56270 31990
rect 56510 31980 56590 31990
rect 56270 31900 56280 31980
rect 56590 31900 56600 31980
rect 56190 31800 56270 31810
rect 56510 31800 56590 31810
rect 56270 31720 56280 31800
rect 56590 31720 56600 31800
rect 56190 31620 56270 31630
rect 56510 31620 56590 31630
rect 56270 31540 56280 31620
rect 56590 31540 56600 31620
rect 56190 31440 56270 31450
rect 56510 31440 56590 31450
rect 56270 31360 56280 31440
rect 56590 31360 56600 31440
rect 56190 31260 56270 31270
rect 56510 31260 56590 31270
rect 56270 31180 56280 31260
rect 56590 31180 56600 31260
rect 56770 31100 56780 37100
rect 56790 31100 56820 37100
rect 56890 37030 56920 37100
rect 57120 37030 57150 37100
rect 56830 37020 56920 37030
rect 56980 37020 57060 37030
rect 57120 37020 57210 37030
rect 57220 37020 57250 37100
rect 56890 36850 56920 37020
rect 57060 36940 57070 37020
rect 57120 36850 57150 37020
rect 57210 36940 57250 37020
rect 56830 36840 56920 36850
rect 56980 36840 57060 36850
rect 57120 36840 57210 36850
rect 57220 36840 57250 36940
rect 56890 36670 56920 36840
rect 57060 36760 57070 36840
rect 57120 36670 57150 36840
rect 57210 36760 57250 36840
rect 56830 36660 56920 36670
rect 56980 36660 57060 36670
rect 57120 36660 57210 36670
rect 57220 36660 57250 36760
rect 56890 36490 56920 36660
rect 57060 36580 57070 36660
rect 57120 36490 57150 36660
rect 57210 36580 57250 36660
rect 56830 36480 56920 36490
rect 56980 36480 57060 36490
rect 57120 36480 57210 36490
rect 57220 36480 57250 36580
rect 56890 36310 56920 36480
rect 57060 36400 57070 36480
rect 57120 36310 57150 36480
rect 57210 36400 57250 36480
rect 56830 36300 56920 36310
rect 56980 36300 57060 36310
rect 57120 36300 57210 36310
rect 57220 36300 57250 36400
rect 56890 36130 56920 36300
rect 57060 36220 57070 36300
rect 57120 36130 57150 36300
rect 57210 36220 57250 36300
rect 56830 36120 56920 36130
rect 56980 36120 57060 36130
rect 57120 36120 57210 36130
rect 57220 36120 57250 36220
rect 56890 35950 56920 36120
rect 57060 36040 57070 36120
rect 57120 35950 57150 36120
rect 57210 36040 57250 36120
rect 56830 35940 56920 35950
rect 56980 35940 57060 35950
rect 57120 35940 57210 35950
rect 57220 35940 57250 36040
rect 56890 35770 56920 35940
rect 57060 35860 57070 35940
rect 57120 35770 57150 35940
rect 57210 35860 57250 35940
rect 56830 35760 56920 35770
rect 56980 35760 57060 35770
rect 57120 35760 57210 35770
rect 57220 35760 57250 35860
rect 56890 35590 56920 35760
rect 57060 35680 57070 35760
rect 57120 35590 57150 35760
rect 57210 35680 57250 35760
rect 56830 35580 56920 35590
rect 56980 35580 57060 35590
rect 57120 35580 57210 35590
rect 57220 35580 57250 35680
rect 56890 35410 56920 35580
rect 57060 35500 57070 35580
rect 57120 35410 57150 35580
rect 57210 35500 57250 35580
rect 56830 35400 56920 35410
rect 56980 35400 57060 35410
rect 57120 35400 57210 35410
rect 57220 35400 57250 35500
rect 56890 35230 56920 35400
rect 57060 35320 57070 35400
rect 57120 35230 57150 35400
rect 57210 35320 57250 35400
rect 56830 35220 56920 35230
rect 56980 35220 57060 35230
rect 57120 35220 57210 35230
rect 57220 35220 57250 35320
rect 56890 35050 56920 35220
rect 57060 35140 57070 35220
rect 57120 35050 57150 35220
rect 57210 35140 57250 35220
rect 56830 35040 56920 35050
rect 56980 35040 57060 35050
rect 57120 35040 57210 35050
rect 57220 35040 57250 35140
rect 56890 34870 56920 35040
rect 57060 34960 57070 35040
rect 57120 34870 57150 35040
rect 57210 34960 57250 35040
rect 56830 34860 56920 34870
rect 56980 34860 57060 34870
rect 57120 34860 57210 34870
rect 57220 34860 57250 34960
rect 56890 34690 56920 34860
rect 57060 34780 57070 34860
rect 57120 34690 57150 34860
rect 57210 34780 57250 34860
rect 56830 34680 56920 34690
rect 56980 34680 57060 34690
rect 57120 34680 57210 34690
rect 57220 34680 57250 34780
rect 56890 34510 56920 34680
rect 57060 34600 57070 34680
rect 57120 34510 57150 34680
rect 57210 34600 57250 34680
rect 56830 34500 56920 34510
rect 56980 34500 57060 34510
rect 57120 34500 57210 34510
rect 57220 34500 57250 34600
rect 56890 34330 56920 34500
rect 57060 34420 57070 34500
rect 57120 34330 57150 34500
rect 57210 34420 57250 34500
rect 56830 34320 56920 34330
rect 56980 34320 57060 34330
rect 57120 34320 57210 34330
rect 57220 34320 57250 34420
rect 56890 34150 56920 34320
rect 57060 34240 57070 34320
rect 57120 34150 57150 34320
rect 57210 34240 57250 34320
rect 56830 34140 56920 34150
rect 56980 34140 57060 34150
rect 57120 34140 57210 34150
rect 57220 34140 57250 34240
rect 56890 33970 56920 34140
rect 57060 34060 57070 34140
rect 57120 33970 57150 34140
rect 57210 34060 57250 34140
rect 56830 33960 56920 33970
rect 56980 33960 57060 33970
rect 57120 33960 57210 33970
rect 57220 33960 57250 34060
rect 56890 33790 56920 33960
rect 57060 33880 57070 33960
rect 57120 33790 57150 33960
rect 57210 33880 57250 33960
rect 56830 33780 56920 33790
rect 56980 33780 57060 33790
rect 57120 33780 57210 33790
rect 57220 33780 57250 33880
rect 56890 33610 56920 33780
rect 57060 33700 57070 33780
rect 57120 33610 57150 33780
rect 57210 33700 57250 33780
rect 56830 33600 56920 33610
rect 56980 33600 57060 33610
rect 57120 33600 57210 33610
rect 57220 33600 57250 33700
rect 56890 33430 56920 33600
rect 57060 33520 57070 33600
rect 57120 33430 57150 33600
rect 57210 33520 57250 33600
rect 56830 33420 56920 33430
rect 56980 33420 57060 33430
rect 57120 33420 57210 33430
rect 57220 33420 57250 33520
rect 56890 33250 56920 33420
rect 57060 33340 57070 33420
rect 57120 33250 57150 33420
rect 57210 33340 57250 33420
rect 56830 33240 56920 33250
rect 56980 33240 57060 33250
rect 57120 33240 57210 33250
rect 57220 33240 57250 33340
rect 56890 33070 56920 33240
rect 57060 33160 57070 33240
rect 57120 33070 57150 33240
rect 57210 33160 57250 33240
rect 56830 33060 56920 33070
rect 56980 33060 57060 33070
rect 57120 33060 57210 33070
rect 57220 33060 57250 33160
rect 56890 32890 56920 33060
rect 57060 32980 57070 33060
rect 57120 32890 57150 33060
rect 57210 32980 57250 33060
rect 56830 32880 56920 32890
rect 56980 32880 57060 32890
rect 57120 32880 57210 32890
rect 57220 32880 57250 32980
rect 56890 32710 56920 32880
rect 57060 32800 57070 32880
rect 57120 32710 57150 32880
rect 57210 32800 57250 32880
rect 56830 32700 56920 32710
rect 56980 32700 57060 32710
rect 57120 32700 57210 32710
rect 57220 32700 57250 32800
rect 56890 32530 56920 32700
rect 57060 32620 57070 32700
rect 57120 32530 57150 32700
rect 57210 32620 57250 32700
rect 56830 32520 56920 32530
rect 56980 32520 57060 32530
rect 57120 32520 57210 32530
rect 57220 32520 57250 32620
rect 56890 32350 56920 32520
rect 57060 32440 57070 32520
rect 57120 32350 57150 32520
rect 57210 32440 57250 32520
rect 56830 32340 56920 32350
rect 56980 32340 57060 32350
rect 57120 32340 57210 32350
rect 57220 32340 57250 32440
rect 56890 32170 56920 32340
rect 57060 32260 57070 32340
rect 57120 32170 57150 32340
rect 57210 32260 57250 32340
rect 56830 32160 56920 32170
rect 56980 32160 57060 32170
rect 57120 32160 57210 32170
rect 57220 32160 57250 32260
rect 56890 31990 56920 32160
rect 57060 32080 57070 32160
rect 57120 31990 57150 32160
rect 57210 32080 57250 32160
rect 56830 31980 56920 31990
rect 56980 31980 57060 31990
rect 57120 31980 57210 31990
rect 57220 31980 57250 32080
rect 56890 31810 56920 31980
rect 57060 31900 57070 31980
rect 57120 31810 57150 31980
rect 57210 31900 57250 31980
rect 56830 31800 56920 31810
rect 56980 31800 57060 31810
rect 57120 31800 57210 31810
rect 57220 31800 57250 31900
rect 56890 31630 56920 31800
rect 57060 31720 57070 31800
rect 57120 31630 57150 31800
rect 57210 31720 57250 31800
rect 56830 31620 56920 31630
rect 56980 31620 57060 31630
rect 57120 31620 57210 31630
rect 57220 31620 57250 31720
rect 56890 31450 56920 31620
rect 57060 31540 57070 31620
rect 57120 31450 57150 31620
rect 57210 31540 57250 31620
rect 56830 31440 56920 31450
rect 56980 31440 57060 31450
rect 57120 31440 57210 31450
rect 57220 31440 57250 31540
rect 56890 31270 56920 31440
rect 57060 31360 57070 31440
rect 57120 31270 57150 31440
rect 57210 31360 57250 31440
rect 56830 31260 56920 31270
rect 56980 31260 57060 31270
rect 57120 31260 57210 31270
rect 57220 31260 57250 31360
rect 56890 31100 56920 31260
rect 57060 31180 57070 31260
rect 57120 31100 57150 31260
rect 57210 31180 57250 31260
rect 57220 31100 57250 31180
rect 57350 31100 57360 37100
rect 57450 37020 57530 37030
rect 57770 37020 57850 37030
rect 57530 36940 57540 37020
rect 57850 36940 57860 37020
rect 57450 36840 57530 36850
rect 57770 36840 57850 36850
rect 57530 36760 57540 36840
rect 57850 36760 57860 36840
rect 57450 36660 57530 36670
rect 57770 36660 57850 36670
rect 57530 36580 57540 36660
rect 57850 36580 57860 36660
rect 57450 36480 57530 36490
rect 57770 36480 57850 36490
rect 57530 36400 57540 36480
rect 57850 36400 57860 36480
rect 57450 36300 57530 36310
rect 57770 36300 57850 36310
rect 57530 36220 57540 36300
rect 57850 36220 57860 36300
rect 57450 36120 57530 36130
rect 57770 36120 57850 36130
rect 57530 36040 57540 36120
rect 57850 36040 57860 36120
rect 57450 35940 57530 35950
rect 57770 35940 57850 35950
rect 57530 35860 57540 35940
rect 57850 35860 57860 35940
rect 57450 35760 57530 35770
rect 57770 35760 57850 35770
rect 57530 35680 57540 35760
rect 57850 35680 57860 35760
rect 57450 35580 57530 35590
rect 57770 35580 57850 35590
rect 57530 35500 57540 35580
rect 57850 35500 57860 35580
rect 57450 35400 57530 35410
rect 57770 35400 57850 35410
rect 57530 35320 57540 35400
rect 57850 35320 57860 35400
rect 57450 35220 57530 35230
rect 57770 35220 57850 35230
rect 57530 35140 57540 35220
rect 57850 35140 57860 35220
rect 57450 35040 57530 35050
rect 57770 35040 57850 35050
rect 57530 34960 57540 35040
rect 57850 34960 57860 35040
rect 57450 34860 57530 34870
rect 57770 34860 57850 34870
rect 57530 34780 57540 34860
rect 57850 34780 57860 34860
rect 57450 34680 57530 34690
rect 57770 34680 57850 34690
rect 57530 34600 57540 34680
rect 57850 34600 57860 34680
rect 57450 34500 57530 34510
rect 57770 34500 57850 34510
rect 57530 34420 57540 34500
rect 57850 34420 57860 34500
rect 57450 34320 57530 34330
rect 57770 34320 57850 34330
rect 57530 34240 57540 34320
rect 57850 34240 57860 34320
rect 57450 34140 57530 34150
rect 57770 34140 57850 34150
rect 57530 34060 57540 34140
rect 57850 34060 57860 34140
rect 57450 33960 57530 33970
rect 57770 33960 57850 33970
rect 57530 33880 57540 33960
rect 57850 33880 57860 33960
rect 57450 33780 57530 33790
rect 57770 33780 57850 33790
rect 57530 33700 57540 33780
rect 57850 33700 57860 33780
rect 57450 33600 57530 33610
rect 57770 33600 57850 33610
rect 57530 33520 57540 33600
rect 57850 33520 57860 33600
rect 57450 33420 57530 33430
rect 57770 33420 57850 33430
rect 57530 33340 57540 33420
rect 57850 33340 57860 33420
rect 57450 33240 57530 33250
rect 57770 33240 57850 33250
rect 57530 33160 57540 33240
rect 57850 33160 57860 33240
rect 57450 33060 57530 33070
rect 57770 33060 57850 33070
rect 57530 32980 57540 33060
rect 57850 32980 57860 33060
rect 57450 32880 57530 32890
rect 57770 32880 57850 32890
rect 57530 32800 57540 32880
rect 57850 32800 57860 32880
rect 57450 32700 57530 32710
rect 57770 32700 57850 32710
rect 57530 32620 57540 32700
rect 57850 32620 57860 32700
rect 57450 32520 57530 32530
rect 57770 32520 57850 32530
rect 57530 32440 57540 32520
rect 57850 32440 57860 32520
rect 57450 32340 57530 32350
rect 57770 32340 57850 32350
rect 57530 32260 57540 32340
rect 57850 32260 57860 32340
rect 57450 32160 57530 32170
rect 57770 32160 57850 32170
rect 57530 32080 57540 32160
rect 57850 32080 57860 32160
rect 57450 31980 57530 31990
rect 57770 31980 57850 31990
rect 57530 31900 57540 31980
rect 57850 31900 57860 31980
rect 57450 31800 57530 31810
rect 57770 31800 57850 31810
rect 57530 31720 57540 31800
rect 57850 31720 57860 31800
rect 57450 31620 57530 31630
rect 57770 31620 57850 31630
rect 57530 31540 57540 31620
rect 57850 31540 57860 31620
rect 57450 31440 57530 31450
rect 57770 31440 57850 31450
rect 57530 31360 57540 31440
rect 57850 31360 57860 31440
rect 57450 31260 57530 31270
rect 57770 31260 57850 31270
rect 57530 31180 57540 31260
rect 57850 31180 57860 31260
rect 58030 31100 58040 37100
rect 58050 31100 58080 37100
rect 58150 37030 58180 37100
rect 58380 37030 58410 37100
rect 58090 37020 58180 37030
rect 58240 37020 58320 37030
rect 58380 37020 58470 37030
rect 58480 37020 58510 37100
rect 58150 36850 58180 37020
rect 58320 36940 58330 37020
rect 58380 36850 58410 37020
rect 58470 36940 58510 37020
rect 58090 36840 58180 36850
rect 58240 36840 58320 36850
rect 58380 36840 58470 36850
rect 58480 36840 58510 36940
rect 58150 36670 58180 36840
rect 58320 36760 58330 36840
rect 58380 36670 58410 36840
rect 58470 36760 58510 36840
rect 58090 36660 58180 36670
rect 58240 36660 58320 36670
rect 58380 36660 58470 36670
rect 58480 36660 58510 36760
rect 58150 36490 58180 36660
rect 58320 36580 58330 36660
rect 58380 36490 58410 36660
rect 58470 36580 58510 36660
rect 58090 36480 58180 36490
rect 58240 36480 58320 36490
rect 58380 36480 58470 36490
rect 58480 36480 58510 36580
rect 58150 36310 58180 36480
rect 58320 36400 58330 36480
rect 58380 36310 58410 36480
rect 58470 36400 58510 36480
rect 58090 36300 58180 36310
rect 58240 36300 58320 36310
rect 58380 36300 58470 36310
rect 58480 36300 58510 36400
rect 58150 36130 58180 36300
rect 58320 36220 58330 36300
rect 58380 36130 58410 36300
rect 58470 36220 58510 36300
rect 58090 36120 58180 36130
rect 58240 36120 58320 36130
rect 58380 36120 58470 36130
rect 58480 36120 58510 36220
rect 58150 35950 58180 36120
rect 58320 36040 58330 36120
rect 58380 35950 58410 36120
rect 58470 36040 58510 36120
rect 58090 35940 58180 35950
rect 58240 35940 58320 35950
rect 58380 35940 58470 35950
rect 58480 35940 58510 36040
rect 58150 35770 58180 35940
rect 58320 35860 58330 35940
rect 58380 35770 58410 35940
rect 58470 35860 58510 35940
rect 58090 35760 58180 35770
rect 58240 35760 58320 35770
rect 58380 35760 58470 35770
rect 58480 35760 58510 35860
rect 58150 35590 58180 35760
rect 58320 35680 58330 35760
rect 58380 35590 58410 35760
rect 58470 35680 58510 35760
rect 58090 35580 58180 35590
rect 58240 35580 58320 35590
rect 58380 35580 58470 35590
rect 58480 35580 58510 35680
rect 58150 35410 58180 35580
rect 58320 35500 58330 35580
rect 58380 35410 58410 35580
rect 58470 35500 58510 35580
rect 58090 35400 58180 35410
rect 58240 35400 58320 35410
rect 58380 35400 58470 35410
rect 58480 35400 58510 35500
rect 58150 35230 58180 35400
rect 58320 35320 58330 35400
rect 58380 35230 58410 35400
rect 58470 35320 58510 35400
rect 58090 35220 58180 35230
rect 58240 35220 58320 35230
rect 58380 35220 58470 35230
rect 58480 35220 58510 35320
rect 58150 35050 58180 35220
rect 58320 35140 58330 35220
rect 58380 35050 58410 35220
rect 58470 35140 58510 35220
rect 58090 35040 58180 35050
rect 58240 35040 58320 35050
rect 58380 35040 58470 35050
rect 58480 35040 58510 35140
rect 58150 34870 58180 35040
rect 58320 34960 58330 35040
rect 58380 34870 58410 35040
rect 58470 34960 58510 35040
rect 58090 34860 58180 34870
rect 58240 34860 58320 34870
rect 58380 34860 58470 34870
rect 58480 34860 58510 34960
rect 58150 34690 58180 34860
rect 58320 34780 58330 34860
rect 58380 34690 58410 34860
rect 58470 34780 58510 34860
rect 58090 34680 58180 34690
rect 58240 34680 58320 34690
rect 58380 34680 58470 34690
rect 58480 34680 58510 34780
rect 58150 34510 58180 34680
rect 58320 34600 58330 34680
rect 58380 34510 58410 34680
rect 58470 34600 58510 34680
rect 58090 34500 58180 34510
rect 58240 34500 58320 34510
rect 58380 34500 58470 34510
rect 58480 34500 58510 34600
rect 58150 34330 58180 34500
rect 58320 34420 58330 34500
rect 58380 34330 58410 34500
rect 58470 34420 58510 34500
rect 58090 34320 58180 34330
rect 58240 34320 58320 34330
rect 58380 34320 58470 34330
rect 58480 34320 58510 34420
rect 58150 34150 58180 34320
rect 58320 34240 58330 34320
rect 58380 34150 58410 34320
rect 58470 34240 58510 34320
rect 58090 34140 58180 34150
rect 58240 34140 58320 34150
rect 58380 34140 58470 34150
rect 58480 34140 58510 34240
rect 58150 33970 58180 34140
rect 58320 34060 58330 34140
rect 58380 33970 58410 34140
rect 58470 34060 58510 34140
rect 58090 33960 58180 33970
rect 58240 33960 58320 33970
rect 58380 33960 58470 33970
rect 58480 33960 58510 34060
rect 58150 33790 58180 33960
rect 58320 33880 58330 33960
rect 58380 33790 58410 33960
rect 58470 33880 58510 33960
rect 58090 33780 58180 33790
rect 58240 33780 58320 33790
rect 58380 33780 58470 33790
rect 58480 33780 58510 33880
rect 58150 33610 58180 33780
rect 58320 33700 58330 33780
rect 58380 33610 58410 33780
rect 58470 33700 58510 33780
rect 58090 33600 58180 33610
rect 58240 33600 58320 33610
rect 58380 33600 58470 33610
rect 58480 33600 58510 33700
rect 58150 33430 58180 33600
rect 58320 33520 58330 33600
rect 58380 33430 58410 33600
rect 58470 33520 58510 33600
rect 58090 33420 58180 33430
rect 58240 33420 58320 33430
rect 58380 33420 58470 33430
rect 58480 33420 58510 33520
rect 58150 33250 58180 33420
rect 58320 33340 58330 33420
rect 58380 33250 58410 33420
rect 58470 33340 58510 33420
rect 58090 33240 58180 33250
rect 58240 33240 58320 33250
rect 58380 33240 58470 33250
rect 58480 33240 58510 33340
rect 58150 33070 58180 33240
rect 58320 33160 58330 33240
rect 58380 33070 58410 33240
rect 58470 33160 58510 33240
rect 58090 33060 58180 33070
rect 58240 33060 58320 33070
rect 58380 33060 58470 33070
rect 58480 33060 58510 33160
rect 58150 32890 58180 33060
rect 58320 32980 58330 33060
rect 58380 32890 58410 33060
rect 58470 32980 58510 33060
rect 58090 32880 58180 32890
rect 58240 32880 58320 32890
rect 58380 32880 58470 32890
rect 58480 32880 58510 32980
rect 58150 32710 58180 32880
rect 58320 32800 58330 32880
rect 58380 32710 58410 32880
rect 58470 32800 58510 32880
rect 58090 32700 58180 32710
rect 58240 32700 58320 32710
rect 58380 32700 58470 32710
rect 58480 32700 58510 32800
rect 58150 32530 58180 32700
rect 58320 32620 58330 32700
rect 58380 32530 58410 32700
rect 58470 32620 58510 32700
rect 58090 32520 58180 32530
rect 58240 32520 58320 32530
rect 58380 32520 58470 32530
rect 58480 32520 58510 32620
rect 58150 32350 58180 32520
rect 58320 32440 58330 32520
rect 58380 32350 58410 32520
rect 58470 32440 58510 32520
rect 58090 32340 58180 32350
rect 58240 32340 58320 32350
rect 58380 32340 58470 32350
rect 58480 32340 58510 32440
rect 58150 32170 58180 32340
rect 58320 32260 58330 32340
rect 58380 32170 58410 32340
rect 58470 32260 58510 32340
rect 58090 32160 58180 32170
rect 58240 32160 58320 32170
rect 58380 32160 58470 32170
rect 58480 32160 58510 32260
rect 58150 31990 58180 32160
rect 58320 32080 58330 32160
rect 58380 31990 58410 32160
rect 58470 32080 58510 32160
rect 58090 31980 58180 31990
rect 58240 31980 58320 31990
rect 58380 31980 58470 31990
rect 58480 31980 58510 32080
rect 58150 31810 58180 31980
rect 58320 31900 58330 31980
rect 58380 31810 58410 31980
rect 58470 31900 58510 31980
rect 58090 31800 58180 31810
rect 58240 31800 58320 31810
rect 58380 31800 58470 31810
rect 58480 31800 58510 31900
rect 58150 31630 58180 31800
rect 58320 31720 58330 31800
rect 58380 31630 58410 31800
rect 58470 31720 58510 31800
rect 58090 31620 58180 31630
rect 58240 31620 58320 31630
rect 58380 31620 58470 31630
rect 58480 31620 58510 31720
rect 58150 31450 58180 31620
rect 58320 31540 58330 31620
rect 58380 31450 58410 31620
rect 58470 31540 58510 31620
rect 58090 31440 58180 31450
rect 58240 31440 58320 31450
rect 58380 31440 58470 31450
rect 58480 31440 58510 31540
rect 58150 31270 58180 31440
rect 58320 31360 58330 31440
rect 58380 31270 58410 31440
rect 58470 31360 58510 31440
rect 58090 31260 58180 31270
rect 58240 31260 58320 31270
rect 58380 31260 58470 31270
rect 58480 31260 58510 31360
rect 58150 31100 58180 31260
rect 58320 31180 58330 31260
rect 58380 31100 58410 31260
rect 58470 31180 58510 31260
rect 58480 31100 58510 31180
rect 58610 31100 58620 37100
rect 58710 37020 58790 37030
rect 59030 37020 59110 37030
rect 58790 36940 58800 37020
rect 59110 36940 59120 37020
rect 58710 36840 58790 36850
rect 59030 36840 59110 36850
rect 58790 36760 58800 36840
rect 59110 36760 59120 36840
rect 58710 36660 58790 36670
rect 59030 36660 59110 36670
rect 58790 36580 58800 36660
rect 59110 36580 59120 36660
rect 58710 36480 58790 36490
rect 59030 36480 59110 36490
rect 58790 36400 58800 36480
rect 59110 36400 59120 36480
rect 58710 36300 58790 36310
rect 59030 36300 59110 36310
rect 58790 36220 58800 36300
rect 59110 36220 59120 36300
rect 58710 36120 58790 36130
rect 59030 36120 59110 36130
rect 58790 36040 58800 36120
rect 59110 36040 59120 36120
rect 58710 35940 58790 35950
rect 59030 35940 59110 35950
rect 58790 35860 58800 35940
rect 59110 35860 59120 35940
rect 58710 35760 58790 35770
rect 59030 35760 59110 35770
rect 58790 35680 58800 35760
rect 59110 35680 59120 35760
rect 58710 35580 58790 35590
rect 59030 35580 59110 35590
rect 58790 35500 58800 35580
rect 59110 35500 59120 35580
rect 58710 35400 58790 35410
rect 59030 35400 59110 35410
rect 58790 35320 58800 35400
rect 59110 35320 59120 35400
rect 58710 35220 58790 35230
rect 59030 35220 59110 35230
rect 58790 35140 58800 35220
rect 59110 35140 59120 35220
rect 58710 35040 58790 35050
rect 59030 35040 59110 35050
rect 58790 34960 58800 35040
rect 59110 34960 59120 35040
rect 58710 34860 58790 34870
rect 59030 34860 59110 34870
rect 58790 34780 58800 34860
rect 59110 34780 59120 34860
rect 58710 34680 58790 34690
rect 59030 34680 59110 34690
rect 58790 34600 58800 34680
rect 59110 34600 59120 34680
rect 58710 34500 58790 34510
rect 59030 34500 59110 34510
rect 58790 34420 58800 34500
rect 59110 34420 59120 34500
rect 58710 34320 58790 34330
rect 59030 34320 59110 34330
rect 58790 34240 58800 34320
rect 59110 34240 59120 34320
rect 58710 34140 58790 34150
rect 59030 34140 59110 34150
rect 58790 34060 58800 34140
rect 59110 34060 59120 34140
rect 58710 33960 58790 33970
rect 59030 33960 59110 33970
rect 58790 33880 58800 33960
rect 59110 33880 59120 33960
rect 58710 33780 58790 33790
rect 59030 33780 59110 33790
rect 58790 33700 58800 33780
rect 59110 33700 59120 33780
rect 58710 33600 58790 33610
rect 59030 33600 59110 33610
rect 58790 33520 58800 33600
rect 59110 33520 59120 33600
rect 58710 33420 58790 33430
rect 59030 33420 59110 33430
rect 58790 33340 58800 33420
rect 59110 33340 59120 33420
rect 58710 33240 58790 33250
rect 59030 33240 59110 33250
rect 58790 33160 58800 33240
rect 59110 33160 59120 33240
rect 58710 33060 58790 33070
rect 59030 33060 59110 33070
rect 58790 32980 58800 33060
rect 59110 32980 59120 33060
rect 58710 32880 58790 32890
rect 59030 32880 59110 32890
rect 58790 32800 58800 32880
rect 59110 32800 59120 32880
rect 58710 32700 58790 32710
rect 59030 32700 59110 32710
rect 58790 32620 58800 32700
rect 59110 32620 59120 32700
rect 58710 32520 58790 32530
rect 59030 32520 59110 32530
rect 58790 32440 58800 32520
rect 59110 32440 59120 32520
rect 58710 32340 58790 32350
rect 59030 32340 59110 32350
rect 58790 32260 58800 32340
rect 59110 32260 59120 32340
rect 58710 32160 58790 32170
rect 59030 32160 59110 32170
rect 58790 32080 58800 32160
rect 59110 32080 59120 32160
rect 58710 31980 58790 31990
rect 59030 31980 59110 31990
rect 58790 31900 58800 31980
rect 59110 31900 59120 31980
rect 58710 31800 58790 31810
rect 59030 31800 59110 31810
rect 58790 31720 58800 31800
rect 59110 31720 59120 31800
rect 58710 31620 58790 31630
rect 59030 31620 59110 31630
rect 58790 31540 58800 31620
rect 59110 31540 59120 31620
rect 58710 31440 58790 31450
rect 59030 31440 59110 31450
rect 58790 31360 58800 31440
rect 59110 31360 59120 31440
rect 58710 31260 58790 31270
rect 59030 31260 59110 31270
rect 58790 31180 58800 31260
rect 59110 31180 59120 31260
rect 59290 31100 59300 37100
rect 59310 31100 59340 37100
rect 59410 37030 59440 37100
rect 59670 37030 59760 37100
rect 60660 37080 60670 37160
rect 60980 37080 60990 37160
rect 61400 37080 61410 37160
rect 61720 37080 61730 37160
rect 62140 37120 62150 37200
rect 62290 37120 62300 37200
rect 62740 37100 68950 37190
rect 63060 37030 63090 37100
rect 59350 37020 59440 37030
rect 59500 37020 59580 37030
rect 59650 37020 59760 37030
rect 60060 37020 60140 37030
rect 60210 37020 60290 37030
rect 60360 37020 60440 37030
rect 62060 37020 62140 37030
rect 62210 37020 62290 37030
rect 62770 37020 62850 37030
rect 62920 37020 63000 37030
rect 63060 37020 63150 37030
rect 63160 37020 63190 37100
rect 59410 36850 59440 37020
rect 59580 36940 59590 37020
rect 59670 36850 59760 37020
rect 60140 36940 60150 37020
rect 60290 36940 60300 37020
rect 60440 36940 60450 37020
rect 60740 37000 60820 37010
rect 61060 37000 61140 37010
rect 61480 37000 61560 37010
rect 61800 37000 61880 37010
rect 60820 36920 60830 37000
rect 61140 36920 61150 37000
rect 61560 36920 61570 37000
rect 61880 36920 61890 37000
rect 62140 36940 62150 37020
rect 62290 36940 62300 37020
rect 62850 36940 62860 37020
rect 63000 36940 63010 37020
rect 63060 36850 63090 37020
rect 63150 36940 63190 37020
rect 59350 36840 59440 36850
rect 59500 36840 59580 36850
rect 59650 36840 59760 36850
rect 60060 36840 60140 36850
rect 60210 36840 60290 36850
rect 60360 36840 60440 36850
rect 60580 36840 60660 36850
rect 60900 36840 60980 36850
rect 61320 36840 61400 36850
rect 61640 36840 61720 36850
rect 62060 36840 62140 36850
rect 62210 36840 62290 36850
rect 62770 36840 62850 36850
rect 62920 36840 63000 36850
rect 63060 36840 63150 36850
rect 63160 36840 63190 36940
rect 59410 36670 59440 36840
rect 59580 36760 59590 36840
rect 59670 36670 59760 36840
rect 60140 36760 60150 36840
rect 60290 36760 60300 36840
rect 60440 36760 60450 36840
rect 60660 36760 60670 36840
rect 60980 36760 60990 36840
rect 61400 36760 61410 36840
rect 61720 36760 61730 36840
rect 62140 36760 62150 36840
rect 62290 36760 62300 36840
rect 62850 36760 62860 36840
rect 63000 36760 63010 36840
rect 60740 36680 60820 36690
rect 61060 36680 61140 36690
rect 61480 36680 61560 36690
rect 61800 36680 61880 36690
rect 59350 36660 59440 36670
rect 59500 36660 59580 36670
rect 59650 36660 59760 36670
rect 60060 36660 60140 36670
rect 60210 36660 60290 36670
rect 60360 36660 60440 36670
rect 59410 36490 59440 36660
rect 59580 36580 59590 36660
rect 59670 36490 59760 36660
rect 60140 36580 60150 36660
rect 60290 36580 60300 36660
rect 60440 36580 60450 36660
rect 60820 36600 60830 36680
rect 61140 36600 61150 36680
rect 61560 36600 61570 36680
rect 61880 36600 61890 36680
rect 63060 36670 63090 36840
rect 63150 36760 63190 36840
rect 62060 36660 62140 36670
rect 62210 36660 62290 36670
rect 62770 36660 62850 36670
rect 62920 36660 63000 36670
rect 63060 36660 63150 36670
rect 63160 36660 63190 36760
rect 62140 36580 62150 36660
rect 62290 36580 62300 36660
rect 62850 36580 62860 36660
rect 63000 36580 63010 36660
rect 60580 36520 60660 36530
rect 60900 36520 60980 36530
rect 61320 36520 61400 36530
rect 61640 36520 61720 36530
rect 59350 36480 59440 36490
rect 59500 36480 59580 36490
rect 59650 36480 59760 36490
rect 60060 36480 60140 36490
rect 60210 36480 60290 36490
rect 60360 36480 60440 36490
rect 59410 36310 59440 36480
rect 59580 36400 59590 36480
rect 59670 36310 59760 36480
rect 60140 36400 60150 36480
rect 60290 36400 60300 36480
rect 60440 36400 60450 36480
rect 60660 36440 60670 36520
rect 60980 36440 60990 36520
rect 61400 36440 61410 36520
rect 61720 36440 61730 36520
rect 63060 36490 63090 36660
rect 63150 36580 63190 36660
rect 62060 36480 62140 36490
rect 62210 36480 62290 36490
rect 62770 36480 62850 36490
rect 62920 36480 63000 36490
rect 63060 36480 63150 36490
rect 63160 36480 63190 36580
rect 62140 36400 62150 36480
rect 62290 36400 62300 36480
rect 62850 36400 62860 36480
rect 63000 36400 63010 36480
rect 60740 36360 60820 36370
rect 61060 36360 61140 36370
rect 61480 36360 61560 36370
rect 61800 36360 61880 36370
rect 59350 36300 59440 36310
rect 59500 36300 59580 36310
rect 59650 36300 59760 36310
rect 60060 36300 60140 36310
rect 60210 36300 60290 36310
rect 60360 36300 60440 36310
rect 59410 36130 59440 36300
rect 59580 36220 59590 36300
rect 59670 36130 59760 36300
rect 60140 36220 60150 36300
rect 60290 36220 60300 36300
rect 60440 36220 60450 36300
rect 60820 36280 60830 36360
rect 61140 36280 61150 36360
rect 61560 36280 61570 36360
rect 61880 36280 61890 36360
rect 63060 36310 63090 36480
rect 63150 36400 63190 36480
rect 62060 36300 62140 36310
rect 62210 36300 62290 36310
rect 62770 36300 62850 36310
rect 62920 36300 63000 36310
rect 63060 36300 63150 36310
rect 63160 36300 63190 36400
rect 62140 36220 62150 36300
rect 62290 36220 62300 36300
rect 62850 36220 62860 36300
rect 63000 36220 63010 36300
rect 60580 36200 60660 36210
rect 60900 36200 60980 36210
rect 61320 36200 61400 36210
rect 61640 36200 61720 36210
rect 59350 36120 59440 36130
rect 59500 36120 59580 36130
rect 59650 36120 59760 36130
rect 60060 36120 60140 36130
rect 60210 36120 60290 36130
rect 60360 36120 60440 36130
rect 60660 36120 60670 36200
rect 60980 36120 60990 36200
rect 61400 36120 61410 36200
rect 61720 36120 61730 36200
rect 63060 36130 63090 36300
rect 63150 36220 63190 36300
rect 62060 36120 62140 36130
rect 62210 36120 62290 36130
rect 62770 36120 62850 36130
rect 62920 36120 63000 36130
rect 63060 36120 63150 36130
rect 63160 36120 63190 36220
rect 59410 35950 59440 36120
rect 59580 36040 59590 36120
rect 59670 35950 59760 36120
rect 60140 36040 60150 36120
rect 60290 36040 60300 36120
rect 60440 36040 60450 36120
rect 60740 36040 60820 36050
rect 61060 36040 61140 36050
rect 61480 36040 61560 36050
rect 61800 36040 61880 36050
rect 62140 36040 62150 36120
rect 62290 36040 62300 36120
rect 62850 36040 62860 36120
rect 63000 36040 63010 36120
rect 60820 35960 60830 36040
rect 61140 35960 61150 36040
rect 61560 35960 61570 36040
rect 61880 35960 61890 36040
rect 63060 36000 63090 36120
rect 63150 36040 63190 36120
rect 63160 36000 63190 36040
rect 63290 36000 63300 37100
rect 63390 37020 63470 37030
rect 63710 37020 63790 37030
rect 63470 36940 63480 37020
rect 63790 36940 63800 37020
rect 63390 36840 63470 36850
rect 63710 36840 63790 36850
rect 63470 36760 63480 36840
rect 63790 36760 63800 36840
rect 63390 36660 63470 36670
rect 63710 36660 63790 36670
rect 63470 36580 63480 36660
rect 63790 36580 63800 36660
rect 63390 36480 63470 36490
rect 63710 36480 63790 36490
rect 63470 36400 63480 36480
rect 63790 36400 63800 36480
rect 63390 36300 63470 36310
rect 63710 36300 63790 36310
rect 63470 36220 63480 36300
rect 63790 36220 63800 36300
rect 63390 36120 63470 36130
rect 63710 36120 63790 36130
rect 63470 36040 63480 36120
rect 63790 36040 63800 36120
rect 63970 36000 63980 37100
rect 63990 36000 64020 37100
rect 64090 37030 64120 37100
rect 64320 37030 64350 37100
rect 64030 37020 64120 37030
rect 64180 37020 64260 37030
rect 64320 37020 64410 37030
rect 64420 37020 64450 37100
rect 64090 36850 64120 37020
rect 64260 36940 64270 37020
rect 64320 36850 64350 37020
rect 64410 36940 64450 37020
rect 64030 36840 64120 36850
rect 64180 36840 64260 36850
rect 64320 36840 64410 36850
rect 64420 36840 64450 36940
rect 64090 36670 64120 36840
rect 64260 36760 64270 36840
rect 64320 36670 64350 36840
rect 64410 36760 64450 36840
rect 64030 36660 64120 36670
rect 64180 36660 64260 36670
rect 64320 36660 64410 36670
rect 64420 36660 64450 36760
rect 64090 36490 64120 36660
rect 64260 36580 64270 36660
rect 64320 36490 64350 36660
rect 64410 36580 64450 36660
rect 64030 36480 64120 36490
rect 64180 36480 64260 36490
rect 64320 36480 64410 36490
rect 64420 36480 64450 36580
rect 64090 36310 64120 36480
rect 64260 36400 64270 36480
rect 64320 36310 64350 36480
rect 64410 36400 64450 36480
rect 64030 36300 64120 36310
rect 64180 36300 64260 36310
rect 64320 36300 64410 36310
rect 64420 36300 64450 36400
rect 64090 36130 64120 36300
rect 64260 36220 64270 36300
rect 64320 36130 64350 36300
rect 64410 36220 64450 36300
rect 64030 36120 64120 36130
rect 64180 36120 64260 36130
rect 64320 36120 64410 36130
rect 64420 36120 64450 36220
rect 64090 36000 64120 36120
rect 64260 36040 64270 36120
rect 64320 36000 64350 36120
rect 64410 36040 64450 36120
rect 64420 36000 64450 36040
rect 64550 36000 64560 37100
rect 64650 37020 64730 37030
rect 64970 37020 65050 37030
rect 64730 36940 64740 37020
rect 65050 36940 65060 37020
rect 64650 36840 64730 36850
rect 64970 36840 65050 36850
rect 64730 36760 64740 36840
rect 65050 36760 65060 36840
rect 64650 36660 64730 36670
rect 64970 36660 65050 36670
rect 64730 36580 64740 36660
rect 65050 36580 65060 36660
rect 64650 36480 64730 36490
rect 64970 36480 65050 36490
rect 64730 36400 64740 36480
rect 65050 36400 65060 36480
rect 64650 36300 64730 36310
rect 64970 36300 65050 36310
rect 64730 36220 64740 36300
rect 65050 36220 65060 36300
rect 64650 36120 64730 36130
rect 64970 36120 65050 36130
rect 64730 36040 64740 36120
rect 65050 36040 65060 36120
rect 65230 36000 65240 37100
rect 65250 36000 65280 37100
rect 65350 37030 65380 37100
rect 65580 37030 65610 37100
rect 65290 37020 65380 37030
rect 65440 37020 65520 37030
rect 65580 37020 65670 37030
rect 65680 37020 65710 37100
rect 65350 36850 65380 37020
rect 65520 36940 65530 37020
rect 65580 36850 65610 37020
rect 65670 36940 65710 37020
rect 65290 36840 65380 36850
rect 65440 36840 65520 36850
rect 65580 36840 65670 36850
rect 65680 36840 65710 36940
rect 65350 36670 65380 36840
rect 65520 36760 65530 36840
rect 65580 36670 65610 36840
rect 65670 36760 65710 36840
rect 65290 36660 65380 36670
rect 65440 36660 65520 36670
rect 65580 36660 65670 36670
rect 65680 36660 65710 36760
rect 65350 36490 65380 36660
rect 65520 36580 65530 36660
rect 65580 36490 65610 36660
rect 65670 36580 65710 36660
rect 65290 36480 65380 36490
rect 65440 36480 65520 36490
rect 65580 36480 65670 36490
rect 65680 36480 65710 36580
rect 65350 36310 65380 36480
rect 65520 36400 65530 36480
rect 65580 36310 65610 36480
rect 65670 36400 65710 36480
rect 65290 36300 65380 36310
rect 65440 36300 65520 36310
rect 65580 36300 65670 36310
rect 65680 36300 65710 36400
rect 65350 36130 65380 36300
rect 65520 36220 65530 36300
rect 65580 36130 65610 36300
rect 65670 36220 65710 36300
rect 65290 36120 65380 36130
rect 65440 36120 65520 36130
rect 65580 36120 65670 36130
rect 65680 36120 65710 36220
rect 65350 36000 65380 36120
rect 65520 36040 65530 36120
rect 65580 36000 65610 36120
rect 65670 36040 65710 36120
rect 65680 36000 65710 36040
rect 65810 36000 65820 37100
rect 65910 37020 65990 37030
rect 66230 37020 66310 37030
rect 65990 36940 66000 37020
rect 66310 36940 66320 37020
rect 65910 36840 65990 36850
rect 66230 36840 66310 36850
rect 65990 36760 66000 36840
rect 66310 36760 66320 36840
rect 65910 36660 65990 36670
rect 66230 36660 66310 36670
rect 65990 36580 66000 36660
rect 66310 36580 66320 36660
rect 65910 36480 65990 36490
rect 66230 36480 66310 36490
rect 65990 36400 66000 36480
rect 66310 36400 66320 36480
rect 65910 36300 65990 36310
rect 66230 36300 66310 36310
rect 65990 36220 66000 36300
rect 66310 36220 66320 36300
rect 65910 36120 65990 36130
rect 66230 36120 66310 36130
rect 65990 36040 66000 36120
rect 66310 36040 66320 36120
rect 66490 36000 66500 37100
rect 66510 36000 66540 37100
rect 66610 37030 66640 37100
rect 66840 37030 66870 37100
rect 66550 37020 66640 37030
rect 66700 37020 66780 37030
rect 66840 37020 66930 37030
rect 66940 37020 66970 37100
rect 66610 36850 66640 37020
rect 66780 36940 66790 37020
rect 66840 36850 66870 37020
rect 66930 36940 66970 37020
rect 66550 36840 66640 36850
rect 66700 36840 66780 36850
rect 66840 36840 66930 36850
rect 66940 36840 66970 36940
rect 66610 36670 66640 36840
rect 66780 36760 66790 36840
rect 66840 36670 66870 36840
rect 66930 36760 66970 36840
rect 66550 36660 66640 36670
rect 66700 36660 66780 36670
rect 66840 36660 66930 36670
rect 66940 36660 66970 36760
rect 66610 36490 66640 36660
rect 66780 36580 66790 36660
rect 66840 36490 66870 36660
rect 66930 36580 66970 36660
rect 66550 36480 66640 36490
rect 66700 36480 66780 36490
rect 66840 36480 66930 36490
rect 66940 36480 66970 36580
rect 66610 36310 66640 36480
rect 66780 36400 66790 36480
rect 66840 36310 66870 36480
rect 66930 36400 66970 36480
rect 66550 36300 66640 36310
rect 66700 36300 66780 36310
rect 66840 36300 66930 36310
rect 66940 36300 66970 36400
rect 66610 36130 66640 36300
rect 66780 36220 66790 36300
rect 66840 36130 66870 36300
rect 66930 36220 66970 36300
rect 66550 36120 66640 36130
rect 66700 36120 66780 36130
rect 66840 36120 66930 36130
rect 66940 36120 66970 36220
rect 66610 36000 66640 36120
rect 66780 36040 66790 36120
rect 66840 36000 66870 36120
rect 66930 36040 66970 36120
rect 66940 36000 66970 36040
rect 67070 36000 67080 37100
rect 67170 37020 67250 37030
rect 67490 37020 67570 37030
rect 67250 36940 67260 37020
rect 67570 36940 67580 37020
rect 67170 36840 67250 36850
rect 67490 36840 67570 36850
rect 67250 36760 67260 36840
rect 67570 36760 67580 36840
rect 67170 36660 67250 36670
rect 67490 36660 67570 36670
rect 67250 36580 67260 36660
rect 67570 36580 67580 36660
rect 67170 36480 67250 36490
rect 67490 36480 67570 36490
rect 67250 36400 67260 36480
rect 67570 36400 67580 36480
rect 67170 36300 67250 36310
rect 67490 36300 67570 36310
rect 67250 36220 67260 36300
rect 67570 36220 67580 36300
rect 67170 36120 67250 36130
rect 67490 36120 67570 36130
rect 67250 36040 67260 36120
rect 67570 36040 67580 36120
rect 67750 36000 67760 37100
rect 67770 36000 67800 37100
rect 67870 37030 67900 37100
rect 68100 37030 68130 37100
rect 67810 37020 67900 37030
rect 67960 37020 68040 37030
rect 68100 37020 68190 37030
rect 68200 37020 68230 37100
rect 67870 36850 67900 37020
rect 68040 36940 68050 37020
rect 68100 36850 68130 37020
rect 68190 36940 68230 37020
rect 67810 36840 67900 36850
rect 67960 36840 68040 36850
rect 68100 36840 68190 36850
rect 68200 36840 68230 36940
rect 67870 36670 67900 36840
rect 68040 36760 68050 36840
rect 68100 36670 68130 36840
rect 68190 36760 68230 36840
rect 67810 36660 67900 36670
rect 67960 36660 68040 36670
rect 68100 36660 68190 36670
rect 68200 36660 68230 36760
rect 67870 36490 67900 36660
rect 68040 36580 68050 36660
rect 68100 36490 68130 36660
rect 68190 36580 68230 36660
rect 67810 36480 67900 36490
rect 67960 36480 68040 36490
rect 68100 36480 68190 36490
rect 68200 36480 68230 36580
rect 67870 36310 67900 36480
rect 68040 36400 68050 36480
rect 68100 36310 68130 36480
rect 68190 36400 68230 36480
rect 67810 36300 67900 36310
rect 67960 36300 68040 36310
rect 68100 36300 68190 36310
rect 68200 36300 68230 36400
rect 67870 36130 67900 36300
rect 68040 36220 68050 36300
rect 68100 36130 68130 36300
rect 68190 36220 68230 36300
rect 67810 36120 67900 36130
rect 67960 36120 68040 36130
rect 68100 36120 68190 36130
rect 68200 36120 68230 36220
rect 67870 36000 67900 36120
rect 68040 36040 68050 36120
rect 68100 36000 68130 36120
rect 68190 36040 68230 36120
rect 68200 36000 68230 36040
rect 68330 36000 68340 37100
rect 68430 37020 68510 37030
rect 68750 37020 68830 37030
rect 68510 36940 68520 37020
rect 68830 36940 68840 37020
rect 68430 36840 68510 36850
rect 68750 36840 68830 36850
rect 68510 36760 68520 36840
rect 68830 36760 68840 36840
rect 68430 36660 68510 36670
rect 68750 36660 68830 36670
rect 68510 36580 68520 36660
rect 68830 36580 68840 36660
rect 68430 36480 68510 36490
rect 68750 36480 68830 36490
rect 68510 36400 68520 36480
rect 68830 36400 68840 36480
rect 68430 36300 68510 36310
rect 68750 36300 68830 36310
rect 68510 36220 68520 36300
rect 68830 36220 68840 36300
rect 68430 36120 68510 36130
rect 68750 36120 68830 36130
rect 68510 36040 68520 36120
rect 68830 36040 68840 36120
rect 59350 35940 59440 35950
rect 59500 35940 59580 35950
rect 59650 35940 59760 35950
rect 60060 35940 60140 35950
rect 60210 35940 60290 35950
rect 60360 35940 60440 35950
rect 62060 35940 62140 35950
rect 62210 35940 62290 35950
rect 59410 35770 59440 35940
rect 59580 35860 59590 35940
rect 59670 35770 59760 35940
rect 60140 35860 60150 35940
rect 60290 35860 60300 35940
rect 60440 35860 60450 35940
rect 60580 35880 60660 35890
rect 60900 35880 60980 35890
rect 61320 35880 61400 35890
rect 61640 35880 61720 35890
rect 60660 35800 60670 35880
rect 60980 35800 60990 35880
rect 61400 35800 61410 35880
rect 61720 35800 61730 35880
rect 62140 35860 62150 35940
rect 62290 35860 62300 35940
rect 59350 35760 59440 35770
rect 59500 35760 59580 35770
rect 59650 35760 59760 35770
rect 60060 35760 60140 35770
rect 60210 35760 60290 35770
rect 60360 35760 60440 35770
rect 62060 35760 62140 35770
rect 62210 35760 62290 35770
rect 59410 35590 59440 35760
rect 59580 35680 59590 35760
rect 59670 35590 59760 35760
rect 60140 35680 60150 35760
rect 60290 35680 60300 35760
rect 60440 35680 60450 35760
rect 60740 35720 60820 35730
rect 61060 35720 61140 35730
rect 61480 35720 61560 35730
rect 61800 35720 61880 35730
rect 60820 35640 60830 35720
rect 61140 35640 61150 35720
rect 61560 35640 61570 35720
rect 61880 35640 61890 35720
rect 62140 35680 62150 35760
rect 62290 35680 62300 35760
rect 59350 35580 59440 35590
rect 59500 35580 59580 35590
rect 59650 35580 59760 35590
rect 60060 35580 60140 35590
rect 60210 35580 60290 35590
rect 60360 35580 60440 35590
rect 62060 35580 62140 35590
rect 62210 35580 62290 35590
rect 59410 35410 59440 35580
rect 59580 35500 59590 35580
rect 59670 35410 59760 35580
rect 60140 35500 60150 35580
rect 60290 35500 60300 35580
rect 60440 35500 60450 35580
rect 60580 35560 60660 35570
rect 60900 35560 60980 35570
rect 61320 35560 61400 35570
rect 61640 35560 61720 35570
rect 60660 35480 60670 35560
rect 60980 35480 60990 35560
rect 61400 35480 61410 35560
rect 61720 35480 61730 35560
rect 62140 35500 62150 35580
rect 62290 35500 62300 35580
rect 59350 35400 59440 35410
rect 59500 35400 59580 35410
rect 59650 35400 59760 35410
rect 60060 35400 60140 35410
rect 60210 35400 60290 35410
rect 60360 35400 60440 35410
rect 60740 35400 60820 35410
rect 61060 35400 61140 35410
rect 61480 35400 61560 35410
rect 61800 35400 61880 35410
rect 62060 35400 62140 35410
rect 62210 35400 62290 35410
rect 59410 35230 59440 35400
rect 59580 35320 59590 35400
rect 59670 35230 59760 35400
rect 60140 35320 60150 35400
rect 60290 35320 60300 35400
rect 60440 35320 60450 35400
rect 60820 35320 60830 35400
rect 61140 35320 61150 35400
rect 61560 35320 61570 35400
rect 61880 35320 61890 35400
rect 62140 35320 62150 35400
rect 62290 35320 62300 35400
rect 60580 35240 60660 35250
rect 60900 35240 60980 35250
rect 61320 35240 61400 35250
rect 61640 35240 61720 35250
rect 59350 35220 59440 35230
rect 59500 35220 59580 35230
rect 59650 35220 59760 35230
rect 60060 35220 60140 35230
rect 60210 35220 60290 35230
rect 60360 35220 60440 35230
rect 59410 35050 59440 35220
rect 59580 35140 59590 35220
rect 59670 35050 59760 35220
rect 60140 35140 60150 35220
rect 60290 35140 60300 35220
rect 60440 35140 60450 35220
rect 60660 35160 60670 35240
rect 60980 35160 60990 35240
rect 61400 35160 61410 35240
rect 61720 35160 61730 35240
rect 62060 35220 62140 35230
rect 62210 35220 62290 35230
rect 62140 35140 62150 35220
rect 62290 35140 62300 35220
rect 60740 35080 60820 35090
rect 61060 35080 61140 35090
rect 61480 35080 61560 35090
rect 61800 35080 61880 35090
rect 59350 35040 59440 35050
rect 59500 35040 59580 35050
rect 59650 35040 59760 35050
rect 60060 35040 60140 35050
rect 60210 35040 60290 35050
rect 60360 35040 60440 35050
rect 59410 34870 59440 35040
rect 59580 34960 59590 35040
rect 59670 34870 59760 35040
rect 60140 34960 60150 35040
rect 60290 34960 60300 35040
rect 60440 34960 60450 35040
rect 60820 35000 60830 35080
rect 61140 35000 61150 35080
rect 61560 35000 61570 35080
rect 61880 35000 61890 35080
rect 62060 35040 62140 35050
rect 62210 35040 62290 35050
rect 62140 34960 62150 35040
rect 62290 34960 62300 35040
rect 60580 34920 60660 34930
rect 60900 34920 60980 34930
rect 61320 34920 61400 34930
rect 61640 34920 61720 34930
rect 59350 34860 59440 34870
rect 59500 34860 59580 34870
rect 59650 34860 59760 34870
rect 60060 34860 60140 34870
rect 60210 34860 60290 34870
rect 60360 34860 60440 34870
rect 59410 34690 59440 34860
rect 59580 34780 59590 34860
rect 59670 34690 59760 34860
rect 60140 34780 60150 34860
rect 60290 34780 60300 34860
rect 60440 34780 60450 34860
rect 60660 34840 60670 34920
rect 60980 34840 60990 34920
rect 61400 34840 61410 34920
rect 61720 34840 61730 34920
rect 62060 34860 62140 34870
rect 62210 34860 62290 34870
rect 62140 34780 62150 34860
rect 62290 34780 62300 34860
rect 60740 34760 60820 34770
rect 61060 34760 61140 34770
rect 61480 34760 61560 34770
rect 61800 34760 61880 34770
rect 59350 34680 59440 34690
rect 59500 34680 59580 34690
rect 59650 34680 59760 34690
rect 60060 34680 60140 34690
rect 60210 34680 60290 34690
rect 60360 34680 60440 34690
rect 60820 34680 60830 34760
rect 61140 34680 61150 34760
rect 61560 34680 61570 34760
rect 61880 34680 61890 34760
rect 62060 34680 62140 34690
rect 62210 34680 62290 34690
rect 59410 34510 59440 34680
rect 59580 34600 59590 34680
rect 59670 34510 59760 34680
rect 60140 34600 60150 34680
rect 60290 34600 60300 34680
rect 60440 34600 60450 34680
rect 60580 34600 60660 34610
rect 60900 34600 60980 34610
rect 61320 34600 61400 34610
rect 61640 34600 61720 34610
rect 62140 34600 62150 34680
rect 62290 34600 62300 34680
rect 60660 34520 60670 34600
rect 60980 34520 60990 34600
rect 61400 34520 61410 34600
rect 61720 34520 61730 34600
rect 59350 34500 59440 34510
rect 59500 34500 59580 34510
rect 59650 34500 59760 34510
rect 60060 34500 60140 34510
rect 60210 34500 60290 34510
rect 60360 34500 60440 34510
rect 62060 34500 62140 34510
rect 62210 34500 62290 34510
rect 59410 34330 59440 34500
rect 59580 34420 59590 34500
rect 59670 34330 59760 34500
rect 60140 34420 60150 34500
rect 60290 34420 60300 34500
rect 60440 34420 60450 34500
rect 60740 34440 60820 34450
rect 61060 34440 61140 34450
rect 61480 34440 61560 34450
rect 61800 34440 61880 34450
rect 60820 34360 60830 34440
rect 61140 34360 61150 34440
rect 61560 34360 61570 34440
rect 61880 34360 61890 34440
rect 62140 34420 62150 34500
rect 62290 34420 62300 34500
rect 59350 34320 59440 34330
rect 59500 34320 59580 34330
rect 59650 34320 59760 34330
rect 60060 34320 60140 34330
rect 60210 34320 60290 34330
rect 60360 34320 60440 34330
rect 62060 34320 62140 34330
rect 62210 34320 62290 34330
rect 59410 34150 59440 34320
rect 59580 34240 59590 34320
rect 59670 34150 59760 34320
rect 60140 34240 60150 34320
rect 60290 34240 60300 34320
rect 60440 34240 60450 34320
rect 60580 34280 60660 34290
rect 60900 34280 60980 34290
rect 61320 34280 61400 34290
rect 61640 34280 61720 34290
rect 60660 34200 60670 34280
rect 60980 34200 60990 34280
rect 61400 34200 61410 34280
rect 61720 34200 61730 34280
rect 62140 34240 62150 34320
rect 62290 34240 62300 34320
rect 59350 34140 59440 34150
rect 59500 34140 59580 34150
rect 59650 34140 59760 34150
rect 60060 34140 60140 34150
rect 60210 34140 60290 34150
rect 60360 34140 60440 34150
rect 62060 34140 62140 34150
rect 62210 34140 62290 34150
rect 59410 33970 59440 34140
rect 59580 34060 59590 34140
rect 59670 33970 59760 34140
rect 60140 34060 60150 34140
rect 60290 34060 60300 34140
rect 60440 34060 60450 34140
rect 60740 34120 60820 34130
rect 61060 34120 61140 34130
rect 61480 34120 61560 34130
rect 61800 34120 61880 34130
rect 60820 34040 60830 34120
rect 61140 34040 61150 34120
rect 61560 34040 61570 34120
rect 61880 34040 61890 34120
rect 62140 34060 62150 34140
rect 62290 34060 62300 34140
rect 59350 33960 59440 33970
rect 59500 33960 59580 33970
rect 59650 33960 59760 33970
rect 60060 33960 60140 33970
rect 60210 33960 60290 33970
rect 60360 33960 60440 33970
rect 60580 33960 60660 33970
rect 60900 33960 60980 33970
rect 61320 33960 61400 33970
rect 61640 33960 61720 33970
rect 62060 33960 62140 33970
rect 62210 33960 62290 33970
rect 59410 33790 59440 33960
rect 59580 33880 59590 33960
rect 59670 33790 59760 33960
rect 60140 33880 60150 33960
rect 60290 33880 60300 33960
rect 60440 33880 60450 33960
rect 60660 33880 60670 33960
rect 60980 33880 60990 33960
rect 61400 33880 61410 33960
rect 61720 33880 61730 33960
rect 62140 33880 62150 33960
rect 62290 33880 62300 33960
rect 60740 33800 60820 33810
rect 61060 33800 61140 33810
rect 61480 33800 61560 33810
rect 61800 33800 61880 33810
rect 59350 33780 59440 33790
rect 59500 33780 59580 33790
rect 59650 33780 59760 33790
rect 60060 33780 60140 33790
rect 60210 33780 60290 33790
rect 60360 33780 60440 33790
rect 59410 33610 59440 33780
rect 59580 33700 59590 33780
rect 59670 33610 59760 33780
rect 60140 33700 60150 33780
rect 60290 33700 60300 33780
rect 60440 33700 60450 33780
rect 60820 33720 60830 33800
rect 61140 33720 61150 33800
rect 61560 33720 61570 33800
rect 61880 33720 61890 33800
rect 62060 33780 62140 33790
rect 62210 33780 62290 33790
rect 62140 33700 62150 33780
rect 62290 33700 62300 33780
rect 60580 33640 60660 33650
rect 60900 33640 60980 33650
rect 61320 33640 61400 33650
rect 61640 33640 61720 33650
rect 59350 33600 59440 33610
rect 59500 33600 59580 33610
rect 59650 33600 59760 33610
rect 60060 33600 60140 33610
rect 60210 33600 60290 33610
rect 60360 33600 60440 33610
rect 59410 33430 59440 33600
rect 59580 33520 59590 33600
rect 59670 33430 59760 33600
rect 60140 33520 60150 33600
rect 60290 33520 60300 33600
rect 60440 33520 60450 33600
rect 60660 33560 60670 33640
rect 60980 33560 60990 33640
rect 61400 33560 61410 33640
rect 61720 33560 61730 33640
rect 62060 33600 62140 33610
rect 62210 33600 62290 33610
rect 62140 33520 62150 33600
rect 62290 33520 62300 33600
rect 60740 33480 60820 33490
rect 61060 33480 61140 33490
rect 61480 33480 61560 33490
rect 61800 33480 61880 33490
rect 59350 33420 59440 33430
rect 59500 33420 59580 33430
rect 59650 33420 59760 33430
rect 60060 33420 60140 33430
rect 60210 33420 60290 33430
rect 60360 33420 60440 33430
rect 59410 33250 59440 33420
rect 59580 33340 59590 33420
rect 59670 33250 59760 33420
rect 60140 33340 60150 33420
rect 60290 33340 60300 33420
rect 60440 33340 60450 33420
rect 60820 33400 60830 33480
rect 61140 33400 61150 33480
rect 61560 33400 61570 33480
rect 61880 33400 61890 33480
rect 62060 33420 62140 33430
rect 62210 33420 62290 33430
rect 62140 33340 62150 33420
rect 62290 33340 62300 33420
rect 60580 33320 60660 33330
rect 60900 33320 60980 33330
rect 61320 33320 61400 33330
rect 61640 33320 61720 33330
rect 59350 33240 59440 33250
rect 59500 33240 59580 33250
rect 59650 33240 59760 33250
rect 60060 33240 60140 33250
rect 60210 33240 60290 33250
rect 60360 33240 60440 33250
rect 60660 33240 60670 33320
rect 60980 33240 60990 33320
rect 61400 33240 61410 33320
rect 61720 33240 61730 33320
rect 62060 33240 62140 33250
rect 62210 33240 62290 33250
rect 59410 33070 59440 33240
rect 59580 33160 59590 33240
rect 59670 33070 59760 33240
rect 60140 33160 60150 33240
rect 60290 33160 60300 33240
rect 60440 33160 60450 33240
rect 60740 33160 60820 33170
rect 61060 33160 61140 33170
rect 61480 33160 61560 33170
rect 61800 33160 61880 33170
rect 62140 33160 62150 33240
rect 62290 33160 62300 33240
rect 60820 33080 60830 33160
rect 61140 33080 61150 33160
rect 61560 33080 61570 33160
rect 61880 33080 61890 33160
rect 59350 33060 59440 33070
rect 59500 33060 59580 33070
rect 59650 33060 59760 33070
rect 60060 33060 60140 33070
rect 60210 33060 60290 33070
rect 60360 33060 60440 33070
rect 62060 33060 62140 33070
rect 62210 33060 62290 33070
rect 59410 32890 59440 33060
rect 59580 32980 59590 33060
rect 59670 32890 59760 33060
rect 60140 32980 60150 33060
rect 60290 32980 60300 33060
rect 60440 32980 60450 33060
rect 60580 33000 60660 33010
rect 60900 33000 60980 33010
rect 61320 33000 61400 33010
rect 61640 33000 61720 33010
rect 60660 32920 60670 33000
rect 60980 32920 60990 33000
rect 61400 32920 61410 33000
rect 61720 32920 61730 33000
rect 62140 32980 62150 33060
rect 62290 32980 62300 33060
rect 59350 32880 59440 32890
rect 59500 32880 59580 32890
rect 59650 32880 59760 32890
rect 60060 32880 60140 32890
rect 60210 32880 60290 32890
rect 60360 32880 60440 32890
rect 62060 32880 62140 32890
rect 62210 32880 62290 32890
rect 59410 32710 59440 32880
rect 59580 32800 59590 32880
rect 59670 32710 59760 32880
rect 60140 32800 60150 32880
rect 60290 32800 60300 32880
rect 60440 32800 60450 32880
rect 60740 32840 60820 32850
rect 61060 32840 61140 32850
rect 61480 32840 61560 32850
rect 61800 32840 61880 32850
rect 60820 32760 60830 32840
rect 61140 32760 61150 32840
rect 61560 32760 61570 32840
rect 61880 32760 61890 32840
rect 62140 32800 62150 32880
rect 62290 32800 62300 32880
rect 59350 32700 59440 32710
rect 59500 32700 59580 32710
rect 59650 32700 59760 32710
rect 60060 32700 60140 32710
rect 60210 32700 60290 32710
rect 60360 32700 60440 32710
rect 62060 32700 62140 32710
rect 62210 32700 62290 32710
rect 59410 32530 59440 32700
rect 59580 32620 59590 32700
rect 59670 32530 59760 32700
rect 60140 32620 60150 32700
rect 60290 32620 60300 32700
rect 60440 32620 60450 32700
rect 60580 32680 60660 32690
rect 60900 32680 60980 32690
rect 61320 32680 61400 32690
rect 61640 32680 61720 32690
rect 60660 32600 60670 32680
rect 60980 32600 60990 32680
rect 61400 32600 61410 32680
rect 61720 32600 61730 32680
rect 62140 32620 62150 32700
rect 62290 32620 62300 32700
rect 59350 32520 59440 32530
rect 59500 32520 59580 32530
rect 59650 32520 59760 32530
rect 60060 32520 60140 32530
rect 60210 32520 60290 32530
rect 60360 32520 60440 32530
rect 60740 32520 60820 32530
rect 61060 32520 61140 32530
rect 61480 32520 61560 32530
rect 61800 32520 61880 32530
rect 62060 32520 62140 32530
rect 62210 32520 62290 32530
rect 59410 32350 59440 32520
rect 59580 32440 59590 32520
rect 59670 32350 59760 32520
rect 60140 32440 60150 32520
rect 60290 32440 60300 32520
rect 60440 32440 60450 32520
rect 60820 32440 60830 32520
rect 61140 32440 61150 32520
rect 61560 32440 61570 32520
rect 61880 32440 61890 32520
rect 62140 32440 62150 32520
rect 62290 32440 62300 32520
rect 60580 32360 60660 32370
rect 60900 32360 60980 32370
rect 61320 32360 61400 32370
rect 61640 32360 61720 32370
rect 59350 32340 59440 32350
rect 59500 32340 59580 32350
rect 59650 32340 59760 32350
rect 60060 32340 60140 32350
rect 60210 32340 60290 32350
rect 60360 32340 60440 32350
rect 59410 32170 59440 32340
rect 59580 32260 59590 32340
rect 59670 32170 59760 32340
rect 60140 32260 60150 32340
rect 60290 32260 60300 32340
rect 60440 32260 60450 32340
rect 60660 32280 60670 32360
rect 60980 32280 60990 32360
rect 61400 32280 61410 32360
rect 61720 32280 61730 32360
rect 62060 32340 62140 32350
rect 62210 32340 62290 32350
rect 62140 32260 62150 32340
rect 62290 32260 62300 32340
rect 60740 32200 60820 32210
rect 61060 32200 61140 32210
rect 61480 32200 61560 32210
rect 61800 32200 61880 32210
rect 59350 32160 59440 32170
rect 59500 32160 59580 32170
rect 59650 32160 59760 32170
rect 60060 32160 60140 32170
rect 60210 32160 60290 32170
rect 60360 32160 60440 32170
rect 59410 31990 59440 32160
rect 59580 32080 59590 32160
rect 59670 31990 59760 32160
rect 60140 32080 60150 32160
rect 60290 32080 60300 32160
rect 60440 32080 60450 32160
rect 60820 32120 60830 32200
rect 61140 32120 61150 32200
rect 61560 32120 61570 32200
rect 61880 32120 61890 32200
rect 62060 32160 62140 32170
rect 62210 32160 62290 32170
rect 62140 32080 62150 32160
rect 62290 32080 62300 32160
rect 60580 32040 60660 32050
rect 60900 32040 60980 32050
rect 61320 32040 61400 32050
rect 61640 32040 61720 32050
rect 59350 31980 59440 31990
rect 59500 31980 59580 31990
rect 59650 31980 59760 31990
rect 60060 31980 60140 31990
rect 60210 31980 60290 31990
rect 60360 31980 60440 31990
rect 59410 31810 59440 31980
rect 59580 31900 59590 31980
rect 59670 31810 59760 31980
rect 60140 31900 60150 31980
rect 60290 31900 60300 31980
rect 60440 31900 60450 31980
rect 60660 31960 60670 32040
rect 60980 31960 60990 32040
rect 61400 31960 61410 32040
rect 61720 31960 61730 32040
rect 62060 31980 62140 31990
rect 62210 31980 62290 31990
rect 62140 31900 62150 31980
rect 62290 31900 62300 31980
rect 60740 31880 60820 31890
rect 61060 31880 61140 31890
rect 61480 31880 61560 31890
rect 61800 31880 61880 31890
rect 59350 31800 59440 31810
rect 59500 31800 59580 31810
rect 59650 31800 59760 31810
rect 60060 31800 60140 31810
rect 60210 31800 60290 31810
rect 60360 31800 60440 31810
rect 60820 31800 60830 31880
rect 61140 31800 61150 31880
rect 61560 31800 61570 31880
rect 61880 31800 61890 31880
rect 62060 31800 62140 31810
rect 62210 31800 62290 31810
rect 59410 31630 59440 31800
rect 59580 31720 59590 31800
rect 59670 31630 59760 31800
rect 60140 31720 60150 31800
rect 60290 31720 60300 31800
rect 60440 31720 60450 31800
rect 60580 31720 60660 31730
rect 60900 31720 60980 31730
rect 61320 31720 61400 31730
rect 61640 31720 61720 31730
rect 62140 31720 62150 31800
rect 62290 31720 62300 31800
rect 60660 31640 60670 31720
rect 60980 31640 60990 31720
rect 61400 31640 61410 31720
rect 61720 31640 61730 31720
rect 59350 31620 59440 31630
rect 59500 31620 59580 31630
rect 59650 31620 59760 31630
rect 60060 31620 60140 31630
rect 60210 31620 60290 31630
rect 60360 31620 60440 31630
rect 62060 31620 62140 31630
rect 62210 31620 62290 31630
rect 59410 31450 59440 31620
rect 59580 31540 59590 31620
rect 59670 31450 59760 31620
rect 60140 31540 60150 31620
rect 60290 31540 60300 31620
rect 60440 31540 60450 31620
rect 60740 31560 60820 31570
rect 61060 31560 61140 31570
rect 61480 31560 61560 31570
rect 61800 31560 61880 31570
rect 60820 31480 60830 31560
rect 61140 31480 61150 31560
rect 61560 31480 61570 31560
rect 61880 31480 61890 31560
rect 62140 31540 62150 31620
rect 62290 31540 62300 31620
rect 59350 31440 59440 31450
rect 59500 31440 59580 31450
rect 59650 31440 59760 31450
rect 60060 31440 60140 31450
rect 60210 31440 60290 31450
rect 60360 31440 60440 31450
rect 62060 31440 62140 31450
rect 62210 31440 62290 31450
rect 59410 31270 59440 31440
rect 59580 31360 59590 31440
rect 59670 31270 59760 31440
rect 60140 31360 60150 31440
rect 60290 31360 60300 31440
rect 60440 31360 60450 31440
rect 60580 31400 60660 31410
rect 60900 31400 60980 31410
rect 61320 31400 61400 31410
rect 61640 31400 61720 31410
rect 60660 31320 60670 31400
rect 60980 31320 60990 31400
rect 61400 31320 61410 31400
rect 61720 31320 61730 31400
rect 62140 31360 62150 31440
rect 62290 31360 62300 31440
rect 59350 31260 59440 31270
rect 59500 31260 59580 31270
rect 59650 31260 59760 31270
rect 60060 31260 60140 31270
rect 60210 31260 60290 31270
rect 60360 31260 60440 31270
rect 62060 31260 62140 31270
rect 62210 31260 62290 31270
rect 59410 31100 59440 31260
rect 59580 31180 59590 31260
rect 59670 31100 59760 31260
rect 60140 31180 60150 31260
rect 60290 31180 60300 31260
rect 60440 31180 60450 31260
rect 60740 31240 60820 31250
rect 61060 31240 61140 31250
rect 61480 31240 61560 31250
rect 61800 31240 61880 31250
rect 60820 31160 60830 31240
rect 61140 31160 61150 31240
rect 61560 31160 61570 31240
rect 61880 31160 61890 31240
rect 62140 31180 62150 31260
rect 62290 31180 62300 31260
rect 73245 31100 73260 37190
rect 73640 37120 73650 37200
rect 73790 37120 73800 37200
rect 73940 37120 73950 37200
rect 74080 37160 74160 37170
rect 74400 37160 74480 37170
rect 74820 37160 74900 37170
rect 75140 37160 75220 37170
rect 74160 37080 74170 37160
rect 74480 37080 74490 37160
rect 74900 37080 74910 37160
rect 75220 37080 75230 37160
rect 75640 37120 75650 37200
rect 75790 37120 75800 37200
rect 76240 37100 76255 37190
rect 73560 37020 73640 37030
rect 73710 37020 73790 37030
rect 73860 37020 73940 37030
rect 75560 37020 75640 37030
rect 75710 37020 75790 37030
rect 73640 36940 73650 37020
rect 73790 36940 73800 37020
rect 73940 36940 73950 37020
rect 74240 37000 74320 37010
rect 74560 37000 74640 37010
rect 74980 37000 75060 37010
rect 75300 37000 75380 37010
rect 74320 36920 74330 37000
rect 74640 36920 74650 37000
rect 75060 36920 75070 37000
rect 75380 36920 75390 37000
rect 75640 36940 75650 37020
rect 75790 36940 75800 37020
rect 73560 36840 73640 36850
rect 73710 36840 73790 36850
rect 73860 36840 73940 36850
rect 74080 36840 74160 36850
rect 74400 36840 74480 36850
rect 74820 36840 74900 36850
rect 75140 36840 75220 36850
rect 75560 36840 75640 36850
rect 75710 36840 75790 36850
rect 73640 36760 73650 36840
rect 73790 36760 73800 36840
rect 73940 36760 73950 36840
rect 74160 36760 74170 36840
rect 74480 36760 74490 36840
rect 74900 36760 74910 36840
rect 75220 36760 75230 36840
rect 75640 36760 75650 36840
rect 75790 36760 75800 36840
rect 74240 36680 74320 36690
rect 74560 36680 74640 36690
rect 74980 36680 75060 36690
rect 75300 36680 75380 36690
rect 73560 36660 73640 36670
rect 73710 36660 73790 36670
rect 73860 36660 73940 36670
rect 73640 36580 73650 36660
rect 73790 36580 73800 36660
rect 73940 36580 73950 36660
rect 74320 36600 74330 36680
rect 74640 36600 74650 36680
rect 75060 36600 75070 36680
rect 75380 36600 75390 36680
rect 75560 36660 75640 36670
rect 75710 36660 75790 36670
rect 75640 36580 75650 36660
rect 75790 36580 75800 36660
rect 74080 36520 74160 36530
rect 74400 36520 74480 36530
rect 74820 36520 74900 36530
rect 75140 36520 75220 36530
rect 73560 36480 73640 36490
rect 73710 36480 73790 36490
rect 73860 36480 73940 36490
rect 73640 36400 73650 36480
rect 73790 36400 73800 36480
rect 73940 36400 73950 36480
rect 74160 36440 74170 36520
rect 74480 36440 74490 36520
rect 74900 36440 74910 36520
rect 75220 36440 75230 36520
rect 75560 36480 75640 36490
rect 75710 36480 75790 36490
rect 75640 36400 75650 36480
rect 75790 36400 75800 36480
rect 74240 36360 74320 36370
rect 74560 36360 74640 36370
rect 74980 36360 75060 36370
rect 75300 36360 75380 36370
rect 73560 36300 73640 36310
rect 73710 36300 73790 36310
rect 73860 36300 73940 36310
rect 73640 36220 73650 36300
rect 73790 36220 73800 36300
rect 73940 36220 73950 36300
rect 74320 36280 74330 36360
rect 74640 36280 74650 36360
rect 75060 36280 75070 36360
rect 75380 36280 75390 36360
rect 75560 36300 75640 36310
rect 75710 36300 75790 36310
rect 75640 36220 75650 36300
rect 75790 36220 75800 36300
rect 74080 36200 74160 36210
rect 74400 36200 74480 36210
rect 74820 36200 74900 36210
rect 75140 36200 75220 36210
rect 73560 36120 73640 36130
rect 73710 36120 73790 36130
rect 73860 36120 73940 36130
rect 74160 36120 74170 36200
rect 74480 36120 74490 36200
rect 74900 36120 74910 36200
rect 75220 36120 75230 36200
rect 75560 36120 75640 36130
rect 75710 36120 75790 36130
rect 73640 36040 73650 36120
rect 73790 36040 73800 36120
rect 73940 36040 73950 36120
rect 74240 36040 74320 36050
rect 74560 36040 74640 36050
rect 74980 36040 75060 36050
rect 75300 36040 75380 36050
rect 75640 36040 75650 36120
rect 75790 36040 75800 36120
rect 74320 35960 74330 36040
rect 74640 35960 74650 36040
rect 75060 35960 75070 36040
rect 75380 35960 75390 36040
rect 73560 35940 73640 35950
rect 73710 35940 73790 35950
rect 73860 35940 73940 35950
rect 75560 35940 75640 35950
rect 75710 35940 75790 35950
rect 73640 35860 73650 35940
rect 73790 35860 73800 35940
rect 73940 35860 73950 35940
rect 74080 35880 74160 35890
rect 74400 35880 74480 35890
rect 74820 35880 74900 35890
rect 75140 35880 75220 35890
rect 74160 35800 74170 35880
rect 74480 35800 74490 35880
rect 74900 35800 74910 35880
rect 75220 35800 75230 35880
rect 75640 35860 75650 35940
rect 75790 35860 75800 35940
rect 73560 35760 73640 35770
rect 73710 35760 73790 35770
rect 73860 35760 73940 35770
rect 75560 35760 75640 35770
rect 75710 35760 75790 35770
rect 73640 35680 73650 35760
rect 73790 35680 73800 35760
rect 73940 35680 73950 35760
rect 74240 35720 74320 35730
rect 74560 35720 74640 35730
rect 74980 35720 75060 35730
rect 75300 35720 75380 35730
rect 74320 35640 74330 35720
rect 74640 35640 74650 35720
rect 75060 35640 75070 35720
rect 75380 35640 75390 35720
rect 75640 35680 75650 35760
rect 75790 35680 75800 35760
rect 73560 35580 73640 35590
rect 73710 35580 73790 35590
rect 73860 35580 73940 35590
rect 75560 35580 75640 35590
rect 75710 35580 75790 35590
rect 73640 35500 73650 35580
rect 73790 35500 73800 35580
rect 73940 35500 73950 35580
rect 74080 35560 74160 35570
rect 74400 35560 74480 35570
rect 74820 35560 74900 35570
rect 75140 35560 75220 35570
rect 74160 35480 74170 35560
rect 74480 35480 74490 35560
rect 74900 35480 74910 35560
rect 75220 35480 75230 35560
rect 75640 35500 75650 35580
rect 75790 35500 75800 35580
rect 73560 35400 73640 35410
rect 73710 35400 73790 35410
rect 73860 35400 73940 35410
rect 74240 35400 74320 35410
rect 74560 35400 74640 35410
rect 74980 35400 75060 35410
rect 75300 35400 75380 35410
rect 75560 35400 75640 35410
rect 75710 35400 75790 35410
rect 73640 35320 73650 35400
rect 73790 35320 73800 35400
rect 73940 35320 73950 35400
rect 74320 35320 74330 35400
rect 74640 35320 74650 35400
rect 75060 35320 75070 35400
rect 75380 35320 75390 35400
rect 75640 35320 75650 35400
rect 75790 35320 75800 35400
rect 74080 35240 74160 35250
rect 74400 35240 74480 35250
rect 74820 35240 74900 35250
rect 75140 35240 75220 35250
rect 73560 35220 73640 35230
rect 73710 35220 73790 35230
rect 73860 35220 73940 35230
rect 73640 35140 73650 35220
rect 73790 35140 73800 35220
rect 73940 35140 73950 35220
rect 74160 35160 74170 35240
rect 74480 35160 74490 35240
rect 74900 35160 74910 35240
rect 75220 35160 75230 35240
rect 75560 35220 75640 35230
rect 75710 35220 75790 35230
rect 75640 35140 75650 35220
rect 75790 35140 75800 35220
rect 74240 35080 74320 35090
rect 74560 35080 74640 35090
rect 74980 35080 75060 35090
rect 75300 35080 75380 35090
rect 73560 35040 73640 35050
rect 73710 35040 73790 35050
rect 73860 35040 73940 35050
rect 73640 34960 73650 35040
rect 73790 34960 73800 35040
rect 73940 34960 73950 35040
rect 74320 35000 74330 35080
rect 74640 35000 74650 35080
rect 75060 35000 75070 35080
rect 75380 35000 75390 35080
rect 75560 35040 75640 35050
rect 75710 35040 75790 35050
rect 75640 34960 75650 35040
rect 75790 34960 75800 35040
rect 74080 34920 74160 34930
rect 74400 34920 74480 34930
rect 74820 34920 74900 34930
rect 75140 34920 75220 34930
rect 73560 34860 73640 34870
rect 73710 34860 73790 34870
rect 73860 34860 73940 34870
rect 73640 34780 73650 34860
rect 73790 34780 73800 34860
rect 73940 34780 73950 34860
rect 74160 34840 74170 34920
rect 74480 34840 74490 34920
rect 74900 34840 74910 34920
rect 75220 34840 75230 34920
rect 75560 34860 75640 34870
rect 75710 34860 75790 34870
rect 75640 34780 75650 34860
rect 75790 34780 75800 34860
rect 74240 34760 74320 34770
rect 74560 34760 74640 34770
rect 74980 34760 75060 34770
rect 75300 34760 75380 34770
rect 73560 34680 73640 34690
rect 73710 34680 73790 34690
rect 73860 34680 73940 34690
rect 74320 34680 74330 34760
rect 74640 34680 74650 34760
rect 75060 34680 75070 34760
rect 75380 34680 75390 34760
rect 75560 34680 75640 34690
rect 75710 34680 75790 34690
rect 73640 34600 73650 34680
rect 73790 34600 73800 34680
rect 73940 34600 73950 34680
rect 74080 34600 74160 34610
rect 74400 34600 74480 34610
rect 74820 34600 74900 34610
rect 75140 34600 75220 34610
rect 75640 34600 75650 34680
rect 75790 34600 75800 34680
rect 74160 34520 74170 34600
rect 74480 34520 74490 34600
rect 74900 34520 74910 34600
rect 75220 34520 75230 34600
rect 73560 34500 73640 34510
rect 73710 34500 73790 34510
rect 73860 34500 73940 34510
rect 75560 34500 75640 34510
rect 75710 34500 75790 34510
rect 73640 34420 73650 34500
rect 73790 34420 73800 34500
rect 73940 34420 73950 34500
rect 74240 34440 74320 34450
rect 74560 34440 74640 34450
rect 74980 34440 75060 34450
rect 75300 34440 75380 34450
rect 74320 34360 74330 34440
rect 74640 34360 74650 34440
rect 75060 34360 75070 34440
rect 75380 34360 75390 34440
rect 75640 34420 75650 34500
rect 75790 34420 75800 34500
rect 73560 34320 73640 34330
rect 73710 34320 73790 34330
rect 73860 34320 73940 34330
rect 75560 34320 75640 34330
rect 75710 34320 75790 34330
rect 73640 34240 73650 34320
rect 73790 34240 73800 34320
rect 73940 34240 73950 34320
rect 74080 34280 74160 34290
rect 74400 34280 74480 34290
rect 74820 34280 74900 34290
rect 75140 34280 75220 34290
rect 74160 34200 74170 34280
rect 74480 34200 74490 34280
rect 74900 34200 74910 34280
rect 75220 34200 75230 34280
rect 75640 34240 75650 34320
rect 75790 34240 75800 34320
rect 73560 34140 73640 34150
rect 73710 34140 73790 34150
rect 73860 34140 73940 34150
rect 75560 34140 75640 34150
rect 75710 34140 75790 34150
rect 73640 34060 73650 34140
rect 73790 34060 73800 34140
rect 73940 34060 73950 34140
rect 74240 34120 74320 34130
rect 74560 34120 74640 34130
rect 74980 34120 75060 34130
rect 75300 34120 75380 34130
rect 74320 34040 74330 34120
rect 74640 34040 74650 34120
rect 75060 34040 75070 34120
rect 75380 34040 75390 34120
rect 75640 34060 75650 34140
rect 75790 34060 75800 34140
rect 73560 33960 73640 33970
rect 73710 33960 73790 33970
rect 73860 33960 73940 33970
rect 74080 33960 74160 33970
rect 74400 33960 74480 33970
rect 74820 33960 74900 33970
rect 75140 33960 75220 33970
rect 75560 33960 75640 33970
rect 75710 33960 75790 33970
rect 73640 33880 73650 33960
rect 73790 33880 73800 33960
rect 73940 33880 73950 33960
rect 74160 33880 74170 33960
rect 74480 33880 74490 33960
rect 74900 33880 74910 33960
rect 75220 33880 75230 33960
rect 75640 33880 75650 33960
rect 75790 33880 75800 33960
rect 74240 33800 74320 33810
rect 74560 33800 74640 33810
rect 74980 33800 75060 33810
rect 75300 33800 75380 33810
rect 73560 33780 73640 33790
rect 73710 33780 73790 33790
rect 73860 33780 73940 33790
rect 73640 33700 73650 33780
rect 73790 33700 73800 33780
rect 73940 33700 73950 33780
rect 74320 33720 74330 33800
rect 74640 33720 74650 33800
rect 75060 33720 75070 33800
rect 75380 33720 75390 33800
rect 75560 33780 75640 33790
rect 75710 33780 75790 33790
rect 75640 33700 75650 33780
rect 75790 33700 75800 33780
rect 74080 33640 74160 33650
rect 74400 33640 74480 33650
rect 74820 33640 74900 33650
rect 75140 33640 75220 33650
rect 73560 33600 73640 33610
rect 73710 33600 73790 33610
rect 73860 33600 73940 33610
rect 73640 33520 73650 33600
rect 73790 33520 73800 33600
rect 73940 33520 73950 33600
rect 74160 33560 74170 33640
rect 74480 33560 74490 33640
rect 74900 33560 74910 33640
rect 75220 33560 75230 33640
rect 75560 33600 75640 33610
rect 75710 33600 75790 33610
rect 75640 33520 75650 33600
rect 75790 33520 75800 33600
rect 74240 33480 74320 33490
rect 74560 33480 74640 33490
rect 74980 33480 75060 33490
rect 75300 33480 75380 33490
rect 73560 33420 73640 33430
rect 73710 33420 73790 33430
rect 73860 33420 73940 33430
rect 73640 33340 73650 33420
rect 73790 33340 73800 33420
rect 73940 33340 73950 33420
rect 74320 33400 74330 33480
rect 74640 33400 74650 33480
rect 75060 33400 75070 33480
rect 75380 33400 75390 33480
rect 75560 33420 75640 33430
rect 75710 33420 75790 33430
rect 75640 33340 75650 33420
rect 75790 33340 75800 33420
rect 74080 33320 74160 33330
rect 74400 33320 74480 33330
rect 74820 33320 74900 33330
rect 75140 33320 75220 33330
rect 73560 33240 73640 33250
rect 73710 33240 73790 33250
rect 73860 33240 73940 33250
rect 74160 33240 74170 33320
rect 74480 33240 74490 33320
rect 74900 33240 74910 33320
rect 75220 33240 75230 33320
rect 75560 33240 75640 33250
rect 75710 33240 75790 33250
rect 73640 33160 73650 33240
rect 73790 33160 73800 33240
rect 73940 33160 73950 33240
rect 74240 33160 74320 33170
rect 74560 33160 74640 33170
rect 74980 33160 75060 33170
rect 75300 33160 75380 33170
rect 75640 33160 75650 33240
rect 75790 33160 75800 33240
rect 74320 33080 74330 33160
rect 74640 33080 74650 33160
rect 75060 33080 75070 33160
rect 75380 33080 75390 33160
rect 73560 33060 73640 33070
rect 73710 33060 73790 33070
rect 73860 33060 73940 33070
rect 75560 33060 75640 33070
rect 75710 33060 75790 33070
rect 73640 32980 73650 33060
rect 73790 32980 73800 33060
rect 73940 32980 73950 33060
rect 74080 33000 74160 33010
rect 74400 33000 74480 33010
rect 74820 33000 74900 33010
rect 75140 33000 75220 33010
rect 74160 32920 74170 33000
rect 74480 32920 74490 33000
rect 74900 32920 74910 33000
rect 75220 32920 75230 33000
rect 75640 32980 75650 33060
rect 75790 32980 75800 33060
rect 73560 32880 73640 32890
rect 73710 32880 73790 32890
rect 73860 32880 73940 32890
rect 75560 32880 75640 32890
rect 75710 32880 75790 32890
rect 73640 32800 73650 32880
rect 73790 32800 73800 32880
rect 73940 32800 73950 32880
rect 74240 32840 74320 32850
rect 74560 32840 74640 32850
rect 74980 32840 75060 32850
rect 75300 32840 75380 32850
rect 74320 32760 74330 32840
rect 74640 32760 74650 32840
rect 75060 32760 75070 32840
rect 75380 32760 75390 32840
rect 75640 32800 75650 32880
rect 75790 32800 75800 32880
rect 73560 32700 73640 32710
rect 73710 32700 73790 32710
rect 73860 32700 73940 32710
rect 75560 32700 75640 32710
rect 75710 32700 75790 32710
rect 73640 32620 73650 32700
rect 73790 32620 73800 32700
rect 73940 32620 73950 32700
rect 74080 32680 74160 32690
rect 74400 32680 74480 32690
rect 74820 32680 74900 32690
rect 75140 32680 75220 32690
rect 74160 32600 74170 32680
rect 74480 32600 74490 32680
rect 74900 32600 74910 32680
rect 75220 32600 75230 32680
rect 75640 32620 75650 32700
rect 75790 32620 75800 32700
rect 73560 32520 73640 32530
rect 73710 32520 73790 32530
rect 73860 32520 73940 32530
rect 74240 32520 74320 32530
rect 74560 32520 74640 32530
rect 74980 32520 75060 32530
rect 75300 32520 75380 32530
rect 75560 32520 75640 32530
rect 75710 32520 75790 32530
rect 73640 32440 73650 32520
rect 73790 32440 73800 32520
rect 73940 32440 73950 32520
rect 74320 32440 74330 32520
rect 74640 32440 74650 32520
rect 75060 32440 75070 32520
rect 75380 32440 75390 32520
rect 75640 32440 75650 32520
rect 75790 32440 75800 32520
rect 74080 32360 74160 32370
rect 74400 32360 74480 32370
rect 74820 32360 74900 32370
rect 75140 32360 75220 32370
rect 73560 32340 73640 32350
rect 73710 32340 73790 32350
rect 73860 32340 73940 32350
rect 73640 32260 73650 32340
rect 73790 32260 73800 32340
rect 73940 32260 73950 32340
rect 74160 32280 74170 32360
rect 74480 32280 74490 32360
rect 74900 32280 74910 32360
rect 75220 32280 75230 32360
rect 75560 32340 75640 32350
rect 75710 32340 75790 32350
rect 75640 32260 75650 32340
rect 75790 32260 75800 32340
rect 74240 32200 74320 32210
rect 74560 32200 74640 32210
rect 74980 32200 75060 32210
rect 75300 32200 75380 32210
rect 73560 32160 73640 32170
rect 73710 32160 73790 32170
rect 73860 32160 73940 32170
rect 73640 32080 73650 32160
rect 73790 32080 73800 32160
rect 73940 32080 73950 32160
rect 74320 32120 74330 32200
rect 74640 32120 74650 32200
rect 75060 32120 75070 32200
rect 75380 32120 75390 32200
rect 75560 32160 75640 32170
rect 75710 32160 75790 32170
rect 75640 32080 75650 32160
rect 75790 32080 75800 32160
rect 74080 32040 74160 32050
rect 74400 32040 74480 32050
rect 74820 32040 74900 32050
rect 75140 32040 75220 32050
rect 73560 31980 73640 31990
rect 73710 31980 73790 31990
rect 73860 31980 73940 31990
rect 73640 31900 73650 31980
rect 73790 31900 73800 31980
rect 73940 31900 73950 31980
rect 74160 31960 74170 32040
rect 74480 31960 74490 32040
rect 74900 31960 74910 32040
rect 75220 31960 75230 32040
rect 75560 31980 75640 31990
rect 75710 31980 75790 31990
rect 75640 31900 75650 31980
rect 75790 31900 75800 31980
rect 74240 31880 74320 31890
rect 74560 31880 74640 31890
rect 74980 31880 75060 31890
rect 75300 31880 75380 31890
rect 73560 31800 73640 31810
rect 73710 31800 73790 31810
rect 73860 31800 73940 31810
rect 74320 31800 74330 31880
rect 74640 31800 74650 31880
rect 75060 31800 75070 31880
rect 75380 31800 75390 31880
rect 75560 31800 75640 31810
rect 75710 31800 75790 31810
rect 73640 31720 73650 31800
rect 73790 31720 73800 31800
rect 73940 31720 73950 31800
rect 74080 31720 74160 31730
rect 74400 31720 74480 31730
rect 74820 31720 74900 31730
rect 75140 31720 75220 31730
rect 75640 31720 75650 31800
rect 75790 31720 75800 31800
rect 74160 31640 74170 31720
rect 74480 31640 74490 31720
rect 74900 31640 74910 31720
rect 75220 31640 75230 31720
rect 73560 31620 73640 31630
rect 73710 31620 73790 31630
rect 73860 31620 73940 31630
rect 75560 31620 75640 31630
rect 75710 31620 75790 31630
rect 73640 31540 73650 31620
rect 73790 31540 73800 31620
rect 73940 31540 73950 31620
rect 74240 31560 74320 31570
rect 74560 31560 74640 31570
rect 74980 31560 75060 31570
rect 75300 31560 75380 31570
rect 74320 31480 74330 31560
rect 74640 31480 74650 31560
rect 75060 31480 75070 31560
rect 75380 31480 75390 31560
rect 75640 31540 75650 31620
rect 75790 31540 75800 31620
rect 73560 31440 73640 31450
rect 73710 31440 73790 31450
rect 73860 31440 73940 31450
rect 75560 31440 75640 31450
rect 75710 31440 75790 31450
rect 73640 31360 73650 31440
rect 73790 31360 73800 31440
rect 73940 31360 73950 31440
rect 74080 31400 74160 31410
rect 74400 31400 74480 31410
rect 74820 31400 74900 31410
rect 75140 31400 75220 31410
rect 74160 31320 74170 31400
rect 74480 31320 74490 31400
rect 74900 31320 74910 31400
rect 75220 31320 75230 31400
rect 75640 31360 75650 31440
rect 75790 31360 75800 31440
rect 73560 31260 73640 31270
rect 73710 31260 73790 31270
rect 73860 31260 73940 31270
rect 75560 31260 75640 31270
rect 75710 31260 75790 31270
rect 73640 31180 73650 31260
rect 73790 31180 73800 31260
rect 73940 31180 73950 31260
rect 74240 31240 74320 31250
rect 74560 31240 74640 31250
rect 74980 31240 75060 31250
rect 75300 31240 75380 31250
rect 74320 31160 74330 31240
rect 74640 31160 74650 31240
rect 75060 31160 75070 31240
rect 75380 31160 75390 31240
rect 75640 31180 75650 31260
rect 75790 31180 75800 31260
rect 86745 31100 86760 37190
rect 87140 37120 87150 37200
rect 87290 37120 87300 37200
rect 87440 37120 87450 37200
rect 87580 37160 87660 37170
rect 87900 37160 87980 37170
rect 88320 37160 88400 37170
rect 88640 37160 88720 37170
rect 87660 37080 87670 37160
rect 87980 37080 87990 37160
rect 88400 37080 88410 37160
rect 88720 37080 88730 37160
rect 89140 37120 89150 37200
rect 89290 37120 89300 37200
rect 89740 37100 89755 37190
rect 87060 37020 87140 37030
rect 87210 37020 87290 37030
rect 87360 37020 87440 37030
rect 89060 37020 89140 37030
rect 89210 37020 89290 37030
rect 87140 36940 87150 37020
rect 87290 36940 87300 37020
rect 87440 36940 87450 37020
rect 87740 37000 87820 37010
rect 88060 37000 88140 37010
rect 88480 37000 88560 37010
rect 88800 37000 88880 37010
rect 87820 36920 87830 37000
rect 88140 36920 88150 37000
rect 88560 36920 88570 37000
rect 88880 36920 88890 37000
rect 89140 36940 89150 37020
rect 89290 36940 89300 37020
rect 87060 36840 87140 36850
rect 87210 36840 87290 36850
rect 87360 36840 87440 36850
rect 87580 36840 87660 36850
rect 87900 36840 87980 36850
rect 88320 36840 88400 36850
rect 88640 36840 88720 36850
rect 89060 36840 89140 36850
rect 89210 36840 89290 36850
rect 87140 36760 87150 36840
rect 87290 36760 87300 36840
rect 87440 36760 87450 36840
rect 87660 36760 87670 36840
rect 87980 36760 87990 36840
rect 88400 36760 88410 36840
rect 88720 36760 88730 36840
rect 89140 36760 89150 36840
rect 89290 36760 89300 36840
rect 87740 36680 87820 36690
rect 88060 36680 88140 36690
rect 88480 36680 88560 36690
rect 88800 36680 88880 36690
rect 87060 36660 87140 36670
rect 87210 36660 87290 36670
rect 87360 36660 87440 36670
rect 87140 36580 87150 36660
rect 87290 36580 87300 36660
rect 87440 36580 87450 36660
rect 87820 36600 87830 36680
rect 88140 36600 88150 36680
rect 88560 36600 88570 36680
rect 88880 36600 88890 36680
rect 89060 36660 89140 36670
rect 89210 36660 89290 36670
rect 89140 36580 89150 36660
rect 89290 36580 89300 36660
rect 87580 36520 87660 36530
rect 87900 36520 87980 36530
rect 88320 36520 88400 36530
rect 88640 36520 88720 36530
rect 87060 36480 87140 36490
rect 87210 36480 87290 36490
rect 87360 36480 87440 36490
rect 87140 36400 87150 36480
rect 87290 36400 87300 36480
rect 87440 36400 87450 36480
rect 87660 36440 87670 36520
rect 87980 36440 87990 36520
rect 88400 36440 88410 36520
rect 88720 36440 88730 36520
rect 89060 36480 89140 36490
rect 89210 36480 89290 36490
rect 89140 36400 89150 36480
rect 89290 36400 89300 36480
rect 87740 36360 87820 36370
rect 88060 36360 88140 36370
rect 88480 36360 88560 36370
rect 88800 36360 88880 36370
rect 87060 36300 87140 36310
rect 87210 36300 87290 36310
rect 87360 36300 87440 36310
rect 87140 36220 87150 36300
rect 87290 36220 87300 36300
rect 87440 36220 87450 36300
rect 87820 36280 87830 36360
rect 88140 36280 88150 36360
rect 88560 36280 88570 36360
rect 88880 36280 88890 36360
rect 89060 36300 89140 36310
rect 89210 36300 89290 36310
rect 89140 36220 89150 36300
rect 89290 36220 89300 36300
rect 87580 36200 87660 36210
rect 87900 36200 87980 36210
rect 88320 36200 88400 36210
rect 88640 36200 88720 36210
rect 87060 36120 87140 36130
rect 87210 36120 87290 36130
rect 87360 36120 87440 36130
rect 87660 36120 87670 36200
rect 87980 36120 87990 36200
rect 88400 36120 88410 36200
rect 88720 36120 88730 36200
rect 89060 36120 89140 36130
rect 89210 36120 89290 36130
rect 87140 36040 87150 36120
rect 87290 36040 87300 36120
rect 87440 36040 87450 36120
rect 87740 36040 87820 36050
rect 88060 36040 88140 36050
rect 88480 36040 88560 36050
rect 88800 36040 88880 36050
rect 89140 36040 89150 36120
rect 89290 36040 89300 36120
rect 87820 35960 87830 36040
rect 88140 35960 88150 36040
rect 88560 35960 88570 36040
rect 88880 35960 88890 36040
rect 87060 35940 87140 35950
rect 87210 35940 87290 35950
rect 87360 35940 87440 35950
rect 89060 35940 89140 35950
rect 89210 35940 89290 35950
rect 87140 35860 87150 35940
rect 87290 35860 87300 35940
rect 87440 35860 87450 35940
rect 87580 35880 87660 35890
rect 87900 35880 87980 35890
rect 88320 35880 88400 35890
rect 88640 35880 88720 35890
rect 87660 35800 87670 35880
rect 87980 35800 87990 35880
rect 88400 35800 88410 35880
rect 88720 35800 88730 35880
rect 89140 35860 89150 35940
rect 89290 35860 89300 35940
rect 87060 35760 87140 35770
rect 87210 35760 87290 35770
rect 87360 35760 87440 35770
rect 89060 35760 89140 35770
rect 89210 35760 89290 35770
rect 87140 35680 87150 35760
rect 87290 35680 87300 35760
rect 87440 35680 87450 35760
rect 87740 35720 87820 35730
rect 88060 35720 88140 35730
rect 88480 35720 88560 35730
rect 88800 35720 88880 35730
rect 87820 35640 87830 35720
rect 88140 35640 88150 35720
rect 88560 35640 88570 35720
rect 88880 35640 88890 35720
rect 89140 35680 89150 35760
rect 89290 35680 89300 35760
rect 87060 35580 87140 35590
rect 87210 35580 87290 35590
rect 87360 35580 87440 35590
rect 89060 35580 89140 35590
rect 89210 35580 89290 35590
rect 87140 35500 87150 35580
rect 87290 35500 87300 35580
rect 87440 35500 87450 35580
rect 87580 35560 87660 35570
rect 87900 35560 87980 35570
rect 88320 35560 88400 35570
rect 88640 35560 88720 35570
rect 87660 35480 87670 35560
rect 87980 35480 87990 35560
rect 88400 35480 88410 35560
rect 88720 35480 88730 35560
rect 89140 35500 89150 35580
rect 89290 35500 89300 35580
rect 87060 35400 87140 35410
rect 87210 35400 87290 35410
rect 87360 35400 87440 35410
rect 87740 35400 87820 35410
rect 88060 35400 88140 35410
rect 88480 35400 88560 35410
rect 88800 35400 88880 35410
rect 89060 35400 89140 35410
rect 89210 35400 89290 35410
rect 87140 35320 87150 35400
rect 87290 35320 87300 35400
rect 87440 35320 87450 35400
rect 87820 35320 87830 35400
rect 88140 35320 88150 35400
rect 88560 35320 88570 35400
rect 88880 35320 88890 35400
rect 89140 35320 89150 35400
rect 89290 35320 89300 35400
rect 87580 35240 87660 35250
rect 87900 35240 87980 35250
rect 88320 35240 88400 35250
rect 88640 35240 88720 35250
rect 87060 35220 87140 35230
rect 87210 35220 87290 35230
rect 87360 35220 87440 35230
rect 87140 35140 87150 35220
rect 87290 35140 87300 35220
rect 87440 35140 87450 35220
rect 87660 35160 87670 35240
rect 87980 35160 87990 35240
rect 88400 35160 88410 35240
rect 88720 35160 88730 35240
rect 89060 35220 89140 35230
rect 89210 35220 89290 35230
rect 89140 35140 89150 35220
rect 89290 35140 89300 35220
rect 87740 35080 87820 35090
rect 88060 35080 88140 35090
rect 88480 35080 88560 35090
rect 88800 35080 88880 35090
rect 87060 35040 87140 35050
rect 87210 35040 87290 35050
rect 87360 35040 87440 35050
rect 87140 34960 87150 35040
rect 87290 34960 87300 35040
rect 87440 34960 87450 35040
rect 87820 35000 87830 35080
rect 88140 35000 88150 35080
rect 88560 35000 88570 35080
rect 88880 35000 88890 35080
rect 89060 35040 89140 35050
rect 89210 35040 89290 35050
rect 89140 34960 89150 35040
rect 89290 34960 89300 35040
rect 87580 34920 87660 34930
rect 87900 34920 87980 34930
rect 88320 34920 88400 34930
rect 88640 34920 88720 34930
rect 87060 34860 87140 34870
rect 87210 34860 87290 34870
rect 87360 34860 87440 34870
rect 87140 34780 87150 34860
rect 87290 34780 87300 34860
rect 87440 34780 87450 34860
rect 87660 34840 87670 34920
rect 87980 34840 87990 34920
rect 88400 34840 88410 34920
rect 88720 34840 88730 34920
rect 89060 34860 89140 34870
rect 89210 34860 89290 34870
rect 89140 34780 89150 34860
rect 89290 34780 89300 34860
rect 87740 34760 87820 34770
rect 88060 34760 88140 34770
rect 88480 34760 88560 34770
rect 88800 34760 88880 34770
rect 87060 34680 87140 34690
rect 87210 34680 87290 34690
rect 87360 34680 87440 34690
rect 87820 34680 87830 34760
rect 88140 34680 88150 34760
rect 88560 34680 88570 34760
rect 88880 34680 88890 34760
rect 89060 34680 89140 34690
rect 89210 34680 89290 34690
rect 87140 34600 87150 34680
rect 87290 34600 87300 34680
rect 87440 34600 87450 34680
rect 87580 34600 87660 34610
rect 87900 34600 87980 34610
rect 88320 34600 88400 34610
rect 88640 34600 88720 34610
rect 89140 34600 89150 34680
rect 89290 34600 89300 34680
rect 87660 34520 87670 34600
rect 87980 34520 87990 34600
rect 88400 34520 88410 34600
rect 88720 34520 88730 34600
rect 87060 34500 87140 34510
rect 87210 34500 87290 34510
rect 87360 34500 87440 34510
rect 89060 34500 89140 34510
rect 89210 34500 89290 34510
rect 87140 34420 87150 34500
rect 87290 34420 87300 34500
rect 87440 34420 87450 34500
rect 87740 34440 87820 34450
rect 88060 34440 88140 34450
rect 88480 34440 88560 34450
rect 88800 34440 88880 34450
rect 87820 34360 87830 34440
rect 88140 34360 88150 34440
rect 88560 34360 88570 34440
rect 88880 34360 88890 34440
rect 89140 34420 89150 34500
rect 89290 34420 89300 34500
rect 87060 34320 87140 34330
rect 87210 34320 87290 34330
rect 87360 34320 87440 34330
rect 89060 34320 89140 34330
rect 89210 34320 89290 34330
rect 87140 34240 87150 34320
rect 87290 34240 87300 34320
rect 87440 34240 87450 34320
rect 87580 34280 87660 34290
rect 87900 34280 87980 34290
rect 88320 34280 88400 34290
rect 88640 34280 88720 34290
rect 87660 34200 87670 34280
rect 87980 34200 87990 34280
rect 88400 34200 88410 34280
rect 88720 34200 88730 34280
rect 89140 34240 89150 34320
rect 89290 34240 89300 34320
rect 87060 34140 87140 34150
rect 87210 34140 87290 34150
rect 87360 34140 87440 34150
rect 89060 34140 89140 34150
rect 89210 34140 89290 34150
rect 87140 34060 87150 34140
rect 87290 34060 87300 34140
rect 87440 34060 87450 34140
rect 87740 34120 87820 34130
rect 88060 34120 88140 34130
rect 88480 34120 88560 34130
rect 88800 34120 88880 34130
rect 87820 34040 87830 34120
rect 88140 34040 88150 34120
rect 88560 34040 88570 34120
rect 88880 34040 88890 34120
rect 89140 34060 89150 34140
rect 89290 34060 89300 34140
rect 87060 33960 87140 33970
rect 87210 33960 87290 33970
rect 87360 33960 87440 33970
rect 87580 33960 87660 33970
rect 87900 33960 87980 33970
rect 88320 33960 88400 33970
rect 88640 33960 88720 33970
rect 89060 33960 89140 33970
rect 89210 33960 89290 33970
rect 87140 33880 87150 33960
rect 87290 33880 87300 33960
rect 87440 33880 87450 33960
rect 87660 33880 87670 33960
rect 87980 33880 87990 33960
rect 88400 33880 88410 33960
rect 88720 33880 88730 33960
rect 89140 33880 89150 33960
rect 89290 33880 89300 33960
rect 87740 33800 87820 33810
rect 88060 33800 88140 33810
rect 88480 33800 88560 33810
rect 88800 33800 88880 33810
rect 87060 33780 87140 33790
rect 87210 33780 87290 33790
rect 87360 33780 87440 33790
rect 87140 33700 87150 33780
rect 87290 33700 87300 33780
rect 87440 33700 87450 33780
rect 87820 33720 87830 33800
rect 88140 33720 88150 33800
rect 88560 33720 88570 33800
rect 88880 33720 88890 33800
rect 89060 33780 89140 33790
rect 89210 33780 89290 33790
rect 89140 33700 89150 33780
rect 89290 33700 89300 33780
rect 87580 33640 87660 33650
rect 87900 33640 87980 33650
rect 88320 33640 88400 33650
rect 88640 33640 88720 33650
rect 87060 33600 87140 33610
rect 87210 33600 87290 33610
rect 87360 33600 87440 33610
rect 87140 33520 87150 33600
rect 87290 33520 87300 33600
rect 87440 33520 87450 33600
rect 87660 33560 87670 33640
rect 87980 33560 87990 33640
rect 88400 33560 88410 33640
rect 88720 33560 88730 33640
rect 89060 33600 89140 33610
rect 89210 33600 89290 33610
rect 89140 33520 89150 33600
rect 89290 33520 89300 33600
rect 87740 33480 87820 33490
rect 88060 33480 88140 33490
rect 88480 33480 88560 33490
rect 88800 33480 88880 33490
rect 87060 33420 87140 33430
rect 87210 33420 87290 33430
rect 87360 33420 87440 33430
rect 87140 33340 87150 33420
rect 87290 33340 87300 33420
rect 87440 33340 87450 33420
rect 87820 33400 87830 33480
rect 88140 33400 88150 33480
rect 88560 33400 88570 33480
rect 88880 33400 88890 33480
rect 89060 33420 89140 33430
rect 89210 33420 89290 33430
rect 89140 33340 89150 33420
rect 89290 33340 89300 33420
rect 87580 33320 87660 33330
rect 87900 33320 87980 33330
rect 88320 33320 88400 33330
rect 88640 33320 88720 33330
rect 87060 33240 87140 33250
rect 87210 33240 87290 33250
rect 87360 33240 87440 33250
rect 87660 33240 87670 33320
rect 87980 33240 87990 33320
rect 88400 33240 88410 33320
rect 88720 33240 88730 33320
rect 89060 33240 89140 33250
rect 89210 33240 89290 33250
rect 87140 33160 87150 33240
rect 87290 33160 87300 33240
rect 87440 33160 87450 33240
rect 87740 33160 87820 33170
rect 88060 33160 88140 33170
rect 88480 33160 88560 33170
rect 88800 33160 88880 33170
rect 89140 33160 89150 33240
rect 89290 33160 89300 33240
rect 87820 33080 87830 33160
rect 88140 33080 88150 33160
rect 88560 33080 88570 33160
rect 88880 33080 88890 33160
rect 87060 33060 87140 33070
rect 87210 33060 87290 33070
rect 87360 33060 87440 33070
rect 89060 33060 89140 33070
rect 89210 33060 89290 33070
rect 87140 32980 87150 33060
rect 87290 32980 87300 33060
rect 87440 32980 87450 33060
rect 87580 33000 87660 33010
rect 87900 33000 87980 33010
rect 88320 33000 88400 33010
rect 88640 33000 88720 33010
rect 87660 32920 87670 33000
rect 87980 32920 87990 33000
rect 88400 32920 88410 33000
rect 88720 32920 88730 33000
rect 89140 32980 89150 33060
rect 89290 32980 89300 33060
rect 87060 32880 87140 32890
rect 87210 32880 87290 32890
rect 87360 32880 87440 32890
rect 89060 32880 89140 32890
rect 89210 32880 89290 32890
rect 87140 32800 87150 32880
rect 87290 32800 87300 32880
rect 87440 32800 87450 32880
rect 87740 32840 87820 32850
rect 88060 32840 88140 32850
rect 88480 32840 88560 32850
rect 88800 32840 88880 32850
rect 87820 32760 87830 32840
rect 88140 32760 88150 32840
rect 88560 32760 88570 32840
rect 88880 32760 88890 32840
rect 89140 32800 89150 32880
rect 89290 32800 89300 32880
rect 87060 32700 87140 32710
rect 87210 32700 87290 32710
rect 87360 32700 87440 32710
rect 89060 32700 89140 32710
rect 89210 32700 89290 32710
rect 87140 32620 87150 32700
rect 87290 32620 87300 32700
rect 87440 32620 87450 32700
rect 87580 32680 87660 32690
rect 87900 32680 87980 32690
rect 88320 32680 88400 32690
rect 88640 32680 88720 32690
rect 87660 32600 87670 32680
rect 87980 32600 87990 32680
rect 88400 32600 88410 32680
rect 88720 32600 88730 32680
rect 89140 32620 89150 32700
rect 89290 32620 89300 32700
rect 87060 32520 87140 32530
rect 87210 32520 87290 32530
rect 87360 32520 87440 32530
rect 87740 32520 87820 32530
rect 88060 32520 88140 32530
rect 88480 32520 88560 32530
rect 88800 32520 88880 32530
rect 89060 32520 89140 32530
rect 89210 32520 89290 32530
rect 87140 32440 87150 32520
rect 87290 32440 87300 32520
rect 87440 32440 87450 32520
rect 87820 32440 87830 32520
rect 88140 32440 88150 32520
rect 88560 32440 88570 32520
rect 88880 32440 88890 32520
rect 89140 32440 89150 32520
rect 89290 32440 89300 32520
rect 87580 32360 87660 32370
rect 87900 32360 87980 32370
rect 88320 32360 88400 32370
rect 88640 32360 88720 32370
rect 87060 32340 87140 32350
rect 87210 32340 87290 32350
rect 87360 32340 87440 32350
rect 87140 32260 87150 32340
rect 87290 32260 87300 32340
rect 87440 32260 87450 32340
rect 87660 32280 87670 32360
rect 87980 32280 87990 32360
rect 88400 32280 88410 32360
rect 88720 32280 88730 32360
rect 89060 32340 89140 32350
rect 89210 32340 89290 32350
rect 89140 32260 89150 32340
rect 89290 32260 89300 32340
rect 87740 32200 87820 32210
rect 88060 32200 88140 32210
rect 88480 32200 88560 32210
rect 88800 32200 88880 32210
rect 87060 32160 87140 32170
rect 87210 32160 87290 32170
rect 87360 32160 87440 32170
rect 87140 32080 87150 32160
rect 87290 32080 87300 32160
rect 87440 32080 87450 32160
rect 87820 32120 87830 32200
rect 88140 32120 88150 32200
rect 88560 32120 88570 32200
rect 88880 32120 88890 32200
rect 89060 32160 89140 32170
rect 89210 32160 89290 32170
rect 89140 32080 89150 32160
rect 89290 32080 89300 32160
rect 87580 32040 87660 32050
rect 87900 32040 87980 32050
rect 88320 32040 88400 32050
rect 88640 32040 88720 32050
rect 87060 31980 87140 31990
rect 87210 31980 87290 31990
rect 87360 31980 87440 31990
rect 87140 31900 87150 31980
rect 87290 31900 87300 31980
rect 87440 31900 87450 31980
rect 87660 31960 87670 32040
rect 87980 31960 87990 32040
rect 88400 31960 88410 32040
rect 88720 31960 88730 32040
rect 89060 31980 89140 31990
rect 89210 31980 89290 31990
rect 89140 31900 89150 31980
rect 89290 31900 89300 31980
rect 87740 31880 87820 31890
rect 88060 31880 88140 31890
rect 88480 31880 88560 31890
rect 88800 31880 88880 31890
rect 87060 31800 87140 31810
rect 87210 31800 87290 31810
rect 87360 31800 87440 31810
rect 87820 31800 87830 31880
rect 88140 31800 88150 31880
rect 88560 31800 88570 31880
rect 88880 31800 88890 31880
rect 89060 31800 89140 31810
rect 89210 31800 89290 31810
rect 87140 31720 87150 31800
rect 87290 31720 87300 31800
rect 87440 31720 87450 31800
rect 87580 31720 87660 31730
rect 87900 31720 87980 31730
rect 88320 31720 88400 31730
rect 88640 31720 88720 31730
rect 89140 31720 89150 31800
rect 89290 31720 89300 31800
rect 87660 31640 87670 31720
rect 87980 31640 87990 31720
rect 88400 31640 88410 31720
rect 88720 31640 88730 31720
rect 87060 31620 87140 31630
rect 87210 31620 87290 31630
rect 87360 31620 87440 31630
rect 89060 31620 89140 31630
rect 89210 31620 89290 31630
rect 87140 31540 87150 31620
rect 87290 31540 87300 31620
rect 87440 31540 87450 31620
rect 87740 31560 87820 31570
rect 88060 31560 88140 31570
rect 88480 31560 88560 31570
rect 88800 31560 88880 31570
rect 87820 31480 87830 31560
rect 88140 31480 88150 31560
rect 88560 31480 88570 31560
rect 88880 31480 88890 31560
rect 89140 31540 89150 31620
rect 89290 31540 89300 31620
rect 87060 31440 87140 31450
rect 87210 31440 87290 31450
rect 87360 31440 87440 31450
rect 89060 31440 89140 31450
rect 89210 31440 89290 31450
rect 87140 31360 87150 31440
rect 87290 31360 87300 31440
rect 87440 31360 87450 31440
rect 87580 31400 87660 31410
rect 87900 31400 87980 31410
rect 88320 31400 88400 31410
rect 88640 31400 88720 31410
rect 87660 31320 87670 31400
rect 87980 31320 87990 31400
rect 88400 31320 88410 31400
rect 88720 31320 88730 31400
rect 89140 31360 89150 31440
rect 89290 31360 89300 31440
rect 87060 31260 87140 31270
rect 87210 31260 87290 31270
rect 87360 31260 87440 31270
rect 89060 31260 89140 31270
rect 89210 31260 89290 31270
rect 87140 31180 87150 31260
rect 87290 31180 87300 31260
rect 87440 31180 87450 31260
rect 87740 31240 87820 31250
rect 88060 31240 88140 31250
rect 88480 31240 88560 31250
rect 88800 31240 88880 31250
rect 87820 31160 87830 31240
rect 88140 31160 88150 31240
rect 88560 31160 88570 31240
rect 88880 31160 88890 31240
rect 89140 31180 89150 31260
rect 89290 31180 89300 31260
rect 100245 31100 100260 37190
rect 100640 37120 100650 37200
rect 100790 37120 100800 37200
rect 100940 37120 100950 37200
rect 101080 37160 101160 37170
rect 101400 37160 101480 37170
rect 101820 37160 101900 37170
rect 102140 37160 102220 37170
rect 101160 37080 101170 37160
rect 101480 37080 101490 37160
rect 101900 37080 101910 37160
rect 102220 37080 102230 37160
rect 102640 37120 102650 37200
rect 102790 37120 102800 37200
rect 103240 37100 103255 37190
rect 100560 37020 100640 37030
rect 100710 37020 100790 37030
rect 100860 37020 100940 37030
rect 102560 37020 102640 37030
rect 102710 37020 102790 37030
rect 100640 36940 100650 37020
rect 100790 36940 100800 37020
rect 100940 36940 100950 37020
rect 101240 37000 101320 37010
rect 101560 37000 101640 37010
rect 101980 37000 102060 37010
rect 102300 37000 102380 37010
rect 101320 36920 101330 37000
rect 101640 36920 101650 37000
rect 102060 36920 102070 37000
rect 102380 36920 102390 37000
rect 102640 36940 102650 37020
rect 102790 36940 102800 37020
rect 100560 36840 100640 36850
rect 100710 36840 100790 36850
rect 100860 36840 100940 36850
rect 101080 36840 101160 36850
rect 101400 36840 101480 36850
rect 101820 36840 101900 36850
rect 102140 36840 102220 36850
rect 102560 36840 102640 36850
rect 102710 36840 102790 36850
rect 100640 36760 100650 36840
rect 100790 36760 100800 36840
rect 100940 36760 100950 36840
rect 101160 36760 101170 36840
rect 101480 36760 101490 36840
rect 101900 36760 101910 36840
rect 102220 36760 102230 36840
rect 102640 36760 102650 36840
rect 102790 36760 102800 36840
rect 101240 36680 101320 36690
rect 101560 36680 101640 36690
rect 101980 36680 102060 36690
rect 102300 36680 102380 36690
rect 100560 36660 100640 36670
rect 100710 36660 100790 36670
rect 100860 36660 100940 36670
rect 100640 36580 100650 36660
rect 100790 36580 100800 36660
rect 100940 36580 100950 36660
rect 101320 36600 101330 36680
rect 101640 36600 101650 36680
rect 102060 36600 102070 36680
rect 102380 36600 102390 36680
rect 102560 36660 102640 36670
rect 102710 36660 102790 36670
rect 102640 36580 102650 36660
rect 102790 36580 102800 36660
rect 101080 36520 101160 36530
rect 101400 36520 101480 36530
rect 101820 36520 101900 36530
rect 102140 36520 102220 36530
rect 100560 36480 100640 36490
rect 100710 36480 100790 36490
rect 100860 36480 100940 36490
rect 100640 36400 100650 36480
rect 100790 36400 100800 36480
rect 100940 36400 100950 36480
rect 101160 36440 101170 36520
rect 101480 36440 101490 36520
rect 101900 36440 101910 36520
rect 102220 36440 102230 36520
rect 102560 36480 102640 36490
rect 102710 36480 102790 36490
rect 102640 36400 102650 36480
rect 102790 36400 102800 36480
rect 101240 36360 101320 36370
rect 101560 36360 101640 36370
rect 101980 36360 102060 36370
rect 102300 36360 102380 36370
rect 100560 36300 100640 36310
rect 100710 36300 100790 36310
rect 100860 36300 100940 36310
rect 100640 36220 100650 36300
rect 100790 36220 100800 36300
rect 100940 36220 100950 36300
rect 101320 36280 101330 36360
rect 101640 36280 101650 36360
rect 102060 36280 102070 36360
rect 102380 36280 102390 36360
rect 102560 36300 102640 36310
rect 102710 36300 102790 36310
rect 102640 36220 102650 36300
rect 102790 36220 102800 36300
rect 101080 36200 101160 36210
rect 101400 36200 101480 36210
rect 101820 36200 101900 36210
rect 102140 36200 102220 36210
rect 100560 36120 100640 36130
rect 100710 36120 100790 36130
rect 100860 36120 100940 36130
rect 101160 36120 101170 36200
rect 101480 36120 101490 36200
rect 101900 36120 101910 36200
rect 102220 36120 102230 36200
rect 102560 36120 102640 36130
rect 102710 36120 102790 36130
rect 100640 36040 100650 36120
rect 100790 36040 100800 36120
rect 100940 36040 100950 36120
rect 101240 36040 101320 36050
rect 101560 36040 101640 36050
rect 101980 36040 102060 36050
rect 102300 36040 102380 36050
rect 102640 36040 102650 36120
rect 102790 36040 102800 36120
rect 101320 35960 101330 36040
rect 101640 35960 101650 36040
rect 102060 35960 102070 36040
rect 102380 35960 102390 36040
rect 100560 35940 100640 35950
rect 100710 35940 100790 35950
rect 100860 35940 100940 35950
rect 102560 35940 102640 35950
rect 102710 35940 102790 35950
rect 100640 35860 100650 35940
rect 100790 35860 100800 35940
rect 100940 35860 100950 35940
rect 101080 35880 101160 35890
rect 101400 35880 101480 35890
rect 101820 35880 101900 35890
rect 102140 35880 102220 35890
rect 101160 35800 101170 35880
rect 101480 35800 101490 35880
rect 101900 35800 101910 35880
rect 102220 35800 102230 35880
rect 102640 35860 102650 35940
rect 102790 35860 102800 35940
rect 100560 35760 100640 35770
rect 100710 35760 100790 35770
rect 100860 35760 100940 35770
rect 102560 35760 102640 35770
rect 102710 35760 102790 35770
rect 100640 35680 100650 35760
rect 100790 35680 100800 35760
rect 100940 35680 100950 35760
rect 101240 35720 101320 35730
rect 101560 35720 101640 35730
rect 101980 35720 102060 35730
rect 102300 35720 102380 35730
rect 101320 35640 101330 35720
rect 101640 35640 101650 35720
rect 102060 35640 102070 35720
rect 102380 35640 102390 35720
rect 102640 35680 102650 35760
rect 102790 35680 102800 35760
rect 100560 35580 100640 35590
rect 100710 35580 100790 35590
rect 100860 35580 100940 35590
rect 102560 35580 102640 35590
rect 102710 35580 102790 35590
rect 100640 35500 100650 35580
rect 100790 35500 100800 35580
rect 100940 35500 100950 35580
rect 101080 35560 101160 35570
rect 101400 35560 101480 35570
rect 101820 35560 101900 35570
rect 102140 35560 102220 35570
rect 101160 35480 101170 35560
rect 101480 35480 101490 35560
rect 101900 35480 101910 35560
rect 102220 35480 102230 35560
rect 102640 35500 102650 35580
rect 102790 35500 102800 35580
rect 100560 35400 100640 35410
rect 100710 35400 100790 35410
rect 100860 35400 100940 35410
rect 101240 35400 101320 35410
rect 101560 35400 101640 35410
rect 101980 35400 102060 35410
rect 102300 35400 102380 35410
rect 102560 35400 102640 35410
rect 102710 35400 102790 35410
rect 100640 35320 100650 35400
rect 100790 35320 100800 35400
rect 100940 35320 100950 35400
rect 101320 35320 101330 35400
rect 101640 35320 101650 35400
rect 102060 35320 102070 35400
rect 102380 35320 102390 35400
rect 102640 35320 102650 35400
rect 102790 35320 102800 35400
rect 101080 35240 101160 35250
rect 101400 35240 101480 35250
rect 101820 35240 101900 35250
rect 102140 35240 102220 35250
rect 100560 35220 100640 35230
rect 100710 35220 100790 35230
rect 100860 35220 100940 35230
rect 100640 35140 100650 35220
rect 100790 35140 100800 35220
rect 100940 35140 100950 35220
rect 101160 35160 101170 35240
rect 101480 35160 101490 35240
rect 101900 35160 101910 35240
rect 102220 35160 102230 35240
rect 102560 35220 102640 35230
rect 102710 35220 102790 35230
rect 102640 35140 102650 35220
rect 102790 35140 102800 35220
rect 101240 35080 101320 35090
rect 101560 35080 101640 35090
rect 101980 35080 102060 35090
rect 102300 35080 102380 35090
rect 100560 35040 100640 35050
rect 100710 35040 100790 35050
rect 100860 35040 100940 35050
rect 100640 34960 100650 35040
rect 100790 34960 100800 35040
rect 100940 34960 100950 35040
rect 101320 35000 101330 35080
rect 101640 35000 101650 35080
rect 102060 35000 102070 35080
rect 102380 35000 102390 35080
rect 102560 35040 102640 35050
rect 102710 35040 102790 35050
rect 102640 34960 102650 35040
rect 102790 34960 102800 35040
rect 101080 34920 101160 34930
rect 101400 34920 101480 34930
rect 101820 34920 101900 34930
rect 102140 34920 102220 34930
rect 100560 34860 100640 34870
rect 100710 34860 100790 34870
rect 100860 34860 100940 34870
rect 100640 34780 100650 34860
rect 100790 34780 100800 34860
rect 100940 34780 100950 34860
rect 101160 34840 101170 34920
rect 101480 34840 101490 34920
rect 101900 34840 101910 34920
rect 102220 34840 102230 34920
rect 102560 34860 102640 34870
rect 102710 34860 102790 34870
rect 102640 34780 102650 34860
rect 102790 34780 102800 34860
rect 101240 34760 101320 34770
rect 101560 34760 101640 34770
rect 101980 34760 102060 34770
rect 102300 34760 102380 34770
rect 100560 34680 100640 34690
rect 100710 34680 100790 34690
rect 100860 34680 100940 34690
rect 101320 34680 101330 34760
rect 101640 34680 101650 34760
rect 102060 34680 102070 34760
rect 102380 34680 102390 34760
rect 102560 34680 102640 34690
rect 102710 34680 102790 34690
rect 100640 34600 100650 34680
rect 100790 34600 100800 34680
rect 100940 34600 100950 34680
rect 101080 34600 101160 34610
rect 101400 34600 101480 34610
rect 101820 34600 101900 34610
rect 102140 34600 102220 34610
rect 102640 34600 102650 34680
rect 102790 34600 102800 34680
rect 101160 34520 101170 34600
rect 101480 34520 101490 34600
rect 101900 34520 101910 34600
rect 102220 34520 102230 34600
rect 100560 34500 100640 34510
rect 100710 34500 100790 34510
rect 100860 34500 100940 34510
rect 102560 34500 102640 34510
rect 102710 34500 102790 34510
rect 100640 34420 100650 34500
rect 100790 34420 100800 34500
rect 100940 34420 100950 34500
rect 101240 34440 101320 34450
rect 101560 34440 101640 34450
rect 101980 34440 102060 34450
rect 102300 34440 102380 34450
rect 101320 34360 101330 34440
rect 101640 34360 101650 34440
rect 102060 34360 102070 34440
rect 102380 34360 102390 34440
rect 102640 34420 102650 34500
rect 102790 34420 102800 34500
rect 100560 34320 100640 34330
rect 100710 34320 100790 34330
rect 100860 34320 100940 34330
rect 102560 34320 102640 34330
rect 102710 34320 102790 34330
rect 100640 34240 100650 34320
rect 100790 34240 100800 34320
rect 100940 34240 100950 34320
rect 101080 34280 101160 34290
rect 101400 34280 101480 34290
rect 101820 34280 101900 34290
rect 102140 34280 102220 34290
rect 101160 34200 101170 34280
rect 101480 34200 101490 34280
rect 101900 34200 101910 34280
rect 102220 34200 102230 34280
rect 102640 34240 102650 34320
rect 102790 34240 102800 34320
rect 100560 34140 100640 34150
rect 100710 34140 100790 34150
rect 100860 34140 100940 34150
rect 102560 34140 102640 34150
rect 102710 34140 102790 34150
rect 100640 34060 100650 34140
rect 100790 34060 100800 34140
rect 100940 34060 100950 34140
rect 101240 34120 101320 34130
rect 101560 34120 101640 34130
rect 101980 34120 102060 34130
rect 102300 34120 102380 34130
rect 101320 34040 101330 34120
rect 101640 34040 101650 34120
rect 102060 34040 102070 34120
rect 102380 34040 102390 34120
rect 102640 34060 102650 34140
rect 102790 34060 102800 34140
rect 100560 33960 100640 33970
rect 100710 33960 100790 33970
rect 100860 33960 100940 33970
rect 101080 33960 101160 33970
rect 101400 33960 101480 33970
rect 101820 33960 101900 33970
rect 102140 33960 102220 33970
rect 102560 33960 102640 33970
rect 102710 33960 102790 33970
rect 100640 33880 100650 33960
rect 100790 33880 100800 33960
rect 100940 33880 100950 33960
rect 101160 33880 101170 33960
rect 101480 33880 101490 33960
rect 101900 33880 101910 33960
rect 102220 33880 102230 33960
rect 102640 33880 102650 33960
rect 102790 33880 102800 33960
rect 101240 33800 101320 33810
rect 101560 33800 101640 33810
rect 101980 33800 102060 33810
rect 102300 33800 102380 33810
rect 100560 33780 100640 33790
rect 100710 33780 100790 33790
rect 100860 33780 100940 33790
rect 100640 33700 100650 33780
rect 100790 33700 100800 33780
rect 100940 33700 100950 33780
rect 101320 33720 101330 33800
rect 101640 33720 101650 33800
rect 102060 33720 102070 33800
rect 102380 33720 102390 33800
rect 102560 33780 102640 33790
rect 102710 33780 102790 33790
rect 102640 33700 102650 33780
rect 102790 33700 102800 33780
rect 101080 33640 101160 33650
rect 101400 33640 101480 33650
rect 101820 33640 101900 33650
rect 102140 33640 102220 33650
rect 100560 33600 100640 33610
rect 100710 33600 100790 33610
rect 100860 33600 100940 33610
rect 100640 33520 100650 33600
rect 100790 33520 100800 33600
rect 100940 33520 100950 33600
rect 101160 33560 101170 33640
rect 101480 33560 101490 33640
rect 101900 33560 101910 33640
rect 102220 33560 102230 33640
rect 102560 33600 102640 33610
rect 102710 33600 102790 33610
rect 102640 33520 102650 33600
rect 102790 33520 102800 33600
rect 101240 33480 101320 33490
rect 101560 33480 101640 33490
rect 101980 33480 102060 33490
rect 102300 33480 102380 33490
rect 100560 33420 100640 33430
rect 100710 33420 100790 33430
rect 100860 33420 100940 33430
rect 100640 33340 100650 33420
rect 100790 33340 100800 33420
rect 100940 33340 100950 33420
rect 101320 33400 101330 33480
rect 101640 33400 101650 33480
rect 102060 33400 102070 33480
rect 102380 33400 102390 33480
rect 102560 33420 102640 33430
rect 102710 33420 102790 33430
rect 102640 33340 102650 33420
rect 102790 33340 102800 33420
rect 101080 33320 101160 33330
rect 101400 33320 101480 33330
rect 101820 33320 101900 33330
rect 102140 33320 102220 33330
rect 100560 33240 100640 33250
rect 100710 33240 100790 33250
rect 100860 33240 100940 33250
rect 101160 33240 101170 33320
rect 101480 33240 101490 33320
rect 101900 33240 101910 33320
rect 102220 33240 102230 33320
rect 102560 33240 102640 33250
rect 102710 33240 102790 33250
rect 100640 33160 100650 33240
rect 100790 33160 100800 33240
rect 100940 33160 100950 33240
rect 101240 33160 101320 33170
rect 101560 33160 101640 33170
rect 101980 33160 102060 33170
rect 102300 33160 102380 33170
rect 102640 33160 102650 33240
rect 102790 33160 102800 33240
rect 101320 33080 101330 33160
rect 101640 33080 101650 33160
rect 102060 33080 102070 33160
rect 102380 33080 102390 33160
rect 100560 33060 100640 33070
rect 100710 33060 100790 33070
rect 100860 33060 100940 33070
rect 102560 33060 102640 33070
rect 102710 33060 102790 33070
rect 100640 32980 100650 33060
rect 100790 32980 100800 33060
rect 100940 32980 100950 33060
rect 101080 33000 101160 33010
rect 101400 33000 101480 33010
rect 101820 33000 101900 33010
rect 102140 33000 102220 33010
rect 101160 32920 101170 33000
rect 101480 32920 101490 33000
rect 101900 32920 101910 33000
rect 102220 32920 102230 33000
rect 102640 32980 102650 33060
rect 102790 32980 102800 33060
rect 100560 32880 100640 32890
rect 100710 32880 100790 32890
rect 100860 32880 100940 32890
rect 102560 32880 102640 32890
rect 102710 32880 102790 32890
rect 100640 32800 100650 32880
rect 100790 32800 100800 32880
rect 100940 32800 100950 32880
rect 101240 32840 101320 32850
rect 101560 32840 101640 32850
rect 101980 32840 102060 32850
rect 102300 32840 102380 32850
rect 101320 32760 101330 32840
rect 101640 32760 101650 32840
rect 102060 32760 102070 32840
rect 102380 32760 102390 32840
rect 102640 32800 102650 32880
rect 102790 32800 102800 32880
rect 100560 32700 100640 32710
rect 100710 32700 100790 32710
rect 100860 32700 100940 32710
rect 102560 32700 102640 32710
rect 102710 32700 102790 32710
rect 100640 32620 100650 32700
rect 100790 32620 100800 32700
rect 100940 32620 100950 32700
rect 101080 32680 101160 32690
rect 101400 32680 101480 32690
rect 101820 32680 101900 32690
rect 102140 32680 102220 32690
rect 101160 32600 101170 32680
rect 101480 32600 101490 32680
rect 101900 32600 101910 32680
rect 102220 32600 102230 32680
rect 102640 32620 102650 32700
rect 102790 32620 102800 32700
rect 100560 32520 100640 32530
rect 100710 32520 100790 32530
rect 100860 32520 100940 32530
rect 101240 32520 101320 32530
rect 101560 32520 101640 32530
rect 101980 32520 102060 32530
rect 102300 32520 102380 32530
rect 102560 32520 102640 32530
rect 102710 32520 102790 32530
rect 100640 32440 100650 32520
rect 100790 32440 100800 32520
rect 100940 32440 100950 32520
rect 101320 32440 101330 32520
rect 101640 32440 101650 32520
rect 102060 32440 102070 32520
rect 102380 32440 102390 32520
rect 102640 32440 102650 32520
rect 102790 32440 102800 32520
rect 101080 32360 101160 32370
rect 101400 32360 101480 32370
rect 101820 32360 101900 32370
rect 102140 32360 102220 32370
rect 100560 32340 100640 32350
rect 100710 32340 100790 32350
rect 100860 32340 100940 32350
rect 100640 32260 100650 32340
rect 100790 32260 100800 32340
rect 100940 32260 100950 32340
rect 101160 32280 101170 32360
rect 101480 32280 101490 32360
rect 101900 32280 101910 32360
rect 102220 32280 102230 32360
rect 102560 32340 102640 32350
rect 102710 32340 102790 32350
rect 102640 32260 102650 32340
rect 102790 32260 102800 32340
rect 101240 32200 101320 32210
rect 101560 32200 101640 32210
rect 101980 32200 102060 32210
rect 102300 32200 102380 32210
rect 100560 32160 100640 32170
rect 100710 32160 100790 32170
rect 100860 32160 100940 32170
rect 100640 32080 100650 32160
rect 100790 32080 100800 32160
rect 100940 32080 100950 32160
rect 101320 32120 101330 32200
rect 101640 32120 101650 32200
rect 102060 32120 102070 32200
rect 102380 32120 102390 32200
rect 102560 32160 102640 32170
rect 102710 32160 102790 32170
rect 102640 32080 102650 32160
rect 102790 32080 102800 32160
rect 101080 32040 101160 32050
rect 101400 32040 101480 32050
rect 101820 32040 101900 32050
rect 102140 32040 102220 32050
rect 100560 31980 100640 31990
rect 100710 31980 100790 31990
rect 100860 31980 100940 31990
rect 100640 31900 100650 31980
rect 100790 31900 100800 31980
rect 100940 31900 100950 31980
rect 101160 31960 101170 32040
rect 101480 31960 101490 32040
rect 101900 31960 101910 32040
rect 102220 31960 102230 32040
rect 102560 31980 102640 31990
rect 102710 31980 102790 31990
rect 102640 31900 102650 31980
rect 102790 31900 102800 31980
rect 101240 31880 101320 31890
rect 101560 31880 101640 31890
rect 101980 31880 102060 31890
rect 102300 31880 102380 31890
rect 100560 31800 100640 31810
rect 100710 31800 100790 31810
rect 100860 31800 100940 31810
rect 101320 31800 101330 31880
rect 101640 31800 101650 31880
rect 102060 31800 102070 31880
rect 102380 31800 102390 31880
rect 102560 31800 102640 31810
rect 102710 31800 102790 31810
rect 100640 31720 100650 31800
rect 100790 31720 100800 31800
rect 100940 31720 100950 31800
rect 101080 31720 101160 31730
rect 101400 31720 101480 31730
rect 101820 31720 101900 31730
rect 102140 31720 102220 31730
rect 102640 31720 102650 31800
rect 102790 31720 102800 31800
rect 101160 31640 101170 31720
rect 101480 31640 101490 31720
rect 101900 31640 101910 31720
rect 102220 31640 102230 31720
rect 100560 31620 100640 31630
rect 100710 31620 100790 31630
rect 100860 31620 100940 31630
rect 102560 31620 102640 31630
rect 102710 31620 102790 31630
rect 100640 31540 100650 31620
rect 100790 31540 100800 31620
rect 100940 31540 100950 31620
rect 101240 31560 101320 31570
rect 101560 31560 101640 31570
rect 101980 31560 102060 31570
rect 102300 31560 102380 31570
rect 101320 31480 101330 31560
rect 101640 31480 101650 31560
rect 102060 31480 102070 31560
rect 102380 31480 102390 31560
rect 102640 31540 102650 31620
rect 102790 31540 102800 31620
rect 100560 31440 100640 31450
rect 100710 31440 100790 31450
rect 100860 31440 100940 31450
rect 102560 31440 102640 31450
rect 102710 31440 102790 31450
rect 100640 31360 100650 31440
rect 100790 31360 100800 31440
rect 100940 31360 100950 31440
rect 101080 31400 101160 31410
rect 101400 31400 101480 31410
rect 101820 31400 101900 31410
rect 102140 31400 102220 31410
rect 101160 31320 101170 31400
rect 101480 31320 101490 31400
rect 101900 31320 101910 31400
rect 102220 31320 102230 31400
rect 102640 31360 102650 31440
rect 102790 31360 102800 31440
rect 100560 31260 100640 31270
rect 100710 31260 100790 31270
rect 100860 31260 100940 31270
rect 102560 31260 102640 31270
rect 102710 31260 102790 31270
rect 100640 31180 100650 31260
rect 100790 31180 100800 31260
rect 100940 31180 100950 31260
rect 101240 31240 101320 31250
rect 101560 31240 101640 31250
rect 101980 31240 102060 31250
rect 102300 31240 102380 31250
rect 101320 31160 101330 31240
rect 101640 31160 101650 31240
rect 102060 31160 102070 31240
rect 102380 31160 102390 31240
rect 102640 31180 102650 31260
rect 102790 31180 102800 31260
rect 113745 31100 113760 37190
rect 114140 37120 114150 37200
rect 114290 37120 114300 37200
rect 114440 37120 114450 37200
rect 114580 37160 114660 37170
rect 114900 37160 114980 37170
rect 115320 37160 115400 37170
rect 115640 37160 115720 37170
rect 114660 37080 114670 37160
rect 114980 37080 114990 37160
rect 115400 37080 115410 37160
rect 115720 37080 115730 37160
rect 116140 37120 116150 37200
rect 116290 37120 116300 37200
rect 116740 37100 116755 37190
rect 114060 37020 114140 37030
rect 114210 37020 114290 37030
rect 114360 37020 114440 37030
rect 116060 37020 116140 37030
rect 116210 37020 116290 37030
rect 114140 36940 114150 37020
rect 114290 36940 114300 37020
rect 114440 36940 114450 37020
rect 114740 37000 114820 37010
rect 115060 37000 115140 37010
rect 115480 37000 115560 37010
rect 115800 37000 115880 37010
rect 114820 36920 114830 37000
rect 115140 36920 115150 37000
rect 115560 36920 115570 37000
rect 115880 36920 115890 37000
rect 116140 36940 116150 37020
rect 116290 36940 116300 37020
rect 114060 36840 114140 36850
rect 114210 36840 114290 36850
rect 114360 36840 114440 36850
rect 114580 36840 114660 36850
rect 114900 36840 114980 36850
rect 115320 36840 115400 36850
rect 115640 36840 115720 36850
rect 116060 36840 116140 36850
rect 116210 36840 116290 36850
rect 114140 36760 114150 36840
rect 114290 36760 114300 36840
rect 114440 36760 114450 36840
rect 114660 36760 114670 36840
rect 114980 36760 114990 36840
rect 115400 36760 115410 36840
rect 115720 36760 115730 36840
rect 116140 36760 116150 36840
rect 116290 36760 116300 36840
rect 114740 36680 114820 36690
rect 115060 36680 115140 36690
rect 115480 36680 115560 36690
rect 115800 36680 115880 36690
rect 114060 36660 114140 36670
rect 114210 36660 114290 36670
rect 114360 36660 114440 36670
rect 114140 36580 114150 36660
rect 114290 36580 114300 36660
rect 114440 36580 114450 36660
rect 114820 36600 114830 36680
rect 115140 36600 115150 36680
rect 115560 36600 115570 36680
rect 115880 36600 115890 36680
rect 116060 36660 116140 36670
rect 116210 36660 116290 36670
rect 116140 36580 116150 36660
rect 116290 36580 116300 36660
rect 114580 36520 114660 36530
rect 114900 36520 114980 36530
rect 115320 36520 115400 36530
rect 115640 36520 115720 36530
rect 114060 36480 114140 36490
rect 114210 36480 114290 36490
rect 114360 36480 114440 36490
rect 114140 36400 114150 36480
rect 114290 36400 114300 36480
rect 114440 36400 114450 36480
rect 114660 36440 114670 36520
rect 114980 36440 114990 36520
rect 115400 36440 115410 36520
rect 115720 36440 115730 36520
rect 116060 36480 116140 36490
rect 116210 36480 116290 36490
rect 116140 36400 116150 36480
rect 116290 36400 116300 36480
rect 114740 36360 114820 36370
rect 115060 36360 115140 36370
rect 115480 36360 115560 36370
rect 115800 36360 115880 36370
rect 114060 36300 114140 36310
rect 114210 36300 114290 36310
rect 114360 36300 114440 36310
rect 114140 36220 114150 36300
rect 114290 36220 114300 36300
rect 114440 36220 114450 36300
rect 114820 36280 114830 36360
rect 115140 36280 115150 36360
rect 115560 36280 115570 36360
rect 115880 36280 115890 36360
rect 116060 36300 116140 36310
rect 116210 36300 116290 36310
rect 116140 36220 116150 36300
rect 116290 36220 116300 36300
rect 114580 36200 114660 36210
rect 114900 36200 114980 36210
rect 115320 36200 115400 36210
rect 115640 36200 115720 36210
rect 114060 36120 114140 36130
rect 114210 36120 114290 36130
rect 114360 36120 114440 36130
rect 114660 36120 114670 36200
rect 114980 36120 114990 36200
rect 115400 36120 115410 36200
rect 115720 36120 115730 36200
rect 116060 36120 116140 36130
rect 116210 36120 116290 36130
rect 114140 36040 114150 36120
rect 114290 36040 114300 36120
rect 114440 36040 114450 36120
rect 114740 36040 114820 36050
rect 115060 36040 115140 36050
rect 115480 36040 115560 36050
rect 115800 36040 115880 36050
rect 116140 36040 116150 36120
rect 116290 36040 116300 36120
rect 114820 35960 114830 36040
rect 115140 35960 115150 36040
rect 115560 35960 115570 36040
rect 115880 35960 115890 36040
rect 114060 35940 114140 35950
rect 114210 35940 114290 35950
rect 114360 35940 114440 35950
rect 116060 35940 116140 35950
rect 116210 35940 116290 35950
rect 114140 35860 114150 35940
rect 114290 35860 114300 35940
rect 114440 35860 114450 35940
rect 114580 35880 114660 35890
rect 114900 35880 114980 35890
rect 115320 35880 115400 35890
rect 115640 35880 115720 35890
rect 114660 35800 114670 35880
rect 114980 35800 114990 35880
rect 115400 35800 115410 35880
rect 115720 35800 115730 35880
rect 116140 35860 116150 35940
rect 116290 35860 116300 35940
rect 114060 35760 114140 35770
rect 114210 35760 114290 35770
rect 114360 35760 114440 35770
rect 116060 35760 116140 35770
rect 116210 35760 116290 35770
rect 114140 35680 114150 35760
rect 114290 35680 114300 35760
rect 114440 35680 114450 35760
rect 114740 35720 114820 35730
rect 115060 35720 115140 35730
rect 115480 35720 115560 35730
rect 115800 35720 115880 35730
rect 114820 35640 114830 35720
rect 115140 35640 115150 35720
rect 115560 35640 115570 35720
rect 115880 35640 115890 35720
rect 116140 35680 116150 35760
rect 116290 35680 116300 35760
rect 114060 35580 114140 35590
rect 114210 35580 114290 35590
rect 114360 35580 114440 35590
rect 116060 35580 116140 35590
rect 116210 35580 116290 35590
rect 114140 35500 114150 35580
rect 114290 35500 114300 35580
rect 114440 35500 114450 35580
rect 114580 35560 114660 35570
rect 114900 35560 114980 35570
rect 115320 35560 115400 35570
rect 115640 35560 115720 35570
rect 114660 35480 114670 35560
rect 114980 35480 114990 35560
rect 115400 35480 115410 35560
rect 115720 35480 115730 35560
rect 116140 35500 116150 35580
rect 116290 35500 116300 35580
rect 114060 35400 114140 35410
rect 114210 35400 114290 35410
rect 114360 35400 114440 35410
rect 114740 35400 114820 35410
rect 115060 35400 115140 35410
rect 115480 35400 115560 35410
rect 115800 35400 115880 35410
rect 116060 35400 116140 35410
rect 116210 35400 116290 35410
rect 114140 35320 114150 35400
rect 114290 35320 114300 35400
rect 114440 35320 114450 35400
rect 114820 35320 114830 35400
rect 115140 35320 115150 35400
rect 115560 35320 115570 35400
rect 115880 35320 115890 35400
rect 116140 35320 116150 35400
rect 116290 35320 116300 35400
rect 114580 35240 114660 35250
rect 114900 35240 114980 35250
rect 115320 35240 115400 35250
rect 115640 35240 115720 35250
rect 114060 35220 114140 35230
rect 114210 35220 114290 35230
rect 114360 35220 114440 35230
rect 114140 35140 114150 35220
rect 114290 35140 114300 35220
rect 114440 35140 114450 35220
rect 114660 35160 114670 35240
rect 114980 35160 114990 35240
rect 115400 35160 115410 35240
rect 115720 35160 115730 35240
rect 116060 35220 116140 35230
rect 116210 35220 116290 35230
rect 116140 35140 116150 35220
rect 116290 35140 116300 35220
rect 114740 35080 114820 35090
rect 115060 35080 115140 35090
rect 115480 35080 115560 35090
rect 115800 35080 115880 35090
rect 114060 35040 114140 35050
rect 114210 35040 114290 35050
rect 114360 35040 114440 35050
rect 114140 34960 114150 35040
rect 114290 34960 114300 35040
rect 114440 34960 114450 35040
rect 114820 35000 114830 35080
rect 115140 35000 115150 35080
rect 115560 35000 115570 35080
rect 115880 35000 115890 35080
rect 116060 35040 116140 35050
rect 116210 35040 116290 35050
rect 116140 34960 116150 35040
rect 116290 34960 116300 35040
rect 114580 34920 114660 34930
rect 114900 34920 114980 34930
rect 115320 34920 115400 34930
rect 115640 34920 115720 34930
rect 114060 34860 114140 34870
rect 114210 34860 114290 34870
rect 114360 34860 114440 34870
rect 114140 34780 114150 34860
rect 114290 34780 114300 34860
rect 114440 34780 114450 34860
rect 114660 34840 114670 34920
rect 114980 34840 114990 34920
rect 115400 34840 115410 34920
rect 115720 34840 115730 34920
rect 116060 34860 116140 34870
rect 116210 34860 116290 34870
rect 116140 34780 116150 34860
rect 116290 34780 116300 34860
rect 114740 34760 114820 34770
rect 115060 34760 115140 34770
rect 115480 34760 115560 34770
rect 115800 34760 115880 34770
rect 114060 34680 114140 34690
rect 114210 34680 114290 34690
rect 114360 34680 114440 34690
rect 114820 34680 114830 34760
rect 115140 34680 115150 34760
rect 115560 34680 115570 34760
rect 115880 34680 115890 34760
rect 116060 34680 116140 34690
rect 116210 34680 116290 34690
rect 114140 34600 114150 34680
rect 114290 34600 114300 34680
rect 114440 34600 114450 34680
rect 114580 34600 114660 34610
rect 114900 34600 114980 34610
rect 115320 34600 115400 34610
rect 115640 34600 115720 34610
rect 116140 34600 116150 34680
rect 116290 34600 116300 34680
rect 114660 34520 114670 34600
rect 114980 34520 114990 34600
rect 115400 34520 115410 34600
rect 115720 34520 115730 34600
rect 114060 34500 114140 34510
rect 114210 34500 114290 34510
rect 114360 34500 114440 34510
rect 116060 34500 116140 34510
rect 116210 34500 116290 34510
rect 114140 34420 114150 34500
rect 114290 34420 114300 34500
rect 114440 34420 114450 34500
rect 114740 34440 114820 34450
rect 115060 34440 115140 34450
rect 115480 34440 115560 34450
rect 115800 34440 115880 34450
rect 114820 34360 114830 34440
rect 115140 34360 115150 34440
rect 115560 34360 115570 34440
rect 115880 34360 115890 34440
rect 116140 34420 116150 34500
rect 116290 34420 116300 34500
rect 114060 34320 114140 34330
rect 114210 34320 114290 34330
rect 114360 34320 114440 34330
rect 116060 34320 116140 34330
rect 116210 34320 116290 34330
rect 114140 34240 114150 34320
rect 114290 34240 114300 34320
rect 114440 34240 114450 34320
rect 114580 34280 114660 34290
rect 114900 34280 114980 34290
rect 115320 34280 115400 34290
rect 115640 34280 115720 34290
rect 114660 34200 114670 34280
rect 114980 34200 114990 34280
rect 115400 34200 115410 34280
rect 115720 34200 115730 34280
rect 116140 34240 116150 34320
rect 116290 34240 116300 34320
rect 114060 34140 114140 34150
rect 114210 34140 114290 34150
rect 114360 34140 114440 34150
rect 116060 34140 116140 34150
rect 116210 34140 116290 34150
rect 114140 34060 114150 34140
rect 114290 34060 114300 34140
rect 114440 34060 114450 34140
rect 114740 34120 114820 34130
rect 115060 34120 115140 34130
rect 115480 34120 115560 34130
rect 115800 34120 115880 34130
rect 114820 34040 114830 34120
rect 115140 34040 115150 34120
rect 115560 34040 115570 34120
rect 115880 34040 115890 34120
rect 116140 34060 116150 34140
rect 116290 34060 116300 34140
rect 114060 33960 114140 33970
rect 114210 33960 114290 33970
rect 114360 33960 114440 33970
rect 114580 33960 114660 33970
rect 114900 33960 114980 33970
rect 115320 33960 115400 33970
rect 115640 33960 115720 33970
rect 116060 33960 116140 33970
rect 116210 33960 116290 33970
rect 114140 33880 114150 33960
rect 114290 33880 114300 33960
rect 114440 33880 114450 33960
rect 114660 33880 114670 33960
rect 114980 33880 114990 33960
rect 115400 33880 115410 33960
rect 115720 33880 115730 33960
rect 116140 33880 116150 33960
rect 116290 33880 116300 33960
rect 114740 33800 114820 33810
rect 115060 33800 115140 33810
rect 115480 33800 115560 33810
rect 115800 33800 115880 33810
rect 114060 33780 114140 33790
rect 114210 33780 114290 33790
rect 114360 33780 114440 33790
rect 114140 33700 114150 33780
rect 114290 33700 114300 33780
rect 114440 33700 114450 33780
rect 114820 33720 114830 33800
rect 115140 33720 115150 33800
rect 115560 33720 115570 33800
rect 115880 33720 115890 33800
rect 116060 33780 116140 33790
rect 116210 33780 116290 33790
rect 116140 33700 116150 33780
rect 116290 33700 116300 33780
rect 114580 33640 114660 33650
rect 114900 33640 114980 33650
rect 115320 33640 115400 33650
rect 115640 33640 115720 33650
rect 114060 33600 114140 33610
rect 114210 33600 114290 33610
rect 114360 33600 114440 33610
rect 114140 33520 114150 33600
rect 114290 33520 114300 33600
rect 114440 33520 114450 33600
rect 114660 33560 114670 33640
rect 114980 33560 114990 33640
rect 115400 33560 115410 33640
rect 115720 33560 115730 33640
rect 116060 33600 116140 33610
rect 116210 33600 116290 33610
rect 116140 33520 116150 33600
rect 116290 33520 116300 33600
rect 114740 33480 114820 33490
rect 115060 33480 115140 33490
rect 115480 33480 115560 33490
rect 115800 33480 115880 33490
rect 114060 33420 114140 33430
rect 114210 33420 114290 33430
rect 114360 33420 114440 33430
rect 114140 33340 114150 33420
rect 114290 33340 114300 33420
rect 114440 33340 114450 33420
rect 114820 33400 114830 33480
rect 115140 33400 115150 33480
rect 115560 33400 115570 33480
rect 115880 33400 115890 33480
rect 116060 33420 116140 33430
rect 116210 33420 116290 33430
rect 116140 33340 116150 33420
rect 116290 33340 116300 33420
rect 114580 33320 114660 33330
rect 114900 33320 114980 33330
rect 115320 33320 115400 33330
rect 115640 33320 115720 33330
rect 114060 33240 114140 33250
rect 114210 33240 114290 33250
rect 114360 33240 114440 33250
rect 114660 33240 114670 33320
rect 114980 33240 114990 33320
rect 115400 33240 115410 33320
rect 115720 33240 115730 33320
rect 116060 33240 116140 33250
rect 116210 33240 116290 33250
rect 114140 33160 114150 33240
rect 114290 33160 114300 33240
rect 114440 33160 114450 33240
rect 114740 33160 114820 33170
rect 115060 33160 115140 33170
rect 115480 33160 115560 33170
rect 115800 33160 115880 33170
rect 116140 33160 116150 33240
rect 116290 33160 116300 33240
rect 114820 33080 114830 33160
rect 115140 33080 115150 33160
rect 115560 33080 115570 33160
rect 115880 33080 115890 33160
rect 114060 33060 114140 33070
rect 114210 33060 114290 33070
rect 114360 33060 114440 33070
rect 116060 33060 116140 33070
rect 116210 33060 116290 33070
rect 114140 32980 114150 33060
rect 114290 32980 114300 33060
rect 114440 32980 114450 33060
rect 114580 33000 114660 33010
rect 114900 33000 114980 33010
rect 115320 33000 115400 33010
rect 115640 33000 115720 33010
rect 114660 32920 114670 33000
rect 114980 32920 114990 33000
rect 115400 32920 115410 33000
rect 115720 32920 115730 33000
rect 116140 32980 116150 33060
rect 116290 32980 116300 33060
rect 114060 32880 114140 32890
rect 114210 32880 114290 32890
rect 114360 32880 114440 32890
rect 116060 32880 116140 32890
rect 116210 32880 116290 32890
rect 114140 32800 114150 32880
rect 114290 32800 114300 32880
rect 114440 32800 114450 32880
rect 114740 32840 114820 32850
rect 115060 32840 115140 32850
rect 115480 32840 115560 32850
rect 115800 32840 115880 32850
rect 114820 32760 114830 32840
rect 115140 32760 115150 32840
rect 115560 32760 115570 32840
rect 115880 32760 115890 32840
rect 116140 32800 116150 32880
rect 116290 32800 116300 32880
rect 114060 32700 114140 32710
rect 114210 32700 114290 32710
rect 114360 32700 114440 32710
rect 116060 32700 116140 32710
rect 116210 32700 116290 32710
rect 114140 32620 114150 32700
rect 114290 32620 114300 32700
rect 114440 32620 114450 32700
rect 114580 32680 114660 32690
rect 114900 32680 114980 32690
rect 115320 32680 115400 32690
rect 115640 32680 115720 32690
rect 114660 32600 114670 32680
rect 114980 32600 114990 32680
rect 115400 32600 115410 32680
rect 115720 32600 115730 32680
rect 116140 32620 116150 32700
rect 116290 32620 116300 32700
rect 114060 32520 114140 32530
rect 114210 32520 114290 32530
rect 114360 32520 114440 32530
rect 114740 32520 114820 32530
rect 115060 32520 115140 32530
rect 115480 32520 115560 32530
rect 115800 32520 115880 32530
rect 116060 32520 116140 32530
rect 116210 32520 116290 32530
rect 114140 32440 114150 32520
rect 114290 32440 114300 32520
rect 114440 32440 114450 32520
rect 114820 32440 114830 32520
rect 115140 32440 115150 32520
rect 115560 32440 115570 32520
rect 115880 32440 115890 32520
rect 116140 32440 116150 32520
rect 116290 32440 116300 32520
rect 114580 32360 114660 32370
rect 114900 32360 114980 32370
rect 115320 32360 115400 32370
rect 115640 32360 115720 32370
rect 114060 32340 114140 32350
rect 114210 32340 114290 32350
rect 114360 32340 114440 32350
rect 114140 32260 114150 32340
rect 114290 32260 114300 32340
rect 114440 32260 114450 32340
rect 114660 32280 114670 32360
rect 114980 32280 114990 32360
rect 115400 32280 115410 32360
rect 115720 32280 115730 32360
rect 116060 32340 116140 32350
rect 116210 32340 116290 32350
rect 116140 32260 116150 32340
rect 116290 32260 116300 32340
rect 114740 32200 114820 32210
rect 115060 32200 115140 32210
rect 115480 32200 115560 32210
rect 115800 32200 115880 32210
rect 114060 32160 114140 32170
rect 114210 32160 114290 32170
rect 114360 32160 114440 32170
rect 114140 32080 114150 32160
rect 114290 32080 114300 32160
rect 114440 32080 114450 32160
rect 114820 32120 114830 32200
rect 115140 32120 115150 32200
rect 115560 32120 115570 32200
rect 115880 32120 115890 32200
rect 116060 32160 116140 32170
rect 116210 32160 116290 32170
rect 116140 32080 116150 32160
rect 116290 32080 116300 32160
rect 114580 32040 114660 32050
rect 114900 32040 114980 32050
rect 115320 32040 115400 32050
rect 115640 32040 115720 32050
rect 114060 31980 114140 31990
rect 114210 31980 114290 31990
rect 114360 31980 114440 31990
rect 114140 31900 114150 31980
rect 114290 31900 114300 31980
rect 114440 31900 114450 31980
rect 114660 31960 114670 32040
rect 114980 31960 114990 32040
rect 115400 31960 115410 32040
rect 115720 31960 115730 32040
rect 116060 31980 116140 31990
rect 116210 31980 116290 31990
rect 116140 31900 116150 31980
rect 116290 31900 116300 31980
rect 114740 31880 114820 31890
rect 115060 31880 115140 31890
rect 115480 31880 115560 31890
rect 115800 31880 115880 31890
rect 114060 31800 114140 31810
rect 114210 31800 114290 31810
rect 114360 31800 114440 31810
rect 114820 31800 114830 31880
rect 115140 31800 115150 31880
rect 115560 31800 115570 31880
rect 115880 31800 115890 31880
rect 116060 31800 116140 31810
rect 116210 31800 116290 31810
rect 114140 31720 114150 31800
rect 114290 31720 114300 31800
rect 114440 31720 114450 31800
rect 114580 31720 114660 31730
rect 114900 31720 114980 31730
rect 115320 31720 115400 31730
rect 115640 31720 115720 31730
rect 116140 31720 116150 31800
rect 116290 31720 116300 31800
rect 114660 31640 114670 31720
rect 114980 31640 114990 31720
rect 115400 31640 115410 31720
rect 115720 31640 115730 31720
rect 114060 31620 114140 31630
rect 114210 31620 114290 31630
rect 114360 31620 114440 31630
rect 116060 31620 116140 31630
rect 116210 31620 116290 31630
rect 114140 31540 114150 31620
rect 114290 31540 114300 31620
rect 114440 31540 114450 31620
rect 114740 31560 114820 31570
rect 115060 31560 115140 31570
rect 115480 31560 115560 31570
rect 115800 31560 115880 31570
rect 114820 31480 114830 31560
rect 115140 31480 115150 31560
rect 115560 31480 115570 31560
rect 115880 31480 115890 31560
rect 116140 31540 116150 31620
rect 116290 31540 116300 31620
rect 114060 31440 114140 31450
rect 114210 31440 114290 31450
rect 114360 31440 114440 31450
rect 116060 31440 116140 31450
rect 116210 31440 116290 31450
rect 114140 31360 114150 31440
rect 114290 31360 114300 31440
rect 114440 31360 114450 31440
rect 114580 31400 114660 31410
rect 114900 31400 114980 31410
rect 115320 31400 115400 31410
rect 115640 31400 115720 31410
rect 114660 31320 114670 31400
rect 114980 31320 114990 31400
rect 115400 31320 115410 31400
rect 115720 31320 115730 31400
rect 116140 31360 116150 31440
rect 116290 31360 116300 31440
rect 114060 31260 114140 31270
rect 114210 31260 114290 31270
rect 114360 31260 114440 31270
rect 116060 31260 116140 31270
rect 116210 31260 116290 31270
rect 114140 31180 114150 31260
rect 114290 31180 114300 31260
rect 114440 31180 114450 31260
rect 114740 31240 114820 31250
rect 115060 31240 115140 31250
rect 115480 31240 115560 31250
rect 115800 31240 115880 31250
rect 114820 31160 114830 31240
rect 115140 31160 115150 31240
rect 115560 31160 115570 31240
rect 115880 31160 115890 31240
rect 116140 31180 116150 31260
rect 116290 31180 116300 31260
rect 127245 31100 127260 37190
rect 127640 37120 127650 37200
rect 127790 37120 127800 37200
rect 127940 37120 127950 37200
rect 128080 37160 128160 37170
rect 128400 37160 128480 37170
rect 128820 37160 128900 37170
rect 129140 37160 129220 37170
rect 128160 37080 128170 37160
rect 128480 37080 128490 37160
rect 128900 37080 128910 37160
rect 129220 37080 129230 37160
rect 129640 37120 129650 37200
rect 129790 37120 129800 37200
rect 130240 37100 130255 37190
rect 141140 37120 141150 37200
rect 141290 37120 141300 37200
rect 141440 37120 141450 37200
rect 127560 37020 127640 37030
rect 127710 37020 127790 37030
rect 127860 37020 127940 37030
rect 129560 37020 129640 37030
rect 129710 37020 129790 37030
rect 141060 37020 141140 37030
rect 141210 37020 141290 37030
rect 141360 37020 141440 37030
rect 127640 36940 127650 37020
rect 127790 36940 127800 37020
rect 127940 36940 127950 37020
rect 128240 37000 128320 37010
rect 128560 37000 128640 37010
rect 128980 37000 129060 37010
rect 129300 37000 129380 37010
rect 128320 36920 128330 37000
rect 128640 36920 128650 37000
rect 129060 36920 129070 37000
rect 129380 36920 129390 37000
rect 129640 36940 129650 37020
rect 129790 36940 129800 37020
rect 141140 36940 141150 37020
rect 141290 36940 141300 37020
rect 141440 36940 141450 37020
rect 127560 36840 127640 36850
rect 127710 36840 127790 36850
rect 127860 36840 127940 36850
rect 128080 36840 128160 36850
rect 128400 36840 128480 36850
rect 128820 36840 128900 36850
rect 129140 36840 129220 36850
rect 129560 36840 129640 36850
rect 129710 36840 129790 36850
rect 141060 36840 141140 36850
rect 141210 36840 141290 36850
rect 141360 36840 141440 36850
rect 127640 36760 127650 36840
rect 127790 36760 127800 36840
rect 127940 36760 127950 36840
rect 128160 36760 128170 36840
rect 128480 36760 128490 36840
rect 128900 36760 128910 36840
rect 129220 36760 129230 36840
rect 129640 36760 129650 36840
rect 129790 36760 129800 36840
rect 141140 36760 141150 36840
rect 141290 36760 141300 36840
rect 141440 36760 141450 36840
rect 128240 36680 128320 36690
rect 128560 36680 128640 36690
rect 128980 36680 129060 36690
rect 129300 36680 129380 36690
rect 127560 36660 127640 36670
rect 127710 36660 127790 36670
rect 127860 36660 127940 36670
rect 127640 36580 127650 36660
rect 127790 36580 127800 36660
rect 127940 36580 127950 36660
rect 128320 36600 128330 36680
rect 128640 36600 128650 36680
rect 129060 36600 129070 36680
rect 129380 36600 129390 36680
rect 129560 36660 129640 36670
rect 129710 36660 129790 36670
rect 141060 36660 141140 36670
rect 141210 36660 141290 36670
rect 141360 36660 141440 36670
rect 129640 36580 129650 36660
rect 129790 36580 129800 36660
rect 141140 36580 141150 36660
rect 141290 36580 141300 36660
rect 141440 36580 141450 36660
rect 128080 36520 128160 36530
rect 128400 36520 128480 36530
rect 128820 36520 128900 36530
rect 129140 36520 129220 36530
rect 127560 36480 127640 36490
rect 127710 36480 127790 36490
rect 127860 36480 127940 36490
rect 127640 36400 127650 36480
rect 127790 36400 127800 36480
rect 127940 36400 127950 36480
rect 128160 36440 128170 36520
rect 128480 36440 128490 36520
rect 128900 36440 128910 36520
rect 129220 36440 129230 36520
rect 129560 36480 129640 36490
rect 129710 36480 129790 36490
rect 141060 36480 141140 36490
rect 141210 36480 141290 36490
rect 141360 36480 141440 36490
rect 129640 36400 129650 36480
rect 129790 36400 129800 36480
rect 141140 36400 141150 36480
rect 141290 36400 141300 36480
rect 141440 36400 141450 36480
rect 128240 36360 128320 36370
rect 128560 36360 128640 36370
rect 128980 36360 129060 36370
rect 129300 36360 129380 36370
rect 127560 36300 127640 36310
rect 127710 36300 127790 36310
rect 127860 36300 127940 36310
rect 127640 36220 127650 36300
rect 127790 36220 127800 36300
rect 127940 36220 127950 36300
rect 128320 36280 128330 36360
rect 128640 36280 128650 36360
rect 129060 36280 129070 36360
rect 129380 36280 129390 36360
rect 129560 36300 129640 36310
rect 129710 36300 129790 36310
rect 141060 36300 141140 36310
rect 141210 36300 141290 36310
rect 141360 36300 141440 36310
rect 129640 36220 129650 36300
rect 129790 36220 129800 36300
rect 141140 36220 141150 36300
rect 141290 36220 141300 36300
rect 141440 36220 141450 36300
rect 128080 36200 128160 36210
rect 128400 36200 128480 36210
rect 128820 36200 128900 36210
rect 129140 36200 129220 36210
rect 127560 36120 127640 36130
rect 127710 36120 127790 36130
rect 127860 36120 127940 36130
rect 128160 36120 128170 36200
rect 128480 36120 128490 36200
rect 128900 36120 128910 36200
rect 129220 36120 129230 36200
rect 129560 36120 129640 36130
rect 129710 36120 129790 36130
rect 141060 36120 141140 36130
rect 141210 36120 141290 36130
rect 141360 36120 141440 36130
rect 127640 36040 127650 36120
rect 127790 36040 127800 36120
rect 127940 36040 127950 36120
rect 128240 36040 128320 36050
rect 128560 36040 128640 36050
rect 128980 36040 129060 36050
rect 129300 36040 129380 36050
rect 129640 36040 129650 36120
rect 129790 36040 129800 36120
rect 141140 36040 141150 36120
rect 141290 36040 141300 36120
rect 141440 36040 141450 36120
rect 128320 35960 128330 36040
rect 128640 35960 128650 36040
rect 129060 35960 129070 36040
rect 129380 35960 129390 36040
rect 127560 35940 127640 35950
rect 127710 35940 127790 35950
rect 127860 35940 127940 35950
rect 129560 35940 129640 35950
rect 129710 35940 129790 35950
rect 141060 35940 141140 35950
rect 141210 35940 141290 35950
rect 141360 35940 141440 35950
rect 127640 35860 127650 35940
rect 127790 35860 127800 35940
rect 127940 35860 127950 35940
rect 128080 35880 128160 35890
rect 128400 35880 128480 35890
rect 128820 35880 128900 35890
rect 129140 35880 129220 35890
rect 128160 35800 128170 35880
rect 128480 35800 128490 35880
rect 128900 35800 128910 35880
rect 129220 35800 129230 35880
rect 129640 35860 129650 35940
rect 129790 35860 129800 35940
rect 141140 35860 141150 35940
rect 141290 35860 141300 35940
rect 141440 35860 141450 35940
rect 127560 35760 127640 35770
rect 127710 35760 127790 35770
rect 127860 35760 127940 35770
rect 129560 35760 129640 35770
rect 129710 35760 129790 35770
rect 141060 35760 141140 35770
rect 141210 35760 141290 35770
rect 141360 35760 141440 35770
rect 127640 35680 127650 35760
rect 127790 35680 127800 35760
rect 127940 35680 127950 35760
rect 128240 35720 128320 35730
rect 128560 35720 128640 35730
rect 128980 35720 129060 35730
rect 129300 35720 129380 35730
rect 128320 35640 128330 35720
rect 128640 35640 128650 35720
rect 129060 35640 129070 35720
rect 129380 35640 129390 35720
rect 129640 35680 129650 35760
rect 129790 35680 129800 35760
rect 141140 35680 141150 35760
rect 141290 35680 141300 35760
rect 141440 35680 141450 35760
rect 127560 35580 127640 35590
rect 127710 35580 127790 35590
rect 127860 35580 127940 35590
rect 129560 35580 129640 35590
rect 129710 35580 129790 35590
rect 141060 35580 141140 35590
rect 141210 35580 141290 35590
rect 141360 35580 141440 35590
rect 127640 35500 127650 35580
rect 127790 35500 127800 35580
rect 127940 35500 127950 35580
rect 128080 35560 128160 35570
rect 128400 35560 128480 35570
rect 128820 35560 128900 35570
rect 129140 35560 129220 35570
rect 128160 35480 128170 35560
rect 128480 35480 128490 35560
rect 128900 35480 128910 35560
rect 129220 35480 129230 35560
rect 129640 35500 129650 35580
rect 129790 35500 129800 35580
rect 141140 35500 141150 35580
rect 141290 35500 141300 35580
rect 141440 35500 141450 35580
rect 127560 35400 127640 35410
rect 127710 35400 127790 35410
rect 127860 35400 127940 35410
rect 128240 35400 128320 35410
rect 128560 35400 128640 35410
rect 128980 35400 129060 35410
rect 129300 35400 129380 35410
rect 129560 35400 129640 35410
rect 129710 35400 129790 35410
rect 141060 35400 141140 35410
rect 141210 35400 141290 35410
rect 141360 35400 141440 35410
rect 127640 35320 127650 35400
rect 127790 35320 127800 35400
rect 127940 35320 127950 35400
rect 128320 35320 128330 35400
rect 128640 35320 128650 35400
rect 129060 35320 129070 35400
rect 129380 35320 129390 35400
rect 129640 35320 129650 35400
rect 129790 35320 129800 35400
rect 141140 35320 141150 35400
rect 141290 35320 141300 35400
rect 141440 35320 141450 35400
rect 128080 35240 128160 35250
rect 128400 35240 128480 35250
rect 128820 35240 128900 35250
rect 129140 35240 129220 35250
rect 127560 35220 127640 35230
rect 127710 35220 127790 35230
rect 127860 35220 127940 35230
rect 127640 35140 127650 35220
rect 127790 35140 127800 35220
rect 127940 35140 127950 35220
rect 128160 35160 128170 35240
rect 128480 35160 128490 35240
rect 128900 35160 128910 35240
rect 129220 35160 129230 35240
rect 129560 35220 129640 35230
rect 129710 35220 129790 35230
rect 141060 35220 141140 35230
rect 141210 35220 141290 35230
rect 141360 35220 141440 35230
rect 129640 35140 129650 35220
rect 129790 35140 129800 35220
rect 141140 35140 141150 35220
rect 141290 35140 141300 35220
rect 141440 35140 141450 35220
rect 128240 35080 128320 35090
rect 128560 35080 128640 35090
rect 128980 35080 129060 35090
rect 129300 35080 129380 35090
rect 127560 35040 127640 35050
rect 127710 35040 127790 35050
rect 127860 35040 127940 35050
rect 127640 34960 127650 35040
rect 127790 34960 127800 35040
rect 127940 34960 127950 35040
rect 128320 35000 128330 35080
rect 128640 35000 128650 35080
rect 129060 35000 129070 35080
rect 129380 35000 129390 35080
rect 129560 35040 129640 35050
rect 129710 35040 129790 35050
rect 141060 35040 141140 35050
rect 141210 35040 141290 35050
rect 141360 35040 141440 35050
rect 129640 34960 129650 35040
rect 129790 34960 129800 35040
rect 141140 34960 141150 35040
rect 141290 34960 141300 35040
rect 141440 34960 141450 35040
rect 128080 34920 128160 34930
rect 128400 34920 128480 34930
rect 128820 34920 128900 34930
rect 129140 34920 129220 34930
rect 127560 34860 127640 34870
rect 127710 34860 127790 34870
rect 127860 34860 127940 34870
rect 127640 34780 127650 34860
rect 127790 34780 127800 34860
rect 127940 34780 127950 34860
rect 128160 34840 128170 34920
rect 128480 34840 128490 34920
rect 128900 34840 128910 34920
rect 129220 34840 129230 34920
rect 129560 34860 129640 34870
rect 129710 34860 129790 34870
rect 141060 34860 141140 34870
rect 141210 34860 141290 34870
rect 141360 34860 141440 34870
rect 129640 34780 129650 34860
rect 129790 34780 129800 34860
rect 141140 34780 141150 34860
rect 141290 34780 141300 34860
rect 141440 34780 141450 34860
rect 128240 34760 128320 34770
rect 128560 34760 128640 34770
rect 128980 34760 129060 34770
rect 129300 34760 129380 34770
rect 127560 34680 127640 34690
rect 127710 34680 127790 34690
rect 127860 34680 127940 34690
rect 128320 34680 128330 34760
rect 128640 34680 128650 34760
rect 129060 34680 129070 34760
rect 129380 34680 129390 34760
rect 129560 34680 129640 34690
rect 129710 34680 129790 34690
rect 141060 34680 141140 34690
rect 141210 34680 141290 34690
rect 141360 34680 141440 34690
rect 127640 34600 127650 34680
rect 127790 34600 127800 34680
rect 127940 34600 127950 34680
rect 128080 34600 128160 34610
rect 128400 34600 128480 34610
rect 128820 34600 128900 34610
rect 129140 34600 129220 34610
rect 129640 34600 129650 34680
rect 129790 34600 129800 34680
rect 141140 34600 141150 34680
rect 141290 34600 141300 34680
rect 141440 34600 141450 34680
rect 128160 34520 128170 34600
rect 128480 34520 128490 34600
rect 128900 34520 128910 34600
rect 129220 34520 129230 34600
rect 127560 34500 127640 34510
rect 127710 34500 127790 34510
rect 127860 34500 127940 34510
rect 129560 34500 129640 34510
rect 129710 34500 129790 34510
rect 141060 34500 141140 34510
rect 141210 34500 141290 34510
rect 141360 34500 141440 34510
rect 127640 34420 127650 34500
rect 127790 34420 127800 34500
rect 127940 34420 127950 34500
rect 128240 34440 128320 34450
rect 128560 34440 128640 34450
rect 128980 34440 129060 34450
rect 129300 34440 129380 34450
rect 128320 34360 128330 34440
rect 128640 34360 128650 34440
rect 129060 34360 129070 34440
rect 129380 34360 129390 34440
rect 129640 34420 129650 34500
rect 129790 34420 129800 34500
rect 141140 34420 141150 34500
rect 141290 34420 141300 34500
rect 141440 34420 141450 34500
rect 127560 34320 127640 34330
rect 127710 34320 127790 34330
rect 127860 34320 127940 34330
rect 129560 34320 129640 34330
rect 129710 34320 129790 34330
rect 141060 34320 141140 34330
rect 141210 34320 141290 34330
rect 141360 34320 141440 34330
rect 127640 34240 127650 34320
rect 127790 34240 127800 34320
rect 127940 34240 127950 34320
rect 128080 34280 128160 34290
rect 128400 34280 128480 34290
rect 128820 34280 128900 34290
rect 129140 34280 129220 34290
rect 128160 34200 128170 34280
rect 128480 34200 128490 34280
rect 128900 34200 128910 34280
rect 129220 34200 129230 34280
rect 129640 34240 129650 34320
rect 129790 34240 129800 34320
rect 141140 34240 141150 34320
rect 141290 34240 141300 34320
rect 141440 34240 141450 34320
rect 127560 34140 127640 34150
rect 127710 34140 127790 34150
rect 127860 34140 127940 34150
rect 129560 34140 129640 34150
rect 129710 34140 129790 34150
rect 141060 34140 141140 34150
rect 141210 34140 141290 34150
rect 141360 34140 141440 34150
rect 127640 34060 127650 34140
rect 127790 34060 127800 34140
rect 127940 34060 127950 34140
rect 128240 34120 128320 34130
rect 128560 34120 128640 34130
rect 128980 34120 129060 34130
rect 129300 34120 129380 34130
rect 128320 34040 128330 34120
rect 128640 34040 128650 34120
rect 129060 34040 129070 34120
rect 129380 34040 129390 34120
rect 129640 34060 129650 34140
rect 129790 34060 129800 34140
rect 141140 34060 141150 34140
rect 141290 34060 141300 34140
rect 141440 34060 141450 34140
rect 127560 33960 127640 33970
rect 127710 33960 127790 33970
rect 127860 33960 127940 33970
rect 128080 33960 128160 33970
rect 128400 33960 128480 33970
rect 128820 33960 128900 33970
rect 129140 33960 129220 33970
rect 129560 33960 129640 33970
rect 129710 33960 129790 33970
rect 141060 33960 141140 33970
rect 141210 33960 141290 33970
rect 141360 33960 141440 33970
rect 127640 33880 127650 33960
rect 127790 33880 127800 33960
rect 127940 33880 127950 33960
rect 128160 33880 128170 33960
rect 128480 33880 128490 33960
rect 128900 33880 128910 33960
rect 129220 33880 129230 33960
rect 129640 33880 129650 33960
rect 129790 33880 129800 33960
rect 141140 33880 141150 33960
rect 141290 33880 141300 33960
rect 141440 33880 141450 33960
rect 128240 33800 128320 33810
rect 128560 33800 128640 33810
rect 128980 33800 129060 33810
rect 129300 33800 129380 33810
rect 127560 33780 127640 33790
rect 127710 33780 127790 33790
rect 127860 33780 127940 33790
rect 127640 33700 127650 33780
rect 127790 33700 127800 33780
rect 127940 33700 127950 33780
rect 128320 33720 128330 33800
rect 128640 33720 128650 33800
rect 129060 33720 129070 33800
rect 129380 33720 129390 33800
rect 129560 33780 129640 33790
rect 129710 33780 129790 33790
rect 141060 33780 141140 33790
rect 141210 33780 141290 33790
rect 141360 33780 141440 33790
rect 129640 33700 129650 33780
rect 129790 33700 129800 33780
rect 141140 33700 141150 33780
rect 141290 33700 141300 33780
rect 141440 33700 141450 33780
rect 128080 33640 128160 33650
rect 128400 33640 128480 33650
rect 128820 33640 128900 33650
rect 129140 33640 129220 33650
rect 127560 33600 127640 33610
rect 127710 33600 127790 33610
rect 127860 33600 127940 33610
rect 127640 33520 127650 33600
rect 127790 33520 127800 33600
rect 127940 33520 127950 33600
rect 128160 33560 128170 33640
rect 128480 33560 128490 33640
rect 128900 33560 128910 33640
rect 129220 33560 129230 33640
rect 129560 33600 129640 33610
rect 129710 33600 129790 33610
rect 141060 33600 141140 33610
rect 141210 33600 141290 33610
rect 141360 33600 141440 33610
rect 129640 33520 129650 33600
rect 129790 33520 129800 33600
rect 141140 33520 141150 33600
rect 141290 33520 141300 33600
rect 141440 33520 141450 33600
rect 128240 33480 128320 33490
rect 128560 33480 128640 33490
rect 128980 33480 129060 33490
rect 129300 33480 129380 33490
rect 127560 33420 127640 33430
rect 127710 33420 127790 33430
rect 127860 33420 127940 33430
rect 127640 33340 127650 33420
rect 127790 33340 127800 33420
rect 127940 33340 127950 33420
rect 128320 33400 128330 33480
rect 128640 33400 128650 33480
rect 129060 33400 129070 33480
rect 129380 33400 129390 33480
rect 129560 33420 129640 33430
rect 129710 33420 129790 33430
rect 141060 33420 141140 33430
rect 141210 33420 141290 33430
rect 141360 33420 141440 33430
rect 129640 33340 129650 33420
rect 129790 33340 129800 33420
rect 141140 33340 141150 33420
rect 141290 33340 141300 33420
rect 141440 33340 141450 33420
rect 128080 33320 128160 33330
rect 128400 33320 128480 33330
rect 128820 33320 128900 33330
rect 129140 33320 129220 33330
rect 127560 33240 127640 33250
rect 127710 33240 127790 33250
rect 127860 33240 127940 33250
rect 128160 33240 128170 33320
rect 128480 33240 128490 33320
rect 128900 33240 128910 33320
rect 129220 33240 129230 33320
rect 129560 33240 129640 33250
rect 129710 33240 129790 33250
rect 141060 33240 141140 33250
rect 141210 33240 141290 33250
rect 141360 33240 141440 33250
rect 127640 33160 127650 33240
rect 127790 33160 127800 33240
rect 127940 33160 127950 33240
rect 128240 33160 128320 33170
rect 128560 33160 128640 33170
rect 128980 33160 129060 33170
rect 129300 33160 129380 33170
rect 129640 33160 129650 33240
rect 129790 33160 129800 33240
rect 141140 33160 141150 33240
rect 141290 33160 141300 33240
rect 141440 33160 141450 33240
rect 128320 33080 128330 33160
rect 128640 33080 128650 33160
rect 129060 33080 129070 33160
rect 129380 33080 129390 33160
rect 127560 33060 127640 33070
rect 127710 33060 127790 33070
rect 127860 33060 127940 33070
rect 129560 33060 129640 33070
rect 129710 33060 129790 33070
rect 141060 33060 141140 33070
rect 141210 33060 141290 33070
rect 141360 33060 141440 33070
rect 127640 32980 127650 33060
rect 127790 32980 127800 33060
rect 127940 32980 127950 33060
rect 128080 33000 128160 33010
rect 128400 33000 128480 33010
rect 128820 33000 128900 33010
rect 129140 33000 129220 33010
rect 128160 32920 128170 33000
rect 128480 32920 128490 33000
rect 128900 32920 128910 33000
rect 129220 32920 129230 33000
rect 129640 32980 129650 33060
rect 129790 32980 129800 33060
rect 141140 32980 141150 33060
rect 141290 32980 141300 33060
rect 141440 32980 141450 33060
rect 127560 32880 127640 32890
rect 127710 32880 127790 32890
rect 127860 32880 127940 32890
rect 129560 32880 129640 32890
rect 129710 32880 129790 32890
rect 141060 32880 141140 32890
rect 141210 32880 141290 32890
rect 141360 32880 141440 32890
rect 127640 32800 127650 32880
rect 127790 32800 127800 32880
rect 127940 32800 127950 32880
rect 128240 32840 128320 32850
rect 128560 32840 128640 32850
rect 128980 32840 129060 32850
rect 129300 32840 129380 32850
rect 128320 32760 128330 32840
rect 128640 32760 128650 32840
rect 129060 32760 129070 32840
rect 129380 32760 129390 32840
rect 129640 32800 129650 32880
rect 129790 32800 129800 32880
rect 141140 32800 141150 32880
rect 141290 32800 141300 32880
rect 141440 32800 141450 32880
rect 127560 32700 127640 32710
rect 127710 32700 127790 32710
rect 127860 32700 127940 32710
rect 129560 32700 129640 32710
rect 129710 32700 129790 32710
rect 141060 32700 141140 32710
rect 141210 32700 141290 32710
rect 141360 32700 141440 32710
rect 127640 32620 127650 32700
rect 127790 32620 127800 32700
rect 127940 32620 127950 32700
rect 128080 32680 128160 32690
rect 128400 32680 128480 32690
rect 128820 32680 128900 32690
rect 129140 32680 129220 32690
rect 128160 32600 128170 32680
rect 128480 32600 128490 32680
rect 128900 32600 128910 32680
rect 129220 32600 129230 32680
rect 129640 32620 129650 32700
rect 129790 32620 129800 32700
rect 141140 32620 141150 32700
rect 141290 32620 141300 32700
rect 141440 32620 141450 32700
rect 127560 32520 127640 32530
rect 127710 32520 127790 32530
rect 127860 32520 127940 32530
rect 128240 32520 128320 32530
rect 128560 32520 128640 32530
rect 128980 32520 129060 32530
rect 129300 32520 129380 32530
rect 129560 32520 129640 32530
rect 129710 32520 129790 32530
rect 141060 32520 141140 32530
rect 141210 32520 141290 32530
rect 141360 32520 141440 32530
rect 127640 32440 127650 32520
rect 127790 32440 127800 32520
rect 127940 32440 127950 32520
rect 128320 32440 128330 32520
rect 128640 32440 128650 32520
rect 129060 32440 129070 32520
rect 129380 32440 129390 32520
rect 129640 32440 129650 32520
rect 129790 32440 129800 32520
rect 141140 32440 141150 32520
rect 141290 32440 141300 32520
rect 141440 32440 141450 32520
rect 128080 32360 128160 32370
rect 128400 32360 128480 32370
rect 128820 32360 128900 32370
rect 129140 32360 129220 32370
rect 127560 32340 127640 32350
rect 127710 32340 127790 32350
rect 127860 32340 127940 32350
rect 127640 32260 127650 32340
rect 127790 32260 127800 32340
rect 127940 32260 127950 32340
rect 128160 32280 128170 32360
rect 128480 32280 128490 32360
rect 128900 32280 128910 32360
rect 129220 32280 129230 32360
rect 129560 32340 129640 32350
rect 129710 32340 129790 32350
rect 141060 32340 141140 32350
rect 141210 32340 141290 32350
rect 141360 32340 141440 32350
rect 129640 32260 129650 32340
rect 129790 32260 129800 32340
rect 141140 32260 141150 32340
rect 141290 32260 141300 32340
rect 141440 32260 141450 32340
rect 128240 32200 128320 32210
rect 128560 32200 128640 32210
rect 128980 32200 129060 32210
rect 129300 32200 129380 32210
rect 127560 32160 127640 32170
rect 127710 32160 127790 32170
rect 127860 32160 127940 32170
rect 127640 32080 127650 32160
rect 127790 32080 127800 32160
rect 127940 32080 127950 32160
rect 128320 32120 128330 32200
rect 128640 32120 128650 32200
rect 129060 32120 129070 32200
rect 129380 32120 129390 32200
rect 129560 32160 129640 32170
rect 129710 32160 129790 32170
rect 141060 32160 141140 32170
rect 141210 32160 141290 32170
rect 141360 32160 141440 32170
rect 129640 32080 129650 32160
rect 129790 32080 129800 32160
rect 141140 32080 141150 32160
rect 141290 32080 141300 32160
rect 141440 32080 141450 32160
rect 128080 32040 128160 32050
rect 128400 32040 128480 32050
rect 128820 32040 128900 32050
rect 129140 32040 129220 32050
rect 127560 31980 127640 31990
rect 127710 31980 127790 31990
rect 127860 31980 127940 31990
rect 127640 31900 127650 31980
rect 127790 31900 127800 31980
rect 127940 31900 127950 31980
rect 128160 31960 128170 32040
rect 128480 31960 128490 32040
rect 128900 31960 128910 32040
rect 129220 31960 129230 32040
rect 129560 31980 129640 31990
rect 129710 31980 129790 31990
rect 141060 31980 141140 31990
rect 141210 31980 141290 31990
rect 141360 31980 141440 31990
rect 129640 31900 129650 31980
rect 129790 31900 129800 31980
rect 141140 31900 141150 31980
rect 141290 31900 141300 31980
rect 141440 31900 141450 31980
rect 128240 31880 128320 31890
rect 128560 31880 128640 31890
rect 128980 31880 129060 31890
rect 129300 31880 129380 31890
rect 127560 31800 127640 31810
rect 127710 31800 127790 31810
rect 127860 31800 127940 31810
rect 128320 31800 128330 31880
rect 128640 31800 128650 31880
rect 129060 31800 129070 31880
rect 129380 31800 129390 31880
rect 129560 31800 129640 31810
rect 129710 31800 129790 31810
rect 141060 31800 141140 31810
rect 141210 31800 141290 31810
rect 141360 31800 141440 31810
rect 127640 31720 127650 31800
rect 127790 31720 127800 31800
rect 127940 31720 127950 31800
rect 128080 31720 128160 31730
rect 128400 31720 128480 31730
rect 128820 31720 128900 31730
rect 129140 31720 129220 31730
rect 129640 31720 129650 31800
rect 129790 31720 129800 31800
rect 141140 31720 141150 31800
rect 141290 31720 141300 31800
rect 141440 31720 141450 31800
rect 128160 31640 128170 31720
rect 128480 31640 128490 31720
rect 128900 31640 128910 31720
rect 129220 31640 129230 31720
rect 127560 31620 127640 31630
rect 127710 31620 127790 31630
rect 127860 31620 127940 31630
rect 129560 31620 129640 31630
rect 129710 31620 129790 31630
rect 141060 31620 141140 31630
rect 141210 31620 141290 31630
rect 141360 31620 141440 31630
rect 127640 31540 127650 31620
rect 127790 31540 127800 31620
rect 127940 31540 127950 31620
rect 128240 31560 128320 31570
rect 128560 31560 128640 31570
rect 128980 31560 129060 31570
rect 129300 31560 129380 31570
rect 128320 31480 128330 31560
rect 128640 31480 128650 31560
rect 129060 31480 129070 31560
rect 129380 31480 129390 31560
rect 129640 31540 129650 31620
rect 129790 31540 129800 31620
rect 141140 31540 141150 31620
rect 141290 31540 141300 31620
rect 141440 31540 141450 31620
rect 127560 31440 127640 31450
rect 127710 31440 127790 31450
rect 127860 31440 127940 31450
rect 129560 31440 129640 31450
rect 129710 31440 129790 31450
rect 141060 31440 141140 31450
rect 141210 31440 141290 31450
rect 141360 31440 141440 31450
rect 127640 31360 127650 31440
rect 127790 31360 127800 31440
rect 127940 31360 127950 31440
rect 128080 31400 128160 31410
rect 128400 31400 128480 31410
rect 128820 31400 128900 31410
rect 129140 31400 129220 31410
rect 128160 31320 128170 31400
rect 128480 31320 128490 31400
rect 128900 31320 128910 31400
rect 129220 31320 129230 31400
rect 129640 31360 129650 31440
rect 129790 31360 129800 31440
rect 141140 31360 141150 31440
rect 141290 31360 141300 31440
rect 141440 31360 141450 31440
rect 127560 31260 127640 31270
rect 127710 31260 127790 31270
rect 127860 31260 127940 31270
rect 129560 31260 129640 31270
rect 129710 31260 129790 31270
rect 141060 31260 141140 31270
rect 141210 31260 141290 31270
rect 141360 31260 141440 31270
rect 127640 31180 127650 31260
rect 127790 31180 127800 31260
rect 127940 31180 127950 31260
rect 128240 31240 128320 31250
rect 128560 31240 128640 31250
rect 128980 31240 129060 31250
rect 129300 31240 129380 31250
rect 128320 31160 128330 31240
rect 128640 31160 128650 31240
rect 129060 31160 129070 31240
rect 129380 31160 129390 31240
rect 129640 31180 129650 31260
rect 129790 31180 129800 31260
rect 141140 31180 141150 31260
rect 141290 31180 141300 31260
rect 141440 31180 141450 31260
rect 43785 31080 43865 31090
rect 44105 31080 44185 31090
rect 44425 31080 44505 31090
rect 44745 31080 44825 31090
rect 45065 31080 45145 31090
rect 45385 31080 45465 31090
rect 45705 31080 45785 31090
rect 46025 31080 46105 31090
rect 46345 31080 46425 31090
rect 46665 31080 46745 31090
rect 46985 31080 47065 31090
rect 47305 31080 47385 31090
rect 47625 31080 47705 31090
rect 47945 31080 48025 31090
rect 48265 31080 48345 31090
rect 48500 31080 48640 31090
rect 48710 31080 48790 31090
rect 60060 31080 60140 31090
rect 60210 31080 60290 31090
rect 60360 31080 60440 31090
rect 60580 31080 60660 31090
rect 60900 31080 60980 31090
rect 61320 31080 61400 31090
rect 61640 31080 61720 31090
rect 62060 31080 62140 31090
rect 62210 31080 62290 31090
rect 73560 31080 73640 31090
rect 73710 31080 73790 31090
rect 73860 31080 73940 31090
rect 74080 31080 74160 31090
rect 74400 31080 74480 31090
rect 74820 31080 74900 31090
rect 75140 31080 75220 31090
rect 75560 31080 75640 31090
rect 75710 31080 75790 31090
rect 87060 31080 87140 31090
rect 87210 31080 87290 31090
rect 87360 31080 87440 31090
rect 87580 31080 87660 31090
rect 87900 31080 87980 31090
rect 88320 31080 88400 31090
rect 88640 31080 88720 31090
rect 89060 31080 89140 31090
rect 89210 31080 89290 31090
rect 100560 31080 100640 31090
rect 100710 31080 100790 31090
rect 100860 31080 100940 31090
rect 101080 31080 101160 31090
rect 101400 31080 101480 31090
rect 101820 31080 101900 31090
rect 102140 31080 102220 31090
rect 102560 31080 102640 31090
rect 102710 31080 102790 31090
rect 114060 31080 114140 31090
rect 114210 31080 114290 31090
rect 114360 31080 114440 31090
rect 114580 31080 114660 31090
rect 114900 31080 114980 31090
rect 115320 31080 115400 31090
rect 115640 31080 115720 31090
rect 116060 31080 116140 31090
rect 116210 31080 116290 31090
rect 127560 31080 127640 31090
rect 127710 31080 127790 31090
rect 127860 31080 127940 31090
rect 128080 31080 128160 31090
rect 128400 31080 128480 31090
rect 128820 31080 128900 31090
rect 129140 31080 129220 31090
rect 129560 31080 129640 31090
rect 129710 31080 129790 31090
rect 141060 31080 141140 31090
rect 141210 31080 141290 31090
rect 141360 31080 141440 31090
rect 43865 31000 43875 31080
rect 44185 31000 44195 31080
rect 44505 31000 44515 31080
rect 44825 31000 44835 31080
rect 45145 31000 45155 31080
rect 45465 31000 45475 31080
rect 45785 31000 45795 31080
rect 46105 31000 46115 31080
rect 46425 31000 46435 31080
rect 46745 31000 46755 31080
rect 47065 31000 47075 31080
rect 47385 31000 47395 31080
rect 47705 31000 47715 31080
rect 48025 31000 48035 31080
rect 48345 31000 48355 31080
rect 43060 30980 43140 30990
rect 43380 30980 43460 30990
rect 43140 30900 43150 30980
rect 43460 30900 43470 30980
rect 43945 30920 44025 30930
rect 44265 30920 44345 30930
rect 44585 30920 44665 30930
rect 44905 30920 44985 30930
rect 45225 30920 45305 30930
rect 45545 30920 45625 30930
rect 45865 30920 45945 30930
rect 46185 30920 46265 30930
rect 46505 30920 46585 30930
rect 46825 30920 46905 30930
rect 47145 30920 47225 30930
rect 47465 30920 47545 30930
rect 47785 30920 47865 30930
rect 48105 30920 48185 30930
rect 44025 30840 44035 30920
rect 44345 30840 44355 30920
rect 44665 30840 44675 30920
rect 44985 30840 44995 30920
rect 45305 30840 45315 30920
rect 45625 30840 45635 30920
rect 45945 30840 45955 30920
rect 46265 30840 46275 30920
rect 46585 30840 46595 30920
rect 46905 30840 46915 30920
rect 47225 30840 47235 30920
rect 47545 30840 47555 30920
rect 47865 30840 47875 30920
rect 48185 30840 48195 30920
rect 48500 30910 48605 31080
rect 48640 31000 48650 31080
rect 48790 31000 48800 31080
rect 60140 31000 60150 31080
rect 60290 31000 60300 31080
rect 60440 31000 60450 31080
rect 60660 31000 60670 31080
rect 60980 31000 60990 31080
rect 61400 31000 61410 31080
rect 61720 31000 61730 31080
rect 62140 31000 62150 31080
rect 62290 31000 62300 31080
rect 73640 31000 73650 31080
rect 73790 31000 73800 31080
rect 73940 31000 73950 31080
rect 74160 31000 74170 31080
rect 74480 31000 74490 31080
rect 74900 31000 74910 31080
rect 75220 31000 75230 31080
rect 75640 31000 75650 31080
rect 75790 31000 75800 31080
rect 87140 31000 87150 31080
rect 87290 31000 87300 31080
rect 87440 31000 87450 31080
rect 87660 31000 87670 31080
rect 87980 31000 87990 31080
rect 88400 31000 88410 31080
rect 88720 31000 88730 31080
rect 89140 31000 89150 31080
rect 89290 31000 89300 31080
rect 100640 31000 100650 31080
rect 100790 31000 100800 31080
rect 100940 31000 100950 31080
rect 101160 31000 101170 31080
rect 101480 31000 101490 31080
rect 101900 31000 101910 31080
rect 102220 31000 102230 31080
rect 102640 31000 102650 31080
rect 102790 31000 102800 31080
rect 114140 31000 114150 31080
rect 114290 31000 114300 31080
rect 114440 31000 114450 31080
rect 114660 31000 114670 31080
rect 114980 31000 114990 31080
rect 115400 31000 115410 31080
rect 115720 31000 115730 31080
rect 116140 31000 116150 31080
rect 116290 31000 116300 31080
rect 127640 31000 127650 31080
rect 127790 31000 127800 31080
rect 127940 31000 127950 31080
rect 128160 31000 128170 31080
rect 128480 31000 128490 31080
rect 128900 31000 128910 31080
rect 129220 31000 129230 31080
rect 129640 31000 129650 31080
rect 129790 31000 129800 31080
rect 141140 31000 141150 31080
rect 141290 31000 141300 31080
rect 141440 31000 141450 31080
rect 60740 30920 60820 30930
rect 61060 30920 61140 30930
rect 61480 30920 61560 30930
rect 61800 30920 61880 30930
rect 74240 30920 74320 30930
rect 74560 30920 74640 30930
rect 74980 30920 75060 30930
rect 75300 30920 75380 30930
rect 87740 30920 87820 30930
rect 88060 30920 88140 30930
rect 88480 30920 88560 30930
rect 88800 30920 88880 30930
rect 101240 30920 101320 30930
rect 101560 30920 101640 30930
rect 101980 30920 102060 30930
rect 102300 30920 102380 30930
rect 114740 30920 114820 30930
rect 115060 30920 115140 30930
rect 115480 30920 115560 30930
rect 115800 30920 115880 30930
rect 128240 30920 128320 30930
rect 128560 30920 128640 30930
rect 128980 30920 129060 30930
rect 129300 30920 129380 30930
rect 48500 30900 48640 30910
rect 48710 30900 48790 30910
rect 60060 30900 60140 30910
rect 60210 30900 60290 30910
rect 60360 30900 60440 30910
rect 42950 30820 42980 30830
rect 43220 30820 43300 30830
rect 42980 30740 42990 30820
rect 43300 30740 43310 30820
rect 43785 30760 43865 30770
rect 44105 30760 44185 30770
rect 44425 30760 44505 30770
rect 44745 30760 44825 30770
rect 45065 30760 45145 30770
rect 45385 30760 45465 30770
rect 45705 30760 45785 30770
rect 46025 30760 46105 30770
rect 46345 30760 46425 30770
rect 46665 30760 46745 30770
rect 46985 30760 47065 30770
rect 47305 30760 47385 30770
rect 47625 30760 47705 30770
rect 47945 30760 48025 30770
rect 48265 30760 48345 30770
rect 43865 30680 43875 30760
rect 44185 30680 44195 30760
rect 44505 30680 44515 30760
rect 44825 30680 44835 30760
rect 45145 30680 45155 30760
rect 45465 30680 45475 30760
rect 45785 30680 45795 30760
rect 46105 30680 46115 30760
rect 46425 30680 46435 30760
rect 46745 30680 46755 30760
rect 47065 30680 47075 30760
rect 47385 30680 47395 30760
rect 47705 30680 47715 30760
rect 48025 30680 48035 30760
rect 48345 30680 48355 30760
rect 48500 30730 48605 30900
rect 48640 30820 48650 30900
rect 48790 30820 48800 30900
rect 60140 30820 60150 30900
rect 60290 30820 60300 30900
rect 60440 30820 60450 30900
rect 60820 30840 60830 30920
rect 61140 30840 61150 30920
rect 61560 30840 61570 30920
rect 61880 30840 61890 30920
rect 62060 30900 62140 30910
rect 62210 30900 62290 30910
rect 73560 30900 73640 30910
rect 73710 30900 73790 30910
rect 73860 30900 73940 30910
rect 62140 30820 62150 30900
rect 62290 30820 62300 30900
rect 73640 30820 73650 30900
rect 73790 30820 73800 30900
rect 73940 30820 73950 30900
rect 74320 30840 74330 30920
rect 74640 30840 74650 30920
rect 75060 30840 75070 30920
rect 75380 30840 75390 30920
rect 75560 30900 75640 30910
rect 75710 30900 75790 30910
rect 87060 30900 87140 30910
rect 87210 30900 87290 30910
rect 87360 30900 87440 30910
rect 75640 30820 75650 30900
rect 75790 30820 75800 30900
rect 87140 30820 87150 30900
rect 87290 30820 87300 30900
rect 87440 30820 87450 30900
rect 87820 30840 87830 30920
rect 88140 30840 88150 30920
rect 88560 30840 88570 30920
rect 88880 30840 88890 30920
rect 89060 30900 89140 30910
rect 89210 30900 89290 30910
rect 100560 30900 100640 30910
rect 100710 30900 100790 30910
rect 100860 30900 100940 30910
rect 89140 30820 89150 30900
rect 89290 30820 89300 30900
rect 100640 30820 100650 30900
rect 100790 30820 100800 30900
rect 100940 30820 100950 30900
rect 101320 30840 101330 30920
rect 101640 30840 101650 30920
rect 102060 30840 102070 30920
rect 102380 30840 102390 30920
rect 102560 30900 102640 30910
rect 102710 30900 102790 30910
rect 114060 30900 114140 30910
rect 114210 30900 114290 30910
rect 114360 30900 114440 30910
rect 102640 30820 102650 30900
rect 102790 30820 102800 30900
rect 114140 30820 114150 30900
rect 114290 30820 114300 30900
rect 114440 30820 114450 30900
rect 114820 30840 114830 30920
rect 115140 30840 115150 30920
rect 115560 30840 115570 30920
rect 115880 30840 115890 30920
rect 116060 30900 116140 30910
rect 116210 30900 116290 30910
rect 127560 30900 127640 30910
rect 127710 30900 127790 30910
rect 127860 30900 127940 30910
rect 116140 30820 116150 30900
rect 116290 30820 116300 30900
rect 127640 30820 127650 30900
rect 127790 30820 127800 30900
rect 127940 30820 127950 30900
rect 128320 30840 128330 30920
rect 128640 30840 128650 30920
rect 129060 30840 129070 30920
rect 129380 30840 129390 30920
rect 129560 30900 129640 30910
rect 129710 30900 129790 30910
rect 141060 30900 141140 30910
rect 141210 30900 141290 30910
rect 141360 30900 141440 30910
rect 129640 30820 129650 30900
rect 129790 30820 129800 30900
rect 141140 30820 141150 30900
rect 141290 30820 141300 30900
rect 141440 30820 141450 30900
rect 60580 30760 60660 30770
rect 60900 30760 60980 30770
rect 61320 30760 61400 30770
rect 61640 30760 61720 30770
rect 74080 30760 74160 30770
rect 74400 30760 74480 30770
rect 74820 30760 74900 30770
rect 75140 30760 75220 30770
rect 87580 30760 87660 30770
rect 87900 30760 87980 30770
rect 88320 30760 88400 30770
rect 88640 30760 88720 30770
rect 101080 30760 101160 30770
rect 101400 30760 101480 30770
rect 101820 30760 101900 30770
rect 102140 30760 102220 30770
rect 114580 30760 114660 30770
rect 114900 30760 114980 30770
rect 115320 30760 115400 30770
rect 115640 30760 115720 30770
rect 128080 30760 128160 30770
rect 128400 30760 128480 30770
rect 128820 30760 128900 30770
rect 129140 30760 129220 30770
rect 48500 30720 48640 30730
rect 48710 30720 48790 30730
rect 60060 30720 60140 30730
rect 60210 30720 60290 30730
rect 60360 30720 60440 30730
rect 43060 30660 43140 30670
rect 43380 30660 43460 30670
rect 43140 30580 43150 30660
rect 43460 30580 43470 30660
rect 43945 30600 44025 30610
rect 44265 30600 44345 30610
rect 44585 30600 44665 30610
rect 44905 30600 44985 30610
rect 45225 30600 45305 30610
rect 45545 30600 45625 30610
rect 45865 30600 45945 30610
rect 46185 30600 46265 30610
rect 46505 30600 46585 30610
rect 46825 30600 46905 30610
rect 47145 30600 47225 30610
rect 47465 30600 47545 30610
rect 47785 30600 47865 30610
rect 48105 30600 48185 30610
rect 44025 30520 44035 30600
rect 44345 30520 44355 30600
rect 44665 30520 44675 30600
rect 44985 30520 44995 30600
rect 45305 30520 45315 30600
rect 45625 30520 45635 30600
rect 45945 30520 45955 30600
rect 46265 30520 46275 30600
rect 46585 30520 46595 30600
rect 46905 30520 46915 30600
rect 47225 30520 47235 30600
rect 47545 30520 47555 30600
rect 47865 30520 47875 30600
rect 48185 30520 48195 30600
rect 48500 30550 48605 30720
rect 48640 30640 48650 30720
rect 48790 30640 48800 30720
rect 60140 30640 60150 30720
rect 60290 30640 60300 30720
rect 60440 30640 60450 30720
rect 60660 30680 60670 30760
rect 60980 30680 60990 30760
rect 61400 30680 61410 30760
rect 61720 30680 61730 30760
rect 62060 30720 62140 30730
rect 62210 30720 62290 30730
rect 73560 30720 73640 30730
rect 73710 30720 73790 30730
rect 73860 30720 73940 30730
rect 62140 30640 62150 30720
rect 62290 30640 62300 30720
rect 73640 30640 73650 30720
rect 73790 30640 73800 30720
rect 73940 30640 73950 30720
rect 74160 30680 74170 30760
rect 74480 30680 74490 30760
rect 74900 30680 74910 30760
rect 75220 30680 75230 30760
rect 75560 30720 75640 30730
rect 75710 30720 75790 30730
rect 87060 30720 87140 30730
rect 87210 30720 87290 30730
rect 87360 30720 87440 30730
rect 75640 30640 75650 30720
rect 75790 30640 75800 30720
rect 87140 30640 87150 30720
rect 87290 30640 87300 30720
rect 87440 30640 87450 30720
rect 87660 30680 87670 30760
rect 87980 30680 87990 30760
rect 88400 30680 88410 30760
rect 88720 30680 88730 30760
rect 89060 30720 89140 30730
rect 89210 30720 89290 30730
rect 100560 30720 100640 30730
rect 100710 30720 100790 30730
rect 100860 30720 100940 30730
rect 89140 30640 89150 30720
rect 89290 30640 89300 30720
rect 100640 30640 100650 30720
rect 100790 30640 100800 30720
rect 100940 30640 100950 30720
rect 101160 30680 101170 30760
rect 101480 30680 101490 30760
rect 101900 30680 101910 30760
rect 102220 30680 102230 30760
rect 102560 30720 102640 30730
rect 102710 30720 102790 30730
rect 114060 30720 114140 30730
rect 114210 30720 114290 30730
rect 114360 30720 114440 30730
rect 102640 30640 102650 30720
rect 102790 30640 102800 30720
rect 114140 30640 114150 30720
rect 114290 30640 114300 30720
rect 114440 30640 114450 30720
rect 114660 30680 114670 30760
rect 114980 30680 114990 30760
rect 115400 30680 115410 30760
rect 115720 30680 115730 30760
rect 116060 30720 116140 30730
rect 116210 30720 116290 30730
rect 127560 30720 127640 30730
rect 127710 30720 127790 30730
rect 127860 30720 127940 30730
rect 116140 30640 116150 30720
rect 116290 30640 116300 30720
rect 127640 30640 127650 30720
rect 127790 30640 127800 30720
rect 127940 30640 127950 30720
rect 128160 30680 128170 30760
rect 128480 30680 128490 30760
rect 128900 30680 128910 30760
rect 129220 30680 129230 30760
rect 129560 30720 129640 30730
rect 129710 30720 129790 30730
rect 141060 30720 141140 30730
rect 141210 30720 141290 30730
rect 141360 30720 141440 30730
rect 129640 30640 129650 30720
rect 129790 30640 129800 30720
rect 141140 30640 141150 30720
rect 141290 30640 141300 30720
rect 141440 30640 141450 30720
rect 60740 30600 60820 30610
rect 61060 30600 61140 30610
rect 61480 30600 61560 30610
rect 61800 30600 61880 30610
rect 74240 30600 74320 30610
rect 74560 30600 74640 30610
rect 74980 30600 75060 30610
rect 75300 30600 75380 30610
rect 87740 30600 87820 30610
rect 88060 30600 88140 30610
rect 88480 30600 88560 30610
rect 88800 30600 88880 30610
rect 101240 30600 101320 30610
rect 101560 30600 101640 30610
rect 101980 30600 102060 30610
rect 102300 30600 102380 30610
rect 114740 30600 114820 30610
rect 115060 30600 115140 30610
rect 115480 30600 115560 30610
rect 115800 30600 115880 30610
rect 128240 30600 128320 30610
rect 128560 30600 128640 30610
rect 128980 30600 129060 30610
rect 129300 30600 129380 30610
rect 49180 30570 49210 30600
rect 49300 30570 49330 30600
rect 49420 30570 49450 30600
rect 49540 30570 49570 30600
rect 49660 30570 49690 30600
rect 49780 30570 49810 30600
rect 49900 30570 49930 30600
rect 50020 30570 50050 30600
rect 50140 30570 50170 30600
rect 50260 30570 50290 30600
rect 50380 30570 50410 30600
rect 50500 30570 50530 30600
rect 50620 30570 50650 30600
rect 50740 30570 50770 30600
rect 50860 30570 50890 30600
rect 50980 30570 51010 30600
rect 51100 30570 51130 30600
rect 51220 30570 51250 30600
rect 51340 30570 51370 30600
rect 51460 30570 51490 30600
rect 51580 30570 51610 30600
rect 51700 30570 51730 30600
rect 51820 30570 51850 30600
rect 51940 30570 51970 30600
rect 52060 30570 52090 30600
rect 52180 30570 52210 30600
rect 52300 30570 52330 30600
rect 52420 30570 52450 30600
rect 52540 30570 52570 30600
rect 52660 30570 52690 30600
rect 52780 30570 52810 30600
rect 52900 30570 52930 30600
rect 53020 30570 53050 30600
rect 53140 30570 53170 30600
rect 53260 30570 53290 30600
rect 53380 30570 53410 30600
rect 53500 30570 53530 30600
rect 53620 30570 53650 30600
rect 53740 30570 53770 30600
rect 53860 30570 53890 30600
rect 53980 30570 54010 30600
rect 54100 30570 54130 30600
rect 54220 30570 54250 30600
rect 54340 30570 54370 30600
rect 54460 30570 54490 30600
rect 54580 30570 54610 30600
rect 54700 30570 54730 30600
rect 54820 30570 54850 30600
rect 54940 30570 54970 30600
rect 55060 30570 55090 30600
rect 55180 30570 55210 30600
rect 55300 30570 55330 30600
rect 55420 30570 55450 30600
rect 55540 30570 55570 30600
rect 55660 30570 55690 30600
rect 55780 30570 55810 30600
rect 55900 30570 55930 30600
rect 56020 30570 56050 30600
rect 56140 30570 56170 30600
rect 56260 30570 56290 30600
rect 56380 30570 56410 30600
rect 56500 30570 56530 30600
rect 56620 30570 56650 30600
rect 56740 30570 56770 30600
rect 56860 30570 56890 30600
rect 56980 30570 57010 30600
rect 57100 30570 57130 30600
rect 57220 30570 57250 30600
rect 57340 30570 57370 30600
rect 57460 30570 57490 30600
rect 57580 30570 57610 30600
rect 57700 30570 57730 30600
rect 57820 30570 57850 30600
rect 57940 30570 57970 30600
rect 58060 30570 58090 30600
rect 58180 30570 58210 30600
rect 58300 30570 58330 30600
rect 58420 30570 58450 30600
rect 58540 30570 58570 30600
rect 58660 30570 58690 30600
rect 58780 30570 58810 30600
rect 58900 30570 58930 30600
rect 59020 30570 59050 30600
rect 59140 30570 59170 30600
rect 59260 30570 59290 30600
rect 59380 30570 59410 30600
rect 59500 30570 59530 30600
rect 59620 30570 59650 30600
rect 59740 30570 59770 30600
rect 59860 30570 59890 30600
rect 48500 30540 48640 30550
rect 48710 30540 48790 30550
rect 49060 30540 49120 30570
rect 49180 30540 49240 30570
rect 49300 30540 49360 30570
rect 49420 30540 49480 30570
rect 49540 30540 49600 30570
rect 49660 30540 49720 30570
rect 49780 30540 49840 30570
rect 49900 30540 49960 30570
rect 50020 30540 50080 30570
rect 50140 30540 50200 30570
rect 50260 30540 50320 30570
rect 50380 30540 50440 30570
rect 50500 30540 50560 30570
rect 50620 30540 50680 30570
rect 50740 30540 50800 30570
rect 50860 30540 50920 30570
rect 50980 30540 51040 30570
rect 51100 30540 51160 30570
rect 51220 30540 51280 30570
rect 51340 30540 51400 30570
rect 51460 30540 51520 30570
rect 51580 30540 51640 30570
rect 51700 30540 51760 30570
rect 51820 30540 51880 30570
rect 51940 30540 52000 30570
rect 52060 30540 52120 30570
rect 52180 30540 52240 30570
rect 52300 30540 52360 30570
rect 52420 30540 52480 30570
rect 52540 30540 52600 30570
rect 52660 30540 52720 30570
rect 52780 30540 52840 30570
rect 52900 30540 52960 30570
rect 53020 30540 53080 30570
rect 53140 30540 53200 30570
rect 53260 30540 53320 30570
rect 53380 30540 53440 30570
rect 53500 30540 53560 30570
rect 53620 30540 53680 30570
rect 53740 30540 53800 30570
rect 53860 30540 53920 30570
rect 53980 30540 54040 30570
rect 54100 30540 54160 30570
rect 54220 30540 54280 30570
rect 54340 30540 54400 30570
rect 54460 30540 54520 30570
rect 54580 30540 54640 30570
rect 54700 30540 54760 30570
rect 54820 30540 54880 30570
rect 54940 30540 55000 30570
rect 55060 30540 55120 30570
rect 55180 30540 55240 30570
rect 55300 30540 55360 30570
rect 55420 30540 55480 30570
rect 55540 30540 55600 30570
rect 55660 30540 55720 30570
rect 55780 30540 55840 30570
rect 55900 30540 55960 30570
rect 56020 30540 56080 30570
rect 56140 30540 56200 30570
rect 56260 30540 56320 30570
rect 56380 30540 56440 30570
rect 56500 30540 56560 30570
rect 56620 30540 56680 30570
rect 56740 30540 56800 30570
rect 56860 30540 56920 30570
rect 56980 30540 57040 30570
rect 57100 30540 57160 30570
rect 57220 30540 57280 30570
rect 57340 30540 57400 30570
rect 57460 30540 57520 30570
rect 57580 30540 57640 30570
rect 57700 30540 57760 30570
rect 57820 30540 57880 30570
rect 57940 30540 58000 30570
rect 58060 30540 58120 30570
rect 58180 30540 58240 30570
rect 58300 30540 58360 30570
rect 58420 30540 58480 30570
rect 58540 30540 58600 30570
rect 58660 30540 58720 30570
rect 58780 30540 58840 30570
rect 58900 30540 58960 30570
rect 59020 30540 59080 30570
rect 59140 30540 59200 30570
rect 59260 30540 59320 30570
rect 59380 30540 59440 30570
rect 59500 30540 59560 30570
rect 59620 30540 59680 30570
rect 59740 30540 59800 30570
rect 59860 30540 59920 30570
rect 60060 30540 60140 30550
rect 60210 30540 60290 30550
rect 60360 30540 60440 30550
rect 42950 30500 42980 30510
rect 43220 30500 43300 30510
rect 42980 30420 42990 30500
rect 43300 30420 43310 30500
rect 43785 30440 43865 30450
rect 44105 30440 44185 30450
rect 44425 30440 44505 30450
rect 44745 30440 44825 30450
rect 45065 30440 45145 30450
rect 45385 30440 45465 30450
rect 45705 30440 45785 30450
rect 46025 30440 46105 30450
rect 46345 30440 46425 30450
rect 46665 30440 46745 30450
rect 46985 30440 47065 30450
rect 47305 30440 47385 30450
rect 47625 30440 47705 30450
rect 47945 30440 48025 30450
rect 48265 30440 48345 30450
rect 43865 30360 43875 30440
rect 44185 30360 44195 30440
rect 44505 30360 44515 30440
rect 44825 30360 44835 30440
rect 45145 30360 45155 30440
rect 45465 30360 45475 30440
rect 45785 30360 45795 30440
rect 46105 30360 46115 30440
rect 46425 30360 46435 30440
rect 46745 30360 46755 30440
rect 47065 30360 47075 30440
rect 47385 30360 47395 30440
rect 47705 30360 47715 30440
rect 48025 30360 48035 30440
rect 48345 30360 48355 30440
rect 48500 30370 48605 30540
rect 48640 30460 48650 30540
rect 48790 30460 48800 30540
rect 49180 30450 49210 30480
rect 49300 30450 49330 30480
rect 49420 30450 49450 30480
rect 49540 30450 49570 30480
rect 49660 30450 49690 30480
rect 49780 30450 49810 30480
rect 49900 30450 49930 30480
rect 50020 30450 50050 30480
rect 50140 30450 50170 30480
rect 50260 30450 50290 30480
rect 50380 30450 50410 30480
rect 50500 30450 50530 30480
rect 50620 30450 50650 30480
rect 50740 30450 50770 30480
rect 50860 30450 50890 30480
rect 50980 30450 51010 30480
rect 51100 30450 51130 30480
rect 51220 30450 51250 30480
rect 51340 30450 51370 30480
rect 51460 30450 51490 30480
rect 51580 30450 51610 30480
rect 51700 30450 51730 30480
rect 51820 30450 51850 30480
rect 51940 30450 51970 30480
rect 52060 30450 52090 30480
rect 52180 30450 52210 30480
rect 52300 30450 52330 30480
rect 52420 30450 52450 30480
rect 52540 30450 52570 30480
rect 52660 30450 52690 30480
rect 52780 30450 52810 30480
rect 52900 30450 52930 30480
rect 53020 30450 53050 30480
rect 53140 30450 53170 30480
rect 53260 30450 53290 30480
rect 53380 30450 53410 30480
rect 53500 30450 53530 30480
rect 53620 30450 53650 30480
rect 53740 30450 53770 30480
rect 53860 30450 53890 30480
rect 53980 30450 54010 30480
rect 54100 30450 54130 30480
rect 54220 30450 54250 30480
rect 54340 30450 54370 30480
rect 54460 30450 54490 30480
rect 54580 30450 54610 30480
rect 54700 30450 54730 30480
rect 54820 30450 54850 30480
rect 54940 30450 54970 30480
rect 55060 30450 55090 30480
rect 55180 30450 55210 30480
rect 55300 30450 55330 30480
rect 55420 30450 55450 30480
rect 55540 30450 55570 30480
rect 55660 30450 55690 30480
rect 55780 30450 55810 30480
rect 55900 30450 55930 30480
rect 56020 30450 56050 30480
rect 56140 30450 56170 30480
rect 56260 30450 56290 30480
rect 56380 30450 56410 30480
rect 56500 30450 56530 30480
rect 56620 30450 56650 30480
rect 56740 30450 56770 30480
rect 56860 30450 56890 30480
rect 56980 30450 57010 30480
rect 57100 30450 57130 30480
rect 57220 30450 57250 30480
rect 57340 30450 57370 30480
rect 57460 30450 57490 30480
rect 57580 30450 57610 30480
rect 57700 30450 57730 30480
rect 57820 30450 57850 30480
rect 57940 30450 57970 30480
rect 58060 30450 58090 30480
rect 58180 30450 58210 30480
rect 58300 30450 58330 30480
rect 58420 30450 58450 30480
rect 58540 30450 58570 30480
rect 58660 30450 58690 30480
rect 58780 30450 58810 30480
rect 58900 30450 58930 30480
rect 59020 30450 59050 30480
rect 59140 30450 59170 30480
rect 59260 30450 59290 30480
rect 59380 30450 59410 30480
rect 59500 30450 59530 30480
rect 59620 30450 59650 30480
rect 59740 30450 59770 30480
rect 59860 30450 59890 30480
rect 60140 30460 60150 30540
rect 60290 30460 60300 30540
rect 60440 30460 60450 30540
rect 60820 30520 60830 30600
rect 61140 30520 61150 30600
rect 61560 30520 61570 30600
rect 61880 30520 61890 30600
rect 62680 30570 62710 30600
rect 73245 30570 73270 30600
rect 73360 30570 73390 30600
rect 62060 30540 62140 30550
rect 62210 30540 62290 30550
rect 62560 30540 62620 30570
rect 62680 30540 62740 30570
rect 73245 30540 73300 30570
rect 73360 30540 73420 30570
rect 73560 30540 73640 30550
rect 73710 30540 73790 30550
rect 73860 30540 73940 30550
rect 62140 30460 62150 30540
rect 62290 30460 62300 30540
rect 62680 30450 62710 30480
rect 73245 30450 73270 30480
rect 73360 30450 73390 30480
rect 73640 30460 73650 30540
rect 73790 30460 73800 30540
rect 73940 30460 73950 30540
rect 74320 30520 74330 30600
rect 74640 30520 74650 30600
rect 75060 30520 75070 30600
rect 75380 30520 75390 30600
rect 76180 30570 76210 30600
rect 86745 30570 86770 30600
rect 86860 30570 86890 30600
rect 75560 30540 75640 30550
rect 75710 30540 75790 30550
rect 76060 30540 76120 30570
rect 76180 30540 76240 30570
rect 86745 30540 86800 30570
rect 86860 30540 86920 30570
rect 87060 30540 87140 30550
rect 87210 30540 87290 30550
rect 87360 30540 87440 30550
rect 75640 30460 75650 30540
rect 75790 30460 75800 30540
rect 76180 30450 76210 30480
rect 86745 30450 86770 30480
rect 86860 30450 86890 30480
rect 87140 30460 87150 30540
rect 87290 30460 87300 30540
rect 87440 30460 87450 30540
rect 87820 30520 87830 30600
rect 88140 30520 88150 30600
rect 88560 30520 88570 30600
rect 88880 30520 88890 30600
rect 89680 30570 89710 30600
rect 100245 30570 100270 30600
rect 100360 30570 100390 30600
rect 89060 30540 89140 30550
rect 89210 30540 89290 30550
rect 89560 30540 89620 30570
rect 89680 30540 89740 30570
rect 100245 30540 100300 30570
rect 100360 30540 100420 30570
rect 100560 30540 100640 30550
rect 100710 30540 100790 30550
rect 100860 30540 100940 30550
rect 89140 30460 89150 30540
rect 89290 30460 89300 30540
rect 89680 30450 89710 30480
rect 100245 30450 100270 30480
rect 100360 30450 100390 30480
rect 100640 30460 100650 30540
rect 100790 30460 100800 30540
rect 100940 30460 100950 30540
rect 101320 30520 101330 30600
rect 101640 30520 101650 30600
rect 102060 30520 102070 30600
rect 102380 30520 102390 30600
rect 103180 30570 103210 30600
rect 113745 30570 113770 30600
rect 113860 30570 113890 30600
rect 102560 30540 102640 30550
rect 102710 30540 102790 30550
rect 103060 30540 103120 30570
rect 103180 30540 103240 30570
rect 113745 30540 113800 30570
rect 113860 30540 113920 30570
rect 114060 30540 114140 30550
rect 114210 30540 114290 30550
rect 114360 30540 114440 30550
rect 102640 30460 102650 30540
rect 102790 30460 102800 30540
rect 103180 30450 103210 30480
rect 113745 30450 113770 30480
rect 113860 30450 113890 30480
rect 114140 30460 114150 30540
rect 114290 30460 114300 30540
rect 114440 30460 114450 30540
rect 114820 30520 114830 30600
rect 115140 30520 115150 30600
rect 115560 30520 115570 30600
rect 115880 30520 115890 30600
rect 116680 30570 116710 30600
rect 127245 30570 127270 30600
rect 127360 30570 127390 30600
rect 116060 30540 116140 30550
rect 116210 30540 116290 30550
rect 116560 30540 116620 30570
rect 116680 30540 116740 30570
rect 127245 30540 127300 30570
rect 127360 30540 127420 30570
rect 127560 30540 127640 30550
rect 127710 30540 127790 30550
rect 127860 30540 127940 30550
rect 116140 30460 116150 30540
rect 116290 30460 116300 30540
rect 116680 30450 116710 30480
rect 127245 30450 127270 30480
rect 127360 30450 127390 30480
rect 127640 30460 127650 30540
rect 127790 30460 127800 30540
rect 127940 30460 127950 30540
rect 128320 30520 128330 30600
rect 128640 30520 128650 30600
rect 129060 30520 129070 30600
rect 129380 30520 129390 30600
rect 130180 30570 130210 30600
rect 140860 30570 140890 30600
rect 129560 30540 129640 30550
rect 129710 30540 129790 30550
rect 130060 30540 130120 30570
rect 130180 30540 130240 30570
rect 140860 30540 140920 30570
rect 141060 30540 141140 30550
rect 141210 30540 141290 30550
rect 141360 30540 141440 30550
rect 129640 30460 129650 30540
rect 129790 30460 129800 30540
rect 130180 30450 130210 30480
rect 140860 30450 140890 30480
rect 141140 30460 141150 30540
rect 141290 30460 141300 30540
rect 141440 30460 141450 30540
rect 49060 30420 49120 30450
rect 49180 30420 49240 30450
rect 49300 30420 49360 30450
rect 49420 30420 49480 30450
rect 49540 30420 49600 30450
rect 49660 30420 49720 30450
rect 49780 30420 49840 30450
rect 49900 30420 49960 30450
rect 50020 30420 50080 30450
rect 50140 30420 50200 30450
rect 50260 30420 50320 30450
rect 50380 30420 50440 30450
rect 50500 30420 50560 30450
rect 50620 30420 50680 30450
rect 50740 30420 50800 30450
rect 50860 30420 50920 30450
rect 50980 30420 51040 30450
rect 51100 30420 51160 30450
rect 51220 30420 51280 30450
rect 51340 30420 51400 30450
rect 51460 30420 51520 30450
rect 51580 30420 51640 30450
rect 51700 30420 51760 30450
rect 51820 30420 51880 30450
rect 51940 30420 52000 30450
rect 52060 30420 52120 30450
rect 52180 30420 52240 30450
rect 52300 30420 52360 30450
rect 52420 30420 52480 30450
rect 52540 30420 52600 30450
rect 52660 30420 52720 30450
rect 52780 30420 52840 30450
rect 52900 30420 52960 30450
rect 53020 30420 53080 30450
rect 53140 30420 53200 30450
rect 53260 30420 53320 30450
rect 53380 30420 53440 30450
rect 53500 30420 53560 30450
rect 53620 30420 53680 30450
rect 53740 30420 53800 30450
rect 53860 30420 53920 30450
rect 53980 30420 54040 30450
rect 54100 30420 54160 30450
rect 54220 30420 54280 30450
rect 54340 30420 54400 30450
rect 54460 30420 54520 30450
rect 54580 30420 54640 30450
rect 54700 30420 54760 30450
rect 54820 30420 54880 30450
rect 54940 30420 55000 30450
rect 55060 30420 55120 30450
rect 55180 30420 55240 30450
rect 55300 30420 55360 30450
rect 55420 30420 55480 30450
rect 55540 30420 55600 30450
rect 55660 30420 55720 30450
rect 55780 30420 55840 30450
rect 55900 30420 55960 30450
rect 56020 30420 56080 30450
rect 56140 30420 56200 30450
rect 56260 30420 56320 30450
rect 56380 30420 56440 30450
rect 56500 30420 56560 30450
rect 56620 30420 56680 30450
rect 56740 30420 56800 30450
rect 56860 30420 56920 30450
rect 56980 30420 57040 30450
rect 57100 30420 57160 30450
rect 57220 30420 57280 30450
rect 57340 30420 57400 30450
rect 57460 30420 57520 30450
rect 57580 30420 57640 30450
rect 57700 30420 57760 30450
rect 57820 30420 57880 30450
rect 57940 30420 58000 30450
rect 58060 30420 58120 30450
rect 58180 30420 58240 30450
rect 58300 30420 58360 30450
rect 58420 30420 58480 30450
rect 58540 30420 58600 30450
rect 58660 30420 58720 30450
rect 58780 30420 58840 30450
rect 58900 30420 58960 30450
rect 59020 30420 59080 30450
rect 59140 30420 59200 30450
rect 59260 30420 59320 30450
rect 59380 30420 59440 30450
rect 59500 30420 59560 30450
rect 59620 30420 59680 30450
rect 59740 30420 59800 30450
rect 59860 30420 59920 30450
rect 60580 30440 60660 30450
rect 60900 30440 60980 30450
rect 61320 30440 61400 30450
rect 61640 30440 61720 30450
rect 48500 30360 48640 30370
rect 48710 30360 48790 30370
rect 60060 30360 60140 30370
rect 60210 30360 60290 30370
rect 60360 30360 60440 30370
rect 60660 30360 60670 30440
rect 60980 30360 60990 30440
rect 61400 30360 61410 30440
rect 61720 30360 61730 30440
rect 62560 30420 62620 30450
rect 62680 30420 62740 30450
rect 73245 30420 73300 30450
rect 73360 30420 73420 30450
rect 74080 30440 74160 30450
rect 74400 30440 74480 30450
rect 74820 30440 74900 30450
rect 75140 30440 75220 30450
rect 62060 30360 62140 30370
rect 62210 30360 62290 30370
rect 73560 30360 73640 30370
rect 73710 30360 73790 30370
rect 73860 30360 73940 30370
rect 74160 30360 74170 30440
rect 74480 30360 74490 30440
rect 74900 30360 74910 30440
rect 75220 30360 75230 30440
rect 76060 30420 76120 30450
rect 76180 30420 76240 30450
rect 86745 30420 86800 30450
rect 86860 30420 86920 30450
rect 87580 30440 87660 30450
rect 87900 30440 87980 30450
rect 88320 30440 88400 30450
rect 88640 30440 88720 30450
rect 75560 30360 75640 30370
rect 75710 30360 75790 30370
rect 87060 30360 87140 30370
rect 87210 30360 87290 30370
rect 87360 30360 87440 30370
rect 87660 30360 87670 30440
rect 87980 30360 87990 30440
rect 88400 30360 88410 30440
rect 88720 30360 88730 30440
rect 89560 30420 89620 30450
rect 89680 30420 89740 30450
rect 100245 30420 100300 30450
rect 100360 30420 100420 30450
rect 101080 30440 101160 30450
rect 101400 30440 101480 30450
rect 101820 30440 101900 30450
rect 102140 30440 102220 30450
rect 89060 30360 89140 30370
rect 89210 30360 89290 30370
rect 100560 30360 100640 30370
rect 100710 30360 100790 30370
rect 100860 30360 100940 30370
rect 101160 30360 101170 30440
rect 101480 30360 101490 30440
rect 101900 30360 101910 30440
rect 102220 30360 102230 30440
rect 103060 30420 103120 30450
rect 103180 30420 103240 30450
rect 113745 30420 113800 30450
rect 113860 30420 113920 30450
rect 114580 30440 114660 30450
rect 114900 30440 114980 30450
rect 115320 30440 115400 30450
rect 115640 30440 115720 30450
rect 102560 30360 102640 30370
rect 102710 30360 102790 30370
rect 114060 30360 114140 30370
rect 114210 30360 114290 30370
rect 114360 30360 114440 30370
rect 114660 30360 114670 30440
rect 114980 30360 114990 30440
rect 115400 30360 115410 30440
rect 115720 30360 115730 30440
rect 116560 30420 116620 30450
rect 116680 30420 116740 30450
rect 127245 30420 127300 30450
rect 127360 30420 127420 30450
rect 128080 30440 128160 30450
rect 128400 30440 128480 30450
rect 128820 30440 128900 30450
rect 129140 30440 129220 30450
rect 116060 30360 116140 30370
rect 116210 30360 116290 30370
rect 127560 30360 127640 30370
rect 127710 30360 127790 30370
rect 127860 30360 127940 30370
rect 128160 30360 128170 30440
rect 128480 30360 128490 30440
rect 128900 30360 128910 30440
rect 129220 30360 129230 30440
rect 130060 30420 130120 30450
rect 130180 30420 130240 30450
rect 140860 30420 140920 30450
rect 129560 30360 129640 30370
rect 129710 30360 129790 30370
rect 141060 30360 141140 30370
rect 141210 30360 141290 30370
rect 141360 30360 141440 30370
rect 48500 30200 48605 30360
rect 48640 30280 48650 30360
rect 48790 30280 48800 30360
rect 49180 30300 49210 30360
rect 49300 30300 49330 30360
rect 49420 30300 49450 30360
rect 49540 30300 49570 30360
rect 49660 30300 49690 30360
rect 49780 30300 49810 30360
rect 49900 30300 49930 30360
rect 50020 30300 50050 30360
rect 50140 30300 50170 30360
rect 50260 30300 50290 30360
rect 50380 30300 50410 30360
rect 50500 30300 50530 30360
rect 50620 30300 50650 30360
rect 50740 30300 50770 30360
rect 50860 30300 50890 30360
rect 50980 30300 51010 30360
rect 51100 30300 51130 30360
rect 51220 30300 51250 30360
rect 51340 30300 51370 30360
rect 51460 30300 51490 30360
rect 51580 30300 51610 30360
rect 51700 30300 51730 30360
rect 51820 30300 51850 30360
rect 51940 30300 51970 30360
rect 52060 30300 52090 30360
rect 52180 30300 52210 30360
rect 52300 30300 52330 30360
rect 52420 30300 52450 30360
rect 52540 30300 52570 30360
rect 52660 30300 52690 30360
rect 52780 30300 52810 30360
rect 52900 30300 52930 30360
rect 53020 30300 53050 30360
rect 53140 30300 53170 30360
rect 53260 30300 53290 30360
rect 53380 30300 53410 30360
rect 53500 30300 53530 30360
rect 53620 30300 53650 30360
rect 53740 30300 53770 30360
rect 53860 30300 53890 30360
rect 53980 30300 54010 30360
rect 54100 30300 54130 30360
rect 54220 30300 54250 30360
rect 54340 30300 54370 30360
rect 54460 30300 54490 30360
rect 54580 30300 54610 30360
rect 54700 30300 54730 30360
rect 54820 30300 54850 30360
rect 54940 30300 54970 30360
rect 55060 30300 55090 30360
rect 55180 30300 55210 30360
rect 55300 30300 55330 30360
rect 55420 30300 55450 30360
rect 55540 30300 55570 30360
rect 55660 30300 55690 30360
rect 55780 30300 55810 30360
rect 55900 30300 55930 30360
rect 56020 30300 56050 30360
rect 56140 30300 56170 30360
rect 56260 30300 56290 30360
rect 56380 30300 56410 30360
rect 56500 30300 56530 30360
rect 56620 30300 56650 30360
rect 56740 30300 56770 30360
rect 56860 30300 56890 30360
rect 56980 30300 57010 30360
rect 57100 30300 57130 30360
rect 57220 30300 57250 30360
rect 57340 30300 57370 30360
rect 57460 30300 57490 30360
rect 57580 30300 57610 30360
rect 57700 30300 57730 30360
rect 57820 30300 57850 30360
rect 57940 30300 57970 30360
rect 58060 30300 58090 30360
rect 58180 30300 58210 30360
rect 58300 30300 58330 30360
rect 58420 30300 58450 30360
rect 58540 30300 58570 30360
rect 58660 30300 58690 30360
rect 58780 30300 58810 30360
rect 58900 30300 58930 30360
rect 59020 30300 59050 30360
rect 59140 30300 59170 30360
rect 59260 30300 59290 30360
rect 59380 30300 59410 30360
rect 59500 30300 59530 30360
rect 59620 30300 59650 30360
rect 59740 30300 59770 30360
rect 59860 30300 59890 30360
rect 60140 30280 60150 30360
rect 60290 30280 60300 30360
rect 60440 30280 60450 30360
rect 62140 30280 62150 30360
rect 62290 30280 62300 30360
rect 62680 30300 62710 30360
rect 73245 30300 73270 30360
rect 73360 30300 73390 30360
rect 73640 30280 73650 30360
rect 73790 30280 73800 30360
rect 73940 30280 73950 30360
rect 75640 30280 75650 30360
rect 75790 30280 75800 30360
rect 76180 30300 76210 30360
rect 86745 30300 86770 30360
rect 86860 30300 86890 30360
rect 87140 30280 87150 30360
rect 87290 30280 87300 30360
rect 87440 30280 87450 30360
rect 89140 30280 89150 30360
rect 89290 30280 89300 30360
rect 89680 30300 89710 30360
rect 100245 30300 100270 30360
rect 100360 30300 100390 30360
rect 100640 30280 100650 30360
rect 100790 30280 100800 30360
rect 100940 30280 100950 30360
rect 102640 30280 102650 30360
rect 102790 30280 102800 30360
rect 103180 30300 103210 30360
rect 113745 30300 113770 30360
rect 113860 30300 113890 30360
rect 114140 30280 114150 30360
rect 114290 30280 114300 30360
rect 114440 30280 114450 30360
rect 116140 30280 116150 30360
rect 116290 30280 116300 30360
rect 116680 30300 116710 30360
rect 127245 30300 127270 30360
rect 127360 30300 127390 30360
rect 127640 30280 127650 30360
rect 127790 30280 127800 30360
rect 127940 30280 127950 30360
rect 129640 30280 129650 30360
rect 129790 30280 129800 30360
rect 130180 30300 130210 30360
rect 140860 30300 140890 30360
rect 141140 30280 141150 30360
rect 141290 30280 141300 30360
rect 141440 30280 141450 30360
rect 141565 30200 141620 38000
rect 150460 37940 150470 38020
rect 150780 37940 150790 38020
rect 151100 37940 151110 38020
rect 151420 37940 151430 38020
rect 151740 37940 151750 38020
rect 152060 37940 152070 38020
rect 152380 37940 152390 38020
rect 152700 37940 152710 38020
rect 153020 37940 153030 38020
rect 153340 37940 153350 38020
rect 153660 37940 153670 38020
rect 153980 37940 153990 38020
rect 154300 37940 154310 38020
rect 154620 37940 154630 38020
rect 154940 37940 154950 38020
rect 155260 37940 155270 38020
rect 155580 37940 155590 38020
rect 155900 37940 155910 38020
rect 150220 37860 150300 37870
rect 150540 37860 150620 37870
rect 150860 37860 150940 37870
rect 151180 37860 151260 37870
rect 151500 37860 151580 37870
rect 151820 37860 151900 37870
rect 152140 37860 152220 37870
rect 152460 37860 152540 37870
rect 152780 37860 152860 37870
rect 153100 37860 153180 37870
rect 153420 37860 153500 37870
rect 153740 37860 153820 37870
rect 154060 37860 154140 37870
rect 154380 37860 154460 37870
rect 154700 37860 154780 37870
rect 155020 37860 155100 37870
rect 155340 37860 155420 37870
rect 155660 37860 155740 37870
rect 155980 37860 156000 37870
rect 141665 37800 141745 37810
rect 141985 37800 142065 37810
rect 145200 37800 145265 37810
rect 145505 37800 145585 37810
rect 145825 37800 145905 37810
rect 146145 37800 146225 37810
rect 141745 37720 141755 37800
rect 142065 37720 142075 37800
rect 145265 37720 145275 37800
rect 145585 37720 145595 37800
rect 145905 37720 145915 37800
rect 146225 37720 146235 37800
rect 150300 37780 150310 37860
rect 150620 37780 150630 37860
rect 150940 37780 150950 37860
rect 151260 37780 151270 37860
rect 151580 37780 151590 37860
rect 151900 37780 151910 37860
rect 152220 37780 152230 37860
rect 152540 37780 152550 37860
rect 152860 37780 152870 37860
rect 153180 37780 153190 37860
rect 153500 37780 153510 37860
rect 153820 37780 153830 37860
rect 154140 37780 154150 37860
rect 154460 37780 154470 37860
rect 154780 37780 154790 37860
rect 155100 37780 155110 37860
rect 155420 37780 155430 37860
rect 155740 37780 155750 37860
rect 146540 37700 146620 37710
rect 146860 37700 146940 37710
rect 147180 37700 147260 37710
rect 147500 37700 147580 37710
rect 147820 37700 147900 37710
rect 148140 37700 148220 37710
rect 148460 37700 148540 37710
rect 148780 37700 148860 37710
rect 149100 37700 149180 37710
rect 149420 37700 149500 37710
rect 149740 37700 149820 37710
rect 150060 37700 150140 37710
rect 150380 37700 150460 37710
rect 150700 37700 150780 37710
rect 151020 37700 151100 37710
rect 151340 37700 151420 37710
rect 151660 37700 151740 37710
rect 151980 37700 152060 37710
rect 152300 37700 152380 37710
rect 152620 37700 152700 37710
rect 152940 37700 153020 37710
rect 153260 37700 153340 37710
rect 153580 37700 153660 37710
rect 153900 37700 153980 37710
rect 154220 37700 154300 37710
rect 154540 37700 154620 37710
rect 154860 37700 154940 37710
rect 155180 37700 155260 37710
rect 155500 37700 155580 37710
rect 155820 37700 155900 37710
rect 141825 37640 141905 37650
rect 142145 37640 142200 37650
rect 145345 37640 145425 37650
rect 145665 37640 145745 37650
rect 145985 37640 146065 37650
rect 141905 37560 141915 37640
rect 145425 37560 145435 37640
rect 145745 37560 145755 37640
rect 146065 37560 146075 37640
rect 146620 37620 146630 37700
rect 146940 37620 146950 37700
rect 147260 37620 147270 37700
rect 147580 37620 147590 37700
rect 147900 37620 147910 37700
rect 148220 37620 148230 37700
rect 148540 37620 148550 37700
rect 148860 37620 148870 37700
rect 149180 37620 149190 37700
rect 149500 37620 149510 37700
rect 149820 37620 149830 37700
rect 150140 37620 150150 37700
rect 150460 37620 150470 37700
rect 150780 37620 150790 37700
rect 151100 37620 151110 37700
rect 151420 37620 151430 37700
rect 151740 37620 151750 37700
rect 152060 37620 152070 37700
rect 152380 37620 152390 37700
rect 152700 37620 152710 37700
rect 153020 37620 153030 37700
rect 153340 37620 153350 37700
rect 153660 37620 153670 37700
rect 153980 37620 153990 37700
rect 154300 37620 154310 37700
rect 154620 37620 154630 37700
rect 154940 37620 154950 37700
rect 155260 37620 155270 37700
rect 155580 37620 155590 37700
rect 155900 37620 155910 37700
rect 146700 37540 146780 37550
rect 147020 37540 147100 37550
rect 147340 37540 147420 37550
rect 147660 37540 147740 37550
rect 147980 37540 148060 37550
rect 148300 37540 148380 37550
rect 148620 37540 148700 37550
rect 148940 37540 149020 37550
rect 149260 37540 149340 37550
rect 149580 37540 149660 37550
rect 149900 37540 149980 37550
rect 150220 37540 150300 37550
rect 150540 37540 150620 37550
rect 150860 37540 150940 37550
rect 151180 37540 151260 37550
rect 151500 37540 151580 37550
rect 151820 37540 151900 37550
rect 152140 37540 152220 37550
rect 152460 37540 152540 37550
rect 152780 37540 152860 37550
rect 153100 37540 153180 37550
rect 153420 37540 153500 37550
rect 153740 37540 153820 37550
rect 154060 37540 154140 37550
rect 154380 37540 154460 37550
rect 154700 37540 154780 37550
rect 155020 37540 155100 37550
rect 155340 37540 155420 37550
rect 155660 37540 155740 37550
rect 155980 37540 156000 37550
rect 141665 37480 141745 37490
rect 141985 37480 142065 37490
rect 145200 37480 145265 37490
rect 145505 37480 145585 37490
rect 145825 37480 145905 37490
rect 146145 37480 146225 37490
rect 141745 37400 141755 37480
rect 142065 37400 142075 37480
rect 145265 37400 145275 37480
rect 145585 37400 145595 37480
rect 145905 37400 145915 37480
rect 146225 37400 146235 37480
rect 146780 37460 146790 37540
rect 147100 37460 147110 37540
rect 147420 37460 147430 37540
rect 147740 37460 147750 37540
rect 148060 37460 148070 37540
rect 148380 37460 148390 37540
rect 148700 37460 148710 37540
rect 149020 37460 149030 37540
rect 149340 37460 149350 37540
rect 149660 37460 149670 37540
rect 149980 37460 149990 37540
rect 150300 37460 150310 37540
rect 150620 37460 150630 37540
rect 150940 37460 150950 37540
rect 151260 37460 151270 37540
rect 151580 37460 151590 37540
rect 151900 37460 151910 37540
rect 152220 37460 152230 37540
rect 152540 37460 152550 37540
rect 152860 37460 152870 37540
rect 153180 37460 153190 37540
rect 153500 37460 153510 37540
rect 153820 37460 153830 37540
rect 154140 37460 154150 37540
rect 154460 37460 154470 37540
rect 154780 37460 154790 37540
rect 155100 37460 155110 37540
rect 155420 37460 155430 37540
rect 155740 37460 155750 37540
rect 146540 37380 146620 37390
rect 146860 37380 146940 37390
rect 147180 37380 147260 37390
rect 147500 37380 147580 37390
rect 147820 37380 147900 37390
rect 148140 37380 148220 37390
rect 148460 37380 148540 37390
rect 148780 37380 148860 37390
rect 149100 37380 149180 37390
rect 149420 37380 149500 37390
rect 149740 37380 149820 37390
rect 150060 37380 150140 37390
rect 150380 37380 150460 37390
rect 150700 37380 150780 37390
rect 151020 37380 151100 37390
rect 151340 37380 151420 37390
rect 151660 37380 151740 37390
rect 151980 37380 152060 37390
rect 152300 37380 152380 37390
rect 152620 37380 152700 37390
rect 152940 37380 153020 37390
rect 153260 37380 153340 37390
rect 153580 37380 153660 37390
rect 153900 37380 153980 37390
rect 154220 37380 154300 37390
rect 154540 37380 154620 37390
rect 154860 37380 154940 37390
rect 155180 37380 155260 37390
rect 155500 37380 155580 37390
rect 155820 37380 155900 37390
rect 141825 37320 141905 37330
rect 142145 37320 142200 37330
rect 145345 37320 145425 37330
rect 145665 37320 145745 37330
rect 145985 37320 146065 37330
rect 141905 37240 141915 37320
rect 145425 37240 145435 37320
rect 145745 37240 145755 37320
rect 146065 37240 146075 37320
rect 146620 37300 146630 37380
rect 146940 37300 146950 37380
rect 147260 37300 147270 37380
rect 147580 37300 147590 37380
rect 147900 37300 147910 37380
rect 148220 37300 148230 37380
rect 148540 37300 148550 37380
rect 148860 37300 148870 37380
rect 149180 37300 149190 37380
rect 149500 37300 149510 37380
rect 149820 37300 149830 37380
rect 150140 37300 150150 37380
rect 150460 37300 150470 37380
rect 150780 37300 150790 37380
rect 151100 37300 151110 37380
rect 151420 37300 151430 37380
rect 151740 37300 151750 37380
rect 152060 37300 152070 37380
rect 152380 37300 152390 37380
rect 152700 37300 152710 37380
rect 153020 37300 153030 37380
rect 153340 37300 153350 37380
rect 153660 37300 153670 37380
rect 153980 37300 153990 37380
rect 154300 37300 154310 37380
rect 154620 37300 154630 37380
rect 154940 37300 154950 37380
rect 155260 37300 155270 37380
rect 155580 37300 155590 37380
rect 155900 37300 155910 37380
rect 146700 37220 146780 37230
rect 147020 37220 147100 37230
rect 147340 37220 147420 37230
rect 147660 37220 147740 37230
rect 147980 37220 148060 37230
rect 148300 37220 148380 37230
rect 148620 37220 148700 37230
rect 148940 37220 149020 37230
rect 149260 37220 149340 37230
rect 149580 37220 149660 37230
rect 149900 37220 149980 37230
rect 150220 37220 150300 37230
rect 150540 37220 150620 37230
rect 150860 37220 150940 37230
rect 151180 37220 151260 37230
rect 151500 37220 151580 37230
rect 151820 37220 151900 37230
rect 152140 37220 152220 37230
rect 152460 37220 152540 37230
rect 152780 37220 152860 37230
rect 153100 37220 153180 37230
rect 153420 37220 153500 37230
rect 153740 37220 153820 37230
rect 154060 37220 154140 37230
rect 154380 37220 154460 37230
rect 154700 37220 154780 37230
rect 155020 37220 155100 37230
rect 155340 37220 155420 37230
rect 155660 37220 155740 37230
rect 155980 37220 156000 37230
rect 141665 37160 141745 37170
rect 141985 37160 142065 37170
rect 145200 37160 145265 37170
rect 145505 37160 145585 37170
rect 145825 37160 145905 37170
rect 146145 37160 146225 37170
rect 141745 37080 141755 37160
rect 142065 37080 142075 37160
rect 145265 37080 145275 37160
rect 145585 37080 145595 37160
rect 145905 37080 145915 37160
rect 146225 37080 146235 37160
rect 146780 37140 146790 37220
rect 147100 37140 147110 37220
rect 147420 37140 147430 37220
rect 147740 37140 147750 37220
rect 148060 37140 148070 37220
rect 148380 37140 148390 37220
rect 148700 37140 148710 37220
rect 149020 37140 149030 37220
rect 149340 37140 149350 37220
rect 149660 37140 149670 37220
rect 149980 37140 149990 37220
rect 150300 37140 150310 37220
rect 150620 37140 150630 37220
rect 150940 37140 150950 37220
rect 151260 37140 151270 37220
rect 151580 37140 151590 37220
rect 151900 37140 151910 37220
rect 152220 37140 152230 37220
rect 152540 37140 152550 37220
rect 152860 37140 152870 37220
rect 153180 37140 153190 37220
rect 153500 37140 153510 37220
rect 153820 37140 153830 37220
rect 154140 37140 154150 37220
rect 154460 37140 154470 37220
rect 154780 37140 154790 37220
rect 155100 37140 155110 37220
rect 155420 37140 155430 37220
rect 155740 37140 155750 37220
rect 146540 37060 146620 37070
rect 146860 37060 146940 37070
rect 147180 37060 147260 37070
rect 147500 37060 147580 37070
rect 147820 37060 147900 37070
rect 148140 37060 148220 37070
rect 148460 37060 148540 37070
rect 148780 37060 148860 37070
rect 149100 37060 149180 37070
rect 149420 37060 149500 37070
rect 149740 37060 149820 37070
rect 150060 37060 150140 37070
rect 150380 37060 150460 37070
rect 150700 37060 150780 37070
rect 151020 37060 151100 37070
rect 151340 37060 151420 37070
rect 151660 37060 151740 37070
rect 151980 37060 152060 37070
rect 152300 37060 152380 37070
rect 152620 37060 152700 37070
rect 152940 37060 153020 37070
rect 153260 37060 153340 37070
rect 153580 37060 153660 37070
rect 153900 37060 153980 37070
rect 154220 37060 154300 37070
rect 154540 37060 154620 37070
rect 154860 37060 154940 37070
rect 155180 37060 155260 37070
rect 155500 37060 155580 37070
rect 155820 37060 155900 37070
rect 141825 37000 141905 37010
rect 142145 37000 142200 37010
rect 145345 37000 145425 37010
rect 145665 37000 145745 37010
rect 145985 37000 146065 37010
rect 141905 36920 141915 37000
rect 145425 36920 145435 37000
rect 145745 36920 145755 37000
rect 146065 36920 146075 37000
rect 146620 36980 146630 37060
rect 146940 36980 146950 37060
rect 147260 36980 147270 37060
rect 147580 36980 147590 37060
rect 147900 36980 147910 37060
rect 148220 36980 148230 37060
rect 148540 36980 148550 37060
rect 148860 36980 148870 37060
rect 149180 36980 149190 37060
rect 149500 36980 149510 37060
rect 149820 36980 149830 37060
rect 150140 36980 150150 37060
rect 150460 36980 150470 37060
rect 150780 36980 150790 37060
rect 151100 36980 151110 37060
rect 151420 36980 151430 37060
rect 151740 36980 151750 37060
rect 152060 36980 152070 37060
rect 152380 36980 152390 37060
rect 152700 36980 152710 37060
rect 153020 36980 153030 37060
rect 153340 36980 153350 37060
rect 153660 36980 153670 37060
rect 153980 36980 153990 37060
rect 154300 36980 154310 37060
rect 154620 36980 154630 37060
rect 154940 36980 154950 37060
rect 155260 36980 155270 37060
rect 155580 36980 155590 37060
rect 155900 36980 155910 37060
rect 146700 36900 146780 36910
rect 147020 36900 147100 36910
rect 147340 36900 147420 36910
rect 147660 36900 147740 36910
rect 147980 36900 148060 36910
rect 148300 36900 148380 36910
rect 148620 36900 148700 36910
rect 148940 36900 149020 36910
rect 149260 36900 149340 36910
rect 149580 36900 149660 36910
rect 149900 36900 149980 36910
rect 150220 36900 150300 36910
rect 150540 36900 150620 36910
rect 150860 36900 150940 36910
rect 151180 36900 151260 36910
rect 151500 36900 151580 36910
rect 151820 36900 151900 36910
rect 152140 36900 152220 36910
rect 152460 36900 152540 36910
rect 152780 36900 152860 36910
rect 153100 36900 153180 36910
rect 153420 36900 153500 36910
rect 153740 36900 153820 36910
rect 154060 36900 154140 36910
rect 154380 36900 154460 36910
rect 154700 36900 154780 36910
rect 155020 36900 155100 36910
rect 155340 36900 155420 36910
rect 155660 36900 155740 36910
rect 155980 36900 156000 36910
rect 141665 36840 141745 36850
rect 141985 36840 142065 36850
rect 145200 36840 145265 36850
rect 145505 36840 145585 36850
rect 145825 36840 145905 36850
rect 146145 36840 146225 36850
rect 141745 36760 141755 36840
rect 142065 36760 142075 36840
rect 145265 36760 145275 36840
rect 145585 36760 145595 36840
rect 145905 36760 145915 36840
rect 146225 36760 146235 36840
rect 146780 36820 146790 36900
rect 147100 36820 147110 36900
rect 147420 36820 147430 36900
rect 147740 36820 147750 36900
rect 148060 36820 148070 36900
rect 148380 36820 148390 36900
rect 148700 36820 148710 36900
rect 149020 36820 149030 36900
rect 149340 36820 149350 36900
rect 149660 36820 149670 36900
rect 149980 36820 149990 36900
rect 150300 36820 150310 36900
rect 150620 36820 150630 36900
rect 150940 36820 150950 36900
rect 151260 36820 151270 36900
rect 151580 36820 151590 36900
rect 151900 36820 151910 36900
rect 152220 36820 152230 36900
rect 152540 36820 152550 36900
rect 152860 36820 152870 36900
rect 153180 36820 153190 36900
rect 153500 36820 153510 36900
rect 153820 36820 153830 36900
rect 154140 36820 154150 36900
rect 154460 36820 154470 36900
rect 154780 36820 154790 36900
rect 155100 36820 155110 36900
rect 155420 36820 155430 36900
rect 155740 36820 155750 36900
rect 146540 36740 146620 36750
rect 146860 36740 146940 36750
rect 147180 36740 147260 36750
rect 147500 36740 147580 36750
rect 147820 36740 147900 36750
rect 148140 36740 148220 36750
rect 148460 36740 148540 36750
rect 148780 36740 148860 36750
rect 149100 36740 149180 36750
rect 149420 36740 149500 36750
rect 149740 36740 149820 36750
rect 150060 36740 150140 36750
rect 150380 36740 150460 36750
rect 150700 36740 150780 36750
rect 151020 36740 151100 36750
rect 151340 36740 151420 36750
rect 151660 36740 151740 36750
rect 151980 36740 152060 36750
rect 152300 36740 152380 36750
rect 152620 36740 152700 36750
rect 152940 36740 153020 36750
rect 153260 36740 153340 36750
rect 153580 36740 153660 36750
rect 153900 36740 153980 36750
rect 154220 36740 154300 36750
rect 154540 36740 154620 36750
rect 154860 36740 154940 36750
rect 155180 36740 155260 36750
rect 155500 36740 155580 36750
rect 155820 36740 155900 36750
rect 141825 36680 141905 36690
rect 142145 36680 142200 36690
rect 145345 36680 145425 36690
rect 145665 36680 145745 36690
rect 145985 36680 146065 36690
rect 141905 36600 141915 36680
rect 145425 36600 145435 36680
rect 145745 36600 145755 36680
rect 146065 36600 146075 36680
rect 146620 36660 146630 36740
rect 146940 36660 146950 36740
rect 147260 36660 147270 36740
rect 147580 36660 147590 36740
rect 147900 36660 147910 36740
rect 148220 36660 148230 36740
rect 148540 36660 148550 36740
rect 148860 36660 148870 36740
rect 149180 36660 149190 36740
rect 149500 36660 149510 36740
rect 149820 36660 149830 36740
rect 150140 36660 150150 36740
rect 150460 36660 150470 36740
rect 150780 36660 150790 36740
rect 151100 36660 151110 36740
rect 151420 36660 151430 36740
rect 151740 36660 151750 36740
rect 152060 36660 152070 36740
rect 152380 36660 152390 36740
rect 152700 36660 152710 36740
rect 153020 36660 153030 36740
rect 153340 36660 153350 36740
rect 153660 36660 153670 36740
rect 153980 36660 153990 36740
rect 154300 36660 154310 36740
rect 154620 36660 154630 36740
rect 154940 36660 154950 36740
rect 155260 36660 155270 36740
rect 155580 36660 155590 36740
rect 155900 36660 155910 36740
rect 146700 36580 146780 36590
rect 147020 36580 147100 36590
rect 147340 36580 147420 36590
rect 147660 36580 147740 36590
rect 147980 36580 148060 36590
rect 148300 36580 148380 36590
rect 148620 36580 148700 36590
rect 148940 36580 149020 36590
rect 149260 36580 149340 36590
rect 149580 36580 149660 36590
rect 149900 36580 149980 36590
rect 150220 36580 150300 36590
rect 150540 36580 150620 36590
rect 150860 36580 150940 36590
rect 151180 36580 151260 36590
rect 151500 36580 151580 36590
rect 151820 36580 151900 36590
rect 152140 36580 152220 36590
rect 152460 36580 152540 36590
rect 152780 36580 152860 36590
rect 153100 36580 153180 36590
rect 153420 36580 153500 36590
rect 153740 36580 153820 36590
rect 154060 36580 154140 36590
rect 154380 36580 154460 36590
rect 154700 36580 154780 36590
rect 155020 36580 155100 36590
rect 155340 36580 155420 36590
rect 155660 36580 155740 36590
rect 155980 36580 156000 36590
rect 141665 36520 141745 36530
rect 141985 36520 142065 36530
rect 145200 36520 145265 36530
rect 145505 36520 145585 36530
rect 145825 36520 145905 36530
rect 146145 36520 146225 36530
rect 141745 36440 141755 36520
rect 142065 36440 142075 36520
rect 145265 36440 145275 36520
rect 145585 36440 145595 36520
rect 145905 36440 145915 36520
rect 146225 36440 146235 36520
rect 146780 36500 146790 36580
rect 147100 36500 147110 36580
rect 147420 36500 147430 36580
rect 147740 36500 147750 36580
rect 148060 36500 148070 36580
rect 148380 36500 148390 36580
rect 148700 36500 148710 36580
rect 149020 36500 149030 36580
rect 149340 36500 149350 36580
rect 149660 36500 149670 36580
rect 149980 36500 149990 36580
rect 150300 36500 150310 36580
rect 150620 36500 150630 36580
rect 150940 36500 150950 36580
rect 151260 36500 151270 36580
rect 151580 36500 151590 36580
rect 151900 36500 151910 36580
rect 152220 36500 152230 36580
rect 152540 36500 152550 36580
rect 152860 36500 152870 36580
rect 153180 36500 153190 36580
rect 153500 36500 153510 36580
rect 153820 36500 153830 36580
rect 154140 36500 154150 36580
rect 154460 36500 154470 36580
rect 154780 36500 154790 36580
rect 155100 36500 155110 36580
rect 155420 36500 155430 36580
rect 155740 36500 155750 36580
rect 146540 36420 146620 36430
rect 146860 36420 146940 36430
rect 147180 36420 147260 36430
rect 147500 36420 147580 36430
rect 147820 36420 147900 36430
rect 148140 36420 148220 36430
rect 148460 36420 148540 36430
rect 148780 36420 148860 36430
rect 149100 36420 149180 36430
rect 149420 36420 149500 36430
rect 149740 36420 149820 36430
rect 150060 36420 150140 36430
rect 150380 36420 150460 36430
rect 150700 36420 150780 36430
rect 151020 36420 151100 36430
rect 151340 36420 151420 36430
rect 151660 36420 151740 36430
rect 151980 36420 152060 36430
rect 152300 36420 152380 36430
rect 152620 36420 152700 36430
rect 152940 36420 153020 36430
rect 153260 36420 153340 36430
rect 153580 36420 153660 36430
rect 153900 36420 153980 36430
rect 154220 36420 154300 36430
rect 154540 36420 154620 36430
rect 154860 36420 154940 36430
rect 155180 36420 155260 36430
rect 155500 36420 155580 36430
rect 155820 36420 155900 36430
rect 141825 36360 141905 36370
rect 142145 36360 142200 36370
rect 145345 36360 145425 36370
rect 145665 36360 145745 36370
rect 145985 36360 146065 36370
rect 141905 36280 141915 36360
rect 145425 36280 145435 36360
rect 145745 36280 145755 36360
rect 146065 36280 146075 36360
rect 146620 36340 146630 36420
rect 146940 36340 146950 36420
rect 147260 36340 147270 36420
rect 147580 36340 147590 36420
rect 147900 36340 147910 36420
rect 148220 36340 148230 36420
rect 148540 36340 148550 36420
rect 148860 36340 148870 36420
rect 149180 36340 149190 36420
rect 149500 36340 149510 36420
rect 149820 36340 149830 36420
rect 150140 36340 150150 36420
rect 150460 36340 150470 36420
rect 150780 36340 150790 36420
rect 151100 36340 151110 36420
rect 151420 36340 151430 36420
rect 151740 36340 151750 36420
rect 152060 36340 152070 36420
rect 152380 36340 152390 36420
rect 152700 36340 152710 36420
rect 153020 36340 153030 36420
rect 153340 36340 153350 36420
rect 153660 36340 153670 36420
rect 153980 36340 153990 36420
rect 154300 36340 154310 36420
rect 154620 36340 154630 36420
rect 154940 36340 154950 36420
rect 155260 36340 155270 36420
rect 155580 36340 155590 36420
rect 155900 36340 155910 36420
rect 146700 36260 146780 36270
rect 147020 36260 147100 36270
rect 147340 36260 147420 36270
rect 147660 36260 147740 36270
rect 147980 36260 148060 36270
rect 148300 36260 148380 36270
rect 148620 36260 148700 36270
rect 148940 36260 149020 36270
rect 149260 36260 149340 36270
rect 149580 36260 149660 36270
rect 149900 36260 149980 36270
rect 150220 36260 150300 36270
rect 150540 36260 150620 36270
rect 150860 36260 150940 36270
rect 151180 36260 151260 36270
rect 151500 36260 151580 36270
rect 151820 36260 151900 36270
rect 152140 36260 152220 36270
rect 152460 36260 152540 36270
rect 152780 36260 152860 36270
rect 153100 36260 153180 36270
rect 153420 36260 153500 36270
rect 153740 36260 153820 36270
rect 154060 36260 154140 36270
rect 154380 36260 154460 36270
rect 154700 36260 154780 36270
rect 155020 36260 155100 36270
rect 155340 36260 155420 36270
rect 155660 36260 155740 36270
rect 155980 36260 156000 36270
rect 141665 36200 141745 36210
rect 141985 36200 142065 36210
rect 145200 36200 145265 36210
rect 145505 36200 145585 36210
rect 145825 36200 145905 36210
rect 146145 36200 146225 36210
rect 141745 36120 141755 36200
rect 142065 36120 142075 36200
rect 145265 36120 145275 36200
rect 145585 36120 145595 36200
rect 145905 36120 145915 36200
rect 146225 36120 146235 36200
rect 146780 36180 146790 36260
rect 147100 36180 147110 36260
rect 147420 36180 147430 36260
rect 147740 36180 147750 36260
rect 148060 36180 148070 36260
rect 148380 36180 148390 36260
rect 148700 36180 148710 36260
rect 149020 36180 149030 36260
rect 149340 36180 149350 36260
rect 149660 36180 149670 36260
rect 149980 36180 149990 36260
rect 150300 36180 150310 36260
rect 150620 36180 150630 36260
rect 150940 36180 150950 36260
rect 151260 36180 151270 36260
rect 151580 36180 151590 36260
rect 151900 36180 151910 36260
rect 152220 36180 152230 36260
rect 152540 36180 152550 36260
rect 152860 36180 152870 36260
rect 153180 36180 153190 36260
rect 153500 36180 153510 36260
rect 153820 36180 153830 36260
rect 154140 36180 154150 36260
rect 154460 36180 154470 36260
rect 154780 36180 154790 36260
rect 155100 36180 155110 36260
rect 155420 36180 155430 36260
rect 155740 36180 155750 36260
rect 146540 36100 146620 36110
rect 146860 36100 146940 36110
rect 147180 36100 147260 36110
rect 147500 36100 147580 36110
rect 147820 36100 147900 36110
rect 148140 36100 148220 36110
rect 148460 36100 148540 36110
rect 148780 36100 148860 36110
rect 149100 36100 149180 36110
rect 149420 36100 149500 36110
rect 149740 36100 149820 36110
rect 150060 36100 150140 36110
rect 150380 36100 150460 36110
rect 150700 36100 150780 36110
rect 151020 36100 151100 36110
rect 151340 36100 151420 36110
rect 151660 36100 151740 36110
rect 151980 36100 152060 36110
rect 152300 36100 152380 36110
rect 152620 36100 152700 36110
rect 152940 36100 153020 36110
rect 153260 36100 153340 36110
rect 153580 36100 153660 36110
rect 153900 36100 153980 36110
rect 154220 36100 154300 36110
rect 154540 36100 154620 36110
rect 154860 36100 154940 36110
rect 155180 36100 155260 36110
rect 155500 36100 155580 36110
rect 155820 36100 155900 36110
rect 141825 36040 141905 36050
rect 142145 36040 142200 36050
rect 145345 36040 145425 36050
rect 145665 36040 145745 36050
rect 145985 36040 146065 36050
rect 141905 35960 141915 36040
rect 145425 35960 145435 36040
rect 145745 35960 145755 36040
rect 146065 35960 146075 36040
rect 146620 36020 146630 36100
rect 146940 36020 146950 36100
rect 147260 36020 147270 36100
rect 147580 36020 147590 36100
rect 147900 36020 147910 36100
rect 148220 36020 148230 36100
rect 148540 36020 148550 36100
rect 148860 36020 148870 36100
rect 149180 36020 149190 36100
rect 149500 36020 149510 36100
rect 149820 36020 149830 36100
rect 150140 36020 150150 36100
rect 150460 36020 150470 36100
rect 150780 36020 150790 36100
rect 151100 36020 151110 36100
rect 151420 36020 151430 36100
rect 151740 36020 151750 36100
rect 152060 36020 152070 36100
rect 152380 36020 152390 36100
rect 152700 36020 152710 36100
rect 153020 36020 153030 36100
rect 153340 36020 153350 36100
rect 153660 36020 153670 36100
rect 153980 36020 153990 36100
rect 154300 36020 154310 36100
rect 154620 36020 154630 36100
rect 154940 36020 154950 36100
rect 155260 36020 155270 36100
rect 155580 36020 155590 36100
rect 155900 36020 155910 36100
rect 146700 35940 146780 35950
rect 147020 35940 147100 35950
rect 141665 35880 141745 35890
rect 141985 35880 142065 35890
rect 145200 35880 145265 35890
rect 145505 35880 145585 35890
rect 145825 35880 145905 35890
rect 146145 35880 146225 35890
rect 141745 35800 141755 35880
rect 142065 35800 142075 35880
rect 145265 35800 145275 35880
rect 145585 35800 145595 35880
rect 145905 35800 145915 35880
rect 146225 35800 146235 35880
rect 146780 35860 146790 35940
rect 146540 35780 146620 35790
rect 146860 35780 146940 35790
rect 141825 35720 141905 35730
rect 142145 35720 142200 35730
rect 145345 35720 145425 35730
rect 145665 35720 145745 35730
rect 145985 35720 146065 35730
rect 141905 35640 141915 35720
rect 145425 35640 145435 35720
rect 145745 35640 145755 35720
rect 146065 35640 146075 35720
rect 146620 35700 146630 35780
rect 146940 35700 146950 35780
rect 146700 35620 146780 35630
rect 147020 35620 147100 35630
rect 141665 35560 141745 35570
rect 141985 35560 142065 35570
rect 145200 35560 145265 35570
rect 145505 35560 145585 35570
rect 145825 35560 145905 35570
rect 146145 35560 146225 35570
rect 141745 35480 141755 35560
rect 142065 35480 142075 35560
rect 145265 35480 145275 35560
rect 145585 35480 145595 35560
rect 145905 35480 145915 35560
rect 146225 35480 146235 35560
rect 146780 35540 146790 35620
rect 146540 35460 146620 35470
rect 146860 35460 146940 35470
rect 141825 35400 141905 35410
rect 142145 35400 142200 35410
rect 145345 35400 145425 35410
rect 145665 35400 145745 35410
rect 145985 35400 146065 35410
rect 141905 35320 141915 35400
rect 145425 35320 145435 35400
rect 145745 35320 145755 35400
rect 146065 35320 146075 35400
rect 146620 35380 146630 35460
rect 146940 35380 146950 35460
rect 146700 35300 146780 35310
rect 147020 35300 147100 35310
rect 141665 35240 141745 35250
rect 141985 35240 142065 35250
rect 145200 35240 145265 35250
rect 145505 35240 145585 35250
rect 145825 35240 145905 35250
rect 146145 35240 146225 35250
rect 141745 35160 141755 35240
rect 142065 35160 142075 35240
rect 145265 35160 145275 35240
rect 145585 35160 145595 35240
rect 145905 35160 145915 35240
rect 146225 35160 146235 35240
rect 146780 35220 146790 35300
rect 146540 35140 146620 35150
rect 146860 35140 146940 35150
rect 141825 35080 141905 35090
rect 142145 35080 142200 35090
rect 145345 35080 145425 35090
rect 145665 35080 145745 35090
rect 145985 35080 146065 35090
rect 141905 35000 141915 35080
rect 145425 35000 145435 35080
rect 145745 35000 145755 35080
rect 146065 35000 146075 35080
rect 146620 35060 146630 35140
rect 146940 35060 146950 35140
rect 146700 34980 146780 34990
rect 147020 34980 147100 34990
rect 141665 34920 141745 34930
rect 141985 34920 142065 34930
rect 145200 34920 145265 34930
rect 145505 34920 145585 34930
rect 145825 34920 145905 34930
rect 146145 34920 146225 34930
rect 141745 34840 141755 34920
rect 142065 34840 142075 34920
rect 145265 34840 145275 34920
rect 145585 34840 145595 34920
rect 145905 34840 145915 34920
rect 146225 34840 146235 34920
rect 146780 34900 146790 34980
rect 146540 34820 146620 34830
rect 146860 34820 146940 34830
rect 141825 34760 141905 34770
rect 142145 34760 142200 34770
rect 145345 34760 145425 34770
rect 145665 34760 145745 34770
rect 145985 34760 146065 34770
rect 141905 34680 141915 34760
rect 145425 34680 145435 34760
rect 145745 34680 145755 34760
rect 146065 34680 146075 34760
rect 146620 34740 146630 34820
rect 146940 34740 146950 34820
rect 146700 34660 146780 34670
rect 147020 34660 147100 34670
rect 141665 34600 141745 34610
rect 141985 34600 142065 34610
rect 145200 34600 145265 34610
rect 145505 34600 145585 34610
rect 145825 34600 145905 34610
rect 146145 34600 146225 34610
rect 141745 34520 141755 34600
rect 142065 34520 142075 34600
rect 145265 34520 145275 34600
rect 145585 34520 145595 34600
rect 145905 34520 145915 34600
rect 146225 34520 146235 34600
rect 146780 34580 146790 34660
rect 146540 34500 146620 34510
rect 146860 34500 146940 34510
rect 141825 34440 141905 34450
rect 142145 34440 142200 34450
rect 145345 34440 145425 34450
rect 145665 34440 145745 34450
rect 145985 34440 146065 34450
rect 141905 34360 141915 34440
rect 145425 34360 145435 34440
rect 145745 34360 145755 34440
rect 146065 34360 146075 34440
rect 146620 34420 146630 34500
rect 146940 34420 146950 34500
rect 146700 34340 146780 34350
rect 147020 34340 147100 34350
rect 141665 34280 141745 34290
rect 141985 34280 142065 34290
rect 145200 34280 145265 34290
rect 145505 34280 145585 34290
rect 145825 34280 145905 34290
rect 146145 34280 146225 34290
rect 141745 34200 141755 34280
rect 142065 34200 142075 34280
rect 145265 34200 145275 34280
rect 145585 34200 145595 34280
rect 145905 34200 145915 34280
rect 146225 34200 146235 34280
rect 146780 34260 146790 34340
rect 146540 34180 146620 34190
rect 146860 34180 146940 34190
rect 141825 34120 141905 34130
rect 142145 34120 142200 34130
rect 145345 34120 145425 34130
rect 145665 34120 145745 34130
rect 145985 34120 146065 34130
rect 141905 34040 141915 34120
rect 145425 34040 145435 34120
rect 145745 34040 145755 34120
rect 146065 34040 146075 34120
rect 146620 34100 146630 34180
rect 146940 34100 146950 34180
rect 146700 34020 146780 34030
rect 147020 34020 147100 34030
rect 141665 33960 141745 33970
rect 141985 33960 142065 33970
rect 145200 33960 145265 33970
rect 145505 33960 145585 33970
rect 145825 33960 145905 33970
rect 146145 33960 146225 33970
rect 141745 33880 141755 33960
rect 142065 33880 142075 33960
rect 145265 33880 145275 33960
rect 145585 33880 145595 33960
rect 145905 33880 145915 33960
rect 146225 33880 146235 33960
rect 146780 33940 146790 34020
rect 146540 33860 146620 33870
rect 146860 33860 146940 33870
rect 141825 33800 141905 33810
rect 142145 33800 142200 33810
rect 145345 33800 145425 33810
rect 145665 33800 145745 33810
rect 145985 33800 146065 33810
rect 141905 33720 141915 33800
rect 145425 33720 145435 33800
rect 145745 33720 145755 33800
rect 146065 33720 146075 33800
rect 146620 33780 146630 33860
rect 146940 33780 146950 33860
rect 146700 33700 146780 33710
rect 147020 33700 147100 33710
rect 141665 33640 141745 33650
rect 141985 33640 142065 33650
rect 145200 33640 145265 33650
rect 145505 33640 145585 33650
rect 145825 33640 145905 33650
rect 146145 33640 146225 33650
rect 141745 33560 141755 33640
rect 142065 33560 142075 33640
rect 145265 33560 145275 33640
rect 145585 33560 145595 33640
rect 145905 33560 145915 33640
rect 146225 33560 146235 33640
rect 146780 33620 146790 33700
rect 146540 33540 146620 33550
rect 146860 33540 146940 33550
rect 141825 33480 141905 33490
rect 142145 33480 142200 33490
rect 145345 33480 145425 33490
rect 145665 33480 145745 33490
rect 145985 33480 146065 33490
rect 141905 33400 141915 33480
rect 145425 33400 145435 33480
rect 145745 33400 145755 33480
rect 146065 33400 146075 33480
rect 146620 33460 146630 33540
rect 146940 33460 146950 33540
rect 146700 33380 146780 33390
rect 147020 33380 147100 33390
rect 141665 33320 141745 33330
rect 141985 33320 142065 33330
rect 145200 33320 145265 33330
rect 145505 33320 145585 33330
rect 145825 33320 145905 33330
rect 146145 33320 146225 33330
rect 141745 33240 141755 33320
rect 142065 33240 142075 33320
rect 145265 33240 145275 33320
rect 145585 33240 145595 33320
rect 145905 33240 145915 33320
rect 146225 33240 146235 33320
rect 146780 33300 146790 33380
rect 146540 33220 146620 33230
rect 146860 33220 146940 33230
rect 141825 33160 141905 33170
rect 142145 33160 142200 33170
rect 145345 33160 145425 33170
rect 145665 33160 145745 33170
rect 145985 33160 146065 33170
rect 141905 33080 141915 33160
rect 145425 33080 145435 33160
rect 145745 33080 145755 33160
rect 146065 33080 146075 33160
rect 146620 33140 146630 33220
rect 146940 33140 146950 33220
rect 146700 33060 146780 33070
rect 147020 33060 147100 33070
rect 141665 33000 141745 33010
rect 141985 33000 142065 33010
rect 145200 33000 145265 33010
rect 145505 33000 145585 33010
rect 145825 33000 145905 33010
rect 146145 33000 146225 33010
rect 141745 32920 141755 33000
rect 142065 32920 142075 33000
rect 145265 32920 145275 33000
rect 145585 32920 145595 33000
rect 145905 32920 145915 33000
rect 146225 32920 146235 33000
rect 146780 32980 146790 33060
rect 146540 32900 146620 32910
rect 146860 32900 146940 32910
rect 141825 32840 141905 32850
rect 142145 32840 142200 32850
rect 145345 32840 145425 32850
rect 145665 32840 145745 32850
rect 145985 32840 146065 32850
rect 141905 32760 141915 32840
rect 145425 32760 145435 32840
rect 145745 32760 145755 32840
rect 146065 32760 146075 32840
rect 146620 32820 146630 32900
rect 146940 32820 146950 32900
rect 146700 32740 146780 32750
rect 147020 32740 147100 32750
rect 141665 32680 141745 32690
rect 141985 32680 142065 32690
rect 145200 32680 145265 32690
rect 145505 32680 145585 32690
rect 145825 32680 145905 32690
rect 146145 32680 146225 32690
rect 141745 32600 141755 32680
rect 142065 32600 142075 32680
rect 145265 32600 145275 32680
rect 145585 32600 145595 32680
rect 145905 32600 145915 32680
rect 146225 32600 146235 32680
rect 146780 32660 146790 32740
rect 146540 32580 146620 32590
rect 146860 32580 146940 32590
rect 141825 32520 141905 32530
rect 142145 32520 142200 32530
rect 145345 32520 145425 32530
rect 145665 32520 145745 32530
rect 145985 32520 146065 32530
rect 141905 32440 141915 32520
rect 145425 32440 145435 32520
rect 145745 32440 145755 32520
rect 146065 32440 146075 32520
rect 146620 32500 146630 32580
rect 146940 32500 146950 32580
rect 146700 32420 146780 32430
rect 147020 32420 147100 32430
rect 141665 32360 141745 32370
rect 141985 32360 142065 32370
rect 145200 32360 145265 32370
rect 145505 32360 145585 32370
rect 145825 32360 145905 32370
rect 146145 32360 146225 32370
rect 141745 32280 141755 32360
rect 142065 32280 142075 32360
rect 145265 32280 145275 32360
rect 145585 32280 145595 32360
rect 145905 32280 145915 32360
rect 146225 32280 146235 32360
rect 146780 32340 146790 32420
rect 146540 32260 146620 32270
rect 146860 32260 146940 32270
rect 141825 32200 141905 32210
rect 142145 32200 142200 32210
rect 145345 32200 145425 32210
rect 145665 32200 145745 32210
rect 145985 32200 146065 32210
rect 141905 32120 141915 32200
rect 145425 32120 145435 32200
rect 145745 32120 145755 32200
rect 146065 32120 146075 32200
rect 146620 32180 146630 32260
rect 146940 32180 146950 32260
rect 146700 32100 146780 32110
rect 147020 32100 147100 32110
rect 141665 32040 141745 32050
rect 141985 32040 142065 32050
rect 145200 32040 145265 32050
rect 145505 32040 145585 32050
rect 145825 32040 145905 32050
rect 146145 32040 146225 32050
rect 141745 31960 141755 32040
rect 142065 31960 142075 32040
rect 145265 31960 145275 32040
rect 145585 31960 145595 32040
rect 145905 31960 145915 32040
rect 146225 31960 146235 32040
rect 146780 32020 146790 32100
rect 146540 31940 146620 31950
rect 146860 31940 146940 31950
rect 141825 31880 141905 31890
rect 142145 31880 142200 31890
rect 145345 31880 145425 31890
rect 145665 31880 145745 31890
rect 145985 31880 146065 31890
rect 141905 31800 141915 31880
rect 145425 31800 145435 31880
rect 145745 31800 145755 31880
rect 146065 31800 146075 31880
rect 146620 31860 146630 31940
rect 146940 31860 146950 31940
rect 146700 31780 146780 31790
rect 147020 31780 147100 31790
rect 141665 31720 141745 31730
rect 141985 31720 142065 31730
rect 145200 31720 145265 31730
rect 145505 31720 145585 31730
rect 145825 31720 145905 31730
rect 146145 31720 146225 31730
rect 141745 31640 141755 31720
rect 142065 31640 142075 31720
rect 145265 31640 145275 31720
rect 145585 31640 145595 31720
rect 145905 31640 145915 31720
rect 146225 31640 146235 31720
rect 146780 31700 146790 31780
rect 146540 31620 146620 31630
rect 146860 31620 146940 31630
rect 141825 31560 141905 31570
rect 142145 31560 142200 31570
rect 145345 31560 145425 31570
rect 145665 31560 145745 31570
rect 145985 31560 146065 31570
rect 141905 31480 141915 31560
rect 145425 31480 145435 31560
rect 145745 31480 145755 31560
rect 146065 31480 146075 31560
rect 146620 31540 146630 31620
rect 146940 31540 146950 31620
rect 146700 31460 146780 31470
rect 147020 31460 147100 31470
rect 141665 31400 141745 31410
rect 141985 31400 142065 31410
rect 145200 31400 145265 31410
rect 145505 31400 145585 31410
rect 145825 31400 145905 31410
rect 146145 31400 146225 31410
rect 141745 31320 141755 31400
rect 142065 31320 142075 31400
rect 145265 31320 145275 31400
rect 145585 31320 145595 31400
rect 145905 31320 145915 31400
rect 146225 31320 146235 31400
rect 146780 31380 146790 31460
rect 146540 31300 146620 31310
rect 146860 31300 146940 31310
rect 141825 31240 141905 31250
rect 142145 31240 142200 31250
rect 145345 31240 145425 31250
rect 145665 31240 145745 31250
rect 145985 31240 146065 31250
rect 141905 31160 141915 31240
rect 145425 31160 145435 31240
rect 145745 31160 145755 31240
rect 146065 31160 146075 31240
rect 146620 31220 146630 31300
rect 146940 31220 146950 31300
rect 146700 31140 146780 31150
rect 147020 31140 147100 31150
rect 141665 31080 141745 31090
rect 141985 31080 142065 31090
rect 145200 31080 145265 31090
rect 145505 31080 145585 31090
rect 145825 31080 145905 31090
rect 146145 31080 146225 31090
rect 141745 31000 141755 31080
rect 142065 31000 142075 31080
rect 145265 31000 145275 31080
rect 145585 31000 145595 31080
rect 145905 31000 145915 31080
rect 146225 31000 146235 31080
rect 146780 31060 146790 31140
rect 146540 30980 146620 30990
rect 146860 30980 146940 30990
rect 141825 30920 141905 30930
rect 142145 30920 142200 30930
rect 145345 30920 145425 30930
rect 145665 30920 145745 30930
rect 145985 30920 146065 30930
rect 141905 30840 141915 30920
rect 145425 30840 145435 30920
rect 145745 30840 145755 30920
rect 146065 30840 146075 30920
rect 146620 30900 146630 30980
rect 146940 30900 146950 30980
rect 146700 30820 146780 30830
rect 147020 30820 147100 30830
rect 141665 30760 141745 30770
rect 141985 30760 142065 30770
rect 145200 30760 145265 30770
rect 145505 30760 145585 30770
rect 145825 30760 145905 30770
rect 146145 30760 146225 30770
rect 141745 30680 141755 30760
rect 142065 30680 142075 30760
rect 145265 30680 145275 30760
rect 145585 30680 145595 30760
rect 145905 30680 145915 30760
rect 146225 30680 146235 30760
rect 146780 30740 146790 30820
rect 146540 30660 146620 30670
rect 146860 30660 146940 30670
rect 141825 30600 141905 30610
rect 142145 30600 142200 30610
rect 145345 30600 145425 30610
rect 145665 30600 145745 30610
rect 145985 30600 146065 30610
rect 141905 30520 141915 30600
rect 145425 30520 145435 30600
rect 145745 30520 145755 30600
rect 146065 30520 146075 30600
rect 146620 30580 146630 30660
rect 146940 30580 146950 30660
rect 146700 30500 146780 30510
rect 147020 30500 147100 30510
rect 141665 30440 141745 30450
rect 141985 30440 142065 30450
rect 145200 30440 145265 30450
rect 145505 30440 145585 30450
rect 145825 30440 145905 30450
rect 146145 30440 146225 30450
rect 141745 30360 141755 30440
rect 142065 30360 142075 30440
rect 145265 30360 145275 30440
rect 145585 30360 145595 30440
rect 145905 30360 145915 30440
rect 146225 30360 146235 30440
rect 146780 30420 146790 30500
rect 48685 29570 48765 29580
rect 62185 29570 62265 29580
rect 75685 29570 75765 29580
rect 89185 29570 89265 29580
rect 102685 29570 102765 29580
rect 116185 29570 116265 29580
rect 129685 29570 129765 29580
rect 48765 29500 48775 29570
rect 62265 29500 62275 29570
rect 75765 29500 75775 29570
rect 89265 29500 89275 29570
rect 102765 29500 102775 29570
rect 116265 29500 116275 29570
rect 129765 29500 129775 29570
rect 48685 29490 48775 29500
rect 62185 29490 62275 29500
rect 75685 29490 75775 29500
rect 89185 29490 89275 29500
rect 102685 29490 102775 29500
rect 116185 29490 116275 29500
rect 129685 29490 129775 29500
rect 48685 29410 48765 29420
rect 62185 29410 62265 29420
rect 75685 29410 75765 29420
rect 89185 29410 89265 29420
rect 102685 29410 102765 29420
rect 116185 29410 116265 29420
rect 129685 29410 129765 29420
rect 48765 29340 48775 29410
rect 62265 29340 62275 29410
rect 75765 29340 75775 29410
rect 89265 29340 89275 29410
rect 102765 29340 102775 29410
rect 116265 29340 116275 29410
rect 129765 29340 129775 29410
rect 48685 29330 48775 29340
rect 62185 29330 62275 29340
rect 75685 29330 75775 29340
rect 89185 29330 89275 29340
rect 102685 29330 102775 29340
rect 116185 29330 116275 29340
rect 129685 29330 129775 29340
rect 48685 29250 48765 29260
rect 62185 29250 62265 29260
rect 75685 29250 75765 29260
rect 89185 29250 89265 29260
rect 102685 29250 102765 29260
rect 116185 29250 116265 29260
rect 129685 29250 129765 29260
rect 48765 29180 48775 29250
rect 62265 29180 62275 29250
rect 75765 29180 75775 29250
rect 89265 29180 89275 29250
rect 102765 29180 102775 29250
rect 116265 29180 116275 29250
rect 129765 29180 129775 29250
rect 48685 29170 48775 29180
rect 62185 29170 62275 29180
rect 75685 29170 75775 29180
rect 89185 29170 89275 29180
rect 102685 29170 102775 29180
rect 116185 29170 116275 29180
rect 129685 29170 129775 29180
rect 48685 29090 48765 29100
rect 62185 29090 62265 29100
rect 75685 29090 75765 29100
rect 89185 29090 89265 29100
rect 102685 29090 102765 29100
rect 116185 29090 116265 29100
rect 129685 29090 129765 29100
rect 48765 29020 48775 29090
rect 62265 29020 62275 29090
rect 75765 29020 75775 29090
rect 89265 29020 89275 29090
rect 102765 29020 102775 29090
rect 116265 29020 116275 29090
rect 129765 29020 129775 29090
rect 48685 29010 48775 29020
rect 62185 29010 62275 29020
rect 75685 29010 75775 29020
rect 89185 29010 89275 29020
rect 102685 29010 102775 29020
rect 116185 29010 116275 29020
rect 129685 29010 129775 29020
rect 48685 28930 48765 28940
rect 62185 28930 62265 28940
rect 75685 28930 75765 28940
rect 89185 28930 89265 28940
rect 102685 28930 102765 28940
rect 116185 28930 116265 28940
rect 129685 28930 129765 28940
rect 48765 28850 48775 28930
rect 62265 28850 62275 28930
rect 75765 28850 75775 28930
rect 89265 28850 89275 28930
rect 102765 28850 102775 28930
rect 116265 28850 116275 28930
rect 129765 28850 129775 28930
rect 60085 28115 60165 28125
rect 60265 28115 60345 28125
rect 73585 28115 73665 28125
rect 73765 28115 73845 28125
rect 87085 28115 87165 28125
rect 87265 28115 87345 28125
rect 100585 28115 100665 28125
rect 100765 28115 100845 28125
rect 114085 28115 114165 28125
rect 114265 28115 114345 28125
rect 127585 28115 127665 28125
rect 127765 28115 127845 28125
rect 141085 28115 141165 28125
rect 141265 28115 141345 28125
rect 60165 28035 60175 28115
rect 60345 28035 60355 28115
rect 73665 28035 73675 28115
rect 73845 28035 73855 28115
rect 87165 28035 87175 28115
rect 87345 28035 87355 28115
rect 100665 28035 100675 28115
rect 100845 28035 100855 28115
rect 114165 28035 114175 28115
rect 114345 28035 114355 28115
rect 127665 28035 127675 28115
rect 127845 28035 127855 28115
rect 141165 28035 141175 28115
rect 141345 28035 141355 28115
rect 60085 27935 60165 27945
rect 60265 27935 60345 27945
rect 73585 27935 73665 27945
rect 73765 27935 73845 27945
rect 87085 27935 87165 27945
rect 87265 27935 87345 27945
rect 100585 27935 100665 27945
rect 100765 27935 100845 27945
rect 114085 27935 114165 27945
rect 114265 27935 114345 27945
rect 127585 27935 127665 27945
rect 127765 27935 127845 27945
rect 141085 27935 141165 27945
rect 141265 27935 141345 27945
rect 60165 27855 60175 27935
rect 60345 27855 60355 27935
rect 73665 27855 73675 27935
rect 73845 27855 73855 27935
rect 87165 27855 87175 27935
rect 87345 27855 87355 27935
rect 100665 27855 100675 27935
rect 100845 27855 100855 27935
rect 114165 27855 114175 27935
rect 114345 27855 114355 27935
rect 127665 27855 127675 27935
rect 127845 27855 127855 27935
rect 141165 27855 141175 27935
rect 141345 27855 141355 27935
rect 60085 27755 60165 27765
rect 60265 27755 60345 27765
rect 73585 27755 73665 27765
rect 73765 27755 73845 27765
rect 87085 27755 87165 27765
rect 87265 27755 87345 27765
rect 100585 27755 100665 27765
rect 100765 27755 100845 27765
rect 114085 27755 114165 27765
rect 114265 27755 114345 27765
rect 127585 27755 127665 27765
rect 127765 27755 127845 27765
rect 141085 27755 141165 27765
rect 141265 27755 141345 27765
rect 60165 27675 60175 27755
rect 60345 27675 60355 27755
rect 73665 27675 73675 27755
rect 73845 27675 73855 27755
rect 87165 27675 87175 27755
rect 87345 27675 87355 27755
rect 100665 27675 100675 27755
rect 100845 27675 100855 27755
rect 114165 27675 114175 27755
rect 114345 27675 114355 27755
rect 127665 27675 127675 27755
rect 127845 27675 127855 27755
rect 141165 27675 141175 27755
rect 141345 27675 141355 27755
rect 60085 27575 60165 27585
rect 60265 27575 60345 27585
rect 73585 27575 73665 27585
rect 73765 27575 73845 27585
rect 87085 27575 87165 27585
rect 87265 27575 87345 27585
rect 100585 27575 100665 27585
rect 100765 27575 100845 27585
rect 114085 27575 114165 27585
rect 114265 27575 114345 27585
rect 127585 27575 127665 27585
rect 127765 27575 127845 27585
rect 141085 27575 141165 27585
rect 141265 27575 141345 27585
rect 60165 27495 60175 27575
rect 60345 27495 60355 27575
rect 73665 27495 73675 27575
rect 73845 27495 73855 27575
rect 87165 27495 87175 27575
rect 87345 27495 87355 27575
rect 100665 27495 100675 27575
rect 100845 27495 100855 27575
rect 114165 27495 114175 27575
rect 114345 27495 114355 27575
rect 127665 27495 127675 27575
rect 127845 27495 127855 27575
rect 141165 27495 141175 27575
rect 141345 27495 141355 27575
rect 60085 27395 60165 27405
rect 60265 27395 60345 27405
rect 73585 27395 73665 27405
rect 73765 27395 73845 27405
rect 87085 27395 87165 27405
rect 87265 27395 87345 27405
rect 100585 27395 100665 27405
rect 100765 27395 100845 27405
rect 114085 27395 114165 27405
rect 114265 27395 114345 27405
rect 127585 27395 127665 27405
rect 127765 27395 127845 27405
rect 141085 27395 141165 27405
rect 141265 27395 141345 27405
rect 60165 27315 60175 27395
rect 60345 27315 60355 27395
rect 73665 27315 73675 27395
rect 73845 27315 73855 27395
rect 87165 27315 87175 27395
rect 87345 27315 87355 27395
rect 100665 27315 100675 27395
rect 100845 27315 100855 27395
rect 114165 27315 114175 27395
rect 114345 27315 114355 27395
rect 127665 27315 127675 27395
rect 127845 27315 127855 27395
rect 141165 27315 141175 27395
rect 141345 27315 141355 27395
rect 48500 26630 48605 26700
rect 48500 26620 48640 26630
rect 48710 26620 48790 26630
rect 60060 26620 60140 26630
rect 60210 26620 60290 26630
rect 60360 26620 60440 26630
rect 62060 26620 62140 26630
rect 62210 26620 62290 26630
rect 73560 26620 73640 26630
rect 73710 26620 73790 26630
rect 73860 26620 73940 26630
rect 75560 26620 75640 26630
rect 75710 26620 75790 26630
rect 87060 26620 87140 26630
rect 87210 26620 87290 26630
rect 87360 26620 87440 26630
rect 89060 26620 89140 26630
rect 89210 26620 89290 26630
rect 100560 26620 100640 26630
rect 100710 26620 100790 26630
rect 100860 26620 100940 26630
rect 102560 26620 102640 26630
rect 102710 26620 102790 26630
rect 114060 26620 114140 26630
rect 114210 26620 114290 26630
rect 114360 26620 114440 26630
rect 116060 26620 116140 26630
rect 116210 26620 116290 26630
rect 127560 26620 127640 26630
rect 127710 26620 127790 26630
rect 127860 26620 127940 26630
rect 129560 26620 129640 26630
rect 129710 26620 129790 26630
rect 141060 26620 141140 26630
rect 141210 26620 141290 26630
rect 141360 26620 141440 26630
rect 43060 26500 43140 26510
rect 43380 26500 43460 26510
rect 43140 26420 43150 26500
rect 43460 26420 43470 26500
rect 48500 26450 48605 26620
rect 48640 26540 48650 26620
rect 48790 26540 48800 26620
rect 49180 26570 49210 26600
rect 49300 26570 49330 26600
rect 49420 26570 49450 26600
rect 49540 26570 49570 26600
rect 49660 26570 49690 26600
rect 49780 26570 49810 26600
rect 49900 26570 49930 26600
rect 50020 26570 50050 26600
rect 50140 26570 50170 26600
rect 50260 26570 50290 26600
rect 50380 26570 50410 26600
rect 50500 26570 50530 26600
rect 50620 26570 50650 26600
rect 50740 26570 50770 26600
rect 50860 26570 50890 26600
rect 50980 26570 51010 26600
rect 51100 26570 51130 26600
rect 51220 26570 51250 26600
rect 51340 26570 51370 26600
rect 51460 26570 51490 26600
rect 51580 26570 51610 26600
rect 51700 26570 51730 26600
rect 51820 26570 51850 26600
rect 51940 26570 51970 26600
rect 52060 26570 52090 26600
rect 52180 26570 52210 26600
rect 52300 26570 52330 26600
rect 52420 26570 52450 26600
rect 52540 26570 52570 26600
rect 52660 26570 52690 26600
rect 52780 26570 52810 26600
rect 52900 26570 52930 26600
rect 53020 26570 53050 26600
rect 53140 26570 53170 26600
rect 53260 26570 53290 26600
rect 53380 26570 53410 26600
rect 53500 26570 53530 26600
rect 53620 26570 53650 26600
rect 53740 26570 53770 26600
rect 53860 26570 53890 26600
rect 53980 26570 54010 26600
rect 54100 26570 54130 26600
rect 54220 26570 54250 26600
rect 54340 26570 54370 26600
rect 54460 26570 54490 26600
rect 54580 26570 54610 26600
rect 54700 26570 54730 26600
rect 54820 26570 54850 26600
rect 54940 26570 54970 26600
rect 55060 26570 55090 26600
rect 55180 26570 55210 26600
rect 55300 26570 55330 26600
rect 55420 26570 55450 26600
rect 55540 26570 55570 26600
rect 55660 26570 55690 26600
rect 55780 26570 55810 26600
rect 55900 26570 55930 26600
rect 56020 26570 56050 26600
rect 56140 26570 56170 26600
rect 56260 26570 56290 26600
rect 56380 26570 56410 26600
rect 56500 26570 56530 26600
rect 56620 26570 56650 26600
rect 56740 26570 56770 26600
rect 56860 26570 56890 26600
rect 56980 26570 57010 26600
rect 57100 26570 57130 26600
rect 57220 26570 57250 26600
rect 57340 26570 57370 26600
rect 57460 26570 57490 26600
rect 57580 26570 57610 26600
rect 57700 26570 57730 26600
rect 57820 26570 57850 26600
rect 57940 26570 57970 26600
rect 58060 26570 58090 26600
rect 58180 26570 58210 26600
rect 58300 26570 58330 26600
rect 58420 26570 58450 26600
rect 58540 26570 58570 26600
rect 58660 26570 58690 26600
rect 58780 26570 58810 26600
rect 58900 26570 58930 26600
rect 59020 26570 59050 26600
rect 59140 26570 59170 26600
rect 59260 26570 59290 26600
rect 59380 26570 59410 26600
rect 59500 26570 59530 26600
rect 59620 26570 59650 26600
rect 59740 26570 59770 26600
rect 49060 26540 49120 26570
rect 49180 26540 49240 26570
rect 49300 26540 49360 26570
rect 49420 26540 49480 26570
rect 49540 26540 49600 26570
rect 49660 26540 49720 26570
rect 49780 26540 49840 26570
rect 49900 26540 49960 26570
rect 50020 26540 50080 26570
rect 50140 26540 50200 26570
rect 50260 26540 50320 26570
rect 50380 26540 50440 26570
rect 50500 26540 50560 26570
rect 50620 26540 50680 26570
rect 50740 26540 50800 26570
rect 50860 26540 50920 26570
rect 50980 26540 51040 26570
rect 51100 26540 51160 26570
rect 51220 26540 51280 26570
rect 51340 26540 51400 26570
rect 51460 26540 51520 26570
rect 51580 26540 51640 26570
rect 51700 26540 51760 26570
rect 51820 26540 51880 26570
rect 51940 26540 52000 26570
rect 52060 26540 52120 26570
rect 52180 26540 52240 26570
rect 52300 26540 52360 26570
rect 52420 26540 52480 26570
rect 52540 26540 52600 26570
rect 52660 26540 52720 26570
rect 52780 26540 52840 26570
rect 52900 26540 52960 26570
rect 53020 26540 53080 26570
rect 53140 26540 53200 26570
rect 53260 26540 53320 26570
rect 53380 26540 53440 26570
rect 53500 26540 53560 26570
rect 53620 26540 53680 26570
rect 53740 26540 53800 26570
rect 53860 26540 53920 26570
rect 53980 26540 54040 26570
rect 54100 26540 54160 26570
rect 54220 26540 54280 26570
rect 54340 26540 54400 26570
rect 54460 26540 54520 26570
rect 54580 26540 54640 26570
rect 54700 26540 54760 26570
rect 54820 26540 54880 26570
rect 54940 26540 55000 26570
rect 55060 26540 55120 26570
rect 55180 26540 55240 26570
rect 55300 26540 55360 26570
rect 55420 26540 55480 26570
rect 55540 26540 55600 26570
rect 55660 26540 55720 26570
rect 55780 26540 55840 26570
rect 55900 26540 55960 26570
rect 56020 26540 56080 26570
rect 56140 26540 56200 26570
rect 56260 26540 56320 26570
rect 56380 26540 56440 26570
rect 56500 26540 56560 26570
rect 56620 26540 56680 26570
rect 56740 26540 56800 26570
rect 56860 26540 56920 26570
rect 56980 26540 57040 26570
rect 57100 26540 57160 26570
rect 57220 26540 57280 26570
rect 57340 26540 57400 26570
rect 57460 26540 57520 26570
rect 57580 26540 57640 26570
rect 57700 26540 57760 26570
rect 57820 26540 57880 26570
rect 57940 26540 58000 26570
rect 58060 26540 58120 26570
rect 58180 26540 58240 26570
rect 58300 26540 58360 26570
rect 58420 26540 58480 26570
rect 58540 26540 58600 26570
rect 58660 26540 58720 26570
rect 58780 26540 58840 26570
rect 58900 26540 58960 26570
rect 59020 26540 59080 26570
rect 59140 26540 59200 26570
rect 59260 26540 59320 26570
rect 59380 26540 59440 26570
rect 59500 26540 59560 26570
rect 59620 26540 59680 26570
rect 59740 26540 59800 26570
rect 60140 26540 60150 26620
rect 60290 26540 60300 26620
rect 60440 26540 60450 26620
rect 62140 26540 62150 26620
rect 62290 26540 62300 26620
rect 62680 26570 62710 26600
rect 73245 26570 73270 26600
rect 62560 26540 62620 26570
rect 62680 26540 62740 26570
rect 73245 26540 73300 26570
rect 73640 26540 73650 26620
rect 73790 26540 73800 26620
rect 73940 26540 73950 26620
rect 75640 26540 75650 26620
rect 75790 26540 75800 26620
rect 76180 26570 76210 26600
rect 86745 26570 86770 26600
rect 76060 26540 76120 26570
rect 76180 26540 76240 26570
rect 86745 26540 86800 26570
rect 87140 26540 87150 26620
rect 87290 26540 87300 26620
rect 87440 26540 87450 26620
rect 89140 26540 89150 26620
rect 89290 26540 89300 26620
rect 89680 26570 89710 26600
rect 100245 26570 100270 26600
rect 89560 26540 89620 26570
rect 89680 26540 89740 26570
rect 100245 26540 100300 26570
rect 100640 26540 100650 26620
rect 100790 26540 100800 26620
rect 100940 26540 100950 26620
rect 102640 26540 102650 26620
rect 102790 26540 102800 26620
rect 103180 26570 103210 26600
rect 113745 26570 113770 26600
rect 103060 26540 103120 26570
rect 103180 26540 103240 26570
rect 113745 26540 113800 26570
rect 114140 26540 114150 26620
rect 114290 26540 114300 26620
rect 114440 26540 114450 26620
rect 116140 26540 116150 26620
rect 116290 26540 116300 26620
rect 116680 26570 116710 26600
rect 127245 26570 127270 26600
rect 116560 26540 116620 26570
rect 116680 26540 116740 26570
rect 127245 26540 127300 26570
rect 127640 26540 127650 26620
rect 127790 26540 127800 26620
rect 127940 26540 127950 26620
rect 129640 26540 129650 26620
rect 129790 26540 129800 26620
rect 130180 26570 130210 26600
rect 130060 26540 130120 26570
rect 130180 26540 130240 26570
rect 141140 26540 141150 26620
rect 141290 26540 141300 26620
rect 141440 26540 141450 26620
rect 49180 26450 49210 26480
rect 49300 26450 49330 26480
rect 49420 26450 49450 26480
rect 49540 26450 49570 26480
rect 49660 26450 49690 26480
rect 49780 26450 49810 26480
rect 49900 26450 49930 26480
rect 50020 26450 50050 26480
rect 50140 26450 50170 26480
rect 50260 26450 50290 26480
rect 50380 26450 50410 26480
rect 50500 26450 50530 26480
rect 50620 26450 50650 26480
rect 50740 26450 50770 26480
rect 50860 26450 50890 26480
rect 50980 26450 51010 26480
rect 51100 26450 51130 26480
rect 51220 26450 51250 26480
rect 51340 26450 51370 26480
rect 51460 26450 51490 26480
rect 51580 26450 51610 26480
rect 51700 26450 51730 26480
rect 51820 26450 51850 26480
rect 51940 26450 51970 26480
rect 52060 26450 52090 26480
rect 52180 26450 52210 26480
rect 52300 26450 52330 26480
rect 52420 26450 52450 26480
rect 52540 26450 52570 26480
rect 52660 26450 52690 26480
rect 52780 26450 52810 26480
rect 52900 26450 52930 26480
rect 53020 26450 53050 26480
rect 53140 26450 53170 26480
rect 53260 26450 53290 26480
rect 53380 26450 53410 26480
rect 53500 26450 53530 26480
rect 53620 26450 53650 26480
rect 53740 26450 53770 26480
rect 53860 26450 53890 26480
rect 53980 26450 54010 26480
rect 54100 26450 54130 26480
rect 54220 26450 54250 26480
rect 54340 26450 54370 26480
rect 54460 26450 54490 26480
rect 54580 26450 54610 26480
rect 54700 26450 54730 26480
rect 54820 26450 54850 26480
rect 54940 26450 54970 26480
rect 55060 26450 55090 26480
rect 55180 26450 55210 26480
rect 55300 26450 55330 26480
rect 55420 26450 55450 26480
rect 55540 26450 55570 26480
rect 55660 26450 55690 26480
rect 55780 26450 55810 26480
rect 55900 26450 55930 26480
rect 56020 26450 56050 26480
rect 56140 26450 56170 26480
rect 56260 26450 56290 26480
rect 56380 26450 56410 26480
rect 56500 26450 56530 26480
rect 56620 26450 56650 26480
rect 56740 26450 56770 26480
rect 56860 26450 56890 26480
rect 56980 26450 57010 26480
rect 57100 26450 57130 26480
rect 57220 26450 57250 26480
rect 57340 26450 57370 26480
rect 57460 26450 57490 26480
rect 57580 26450 57610 26480
rect 57700 26450 57730 26480
rect 57820 26450 57850 26480
rect 57940 26450 57970 26480
rect 58060 26450 58090 26480
rect 58180 26450 58210 26480
rect 58300 26450 58330 26480
rect 58420 26450 58450 26480
rect 58540 26450 58570 26480
rect 58660 26450 58690 26480
rect 58780 26450 58810 26480
rect 58900 26450 58930 26480
rect 59020 26450 59050 26480
rect 59140 26450 59170 26480
rect 59260 26450 59290 26480
rect 59380 26450 59410 26480
rect 59500 26450 59530 26480
rect 59620 26450 59650 26480
rect 59740 26450 59770 26480
rect 62680 26450 62710 26480
rect 73245 26450 73270 26480
rect 76180 26450 76210 26480
rect 86745 26450 86770 26480
rect 89680 26450 89710 26480
rect 100245 26450 100270 26480
rect 103180 26450 103210 26480
rect 113745 26450 113770 26480
rect 116680 26450 116710 26480
rect 127245 26450 127270 26480
rect 130180 26450 130210 26480
rect 48500 26440 48640 26450
rect 48710 26440 48790 26450
rect 44065 26410 44145 26420
rect 44385 26410 44465 26420
rect 44705 26410 44785 26420
rect 45025 26410 45105 26420
rect 45345 26410 45425 26420
rect 45665 26410 45745 26420
rect 45985 26410 46065 26420
rect 46305 26410 46385 26420
rect 46625 26410 46705 26420
rect 46945 26410 47025 26420
rect 47265 26410 47345 26420
rect 47585 26410 47665 26420
rect 47905 26410 47985 26420
rect 48225 26410 48305 26420
rect 42950 26340 42980 26350
rect 43220 26340 43300 26350
rect 42980 26260 42990 26340
rect 43300 26260 43310 26340
rect 44145 26330 44155 26410
rect 44465 26330 44475 26410
rect 44785 26330 44795 26410
rect 45105 26330 45115 26410
rect 45425 26330 45435 26410
rect 45745 26330 45755 26410
rect 46065 26330 46075 26410
rect 46385 26330 46395 26410
rect 46705 26330 46715 26410
rect 47025 26330 47035 26410
rect 47345 26330 47355 26410
rect 47665 26330 47675 26410
rect 47985 26330 47995 26410
rect 48305 26330 48315 26410
rect 48500 26270 48605 26440
rect 48640 26360 48650 26440
rect 48790 26360 48800 26440
rect 49060 26420 49120 26450
rect 49180 26420 49240 26450
rect 49300 26420 49360 26450
rect 49420 26420 49480 26450
rect 49540 26420 49600 26450
rect 49660 26420 49720 26450
rect 49780 26420 49840 26450
rect 49900 26420 49960 26450
rect 50020 26420 50080 26450
rect 50140 26420 50200 26450
rect 50260 26420 50320 26450
rect 50380 26420 50440 26450
rect 50500 26420 50560 26450
rect 50620 26420 50680 26450
rect 50740 26420 50800 26450
rect 50860 26420 50920 26450
rect 50980 26420 51040 26450
rect 51100 26420 51160 26450
rect 51220 26420 51280 26450
rect 51340 26420 51400 26450
rect 51460 26420 51520 26450
rect 51580 26420 51640 26450
rect 51700 26420 51760 26450
rect 51820 26420 51880 26450
rect 51940 26420 52000 26450
rect 52060 26420 52120 26450
rect 52180 26420 52240 26450
rect 52300 26420 52360 26450
rect 52420 26420 52480 26450
rect 52540 26420 52600 26450
rect 52660 26420 52720 26450
rect 52780 26420 52840 26450
rect 52900 26420 52960 26450
rect 53020 26420 53080 26450
rect 53140 26420 53200 26450
rect 53260 26420 53320 26450
rect 53380 26420 53440 26450
rect 53500 26420 53560 26450
rect 53620 26420 53680 26450
rect 53740 26420 53800 26450
rect 53860 26420 53920 26450
rect 53980 26420 54040 26450
rect 54100 26420 54160 26450
rect 54220 26420 54280 26450
rect 54340 26420 54400 26450
rect 54460 26420 54520 26450
rect 54580 26420 54640 26450
rect 54700 26420 54760 26450
rect 54820 26420 54880 26450
rect 54940 26420 55000 26450
rect 55060 26420 55120 26450
rect 55180 26420 55240 26450
rect 55300 26420 55360 26450
rect 55420 26420 55480 26450
rect 55540 26420 55600 26450
rect 55660 26420 55720 26450
rect 55780 26420 55840 26450
rect 55900 26420 55960 26450
rect 56020 26420 56080 26450
rect 56140 26420 56200 26450
rect 56260 26420 56320 26450
rect 56380 26420 56440 26450
rect 56500 26420 56560 26450
rect 56620 26420 56680 26450
rect 56740 26420 56800 26450
rect 56860 26420 56920 26450
rect 56980 26420 57040 26450
rect 57100 26420 57160 26450
rect 57220 26420 57280 26450
rect 57340 26420 57400 26450
rect 57460 26420 57520 26450
rect 57580 26420 57640 26450
rect 57700 26420 57760 26450
rect 57820 26420 57880 26450
rect 57940 26420 58000 26450
rect 58060 26420 58120 26450
rect 58180 26420 58240 26450
rect 58300 26420 58360 26450
rect 58420 26420 58480 26450
rect 58540 26420 58600 26450
rect 58660 26420 58720 26450
rect 58780 26420 58840 26450
rect 58900 26420 58960 26450
rect 59020 26420 59080 26450
rect 59140 26420 59200 26450
rect 59260 26420 59320 26450
rect 59380 26420 59440 26450
rect 59500 26420 59560 26450
rect 59620 26420 59680 26450
rect 59740 26420 59800 26450
rect 60060 26440 60140 26450
rect 60210 26440 60290 26450
rect 60360 26440 60440 26450
rect 62060 26440 62140 26450
rect 62210 26440 62290 26450
rect 60140 26360 60150 26440
rect 60290 26360 60300 26440
rect 60440 26360 60450 26440
rect 60610 26410 60690 26420
rect 60930 26410 61010 26420
rect 61350 26410 61430 26420
rect 61670 26410 61750 26420
rect 49180 26300 49210 26360
rect 49300 26300 49330 26360
rect 49420 26300 49450 26360
rect 49540 26300 49570 26360
rect 49660 26300 49690 26360
rect 49780 26300 49810 26360
rect 49900 26300 49930 26360
rect 50020 26300 50050 26360
rect 50140 26300 50170 26360
rect 50260 26300 50290 26360
rect 50380 26300 50410 26360
rect 50500 26300 50530 26360
rect 50620 26300 50650 26360
rect 50740 26300 50770 26360
rect 50860 26300 50890 26360
rect 50980 26300 51010 26360
rect 51100 26300 51130 26360
rect 51220 26300 51250 26360
rect 51340 26300 51370 26360
rect 51460 26300 51490 26360
rect 51580 26300 51610 26360
rect 51700 26300 51730 26360
rect 51820 26300 51850 26360
rect 51940 26300 51970 26360
rect 52060 26300 52090 26360
rect 52180 26300 52210 26360
rect 52300 26300 52330 26360
rect 52420 26300 52450 26360
rect 52540 26300 52570 26360
rect 52660 26300 52690 26360
rect 52780 26300 52810 26360
rect 52900 26300 52930 26360
rect 53020 26300 53050 26360
rect 53140 26300 53170 26360
rect 53260 26300 53290 26360
rect 53380 26300 53410 26360
rect 53500 26300 53530 26360
rect 53620 26300 53650 26360
rect 53740 26300 53770 26360
rect 53860 26300 53890 26360
rect 53980 26300 54010 26360
rect 54100 26300 54130 26360
rect 54220 26300 54250 26360
rect 54340 26300 54370 26360
rect 54460 26300 54490 26360
rect 54580 26300 54610 26360
rect 54700 26300 54730 26360
rect 54820 26300 54850 26360
rect 54940 26300 54970 26360
rect 55060 26300 55090 26360
rect 55180 26300 55210 26360
rect 55300 26300 55330 26360
rect 55420 26300 55450 26360
rect 55540 26300 55570 26360
rect 55660 26300 55690 26360
rect 55780 26300 55810 26360
rect 55900 26300 55930 26360
rect 56020 26300 56050 26360
rect 56140 26300 56170 26360
rect 56260 26300 56290 26360
rect 56380 26300 56410 26360
rect 56500 26300 56530 26360
rect 56620 26300 56650 26360
rect 56740 26300 56770 26360
rect 56860 26300 56890 26360
rect 56980 26300 57010 26360
rect 57100 26300 57130 26360
rect 57220 26300 57250 26360
rect 57340 26300 57370 26360
rect 57460 26300 57490 26360
rect 57580 26300 57610 26360
rect 57700 26300 57730 26360
rect 57820 26300 57850 26360
rect 57940 26300 57970 26360
rect 58060 26300 58090 26360
rect 58180 26300 58210 26360
rect 58300 26300 58330 26360
rect 58420 26300 58450 26360
rect 58540 26300 58570 26360
rect 58660 26300 58690 26360
rect 58780 26300 58810 26360
rect 58900 26300 58930 26360
rect 59020 26300 59050 26360
rect 59140 26300 59170 26360
rect 59260 26300 59290 26360
rect 59380 26300 59410 26360
rect 59500 26300 59530 26360
rect 59620 26300 59650 26360
rect 59740 26300 59770 26360
rect 60690 26330 60700 26410
rect 61010 26330 61020 26410
rect 61430 26330 61440 26410
rect 61750 26330 61760 26410
rect 62140 26360 62150 26440
rect 62290 26360 62300 26440
rect 62560 26420 62620 26450
rect 62680 26420 62740 26450
rect 73245 26420 73300 26450
rect 73560 26440 73640 26450
rect 73710 26440 73790 26450
rect 73860 26440 73940 26450
rect 75560 26440 75640 26450
rect 75710 26440 75790 26450
rect 73640 26360 73650 26440
rect 73790 26360 73800 26440
rect 73940 26360 73950 26440
rect 74110 26410 74190 26420
rect 74430 26410 74510 26420
rect 74850 26410 74930 26420
rect 75170 26410 75250 26420
rect 62680 26300 62710 26360
rect 73245 26300 73270 26360
rect 74190 26330 74200 26410
rect 74510 26330 74520 26410
rect 74930 26330 74940 26410
rect 75250 26330 75260 26410
rect 75640 26360 75650 26440
rect 75790 26360 75800 26440
rect 76060 26420 76120 26450
rect 76180 26420 76240 26450
rect 86745 26420 86800 26450
rect 87060 26440 87140 26450
rect 87210 26440 87290 26450
rect 87360 26440 87440 26450
rect 89060 26440 89140 26450
rect 89210 26440 89290 26450
rect 87140 26360 87150 26440
rect 87290 26360 87300 26440
rect 87440 26360 87450 26440
rect 87610 26410 87690 26420
rect 87930 26410 88010 26420
rect 88350 26410 88430 26420
rect 88670 26410 88750 26420
rect 76180 26300 76210 26360
rect 86745 26300 86770 26360
rect 87690 26330 87700 26410
rect 88010 26330 88020 26410
rect 88430 26330 88440 26410
rect 88750 26330 88760 26410
rect 89140 26360 89150 26440
rect 89290 26360 89300 26440
rect 89560 26420 89620 26450
rect 89680 26420 89740 26450
rect 100245 26420 100300 26450
rect 100560 26440 100640 26450
rect 100710 26440 100790 26450
rect 100860 26440 100940 26450
rect 102560 26440 102640 26450
rect 102710 26440 102790 26450
rect 100640 26360 100650 26440
rect 100790 26360 100800 26440
rect 100940 26360 100950 26440
rect 101110 26410 101190 26420
rect 101430 26410 101510 26420
rect 101850 26410 101930 26420
rect 102170 26410 102250 26420
rect 89680 26300 89710 26360
rect 100245 26300 100270 26360
rect 101190 26330 101200 26410
rect 101510 26330 101520 26410
rect 101930 26330 101940 26410
rect 102250 26330 102260 26410
rect 102640 26360 102650 26440
rect 102790 26360 102800 26440
rect 103060 26420 103120 26450
rect 103180 26420 103240 26450
rect 113745 26420 113800 26450
rect 114060 26440 114140 26450
rect 114210 26440 114290 26450
rect 114360 26440 114440 26450
rect 116060 26440 116140 26450
rect 116210 26440 116290 26450
rect 114140 26360 114150 26440
rect 114290 26360 114300 26440
rect 114440 26360 114450 26440
rect 114610 26410 114690 26420
rect 114930 26410 115010 26420
rect 115350 26410 115430 26420
rect 115670 26410 115750 26420
rect 103180 26300 103210 26360
rect 113745 26300 113770 26360
rect 114690 26330 114700 26410
rect 115010 26330 115020 26410
rect 115430 26330 115440 26410
rect 115750 26330 115760 26410
rect 116140 26360 116150 26440
rect 116290 26360 116300 26440
rect 116560 26420 116620 26450
rect 116680 26420 116740 26450
rect 127245 26420 127300 26450
rect 127560 26440 127640 26450
rect 127710 26440 127790 26450
rect 127860 26440 127940 26450
rect 129560 26440 129640 26450
rect 129710 26440 129790 26450
rect 127640 26360 127650 26440
rect 127790 26360 127800 26440
rect 127940 26360 127950 26440
rect 128110 26410 128190 26420
rect 128430 26410 128510 26420
rect 128850 26410 128930 26420
rect 129170 26410 129250 26420
rect 116680 26300 116710 26360
rect 127245 26300 127270 26360
rect 128190 26330 128200 26410
rect 128510 26330 128520 26410
rect 128930 26330 128940 26410
rect 129250 26330 129260 26410
rect 129640 26360 129650 26440
rect 129790 26360 129800 26440
rect 130060 26420 130120 26450
rect 130180 26420 130240 26450
rect 141060 26440 141140 26450
rect 141210 26440 141290 26450
rect 141360 26440 141440 26450
rect 141140 26360 141150 26440
rect 141290 26360 141300 26440
rect 141440 26360 141450 26440
rect 130180 26300 130210 26360
rect 48500 26260 48640 26270
rect 48710 26260 48790 26270
rect 60060 26260 60140 26270
rect 60210 26260 60290 26270
rect 60360 26260 60440 26270
rect 62060 26260 62140 26270
rect 62210 26260 62290 26270
rect 73560 26260 73640 26270
rect 73710 26260 73790 26270
rect 73860 26260 73940 26270
rect 75560 26260 75640 26270
rect 75710 26260 75790 26270
rect 87060 26260 87140 26270
rect 87210 26260 87290 26270
rect 87360 26260 87440 26270
rect 89060 26260 89140 26270
rect 89210 26260 89290 26270
rect 100560 26260 100640 26270
rect 100710 26260 100790 26270
rect 100860 26260 100940 26270
rect 102560 26260 102640 26270
rect 102710 26260 102790 26270
rect 114060 26260 114140 26270
rect 114210 26260 114290 26270
rect 114360 26260 114440 26270
rect 116060 26260 116140 26270
rect 116210 26260 116290 26270
rect 127560 26260 127640 26270
rect 127710 26260 127790 26270
rect 127860 26260 127940 26270
rect 129560 26260 129640 26270
rect 129710 26260 129790 26270
rect 141060 26260 141140 26270
rect 141210 26260 141290 26270
rect 141360 26260 141440 26270
rect 43905 26250 43985 26260
rect 44225 26250 44305 26260
rect 44545 26250 44625 26260
rect 44865 26250 44945 26260
rect 45185 26250 45265 26260
rect 45505 26250 45585 26260
rect 45825 26250 45905 26260
rect 46145 26250 46225 26260
rect 46465 26250 46545 26260
rect 46785 26250 46865 26260
rect 47105 26250 47185 26260
rect 47425 26250 47505 26260
rect 47745 26250 47825 26260
rect 48065 26250 48145 26260
rect 43060 26180 43140 26190
rect 43380 26180 43460 26190
rect 43140 26100 43150 26180
rect 43460 26100 43470 26180
rect 43985 26170 43995 26250
rect 44305 26170 44315 26250
rect 44625 26170 44635 26250
rect 44945 26170 44955 26250
rect 45265 26170 45275 26250
rect 45585 26170 45595 26250
rect 45905 26170 45915 26250
rect 46225 26170 46235 26250
rect 46545 26170 46555 26250
rect 46865 26170 46875 26250
rect 47185 26170 47195 26250
rect 47505 26170 47515 26250
rect 47825 26170 47835 26250
rect 48145 26170 48155 26250
rect 44065 26090 44145 26100
rect 44385 26090 44465 26100
rect 44705 26090 44785 26100
rect 45025 26090 45105 26100
rect 45345 26090 45425 26100
rect 45665 26090 45745 26100
rect 45985 26090 46065 26100
rect 46305 26090 46385 26100
rect 46625 26090 46705 26100
rect 46945 26090 47025 26100
rect 47265 26090 47345 26100
rect 47585 26090 47665 26100
rect 47905 26090 47985 26100
rect 48225 26090 48305 26100
rect 48500 26090 48605 26260
rect 48640 26180 48650 26260
rect 48790 26180 48800 26260
rect 60140 26180 60150 26260
rect 60290 26180 60300 26260
rect 60440 26180 60450 26260
rect 60770 26250 60850 26260
rect 61090 26250 61170 26260
rect 61510 26250 61590 26260
rect 61830 26250 61910 26260
rect 60850 26170 60860 26250
rect 61170 26170 61180 26250
rect 61590 26170 61600 26250
rect 61910 26170 61920 26250
rect 62140 26180 62150 26260
rect 62290 26180 62300 26260
rect 73640 26180 73650 26260
rect 73790 26180 73800 26260
rect 73940 26180 73950 26260
rect 74270 26250 74350 26260
rect 74590 26250 74670 26260
rect 75010 26250 75090 26260
rect 75330 26250 75410 26260
rect 74350 26170 74360 26250
rect 74670 26170 74680 26250
rect 75090 26170 75100 26250
rect 75410 26170 75420 26250
rect 75640 26180 75650 26260
rect 75790 26180 75800 26260
rect 87140 26180 87150 26260
rect 87290 26180 87300 26260
rect 87440 26180 87450 26260
rect 87770 26250 87850 26260
rect 88090 26250 88170 26260
rect 88510 26250 88590 26260
rect 88830 26250 88910 26260
rect 87850 26170 87860 26250
rect 88170 26170 88180 26250
rect 88590 26170 88600 26250
rect 88910 26170 88920 26250
rect 89140 26180 89150 26260
rect 89290 26180 89300 26260
rect 100640 26180 100650 26260
rect 100790 26180 100800 26260
rect 100940 26180 100950 26260
rect 101270 26250 101350 26260
rect 101590 26250 101670 26260
rect 102010 26250 102090 26260
rect 102330 26250 102410 26260
rect 101350 26170 101360 26250
rect 101670 26170 101680 26250
rect 102090 26170 102100 26250
rect 102410 26170 102420 26250
rect 102640 26180 102650 26260
rect 102790 26180 102800 26260
rect 114140 26180 114150 26260
rect 114290 26180 114300 26260
rect 114440 26180 114450 26260
rect 114770 26250 114850 26260
rect 115090 26250 115170 26260
rect 115510 26250 115590 26260
rect 115830 26250 115910 26260
rect 114850 26170 114860 26250
rect 115170 26170 115180 26250
rect 115590 26170 115600 26250
rect 115910 26170 115920 26250
rect 116140 26180 116150 26260
rect 116290 26180 116300 26260
rect 127640 26180 127650 26260
rect 127790 26180 127800 26260
rect 127940 26180 127950 26260
rect 128270 26250 128350 26260
rect 128590 26250 128670 26260
rect 129010 26250 129090 26260
rect 129330 26250 129410 26260
rect 128350 26170 128360 26250
rect 128670 26170 128680 26250
rect 129090 26170 129100 26250
rect 129410 26170 129420 26250
rect 129640 26180 129650 26260
rect 129790 26180 129800 26260
rect 141140 26180 141150 26260
rect 141290 26180 141300 26260
rect 141440 26180 141450 26260
rect 60610 26090 60690 26100
rect 60930 26090 61010 26100
rect 61350 26090 61430 26100
rect 61670 26090 61750 26100
rect 74110 26090 74190 26100
rect 74430 26090 74510 26100
rect 74850 26090 74930 26100
rect 75170 26090 75250 26100
rect 87610 26090 87690 26100
rect 87930 26090 88010 26100
rect 88350 26090 88430 26100
rect 88670 26090 88750 26100
rect 101110 26090 101190 26100
rect 101430 26090 101510 26100
rect 101850 26090 101930 26100
rect 102170 26090 102250 26100
rect 114610 26090 114690 26100
rect 114930 26090 115010 26100
rect 115350 26090 115430 26100
rect 115670 26090 115750 26100
rect 128110 26090 128190 26100
rect 128430 26090 128510 26100
rect 128850 26090 128930 26100
rect 129170 26090 129250 26100
rect 42950 26020 42980 26030
rect 43220 26020 43300 26030
rect 42980 25940 42990 26020
rect 43300 25940 43310 26020
rect 44145 26010 44155 26090
rect 44465 26010 44475 26090
rect 44785 26010 44795 26090
rect 45105 26010 45115 26090
rect 45425 26010 45435 26090
rect 45745 26010 45755 26090
rect 46065 26010 46075 26090
rect 46385 26010 46395 26090
rect 46705 26010 46715 26090
rect 47025 26010 47035 26090
rect 47345 26010 47355 26090
rect 47665 26010 47675 26090
rect 47985 26010 47995 26090
rect 48305 26010 48315 26090
rect 48500 26080 48640 26090
rect 48710 26080 48790 26090
rect 60060 26080 60140 26090
rect 60210 26080 60290 26090
rect 60360 26080 60440 26090
rect 43905 25930 43985 25940
rect 44225 25930 44305 25940
rect 44545 25930 44625 25940
rect 44865 25930 44945 25940
rect 45185 25930 45265 25940
rect 45505 25930 45585 25940
rect 45825 25930 45905 25940
rect 46145 25930 46225 25940
rect 46465 25930 46545 25940
rect 46785 25930 46865 25940
rect 47105 25930 47185 25940
rect 47425 25930 47505 25940
rect 47745 25930 47825 25940
rect 48065 25930 48145 25940
rect 43060 25860 43140 25870
rect 43380 25860 43460 25870
rect 43140 25780 43150 25860
rect 43460 25780 43470 25860
rect 43985 25850 43995 25930
rect 44305 25850 44315 25930
rect 44625 25850 44635 25930
rect 44945 25850 44955 25930
rect 45265 25850 45275 25930
rect 45585 25850 45595 25930
rect 45905 25850 45915 25930
rect 46225 25850 46235 25930
rect 46545 25850 46555 25930
rect 46865 25850 46875 25930
rect 47185 25850 47195 25930
rect 47505 25850 47515 25930
rect 47825 25850 47835 25930
rect 48145 25850 48155 25930
rect 48500 25910 48605 26080
rect 48640 26000 48650 26080
rect 48790 26000 48800 26080
rect 60140 26000 60150 26080
rect 60290 26000 60300 26080
rect 60440 26000 60450 26080
rect 60690 26010 60700 26090
rect 61010 26010 61020 26090
rect 61430 26010 61440 26090
rect 61750 26010 61760 26090
rect 62060 26080 62140 26090
rect 62210 26080 62290 26090
rect 73560 26080 73640 26090
rect 73710 26080 73790 26090
rect 73860 26080 73940 26090
rect 62140 26000 62150 26080
rect 62290 26000 62300 26080
rect 73640 26000 73650 26080
rect 73790 26000 73800 26080
rect 73940 26000 73950 26080
rect 74190 26010 74200 26090
rect 74510 26010 74520 26090
rect 74930 26010 74940 26090
rect 75250 26010 75260 26090
rect 75560 26080 75640 26090
rect 75710 26080 75790 26090
rect 87060 26080 87140 26090
rect 87210 26080 87290 26090
rect 87360 26080 87440 26090
rect 75640 26000 75650 26080
rect 75790 26000 75800 26080
rect 87140 26000 87150 26080
rect 87290 26000 87300 26080
rect 87440 26000 87450 26080
rect 87690 26010 87700 26090
rect 88010 26010 88020 26090
rect 88430 26010 88440 26090
rect 88750 26010 88760 26090
rect 89060 26080 89140 26090
rect 89210 26080 89290 26090
rect 100560 26080 100640 26090
rect 100710 26080 100790 26090
rect 100860 26080 100940 26090
rect 89140 26000 89150 26080
rect 89290 26000 89300 26080
rect 100640 26000 100650 26080
rect 100790 26000 100800 26080
rect 100940 26000 100950 26080
rect 101190 26010 101200 26090
rect 101510 26010 101520 26090
rect 101930 26010 101940 26090
rect 102250 26010 102260 26090
rect 102560 26080 102640 26090
rect 102710 26080 102790 26090
rect 114060 26080 114140 26090
rect 114210 26080 114290 26090
rect 114360 26080 114440 26090
rect 102640 26000 102650 26080
rect 102790 26000 102800 26080
rect 114140 26000 114150 26080
rect 114290 26000 114300 26080
rect 114440 26000 114450 26080
rect 114690 26010 114700 26090
rect 115010 26010 115020 26090
rect 115430 26010 115440 26090
rect 115750 26010 115760 26090
rect 116060 26080 116140 26090
rect 116210 26080 116290 26090
rect 127560 26080 127640 26090
rect 127710 26080 127790 26090
rect 127860 26080 127940 26090
rect 116140 26000 116150 26080
rect 116290 26000 116300 26080
rect 127640 26000 127650 26080
rect 127790 26000 127800 26080
rect 127940 26000 127950 26080
rect 128190 26010 128200 26090
rect 128510 26010 128520 26090
rect 128930 26010 128940 26090
rect 129250 26010 129260 26090
rect 129560 26080 129640 26090
rect 129710 26080 129790 26090
rect 141060 26080 141140 26090
rect 141210 26080 141290 26090
rect 141360 26080 141440 26090
rect 129640 26000 129650 26080
rect 129790 26000 129800 26080
rect 141140 26000 141150 26080
rect 141290 26000 141300 26080
rect 141440 26000 141450 26080
rect 60770 25930 60850 25940
rect 61090 25930 61170 25940
rect 61510 25930 61590 25940
rect 61830 25930 61910 25940
rect 74270 25930 74350 25940
rect 74590 25930 74670 25940
rect 75010 25930 75090 25940
rect 75330 25930 75410 25940
rect 87770 25930 87850 25940
rect 88090 25930 88170 25940
rect 88510 25930 88590 25940
rect 88830 25930 88910 25940
rect 101270 25930 101350 25940
rect 101590 25930 101670 25940
rect 102010 25930 102090 25940
rect 102330 25930 102410 25940
rect 114770 25930 114850 25940
rect 115090 25930 115170 25940
rect 115510 25930 115590 25940
rect 115830 25930 115910 25940
rect 128270 25930 128350 25940
rect 128590 25930 128670 25940
rect 129010 25930 129090 25940
rect 129330 25930 129410 25940
rect 48500 25900 48640 25910
rect 48710 25900 48790 25910
rect 60060 25900 60140 25910
rect 60210 25900 60290 25910
rect 60360 25900 60440 25910
rect 44065 25770 44145 25780
rect 44385 25770 44465 25780
rect 44705 25770 44785 25780
rect 45025 25770 45105 25780
rect 45345 25770 45425 25780
rect 45665 25770 45745 25780
rect 45985 25770 46065 25780
rect 46305 25770 46385 25780
rect 46625 25770 46705 25780
rect 46945 25770 47025 25780
rect 47265 25770 47345 25780
rect 47585 25770 47665 25780
rect 47905 25770 47985 25780
rect 48225 25770 48305 25780
rect 42950 25700 42980 25710
rect 43220 25700 43300 25710
rect 42980 25620 42990 25700
rect 43300 25620 43310 25700
rect 44145 25690 44155 25770
rect 44465 25690 44475 25770
rect 44785 25690 44795 25770
rect 45105 25690 45115 25770
rect 45425 25690 45435 25770
rect 45745 25690 45755 25770
rect 46065 25690 46075 25770
rect 46385 25690 46395 25770
rect 46705 25690 46715 25770
rect 47025 25690 47035 25770
rect 47345 25690 47355 25770
rect 47665 25690 47675 25770
rect 47985 25690 47995 25770
rect 48305 25690 48315 25770
rect 48500 25730 48605 25900
rect 48640 25820 48650 25900
rect 48790 25820 48800 25900
rect 60140 25820 60150 25900
rect 60290 25820 60300 25900
rect 60440 25820 60450 25900
rect 60850 25850 60860 25930
rect 61170 25850 61180 25930
rect 61590 25850 61600 25930
rect 61910 25850 61920 25930
rect 62060 25900 62140 25910
rect 62210 25900 62290 25910
rect 73560 25900 73640 25910
rect 73710 25900 73790 25910
rect 73860 25900 73940 25910
rect 62140 25820 62150 25900
rect 62290 25820 62300 25900
rect 73640 25820 73650 25900
rect 73790 25820 73800 25900
rect 73940 25820 73950 25900
rect 74350 25850 74360 25930
rect 74670 25850 74680 25930
rect 75090 25850 75100 25930
rect 75410 25850 75420 25930
rect 75560 25900 75640 25910
rect 75710 25900 75790 25910
rect 87060 25900 87140 25910
rect 87210 25900 87290 25910
rect 87360 25900 87440 25910
rect 75640 25820 75650 25900
rect 75790 25820 75800 25900
rect 87140 25820 87150 25900
rect 87290 25820 87300 25900
rect 87440 25820 87450 25900
rect 87850 25850 87860 25930
rect 88170 25850 88180 25930
rect 88590 25850 88600 25930
rect 88910 25850 88920 25930
rect 89060 25900 89140 25910
rect 89210 25900 89290 25910
rect 100560 25900 100640 25910
rect 100710 25900 100790 25910
rect 100860 25900 100940 25910
rect 89140 25820 89150 25900
rect 89290 25820 89300 25900
rect 100640 25820 100650 25900
rect 100790 25820 100800 25900
rect 100940 25820 100950 25900
rect 101350 25850 101360 25930
rect 101670 25850 101680 25930
rect 102090 25850 102100 25930
rect 102410 25850 102420 25930
rect 102560 25900 102640 25910
rect 102710 25900 102790 25910
rect 114060 25900 114140 25910
rect 114210 25900 114290 25910
rect 114360 25900 114440 25910
rect 102640 25820 102650 25900
rect 102790 25820 102800 25900
rect 114140 25820 114150 25900
rect 114290 25820 114300 25900
rect 114440 25820 114450 25900
rect 114850 25850 114860 25930
rect 115170 25850 115180 25930
rect 115590 25850 115600 25930
rect 115910 25850 115920 25930
rect 116060 25900 116140 25910
rect 116210 25900 116290 25910
rect 127560 25900 127640 25910
rect 127710 25900 127790 25910
rect 127860 25900 127940 25910
rect 116140 25820 116150 25900
rect 116290 25820 116300 25900
rect 127640 25820 127650 25900
rect 127790 25820 127800 25900
rect 127940 25820 127950 25900
rect 128350 25850 128360 25930
rect 128670 25850 128680 25930
rect 129090 25850 129100 25930
rect 129410 25850 129420 25930
rect 129560 25900 129640 25910
rect 129710 25900 129790 25910
rect 141060 25900 141140 25910
rect 141210 25900 141290 25910
rect 141360 25900 141440 25910
rect 129640 25820 129650 25900
rect 129790 25820 129800 25900
rect 141140 25820 141150 25900
rect 141290 25820 141300 25900
rect 141440 25820 141450 25900
rect 48500 25720 48640 25730
rect 48710 25720 48790 25730
rect 49270 25720 49350 25730
rect 49420 25720 49500 25730
rect 49570 25720 49650 25730
rect 43905 25610 43985 25620
rect 44225 25610 44305 25620
rect 44545 25610 44625 25620
rect 44865 25610 44945 25620
rect 45185 25610 45265 25620
rect 45505 25610 45585 25620
rect 45825 25610 45905 25620
rect 46145 25610 46225 25620
rect 46465 25610 46545 25620
rect 46785 25610 46865 25620
rect 47105 25610 47185 25620
rect 47425 25610 47505 25620
rect 47745 25610 47825 25620
rect 48065 25610 48145 25620
rect 43060 25540 43140 25550
rect 43380 25540 43460 25550
rect 43140 25460 43150 25540
rect 43460 25460 43470 25540
rect 43985 25530 43995 25610
rect 44305 25530 44315 25610
rect 44625 25530 44635 25610
rect 44945 25530 44955 25610
rect 45265 25530 45275 25610
rect 45585 25530 45595 25610
rect 45905 25530 45915 25610
rect 46225 25530 46235 25610
rect 46545 25530 46555 25610
rect 46865 25530 46875 25610
rect 47185 25530 47195 25610
rect 47505 25530 47515 25610
rect 47825 25530 47835 25610
rect 48145 25530 48155 25610
rect 48500 25550 48605 25720
rect 48640 25640 48650 25720
rect 48790 25640 48800 25720
rect 49350 25640 49360 25720
rect 49500 25640 49510 25720
rect 49650 25640 49660 25720
rect 48500 25540 48640 25550
rect 48710 25540 48790 25550
rect 49270 25540 49350 25550
rect 49420 25540 49500 25550
rect 49570 25540 49650 25550
rect 44065 25450 44145 25460
rect 44385 25450 44465 25460
rect 44705 25450 44785 25460
rect 45025 25450 45105 25460
rect 45345 25450 45425 25460
rect 45665 25450 45745 25460
rect 45985 25450 46065 25460
rect 46305 25450 46385 25460
rect 46625 25450 46705 25460
rect 46945 25450 47025 25460
rect 47265 25450 47345 25460
rect 47585 25450 47665 25460
rect 47905 25450 47985 25460
rect 48225 25450 48305 25460
rect 42950 25380 42980 25390
rect 43220 25380 43300 25390
rect 42980 25300 42990 25380
rect 43300 25300 43310 25380
rect 44145 25370 44155 25450
rect 44465 25370 44475 25450
rect 44785 25370 44795 25450
rect 45105 25370 45115 25450
rect 45425 25370 45435 25450
rect 45745 25370 45755 25450
rect 46065 25370 46075 25450
rect 46385 25370 46395 25450
rect 46705 25370 46715 25450
rect 47025 25370 47035 25450
rect 47345 25370 47355 25450
rect 47665 25370 47675 25450
rect 47985 25370 47995 25450
rect 48305 25370 48315 25450
rect 48500 25370 48605 25540
rect 48640 25460 48650 25540
rect 48790 25460 48800 25540
rect 49350 25460 49360 25540
rect 49500 25460 49510 25540
rect 49650 25460 49660 25540
rect 48500 25360 48640 25370
rect 48710 25360 48790 25370
rect 49270 25360 49350 25370
rect 49420 25360 49500 25370
rect 49570 25360 49650 25370
rect 43905 25290 43985 25300
rect 44225 25290 44305 25300
rect 44545 25290 44625 25300
rect 44865 25290 44945 25300
rect 45185 25290 45265 25300
rect 45505 25290 45585 25300
rect 45825 25290 45905 25300
rect 46145 25290 46225 25300
rect 46465 25290 46545 25300
rect 46785 25290 46865 25300
rect 47105 25290 47185 25300
rect 47425 25290 47505 25300
rect 47745 25290 47825 25300
rect 48065 25290 48145 25300
rect 43060 25220 43140 25230
rect 43380 25220 43460 25230
rect 43140 25140 43150 25220
rect 43460 25140 43470 25220
rect 43985 25210 43995 25290
rect 44305 25210 44315 25290
rect 44625 25210 44635 25290
rect 44945 25210 44955 25290
rect 45265 25210 45275 25290
rect 45585 25210 45595 25290
rect 45905 25210 45915 25290
rect 46225 25210 46235 25290
rect 46545 25210 46555 25290
rect 46865 25210 46875 25290
rect 47185 25210 47195 25290
rect 47505 25210 47515 25290
rect 47825 25210 47835 25290
rect 48145 25210 48155 25290
rect 48500 25190 48605 25360
rect 48640 25280 48650 25360
rect 48790 25280 48800 25360
rect 49350 25280 49360 25360
rect 49500 25280 49510 25360
rect 49650 25280 49660 25360
rect 48500 25180 48640 25190
rect 48710 25180 48790 25190
rect 49270 25180 49350 25190
rect 49420 25180 49500 25190
rect 49570 25180 49650 25190
rect 44065 25130 44145 25140
rect 44385 25130 44465 25140
rect 44705 25130 44785 25140
rect 45025 25130 45105 25140
rect 45345 25130 45425 25140
rect 45665 25130 45745 25140
rect 45985 25130 46065 25140
rect 46305 25130 46385 25140
rect 46625 25130 46705 25140
rect 46945 25130 47025 25140
rect 47265 25130 47345 25140
rect 47585 25130 47665 25140
rect 47905 25130 47985 25140
rect 48225 25130 48305 25140
rect 42950 25060 42980 25070
rect 43220 25060 43300 25070
rect 42980 24980 42990 25060
rect 43300 24980 43310 25060
rect 44145 25050 44155 25130
rect 44465 25050 44475 25130
rect 44785 25050 44795 25130
rect 45105 25050 45115 25130
rect 45425 25050 45435 25130
rect 45745 25050 45755 25130
rect 46065 25050 46075 25130
rect 46385 25050 46395 25130
rect 46705 25050 46715 25130
rect 47025 25050 47035 25130
rect 47345 25050 47355 25130
rect 47665 25050 47675 25130
rect 47985 25050 47995 25130
rect 48305 25050 48315 25130
rect 48500 25010 48605 25180
rect 48640 25100 48650 25180
rect 48790 25100 48800 25180
rect 49350 25100 49360 25180
rect 49500 25100 49510 25180
rect 49650 25100 49660 25180
rect 48500 25000 48640 25010
rect 48710 25000 48790 25010
rect 49270 25000 49350 25010
rect 49420 25000 49500 25010
rect 49570 25000 49650 25010
rect 43905 24970 43985 24980
rect 44225 24970 44305 24980
rect 44545 24970 44625 24980
rect 44865 24970 44945 24980
rect 45185 24970 45265 24980
rect 45505 24970 45585 24980
rect 45825 24970 45905 24980
rect 46145 24970 46225 24980
rect 46465 24970 46545 24980
rect 46785 24970 46865 24980
rect 47105 24970 47185 24980
rect 47425 24970 47505 24980
rect 47745 24970 47825 24980
rect 48065 24970 48145 24980
rect 43060 24900 43140 24910
rect 43380 24900 43460 24910
rect 43140 24820 43150 24900
rect 43460 24820 43470 24900
rect 43985 24890 43995 24970
rect 44305 24890 44315 24970
rect 44625 24890 44635 24970
rect 44945 24890 44955 24970
rect 45265 24890 45275 24970
rect 45585 24890 45595 24970
rect 45905 24890 45915 24970
rect 46225 24890 46235 24970
rect 46545 24890 46555 24970
rect 46865 24890 46875 24970
rect 47185 24890 47195 24970
rect 47505 24890 47515 24970
rect 47825 24890 47835 24970
rect 48145 24890 48155 24970
rect 48500 24830 48605 25000
rect 48640 24920 48650 25000
rect 48790 24920 48800 25000
rect 49350 24920 49360 25000
rect 49500 24920 49510 25000
rect 49650 24920 49660 25000
rect 48500 24820 48640 24830
rect 48710 24820 48790 24830
rect 49270 24820 49350 24830
rect 49420 24820 49500 24830
rect 49570 24820 49650 24830
rect 44065 24810 44145 24820
rect 44385 24810 44465 24820
rect 44705 24810 44785 24820
rect 45025 24810 45105 24820
rect 45345 24810 45425 24820
rect 45665 24810 45745 24820
rect 45985 24810 46065 24820
rect 46305 24810 46385 24820
rect 46625 24810 46705 24820
rect 46945 24810 47025 24820
rect 47265 24810 47345 24820
rect 47585 24810 47665 24820
rect 47905 24810 47985 24820
rect 48225 24810 48305 24820
rect 42950 24740 42980 24750
rect 43220 24740 43300 24750
rect 42980 24660 42990 24740
rect 43300 24660 43310 24740
rect 44145 24730 44155 24810
rect 44465 24730 44475 24810
rect 44785 24730 44795 24810
rect 45105 24730 45115 24810
rect 45425 24730 45435 24810
rect 45745 24730 45755 24810
rect 46065 24730 46075 24810
rect 46385 24730 46395 24810
rect 46705 24730 46715 24810
rect 47025 24730 47035 24810
rect 47345 24730 47355 24810
rect 47665 24730 47675 24810
rect 47985 24730 47995 24810
rect 48305 24730 48315 24810
rect 43905 24650 43985 24660
rect 44225 24650 44305 24660
rect 44545 24650 44625 24660
rect 44865 24650 44945 24660
rect 45185 24650 45265 24660
rect 45505 24650 45585 24660
rect 45825 24650 45905 24660
rect 46145 24650 46225 24660
rect 46465 24650 46545 24660
rect 46785 24650 46865 24660
rect 47105 24650 47185 24660
rect 47425 24650 47505 24660
rect 47745 24650 47825 24660
rect 48065 24650 48145 24660
rect 48500 24650 48605 24820
rect 48640 24740 48650 24820
rect 48790 24740 48800 24820
rect 49350 24740 49360 24820
rect 49500 24740 49510 24820
rect 49650 24740 49660 24820
rect 43060 24580 43140 24590
rect 43380 24580 43460 24590
rect 43140 24500 43150 24580
rect 43460 24500 43470 24580
rect 43985 24570 43995 24650
rect 44305 24570 44315 24650
rect 44625 24570 44635 24650
rect 44945 24570 44955 24650
rect 45265 24570 45275 24650
rect 45585 24570 45595 24650
rect 45905 24570 45915 24650
rect 46225 24570 46235 24650
rect 46545 24570 46555 24650
rect 46865 24570 46875 24650
rect 47185 24570 47195 24650
rect 47505 24570 47515 24650
rect 47825 24570 47835 24650
rect 48145 24570 48155 24650
rect 48500 24640 48640 24650
rect 48710 24640 48790 24650
rect 49270 24640 49350 24650
rect 49420 24640 49500 24650
rect 49570 24640 49650 24650
rect 44065 24490 44145 24500
rect 44385 24490 44465 24500
rect 44705 24490 44785 24500
rect 45025 24490 45105 24500
rect 45345 24490 45425 24500
rect 45665 24490 45745 24500
rect 45985 24490 46065 24500
rect 46305 24490 46385 24500
rect 46625 24490 46705 24500
rect 46945 24490 47025 24500
rect 47265 24490 47345 24500
rect 47585 24490 47665 24500
rect 47905 24490 47985 24500
rect 48225 24490 48305 24500
rect 42950 24420 42980 24430
rect 43220 24420 43300 24430
rect 42980 24340 42990 24420
rect 43300 24340 43310 24420
rect 44145 24410 44155 24490
rect 44465 24410 44475 24490
rect 44785 24410 44795 24490
rect 45105 24410 45115 24490
rect 45425 24410 45435 24490
rect 45745 24410 45755 24490
rect 46065 24410 46075 24490
rect 46385 24410 46395 24490
rect 46705 24410 46715 24490
rect 47025 24410 47035 24490
rect 47345 24410 47355 24490
rect 47665 24410 47675 24490
rect 47985 24410 47995 24490
rect 48305 24410 48315 24490
rect 48500 24470 48605 24640
rect 48640 24560 48650 24640
rect 48790 24560 48800 24640
rect 49350 24560 49360 24640
rect 49500 24560 49510 24640
rect 49650 24560 49660 24640
rect 48500 24460 48640 24470
rect 48710 24460 48790 24470
rect 49270 24460 49350 24470
rect 49420 24460 49500 24470
rect 49570 24460 49650 24470
rect 43905 24330 43985 24340
rect 44225 24330 44305 24340
rect 44545 24330 44625 24340
rect 44865 24330 44945 24340
rect 45185 24330 45265 24340
rect 45505 24330 45585 24340
rect 45825 24330 45905 24340
rect 46145 24330 46225 24340
rect 46465 24330 46545 24340
rect 46785 24330 46865 24340
rect 47105 24330 47185 24340
rect 47425 24330 47505 24340
rect 47745 24330 47825 24340
rect 48065 24330 48145 24340
rect 43060 24260 43140 24270
rect 43380 24260 43460 24270
rect 43140 24180 43150 24260
rect 43460 24180 43470 24260
rect 43985 24250 43995 24330
rect 44305 24250 44315 24330
rect 44625 24250 44635 24330
rect 44945 24250 44955 24330
rect 45265 24250 45275 24330
rect 45585 24250 45595 24330
rect 45905 24250 45915 24330
rect 46225 24250 46235 24330
rect 46545 24250 46555 24330
rect 46865 24250 46875 24330
rect 47185 24250 47195 24330
rect 47505 24250 47515 24330
rect 47825 24250 47835 24330
rect 48145 24250 48155 24330
rect 48500 24290 48605 24460
rect 48640 24380 48650 24460
rect 48790 24380 48800 24460
rect 49350 24380 49360 24460
rect 49500 24380 49510 24460
rect 49650 24380 49660 24460
rect 48500 24280 48640 24290
rect 48710 24280 48790 24290
rect 49270 24280 49350 24290
rect 49420 24280 49500 24290
rect 49570 24280 49650 24290
rect 44065 24170 44145 24180
rect 44385 24170 44465 24180
rect 44705 24170 44785 24180
rect 45025 24170 45105 24180
rect 45345 24170 45425 24180
rect 45665 24170 45745 24180
rect 45985 24170 46065 24180
rect 46305 24170 46385 24180
rect 46625 24170 46705 24180
rect 46945 24170 47025 24180
rect 47265 24170 47345 24180
rect 47585 24170 47665 24180
rect 47905 24170 47985 24180
rect 48225 24170 48305 24180
rect 42950 24100 42980 24110
rect 43220 24100 43300 24110
rect 42980 24020 42990 24100
rect 43300 24020 43310 24100
rect 44145 24090 44155 24170
rect 44465 24090 44475 24170
rect 44785 24090 44795 24170
rect 45105 24090 45115 24170
rect 45425 24090 45435 24170
rect 45745 24090 45755 24170
rect 46065 24090 46075 24170
rect 46385 24090 46395 24170
rect 46705 24090 46715 24170
rect 47025 24090 47035 24170
rect 47345 24090 47355 24170
rect 47665 24090 47675 24170
rect 47985 24090 47995 24170
rect 48305 24090 48315 24170
rect 48500 24110 48605 24280
rect 48640 24200 48650 24280
rect 48790 24200 48800 24280
rect 49350 24200 49360 24280
rect 49500 24200 49510 24280
rect 49650 24200 49660 24280
rect 48500 24100 48640 24110
rect 48710 24100 48790 24110
rect 49270 24100 49350 24110
rect 49420 24100 49500 24110
rect 49570 24100 49650 24110
rect 43905 24010 43985 24020
rect 44225 24010 44305 24020
rect 44545 24010 44625 24020
rect 44865 24010 44945 24020
rect 45185 24010 45265 24020
rect 45505 24010 45585 24020
rect 45825 24010 45905 24020
rect 46145 24010 46225 24020
rect 46465 24010 46545 24020
rect 46785 24010 46865 24020
rect 47105 24010 47185 24020
rect 47425 24010 47505 24020
rect 47745 24010 47825 24020
rect 48065 24010 48145 24020
rect 43060 23940 43140 23950
rect 43380 23940 43460 23950
rect 43140 23860 43150 23940
rect 43460 23860 43470 23940
rect 43985 23930 43995 24010
rect 44305 23930 44315 24010
rect 44625 23930 44635 24010
rect 44945 23930 44955 24010
rect 45265 23930 45275 24010
rect 45585 23930 45595 24010
rect 45905 23930 45915 24010
rect 46225 23930 46235 24010
rect 46545 23930 46555 24010
rect 46865 23930 46875 24010
rect 47185 23930 47195 24010
rect 47505 23930 47515 24010
rect 47825 23930 47835 24010
rect 48145 23930 48155 24010
rect 48500 23930 48605 24100
rect 48640 24020 48650 24100
rect 48790 24020 48800 24100
rect 49350 24020 49360 24100
rect 49500 24020 49510 24100
rect 49650 24020 49660 24100
rect 48500 23920 48640 23930
rect 48710 23920 48790 23930
rect 49270 23920 49350 23930
rect 49420 23920 49500 23930
rect 49570 23920 49650 23930
rect 44065 23850 44145 23860
rect 44385 23850 44465 23860
rect 44705 23850 44785 23860
rect 45025 23850 45105 23860
rect 45345 23850 45425 23860
rect 45665 23850 45745 23860
rect 45985 23850 46065 23860
rect 46305 23850 46385 23860
rect 46625 23850 46705 23860
rect 46945 23850 47025 23860
rect 47265 23850 47345 23860
rect 47585 23850 47665 23860
rect 47905 23850 47985 23860
rect 48225 23850 48305 23860
rect 42950 23780 42980 23790
rect 43220 23780 43300 23790
rect 42980 23700 42990 23780
rect 43300 23700 43310 23780
rect 44145 23770 44155 23850
rect 44465 23770 44475 23850
rect 44785 23770 44795 23850
rect 45105 23770 45115 23850
rect 45425 23770 45435 23850
rect 45745 23770 45755 23850
rect 46065 23770 46075 23850
rect 46385 23770 46395 23850
rect 46705 23770 46715 23850
rect 47025 23770 47035 23850
rect 47345 23770 47355 23850
rect 47665 23770 47675 23850
rect 47985 23770 47995 23850
rect 48305 23770 48315 23850
rect 48500 23750 48605 23920
rect 48640 23840 48650 23920
rect 48790 23840 48800 23920
rect 49350 23840 49360 23920
rect 49500 23840 49510 23920
rect 49650 23840 49660 23920
rect 48500 23740 48640 23750
rect 48710 23740 48790 23750
rect 49270 23740 49350 23750
rect 49420 23740 49500 23750
rect 49570 23740 49650 23750
rect 43905 23690 43985 23700
rect 44225 23690 44305 23700
rect 44545 23690 44625 23700
rect 44865 23690 44945 23700
rect 45185 23690 45265 23700
rect 45505 23690 45585 23700
rect 45825 23690 45905 23700
rect 46145 23690 46225 23700
rect 46465 23690 46545 23700
rect 46785 23690 46865 23700
rect 47105 23690 47185 23700
rect 47425 23690 47505 23700
rect 47745 23690 47825 23700
rect 48065 23690 48145 23700
rect 43060 23620 43140 23630
rect 43380 23620 43460 23630
rect 43140 23540 43150 23620
rect 43460 23540 43470 23620
rect 43985 23610 43995 23690
rect 44305 23610 44315 23690
rect 44625 23610 44635 23690
rect 44945 23610 44955 23690
rect 45265 23610 45275 23690
rect 45585 23610 45595 23690
rect 45905 23610 45915 23690
rect 46225 23610 46235 23690
rect 46545 23610 46555 23690
rect 46865 23610 46875 23690
rect 47185 23610 47195 23690
rect 47505 23610 47515 23690
rect 47825 23610 47835 23690
rect 48145 23610 48155 23690
rect 48500 23570 48605 23740
rect 48640 23660 48650 23740
rect 48790 23660 48800 23740
rect 49350 23660 49360 23740
rect 49500 23660 49510 23740
rect 49650 23660 49660 23740
rect 48500 23560 48640 23570
rect 48710 23560 48790 23570
rect 49270 23560 49350 23570
rect 49420 23560 49500 23570
rect 49570 23560 49650 23570
rect 44065 23530 44145 23540
rect 44385 23530 44465 23540
rect 44705 23530 44785 23540
rect 45025 23530 45105 23540
rect 45345 23530 45425 23540
rect 45665 23530 45745 23540
rect 45985 23530 46065 23540
rect 46305 23530 46385 23540
rect 46625 23530 46705 23540
rect 46945 23530 47025 23540
rect 47265 23530 47345 23540
rect 47585 23530 47665 23540
rect 47905 23530 47985 23540
rect 48225 23530 48305 23540
rect 42950 23460 42980 23470
rect 43220 23460 43300 23470
rect 42980 23380 42990 23460
rect 43300 23380 43310 23460
rect 44145 23450 44155 23530
rect 44465 23450 44475 23530
rect 44785 23450 44795 23530
rect 45105 23450 45115 23530
rect 45425 23450 45435 23530
rect 45745 23450 45755 23530
rect 46065 23450 46075 23530
rect 46385 23450 46395 23530
rect 46705 23450 46715 23530
rect 47025 23450 47035 23530
rect 47345 23450 47355 23530
rect 47665 23450 47675 23530
rect 47985 23450 47995 23530
rect 48305 23450 48315 23530
rect 48500 23390 48605 23560
rect 48640 23480 48650 23560
rect 48790 23480 48800 23560
rect 49350 23480 49360 23560
rect 49500 23480 49510 23560
rect 49650 23480 49660 23560
rect 48500 23380 48640 23390
rect 48710 23380 48790 23390
rect 49270 23380 49350 23390
rect 49420 23380 49500 23390
rect 49570 23380 49650 23390
rect 43905 23370 43985 23380
rect 44225 23370 44305 23380
rect 44545 23370 44625 23380
rect 44865 23370 44945 23380
rect 45185 23370 45265 23380
rect 45505 23370 45585 23380
rect 45825 23370 45905 23380
rect 46145 23370 46225 23380
rect 46465 23370 46545 23380
rect 46785 23370 46865 23380
rect 47105 23370 47185 23380
rect 47425 23370 47505 23380
rect 47745 23370 47825 23380
rect 48065 23370 48145 23380
rect 43060 23300 43140 23310
rect 43380 23300 43460 23310
rect 43140 23220 43150 23300
rect 43460 23220 43470 23300
rect 43985 23290 43995 23370
rect 44305 23290 44315 23370
rect 44625 23290 44635 23370
rect 44945 23290 44955 23370
rect 45265 23290 45275 23370
rect 45585 23290 45595 23370
rect 45905 23290 45915 23370
rect 46225 23290 46235 23370
rect 46545 23290 46555 23370
rect 46865 23290 46875 23370
rect 47185 23290 47195 23370
rect 47505 23290 47515 23370
rect 47825 23290 47835 23370
rect 48145 23290 48155 23370
rect 44065 23210 44145 23220
rect 44385 23210 44465 23220
rect 44705 23210 44785 23220
rect 45025 23210 45105 23220
rect 45345 23210 45425 23220
rect 45665 23210 45745 23220
rect 45985 23210 46065 23220
rect 46305 23210 46385 23220
rect 46625 23210 46705 23220
rect 46945 23210 47025 23220
rect 47265 23210 47345 23220
rect 47585 23210 47665 23220
rect 47905 23210 47985 23220
rect 48225 23210 48305 23220
rect 48500 23210 48605 23380
rect 48640 23300 48650 23380
rect 48790 23300 48800 23380
rect 49350 23300 49360 23380
rect 49500 23300 49510 23380
rect 49650 23300 49660 23380
rect 42950 23140 42980 23150
rect 43220 23140 43300 23150
rect 42980 23060 42990 23140
rect 43300 23060 43310 23140
rect 44145 23130 44155 23210
rect 44465 23130 44475 23210
rect 44785 23130 44795 23210
rect 45105 23130 45115 23210
rect 45425 23130 45435 23210
rect 45745 23130 45755 23210
rect 46065 23130 46075 23210
rect 46385 23130 46395 23210
rect 46705 23130 46715 23210
rect 47025 23130 47035 23210
rect 47345 23130 47355 23210
rect 47665 23130 47675 23210
rect 47985 23130 47995 23210
rect 48305 23130 48315 23210
rect 48500 23200 48640 23210
rect 48710 23200 48790 23210
rect 49270 23200 49350 23210
rect 49420 23200 49500 23210
rect 49570 23200 49650 23210
rect 43905 23050 43985 23060
rect 44225 23050 44305 23060
rect 44545 23050 44625 23060
rect 44865 23050 44945 23060
rect 45185 23050 45265 23060
rect 45505 23050 45585 23060
rect 45825 23050 45905 23060
rect 46145 23050 46225 23060
rect 46465 23050 46545 23060
rect 46785 23050 46865 23060
rect 47105 23050 47185 23060
rect 47425 23050 47505 23060
rect 47745 23050 47825 23060
rect 48065 23050 48145 23060
rect 43060 22980 43140 22990
rect 43380 22980 43460 22990
rect 43140 22900 43150 22980
rect 43460 22900 43470 22980
rect 43985 22970 43995 23050
rect 44305 22970 44315 23050
rect 44625 22970 44635 23050
rect 44945 22970 44955 23050
rect 45265 22970 45275 23050
rect 45585 22970 45595 23050
rect 45905 22970 45915 23050
rect 46225 22970 46235 23050
rect 46545 22970 46555 23050
rect 46865 22970 46875 23050
rect 47185 22970 47195 23050
rect 47505 22970 47515 23050
rect 47825 22970 47835 23050
rect 48145 22970 48155 23050
rect 48500 23030 48605 23200
rect 48640 23120 48650 23200
rect 48790 23120 48800 23200
rect 49350 23120 49360 23200
rect 49500 23120 49510 23200
rect 49650 23120 49660 23200
rect 48500 23020 48640 23030
rect 48710 23020 48790 23030
rect 49270 23020 49350 23030
rect 49420 23020 49500 23030
rect 49570 23020 49650 23030
rect 44065 22890 44145 22900
rect 44385 22890 44465 22900
rect 44705 22890 44785 22900
rect 45025 22890 45105 22900
rect 45345 22890 45425 22900
rect 45665 22890 45745 22900
rect 45985 22890 46065 22900
rect 46305 22890 46385 22900
rect 46625 22890 46705 22900
rect 46945 22890 47025 22900
rect 47265 22890 47345 22900
rect 47585 22890 47665 22900
rect 47905 22890 47985 22900
rect 48225 22890 48305 22900
rect 42950 22820 42980 22830
rect 43220 22820 43300 22830
rect 42980 22740 42990 22820
rect 43300 22740 43310 22820
rect 44145 22810 44155 22890
rect 44465 22810 44475 22890
rect 44785 22810 44795 22890
rect 45105 22810 45115 22890
rect 45425 22810 45435 22890
rect 45745 22810 45755 22890
rect 46065 22810 46075 22890
rect 46385 22810 46395 22890
rect 46705 22810 46715 22890
rect 47025 22810 47035 22890
rect 47345 22810 47355 22890
rect 47665 22810 47675 22890
rect 47985 22810 47995 22890
rect 48305 22810 48315 22890
rect 48500 22850 48605 23020
rect 48640 22940 48650 23020
rect 48790 22940 48800 23020
rect 49350 22940 49360 23020
rect 49500 22940 49510 23020
rect 49650 22940 49660 23020
rect 48500 22840 48640 22850
rect 48710 22840 48790 22850
rect 49270 22840 49350 22850
rect 49420 22840 49500 22850
rect 49570 22840 49650 22850
rect 43905 22730 43985 22740
rect 44225 22730 44305 22740
rect 44545 22730 44625 22740
rect 44865 22730 44945 22740
rect 45185 22730 45265 22740
rect 45505 22730 45585 22740
rect 45825 22730 45905 22740
rect 46145 22730 46225 22740
rect 46465 22730 46545 22740
rect 46785 22730 46865 22740
rect 47105 22730 47185 22740
rect 47425 22730 47505 22740
rect 47745 22730 47825 22740
rect 48065 22730 48145 22740
rect 43060 22660 43140 22670
rect 43380 22660 43460 22670
rect 43140 22580 43150 22660
rect 43460 22580 43470 22660
rect 43985 22650 43995 22730
rect 44305 22650 44315 22730
rect 44625 22650 44635 22730
rect 44945 22650 44955 22730
rect 45265 22650 45275 22730
rect 45585 22650 45595 22730
rect 45905 22650 45915 22730
rect 46225 22650 46235 22730
rect 46545 22650 46555 22730
rect 46865 22650 46875 22730
rect 47185 22650 47195 22730
rect 47505 22650 47515 22730
rect 47825 22650 47835 22730
rect 48145 22650 48155 22730
rect 48500 22670 48605 22840
rect 48640 22760 48650 22840
rect 48790 22760 48800 22840
rect 49350 22760 49360 22840
rect 49500 22760 49510 22840
rect 49650 22760 49660 22840
rect 48500 22660 48640 22670
rect 48710 22660 48790 22670
rect 49270 22660 49350 22670
rect 49420 22660 49500 22670
rect 49570 22660 49650 22670
rect 44065 22570 44145 22580
rect 44385 22570 44465 22580
rect 44705 22570 44785 22580
rect 45025 22570 45105 22580
rect 45345 22570 45425 22580
rect 45665 22570 45745 22580
rect 45985 22570 46065 22580
rect 46305 22570 46385 22580
rect 46625 22570 46705 22580
rect 46945 22570 47025 22580
rect 47265 22570 47345 22580
rect 47585 22570 47665 22580
rect 47905 22570 47985 22580
rect 48225 22570 48305 22580
rect 42950 22500 42980 22510
rect 43220 22500 43300 22510
rect 42980 22420 42990 22500
rect 43300 22420 43310 22500
rect 44145 22490 44155 22570
rect 44465 22490 44475 22570
rect 44785 22490 44795 22570
rect 45105 22490 45115 22570
rect 45425 22490 45435 22570
rect 45745 22490 45755 22570
rect 46065 22490 46075 22570
rect 46385 22490 46395 22570
rect 46705 22490 46715 22570
rect 47025 22490 47035 22570
rect 47345 22490 47355 22570
rect 47665 22490 47675 22570
rect 47985 22490 47995 22570
rect 48305 22490 48315 22570
rect 48500 22490 48605 22660
rect 48640 22580 48650 22660
rect 48790 22580 48800 22660
rect 49350 22580 49360 22660
rect 49500 22580 49510 22660
rect 49650 22580 49660 22660
rect 48500 22480 48640 22490
rect 48710 22480 48790 22490
rect 49270 22480 49350 22490
rect 49420 22480 49500 22490
rect 49570 22480 49650 22490
rect 43905 22410 43985 22420
rect 44225 22410 44305 22420
rect 44545 22410 44625 22420
rect 44865 22410 44945 22420
rect 45185 22410 45265 22420
rect 45505 22410 45585 22420
rect 45825 22410 45905 22420
rect 46145 22410 46225 22420
rect 46465 22410 46545 22420
rect 46785 22410 46865 22420
rect 47105 22410 47185 22420
rect 47425 22410 47505 22420
rect 47745 22410 47825 22420
rect 48065 22410 48145 22420
rect 43060 22340 43140 22350
rect 43380 22340 43460 22350
rect 43140 22260 43150 22340
rect 43460 22260 43470 22340
rect 43985 22330 43995 22410
rect 44305 22330 44315 22410
rect 44625 22330 44635 22410
rect 44945 22330 44955 22410
rect 45265 22330 45275 22410
rect 45585 22330 45595 22410
rect 45905 22330 45915 22410
rect 46225 22330 46235 22410
rect 46545 22330 46555 22410
rect 46865 22330 46875 22410
rect 47185 22330 47195 22410
rect 47505 22330 47515 22410
rect 47825 22330 47835 22410
rect 48145 22330 48155 22410
rect 48500 22310 48605 22480
rect 48640 22400 48650 22480
rect 48790 22400 48800 22480
rect 49350 22400 49360 22480
rect 49500 22400 49510 22480
rect 49650 22400 49660 22480
rect 48500 22300 48640 22310
rect 48710 22300 48790 22310
rect 49270 22300 49350 22310
rect 49420 22300 49500 22310
rect 49570 22300 49650 22310
rect 44065 22250 44145 22260
rect 44385 22250 44465 22260
rect 44705 22250 44785 22260
rect 45025 22250 45105 22260
rect 45345 22250 45425 22260
rect 45665 22250 45745 22260
rect 45985 22250 46065 22260
rect 46305 22250 46385 22260
rect 46625 22250 46705 22260
rect 46945 22250 47025 22260
rect 47265 22250 47345 22260
rect 47585 22250 47665 22260
rect 47905 22250 47985 22260
rect 48225 22250 48305 22260
rect 42950 22180 42980 22190
rect 43220 22180 43300 22190
rect 42980 22100 42990 22180
rect 43300 22100 43310 22180
rect 44145 22170 44155 22250
rect 44465 22170 44475 22250
rect 44785 22170 44795 22250
rect 45105 22170 45115 22250
rect 45425 22170 45435 22250
rect 45745 22170 45755 22250
rect 46065 22170 46075 22250
rect 46385 22170 46395 22250
rect 46705 22170 46715 22250
rect 47025 22170 47035 22250
rect 47345 22170 47355 22250
rect 47665 22170 47675 22250
rect 47985 22170 47995 22250
rect 48305 22170 48315 22250
rect 48500 22130 48605 22300
rect 48640 22220 48650 22300
rect 48790 22220 48800 22300
rect 49350 22220 49360 22300
rect 49500 22220 49510 22300
rect 49650 22220 49660 22300
rect 48500 22120 48640 22130
rect 48710 22120 48790 22130
rect 49270 22120 49350 22130
rect 49420 22120 49500 22130
rect 49570 22120 49650 22130
rect 43905 22090 43985 22100
rect 44225 22090 44305 22100
rect 44545 22090 44625 22100
rect 44865 22090 44945 22100
rect 45185 22090 45265 22100
rect 45505 22090 45585 22100
rect 45825 22090 45905 22100
rect 46145 22090 46225 22100
rect 46465 22090 46545 22100
rect 46785 22090 46865 22100
rect 47105 22090 47185 22100
rect 47425 22090 47505 22100
rect 47745 22090 47825 22100
rect 48065 22090 48145 22100
rect 43060 22020 43140 22030
rect 43380 22020 43460 22030
rect 43140 21940 43150 22020
rect 43460 21940 43470 22020
rect 43985 22010 43995 22090
rect 44305 22010 44315 22090
rect 44625 22010 44635 22090
rect 44945 22010 44955 22090
rect 45265 22010 45275 22090
rect 45585 22010 45595 22090
rect 45905 22010 45915 22090
rect 46225 22010 46235 22090
rect 46545 22010 46555 22090
rect 46865 22010 46875 22090
rect 47185 22010 47195 22090
rect 47505 22010 47515 22090
rect 47825 22010 47835 22090
rect 48145 22010 48155 22090
rect 48500 21950 48605 22120
rect 48640 22040 48650 22120
rect 48790 22040 48800 22120
rect 49350 22040 49360 22120
rect 49500 22040 49510 22120
rect 49650 22040 49660 22120
rect 48500 21940 48640 21950
rect 48710 21940 48790 21950
rect 49270 21940 49350 21950
rect 49420 21940 49500 21950
rect 49570 21940 49650 21950
rect 44065 21930 44145 21940
rect 44385 21930 44465 21940
rect 44705 21930 44785 21940
rect 45025 21930 45105 21940
rect 45345 21930 45425 21940
rect 45665 21930 45745 21940
rect 45985 21930 46065 21940
rect 46305 21930 46385 21940
rect 46625 21930 46705 21940
rect 46945 21930 47025 21940
rect 47265 21930 47345 21940
rect 47585 21930 47665 21940
rect 47905 21930 47985 21940
rect 48225 21930 48305 21940
rect 42950 21860 42980 21870
rect 43220 21860 43300 21870
rect 42980 21780 42990 21860
rect 43300 21780 43310 21860
rect 44145 21850 44155 21930
rect 44465 21850 44475 21930
rect 44785 21850 44795 21930
rect 45105 21850 45115 21930
rect 45425 21850 45435 21930
rect 45745 21850 45755 21930
rect 46065 21850 46075 21930
rect 46385 21850 46395 21930
rect 46705 21850 46715 21930
rect 47025 21850 47035 21930
rect 47345 21850 47355 21930
rect 47665 21850 47675 21930
rect 47985 21850 47995 21930
rect 48305 21850 48315 21930
rect 43905 21770 43985 21780
rect 44225 21770 44305 21780
rect 44545 21770 44625 21780
rect 44865 21770 44945 21780
rect 45185 21770 45265 21780
rect 45505 21770 45585 21780
rect 45825 21770 45905 21780
rect 46145 21770 46225 21780
rect 46465 21770 46545 21780
rect 46785 21770 46865 21780
rect 47105 21770 47185 21780
rect 47425 21770 47505 21780
rect 47745 21770 47825 21780
rect 48065 21770 48145 21780
rect 48500 21770 48605 21940
rect 48640 21860 48650 21940
rect 48790 21860 48800 21940
rect 49350 21860 49360 21940
rect 49500 21860 49510 21940
rect 49650 21860 49660 21940
rect 43060 21700 43140 21710
rect 43380 21700 43460 21710
rect 43140 21620 43150 21700
rect 43460 21620 43470 21700
rect 43985 21690 43995 21770
rect 44305 21690 44315 21770
rect 44625 21690 44635 21770
rect 44945 21690 44955 21770
rect 45265 21690 45275 21770
rect 45585 21690 45595 21770
rect 45905 21690 45915 21770
rect 46225 21690 46235 21770
rect 46545 21690 46555 21770
rect 46865 21690 46875 21770
rect 47185 21690 47195 21770
rect 47505 21690 47515 21770
rect 47825 21690 47835 21770
rect 48145 21690 48155 21770
rect 48500 21760 48640 21770
rect 48710 21760 48790 21770
rect 49270 21760 49350 21770
rect 49420 21760 49500 21770
rect 49570 21760 49650 21770
rect 44065 21610 44145 21620
rect 44385 21610 44465 21620
rect 44705 21610 44785 21620
rect 45025 21610 45105 21620
rect 45345 21610 45425 21620
rect 45665 21610 45745 21620
rect 45985 21610 46065 21620
rect 46305 21610 46385 21620
rect 46625 21610 46705 21620
rect 46945 21610 47025 21620
rect 47265 21610 47345 21620
rect 47585 21610 47665 21620
rect 47905 21610 47985 21620
rect 48225 21610 48305 21620
rect 42950 21540 42980 21550
rect 43220 21540 43300 21550
rect 42980 21460 42990 21540
rect 43300 21460 43310 21540
rect 44145 21530 44155 21610
rect 44465 21530 44475 21610
rect 44785 21530 44795 21610
rect 45105 21530 45115 21610
rect 45425 21530 45435 21610
rect 45745 21530 45755 21610
rect 46065 21530 46075 21610
rect 46385 21530 46395 21610
rect 46705 21530 46715 21610
rect 47025 21530 47035 21610
rect 47345 21530 47355 21610
rect 47665 21530 47675 21610
rect 47985 21530 47995 21610
rect 48305 21530 48315 21610
rect 48500 21590 48605 21760
rect 48640 21680 48650 21760
rect 48790 21680 48800 21760
rect 49350 21680 49360 21760
rect 49500 21680 49510 21760
rect 49650 21680 49660 21760
rect 48500 21580 48640 21590
rect 48710 21580 48790 21590
rect 49270 21580 49350 21590
rect 49420 21580 49500 21590
rect 49570 21580 49650 21590
rect 43905 21450 43985 21460
rect 44225 21450 44305 21460
rect 44545 21450 44625 21460
rect 44865 21450 44945 21460
rect 45185 21450 45265 21460
rect 45505 21450 45585 21460
rect 45825 21450 45905 21460
rect 46145 21450 46225 21460
rect 46465 21450 46545 21460
rect 46785 21450 46865 21460
rect 47105 21450 47185 21460
rect 47425 21450 47505 21460
rect 47745 21450 47825 21460
rect 48065 21450 48145 21460
rect 43060 21380 43140 21390
rect 43380 21380 43460 21390
rect 43140 21300 43150 21380
rect 43460 21300 43470 21380
rect 43985 21370 43995 21450
rect 44305 21370 44315 21450
rect 44625 21370 44635 21450
rect 44945 21370 44955 21450
rect 45265 21370 45275 21450
rect 45585 21370 45595 21450
rect 45905 21370 45915 21450
rect 46225 21370 46235 21450
rect 46545 21370 46555 21450
rect 46865 21370 46875 21450
rect 47185 21370 47195 21450
rect 47505 21370 47515 21450
rect 47825 21370 47835 21450
rect 48145 21370 48155 21450
rect 48500 21410 48605 21580
rect 48640 21500 48650 21580
rect 48790 21500 48800 21580
rect 49350 21500 49360 21580
rect 49500 21500 49510 21580
rect 49650 21500 49660 21580
rect 48500 21400 48640 21410
rect 48710 21400 48790 21410
rect 49270 21400 49350 21410
rect 49420 21400 49500 21410
rect 49570 21400 49650 21410
rect 44065 21290 44145 21300
rect 44385 21290 44465 21300
rect 44705 21290 44785 21300
rect 45025 21290 45105 21300
rect 45345 21290 45425 21300
rect 45665 21290 45745 21300
rect 45985 21290 46065 21300
rect 46305 21290 46385 21300
rect 46625 21290 46705 21300
rect 46945 21290 47025 21300
rect 47265 21290 47345 21300
rect 47585 21290 47665 21300
rect 47905 21290 47985 21300
rect 48225 21290 48305 21300
rect 42950 21220 42980 21230
rect 43220 21220 43300 21230
rect 42980 21140 42990 21220
rect 43300 21140 43310 21220
rect 44145 21210 44155 21290
rect 44465 21210 44475 21290
rect 44785 21210 44795 21290
rect 45105 21210 45115 21290
rect 45425 21210 45435 21290
rect 45745 21210 45755 21290
rect 46065 21210 46075 21290
rect 46385 21210 46395 21290
rect 46705 21210 46715 21290
rect 47025 21210 47035 21290
rect 47345 21210 47355 21290
rect 47665 21210 47675 21290
rect 47985 21210 47995 21290
rect 48305 21210 48315 21290
rect 48500 21230 48605 21400
rect 48640 21320 48650 21400
rect 48790 21320 48800 21400
rect 49350 21320 49360 21400
rect 49500 21320 49510 21400
rect 49650 21320 49660 21400
rect 48500 21220 48640 21230
rect 48710 21220 48790 21230
rect 49270 21220 49350 21230
rect 49420 21220 49500 21230
rect 49570 21220 49650 21230
rect 43905 21130 43985 21140
rect 44225 21130 44305 21140
rect 44545 21130 44625 21140
rect 44865 21130 44945 21140
rect 45185 21130 45265 21140
rect 45505 21130 45585 21140
rect 45825 21130 45905 21140
rect 46145 21130 46225 21140
rect 46465 21130 46545 21140
rect 46785 21130 46865 21140
rect 47105 21130 47185 21140
rect 47425 21130 47505 21140
rect 47745 21130 47825 21140
rect 48065 21130 48145 21140
rect 43060 21060 43140 21070
rect 43380 21060 43460 21070
rect 43140 20980 43150 21060
rect 43460 20980 43470 21060
rect 43985 21050 43995 21130
rect 44305 21050 44315 21130
rect 44625 21050 44635 21130
rect 44945 21050 44955 21130
rect 45265 21050 45275 21130
rect 45585 21050 45595 21130
rect 45905 21050 45915 21130
rect 46225 21050 46235 21130
rect 46545 21050 46555 21130
rect 46865 21050 46875 21130
rect 47185 21050 47195 21130
rect 47505 21050 47515 21130
rect 47825 21050 47835 21130
rect 48145 21050 48155 21130
rect 48500 21050 48605 21220
rect 48640 21140 48650 21220
rect 48790 21140 48800 21220
rect 49350 21140 49360 21220
rect 49500 21140 49510 21220
rect 49650 21140 49660 21220
rect 48500 21040 48640 21050
rect 48710 21040 48790 21050
rect 49270 21040 49350 21050
rect 49420 21040 49500 21050
rect 49570 21040 49650 21050
rect 44065 20970 44145 20980
rect 44385 20970 44465 20980
rect 44705 20970 44785 20980
rect 45025 20970 45105 20980
rect 45345 20970 45425 20980
rect 45665 20970 45745 20980
rect 45985 20970 46065 20980
rect 46305 20970 46385 20980
rect 46625 20970 46705 20980
rect 46945 20970 47025 20980
rect 47265 20970 47345 20980
rect 47585 20970 47665 20980
rect 47905 20970 47985 20980
rect 48225 20970 48305 20980
rect 42950 20900 42980 20910
rect 43220 20900 43300 20910
rect 42980 20820 42990 20900
rect 43300 20820 43310 20900
rect 44145 20890 44155 20970
rect 44465 20890 44475 20970
rect 44785 20890 44795 20970
rect 45105 20890 45115 20970
rect 45425 20890 45435 20970
rect 45745 20890 45755 20970
rect 46065 20890 46075 20970
rect 46385 20890 46395 20970
rect 46705 20890 46715 20970
rect 47025 20890 47035 20970
rect 47345 20890 47355 20970
rect 47665 20890 47675 20970
rect 47985 20890 47995 20970
rect 48305 20890 48315 20970
rect 48500 20870 48605 21040
rect 48640 20960 48650 21040
rect 48790 20960 48800 21040
rect 49350 20960 49360 21040
rect 49500 20960 49510 21040
rect 49650 20960 49660 21040
rect 48500 20860 48640 20870
rect 48710 20860 48790 20870
rect 49270 20860 49350 20870
rect 49420 20860 49500 20870
rect 49570 20860 49650 20870
rect 43905 20810 43985 20820
rect 44225 20810 44305 20820
rect 44545 20810 44625 20820
rect 44865 20810 44945 20820
rect 45185 20810 45265 20820
rect 45505 20810 45585 20820
rect 45825 20810 45905 20820
rect 46145 20810 46225 20820
rect 46465 20810 46545 20820
rect 46785 20810 46865 20820
rect 47105 20810 47185 20820
rect 47425 20810 47505 20820
rect 47745 20810 47825 20820
rect 48065 20810 48145 20820
rect 43060 20740 43140 20750
rect 43380 20740 43460 20750
rect 43140 20660 43150 20740
rect 43460 20660 43470 20740
rect 43985 20730 43995 20810
rect 44305 20730 44315 20810
rect 44625 20730 44635 20810
rect 44945 20730 44955 20810
rect 45265 20730 45275 20810
rect 45585 20730 45595 20810
rect 45905 20730 45915 20810
rect 46225 20730 46235 20810
rect 46545 20730 46555 20810
rect 46865 20730 46875 20810
rect 47185 20730 47195 20810
rect 47505 20730 47515 20810
rect 47825 20730 47835 20810
rect 48145 20730 48155 20810
rect 48500 20690 48605 20860
rect 48640 20780 48650 20860
rect 48790 20780 48800 20860
rect 49350 20780 49360 20860
rect 49500 20780 49510 20860
rect 49650 20780 49660 20860
rect 48500 20680 48640 20690
rect 48710 20680 48790 20690
rect 49270 20680 49350 20690
rect 49420 20680 49500 20690
rect 49570 20680 49650 20690
rect 44065 20650 44145 20660
rect 44385 20650 44465 20660
rect 44705 20650 44785 20660
rect 45025 20650 45105 20660
rect 45345 20650 45425 20660
rect 45665 20650 45745 20660
rect 45985 20650 46065 20660
rect 46305 20650 46385 20660
rect 46625 20650 46705 20660
rect 46945 20650 47025 20660
rect 47265 20650 47345 20660
rect 47585 20650 47665 20660
rect 47905 20650 47985 20660
rect 48225 20650 48305 20660
rect 42950 20580 42980 20590
rect 43220 20580 43300 20590
rect 42980 20500 42990 20580
rect 43300 20500 43310 20580
rect 44145 20570 44155 20650
rect 44465 20570 44475 20650
rect 44785 20570 44795 20650
rect 45105 20570 45115 20650
rect 45425 20570 45435 20650
rect 45745 20570 45755 20650
rect 46065 20570 46075 20650
rect 46385 20570 46395 20650
rect 46705 20570 46715 20650
rect 47025 20570 47035 20650
rect 47345 20570 47355 20650
rect 47665 20570 47675 20650
rect 47985 20570 47995 20650
rect 48305 20570 48315 20650
rect 48500 20510 48605 20680
rect 48640 20600 48650 20680
rect 48790 20600 48800 20680
rect 49350 20600 49360 20680
rect 49500 20600 49510 20680
rect 49650 20600 49660 20680
rect 48500 20500 48640 20510
rect 48710 20500 48790 20510
rect 49270 20500 49350 20510
rect 49420 20500 49500 20510
rect 49570 20500 49650 20510
rect 43905 20490 43985 20500
rect 44225 20490 44305 20500
rect 44545 20490 44625 20500
rect 44865 20490 44945 20500
rect 45185 20490 45265 20500
rect 45505 20490 45585 20500
rect 45825 20490 45905 20500
rect 46145 20490 46225 20500
rect 46465 20490 46545 20500
rect 46785 20490 46865 20500
rect 47105 20490 47185 20500
rect 47425 20490 47505 20500
rect 47745 20490 47825 20500
rect 48065 20490 48145 20500
rect 43060 20420 43140 20430
rect 43380 20420 43460 20430
rect 43140 20340 43150 20420
rect 43460 20340 43470 20420
rect 43985 20410 43995 20490
rect 44305 20410 44315 20490
rect 44625 20410 44635 20490
rect 44945 20410 44955 20490
rect 45265 20410 45275 20490
rect 45585 20410 45595 20490
rect 45905 20410 45915 20490
rect 46225 20410 46235 20490
rect 46545 20410 46555 20490
rect 46865 20410 46875 20490
rect 47185 20410 47195 20490
rect 47505 20410 47515 20490
rect 47825 20410 47835 20490
rect 48145 20410 48155 20490
rect 44065 20330 44145 20340
rect 44385 20330 44465 20340
rect 44705 20330 44785 20340
rect 45025 20330 45105 20340
rect 45345 20330 45425 20340
rect 45665 20330 45745 20340
rect 45985 20330 46065 20340
rect 46305 20330 46385 20340
rect 46625 20330 46705 20340
rect 46945 20330 47025 20340
rect 47265 20330 47345 20340
rect 47585 20330 47665 20340
rect 47905 20330 47985 20340
rect 48225 20330 48305 20340
rect 48500 20330 48605 20500
rect 48640 20420 48650 20500
rect 48790 20420 48800 20500
rect 49350 20420 49360 20500
rect 49500 20420 49510 20500
rect 49650 20420 49660 20500
rect 42950 20260 42980 20270
rect 43220 20260 43300 20270
rect 42980 20180 42990 20260
rect 43300 20180 43310 20260
rect 44145 20250 44155 20330
rect 44465 20250 44475 20330
rect 44785 20250 44795 20330
rect 45105 20250 45115 20330
rect 45425 20250 45435 20330
rect 45745 20250 45755 20330
rect 46065 20250 46075 20330
rect 46385 20250 46395 20330
rect 46705 20250 46715 20330
rect 47025 20250 47035 20330
rect 47345 20250 47355 20330
rect 47665 20250 47675 20330
rect 47985 20250 47995 20330
rect 48305 20250 48315 20330
rect 48500 20320 48640 20330
rect 48710 20320 48790 20330
rect 49270 20320 49350 20330
rect 49420 20320 49500 20330
rect 49570 20320 49650 20330
rect 43905 20170 43985 20180
rect 44225 20170 44305 20180
rect 44545 20170 44625 20180
rect 44865 20170 44945 20180
rect 45185 20170 45265 20180
rect 45505 20170 45585 20180
rect 45825 20170 45905 20180
rect 46145 20170 46225 20180
rect 46465 20170 46545 20180
rect 46785 20170 46865 20180
rect 47105 20170 47185 20180
rect 47425 20170 47505 20180
rect 47745 20170 47825 20180
rect 48065 20170 48145 20180
rect 43060 20100 43140 20110
rect 43380 20100 43460 20110
rect 43140 20020 43150 20100
rect 43460 20020 43470 20100
rect 43985 20090 43995 20170
rect 44305 20090 44315 20170
rect 44625 20090 44635 20170
rect 44945 20090 44955 20170
rect 45265 20090 45275 20170
rect 45585 20090 45595 20170
rect 45905 20090 45915 20170
rect 46225 20090 46235 20170
rect 46545 20090 46555 20170
rect 46865 20090 46875 20170
rect 47185 20090 47195 20170
rect 47505 20090 47515 20170
rect 47825 20090 47835 20170
rect 48145 20090 48155 20170
rect 48500 20150 48605 20320
rect 48640 20240 48650 20320
rect 48790 20240 48800 20320
rect 49350 20240 49360 20320
rect 49500 20240 49510 20320
rect 49650 20240 49660 20320
rect 48500 20140 48640 20150
rect 48710 20140 48790 20150
rect 49270 20140 49350 20150
rect 49420 20140 49500 20150
rect 49570 20140 49650 20150
rect 44065 20010 44145 20020
rect 44385 20010 44465 20020
rect 44705 20010 44785 20020
rect 45025 20010 45105 20020
rect 45345 20010 45425 20020
rect 45665 20010 45745 20020
rect 45985 20010 46065 20020
rect 46305 20010 46385 20020
rect 46625 20010 46705 20020
rect 46945 20010 47025 20020
rect 47265 20010 47345 20020
rect 47585 20010 47665 20020
rect 47905 20010 47985 20020
rect 48225 20010 48305 20020
rect 42950 19940 42980 19950
rect 43220 19940 43300 19950
rect 42980 19860 42990 19940
rect 43300 19860 43310 19940
rect 44145 19930 44155 20010
rect 44465 19930 44475 20010
rect 44785 19930 44795 20010
rect 45105 19930 45115 20010
rect 45425 19930 45435 20010
rect 45745 19930 45755 20010
rect 46065 19930 46075 20010
rect 46385 19930 46395 20010
rect 46705 19930 46715 20010
rect 47025 19930 47035 20010
rect 47345 19930 47355 20010
rect 47665 19930 47675 20010
rect 47985 19930 47995 20010
rect 48305 19930 48315 20010
rect 48500 19970 48605 20140
rect 48640 20060 48650 20140
rect 48790 20060 48800 20140
rect 49350 20060 49360 20140
rect 49500 20060 49510 20140
rect 49650 20060 49660 20140
rect 48500 19960 48640 19970
rect 48710 19960 48790 19970
rect 49270 19960 49350 19970
rect 49420 19960 49500 19970
rect 49570 19960 49650 19970
rect 43905 19850 43985 19860
rect 44225 19850 44305 19860
rect 44545 19850 44625 19860
rect 44865 19850 44945 19860
rect 45185 19850 45265 19860
rect 45505 19850 45585 19860
rect 45825 19850 45905 19860
rect 46145 19850 46225 19860
rect 46465 19850 46545 19860
rect 46785 19850 46865 19860
rect 47105 19850 47185 19860
rect 47425 19850 47505 19860
rect 47745 19850 47825 19860
rect 48065 19850 48145 19860
rect 43060 19780 43140 19790
rect 43380 19780 43460 19790
rect 43140 19700 43150 19780
rect 43460 19700 43470 19780
rect 43985 19770 43995 19850
rect 44305 19770 44315 19850
rect 44625 19770 44635 19850
rect 44945 19770 44955 19850
rect 45265 19770 45275 19850
rect 45585 19770 45595 19850
rect 45905 19770 45915 19850
rect 46225 19770 46235 19850
rect 46545 19770 46555 19850
rect 46865 19770 46875 19850
rect 47185 19770 47195 19850
rect 47505 19770 47515 19850
rect 47825 19770 47835 19850
rect 48145 19770 48155 19850
rect 48500 19790 48605 19960
rect 48640 19880 48650 19960
rect 48790 19880 48800 19960
rect 49350 19880 49360 19960
rect 49500 19880 49510 19960
rect 49650 19880 49660 19960
rect 49790 19800 49800 25800
rect 49910 25720 49990 25730
rect 50210 25720 50290 25730
rect 49990 25640 50000 25720
rect 50290 25640 50300 25720
rect 49910 25540 49990 25550
rect 50210 25540 50290 25550
rect 49990 25460 50000 25540
rect 50290 25460 50300 25540
rect 49910 25360 49990 25370
rect 50210 25360 50290 25370
rect 49990 25280 50000 25360
rect 50290 25280 50300 25360
rect 49910 25180 49990 25190
rect 50210 25180 50290 25190
rect 49990 25100 50000 25180
rect 50290 25100 50300 25180
rect 49910 25000 49990 25010
rect 50210 25000 50290 25010
rect 49990 24920 50000 25000
rect 50290 24920 50300 25000
rect 49910 24820 49990 24830
rect 50210 24820 50290 24830
rect 49990 24740 50000 24820
rect 50290 24740 50300 24820
rect 49910 24640 49990 24650
rect 50210 24640 50290 24650
rect 49990 24560 50000 24640
rect 50290 24560 50300 24640
rect 49910 24460 49990 24470
rect 50210 24460 50290 24470
rect 49990 24380 50000 24460
rect 50290 24380 50300 24460
rect 49910 24280 49990 24290
rect 50210 24280 50290 24290
rect 49990 24200 50000 24280
rect 50290 24200 50300 24280
rect 49910 24100 49990 24110
rect 50210 24100 50290 24110
rect 49990 24020 50000 24100
rect 50290 24020 50300 24100
rect 49910 23920 49990 23930
rect 50210 23920 50290 23930
rect 49990 23840 50000 23920
rect 50290 23840 50300 23920
rect 49910 23740 49990 23750
rect 50210 23740 50290 23750
rect 49990 23660 50000 23740
rect 50290 23660 50300 23740
rect 49910 23560 49990 23570
rect 50210 23560 50290 23570
rect 49990 23480 50000 23560
rect 50290 23480 50300 23560
rect 49910 23380 49990 23390
rect 50210 23380 50290 23390
rect 49990 23300 50000 23380
rect 50290 23300 50300 23380
rect 49910 23200 49990 23210
rect 50210 23200 50290 23210
rect 49990 23120 50000 23200
rect 50290 23120 50300 23200
rect 49910 23020 49990 23030
rect 50210 23020 50290 23030
rect 49990 22940 50000 23020
rect 50290 22940 50300 23020
rect 49910 22840 49990 22850
rect 50210 22840 50290 22850
rect 49990 22760 50000 22840
rect 50290 22760 50300 22840
rect 49910 22660 49990 22670
rect 50210 22660 50290 22670
rect 49990 22580 50000 22660
rect 50290 22580 50300 22660
rect 49910 22480 49990 22490
rect 50210 22480 50290 22490
rect 49990 22400 50000 22480
rect 50290 22400 50300 22480
rect 49910 22300 49990 22310
rect 50210 22300 50290 22310
rect 49990 22220 50000 22300
rect 50290 22220 50300 22300
rect 49910 22120 49990 22130
rect 50210 22120 50290 22130
rect 49990 22040 50000 22120
rect 50290 22040 50300 22120
rect 49910 21940 49990 21950
rect 50210 21940 50290 21950
rect 49990 21860 50000 21940
rect 50290 21860 50300 21940
rect 49910 21760 49990 21770
rect 50210 21760 50290 21770
rect 49990 21680 50000 21760
rect 50290 21680 50300 21760
rect 49910 21580 49990 21590
rect 50210 21580 50290 21590
rect 49990 21500 50000 21580
rect 50290 21500 50300 21580
rect 49910 21400 49990 21410
rect 50210 21400 50290 21410
rect 49990 21320 50000 21400
rect 50290 21320 50300 21400
rect 49910 21220 49990 21230
rect 50210 21220 50290 21230
rect 49990 21140 50000 21220
rect 50290 21140 50300 21220
rect 49910 21040 49990 21050
rect 50210 21040 50290 21050
rect 49990 20960 50000 21040
rect 50290 20960 50300 21040
rect 49910 20860 49990 20870
rect 50210 20860 50290 20870
rect 49990 20780 50000 20860
rect 50290 20780 50300 20860
rect 49910 20680 49990 20690
rect 50210 20680 50290 20690
rect 49990 20600 50000 20680
rect 50290 20600 50300 20680
rect 49910 20500 49990 20510
rect 50210 20500 50290 20510
rect 49990 20420 50000 20500
rect 50290 20420 50300 20500
rect 49910 20320 49990 20330
rect 50210 20320 50290 20330
rect 49990 20240 50000 20320
rect 50290 20240 50300 20320
rect 49910 20140 49990 20150
rect 50210 20140 50290 20150
rect 49990 20060 50000 20140
rect 50290 20060 50300 20140
rect 49910 19960 49990 19970
rect 50210 19960 50290 19970
rect 49990 19880 50000 19960
rect 50290 19880 50300 19960
rect 50470 19800 50480 25800
rect 50530 25720 50610 25730
rect 50680 25720 50760 25730
rect 50830 25720 50910 25730
rect 50610 25640 50620 25720
rect 50760 25640 50770 25720
rect 50910 25640 50920 25720
rect 50530 25540 50610 25550
rect 50680 25540 50760 25550
rect 50830 25540 50910 25550
rect 50610 25460 50620 25540
rect 50760 25460 50770 25540
rect 50910 25460 50920 25540
rect 50530 25360 50610 25370
rect 50680 25360 50760 25370
rect 50830 25360 50910 25370
rect 50610 25280 50620 25360
rect 50760 25280 50770 25360
rect 50910 25280 50920 25360
rect 50530 25180 50610 25190
rect 50680 25180 50760 25190
rect 50830 25180 50910 25190
rect 50610 25100 50620 25180
rect 50760 25100 50770 25180
rect 50910 25100 50920 25180
rect 50530 25000 50610 25010
rect 50680 25000 50760 25010
rect 50830 25000 50910 25010
rect 50610 24920 50620 25000
rect 50760 24920 50770 25000
rect 50910 24920 50920 25000
rect 50530 24820 50610 24830
rect 50680 24820 50760 24830
rect 50830 24820 50910 24830
rect 50610 24740 50620 24820
rect 50760 24740 50770 24820
rect 50910 24740 50920 24820
rect 50530 24640 50610 24650
rect 50680 24640 50760 24650
rect 50830 24640 50910 24650
rect 50610 24560 50620 24640
rect 50760 24560 50770 24640
rect 50910 24560 50920 24640
rect 50530 24460 50610 24470
rect 50680 24460 50760 24470
rect 50830 24460 50910 24470
rect 50610 24380 50620 24460
rect 50760 24380 50770 24460
rect 50910 24380 50920 24460
rect 50530 24280 50610 24290
rect 50680 24280 50760 24290
rect 50830 24280 50910 24290
rect 50610 24200 50620 24280
rect 50760 24200 50770 24280
rect 50910 24200 50920 24280
rect 50530 24100 50610 24110
rect 50680 24100 50760 24110
rect 50830 24100 50910 24110
rect 50610 24020 50620 24100
rect 50760 24020 50770 24100
rect 50910 24020 50920 24100
rect 50530 23920 50610 23930
rect 50680 23920 50760 23930
rect 50830 23920 50910 23930
rect 50610 23840 50620 23920
rect 50760 23840 50770 23920
rect 50910 23840 50920 23920
rect 50530 23740 50610 23750
rect 50680 23740 50760 23750
rect 50830 23740 50910 23750
rect 50610 23660 50620 23740
rect 50760 23660 50770 23740
rect 50910 23660 50920 23740
rect 50530 23560 50610 23570
rect 50680 23560 50760 23570
rect 50830 23560 50910 23570
rect 50610 23480 50620 23560
rect 50760 23480 50770 23560
rect 50910 23480 50920 23560
rect 50530 23380 50610 23390
rect 50680 23380 50760 23390
rect 50830 23380 50910 23390
rect 50610 23300 50620 23380
rect 50760 23300 50770 23380
rect 50910 23300 50920 23380
rect 50530 23200 50610 23210
rect 50680 23200 50760 23210
rect 50830 23200 50910 23210
rect 50610 23120 50620 23200
rect 50760 23120 50770 23200
rect 50910 23120 50920 23200
rect 50530 23020 50610 23030
rect 50680 23020 50760 23030
rect 50830 23020 50910 23030
rect 50610 22940 50620 23020
rect 50760 22940 50770 23020
rect 50910 22940 50920 23020
rect 50530 22840 50610 22850
rect 50680 22840 50760 22850
rect 50830 22840 50910 22850
rect 50610 22760 50620 22840
rect 50760 22760 50770 22840
rect 50910 22760 50920 22840
rect 50530 22660 50610 22670
rect 50680 22660 50760 22670
rect 50830 22660 50910 22670
rect 50610 22580 50620 22660
rect 50760 22580 50770 22660
rect 50910 22580 50920 22660
rect 50530 22480 50610 22490
rect 50680 22480 50760 22490
rect 50830 22480 50910 22490
rect 50610 22400 50620 22480
rect 50760 22400 50770 22480
rect 50910 22400 50920 22480
rect 50530 22300 50610 22310
rect 50680 22300 50760 22310
rect 50830 22300 50910 22310
rect 50610 22220 50620 22300
rect 50760 22220 50770 22300
rect 50910 22220 50920 22300
rect 50530 22120 50610 22130
rect 50680 22120 50760 22130
rect 50830 22120 50910 22130
rect 50610 22040 50620 22120
rect 50760 22040 50770 22120
rect 50910 22040 50920 22120
rect 50530 21940 50610 21950
rect 50680 21940 50760 21950
rect 50830 21940 50910 21950
rect 50610 21860 50620 21940
rect 50760 21860 50770 21940
rect 50910 21860 50920 21940
rect 50530 21760 50610 21770
rect 50680 21760 50760 21770
rect 50830 21760 50910 21770
rect 50610 21680 50620 21760
rect 50760 21680 50770 21760
rect 50910 21680 50920 21760
rect 50530 21580 50610 21590
rect 50680 21580 50760 21590
rect 50830 21580 50910 21590
rect 50610 21500 50620 21580
rect 50760 21500 50770 21580
rect 50910 21500 50920 21580
rect 50530 21400 50610 21410
rect 50680 21400 50760 21410
rect 50830 21400 50910 21410
rect 50610 21320 50620 21400
rect 50760 21320 50770 21400
rect 50910 21320 50920 21400
rect 50530 21220 50610 21230
rect 50680 21220 50760 21230
rect 50830 21220 50910 21230
rect 50610 21140 50620 21220
rect 50760 21140 50770 21220
rect 50910 21140 50920 21220
rect 50530 21040 50610 21050
rect 50680 21040 50760 21050
rect 50830 21040 50910 21050
rect 50610 20960 50620 21040
rect 50760 20960 50770 21040
rect 50910 20960 50920 21040
rect 50530 20860 50610 20870
rect 50680 20860 50760 20870
rect 50830 20860 50910 20870
rect 50610 20780 50620 20860
rect 50760 20780 50770 20860
rect 50910 20780 50920 20860
rect 50530 20680 50610 20690
rect 50680 20680 50760 20690
rect 50830 20680 50910 20690
rect 50610 20600 50620 20680
rect 50760 20600 50770 20680
rect 50910 20600 50920 20680
rect 50530 20500 50610 20510
rect 50680 20500 50760 20510
rect 50830 20500 50910 20510
rect 50610 20420 50620 20500
rect 50760 20420 50770 20500
rect 50910 20420 50920 20500
rect 50530 20320 50610 20330
rect 50680 20320 50760 20330
rect 50830 20320 50910 20330
rect 50610 20240 50620 20320
rect 50760 20240 50770 20320
rect 50910 20240 50920 20320
rect 50530 20140 50610 20150
rect 50680 20140 50760 20150
rect 50830 20140 50910 20150
rect 50610 20060 50620 20140
rect 50760 20060 50770 20140
rect 50910 20060 50920 20140
rect 50530 19960 50610 19970
rect 50680 19960 50760 19970
rect 50830 19960 50910 19970
rect 50610 19880 50620 19960
rect 50760 19880 50770 19960
rect 50910 19880 50920 19960
rect 51050 19800 51060 25800
rect 51170 25720 51250 25730
rect 51470 25720 51550 25730
rect 51250 25640 51260 25720
rect 51550 25640 51560 25720
rect 51170 25540 51250 25550
rect 51470 25540 51550 25550
rect 51250 25460 51260 25540
rect 51550 25460 51560 25540
rect 51170 25360 51250 25370
rect 51470 25360 51550 25370
rect 51250 25280 51260 25360
rect 51550 25280 51560 25360
rect 51170 25180 51250 25190
rect 51470 25180 51550 25190
rect 51250 25100 51260 25180
rect 51550 25100 51560 25180
rect 51170 25000 51250 25010
rect 51470 25000 51550 25010
rect 51250 24920 51260 25000
rect 51550 24920 51560 25000
rect 51170 24820 51250 24830
rect 51470 24820 51550 24830
rect 51250 24740 51260 24820
rect 51550 24740 51560 24820
rect 51170 24640 51250 24650
rect 51470 24640 51550 24650
rect 51250 24560 51260 24640
rect 51550 24560 51560 24640
rect 51170 24460 51250 24470
rect 51470 24460 51550 24470
rect 51250 24380 51260 24460
rect 51550 24380 51560 24460
rect 51170 24280 51250 24290
rect 51470 24280 51550 24290
rect 51250 24200 51260 24280
rect 51550 24200 51560 24280
rect 51170 24100 51250 24110
rect 51470 24100 51550 24110
rect 51250 24020 51260 24100
rect 51550 24020 51560 24100
rect 51170 23920 51250 23930
rect 51470 23920 51550 23930
rect 51250 23840 51260 23920
rect 51550 23840 51560 23920
rect 51170 23740 51250 23750
rect 51470 23740 51550 23750
rect 51250 23660 51260 23740
rect 51550 23660 51560 23740
rect 51170 23560 51250 23570
rect 51470 23560 51550 23570
rect 51250 23480 51260 23560
rect 51550 23480 51560 23560
rect 51170 23380 51250 23390
rect 51470 23380 51550 23390
rect 51250 23300 51260 23380
rect 51550 23300 51560 23380
rect 51170 23200 51250 23210
rect 51470 23200 51550 23210
rect 51250 23120 51260 23200
rect 51550 23120 51560 23200
rect 51170 23020 51250 23030
rect 51470 23020 51550 23030
rect 51250 22940 51260 23020
rect 51550 22940 51560 23020
rect 51170 22840 51250 22850
rect 51470 22840 51550 22850
rect 51250 22760 51260 22840
rect 51550 22760 51560 22840
rect 51170 22660 51250 22670
rect 51470 22660 51550 22670
rect 51250 22580 51260 22660
rect 51550 22580 51560 22660
rect 51170 22480 51250 22490
rect 51470 22480 51550 22490
rect 51250 22400 51260 22480
rect 51550 22400 51560 22480
rect 51170 22300 51250 22310
rect 51470 22300 51550 22310
rect 51250 22220 51260 22300
rect 51550 22220 51560 22300
rect 51170 22120 51250 22130
rect 51470 22120 51550 22130
rect 51250 22040 51260 22120
rect 51550 22040 51560 22120
rect 51170 21940 51250 21950
rect 51470 21940 51550 21950
rect 51250 21860 51260 21940
rect 51550 21860 51560 21940
rect 51170 21760 51250 21770
rect 51470 21760 51550 21770
rect 51250 21680 51260 21760
rect 51550 21680 51560 21760
rect 51170 21580 51250 21590
rect 51470 21580 51550 21590
rect 51250 21500 51260 21580
rect 51550 21500 51560 21580
rect 51170 21400 51250 21410
rect 51470 21400 51550 21410
rect 51250 21320 51260 21400
rect 51550 21320 51560 21400
rect 51170 21220 51250 21230
rect 51470 21220 51550 21230
rect 51250 21140 51260 21220
rect 51550 21140 51560 21220
rect 51170 21040 51250 21050
rect 51470 21040 51550 21050
rect 51250 20960 51260 21040
rect 51550 20960 51560 21040
rect 51170 20860 51250 20870
rect 51470 20860 51550 20870
rect 51250 20780 51260 20860
rect 51550 20780 51560 20860
rect 51170 20680 51250 20690
rect 51470 20680 51550 20690
rect 51250 20600 51260 20680
rect 51550 20600 51560 20680
rect 51170 20500 51250 20510
rect 51470 20500 51550 20510
rect 51250 20420 51260 20500
rect 51550 20420 51560 20500
rect 51170 20320 51250 20330
rect 51470 20320 51550 20330
rect 51250 20240 51260 20320
rect 51550 20240 51560 20320
rect 51170 20140 51250 20150
rect 51470 20140 51550 20150
rect 51250 20060 51260 20140
rect 51550 20060 51560 20140
rect 51170 19960 51250 19970
rect 51470 19960 51550 19970
rect 51250 19880 51260 19960
rect 51550 19880 51560 19960
rect 51730 19800 51740 25800
rect 51790 25720 51870 25730
rect 51940 25720 52020 25730
rect 52090 25720 52170 25730
rect 51870 25640 51880 25720
rect 52020 25640 52030 25720
rect 52170 25640 52180 25720
rect 51790 25540 51870 25550
rect 51940 25540 52020 25550
rect 52090 25540 52170 25550
rect 51870 25460 51880 25540
rect 52020 25460 52030 25540
rect 52170 25460 52180 25540
rect 51790 25360 51870 25370
rect 51940 25360 52020 25370
rect 52090 25360 52170 25370
rect 51870 25280 51880 25360
rect 52020 25280 52030 25360
rect 52170 25280 52180 25360
rect 51790 25180 51870 25190
rect 51940 25180 52020 25190
rect 52090 25180 52170 25190
rect 51870 25100 51880 25180
rect 52020 25100 52030 25180
rect 52170 25100 52180 25180
rect 51790 25000 51870 25010
rect 51940 25000 52020 25010
rect 52090 25000 52170 25010
rect 51870 24920 51880 25000
rect 52020 24920 52030 25000
rect 52170 24920 52180 25000
rect 51790 24820 51870 24830
rect 51940 24820 52020 24830
rect 52090 24820 52170 24830
rect 51870 24740 51880 24820
rect 52020 24740 52030 24820
rect 52170 24740 52180 24820
rect 51790 24640 51870 24650
rect 51940 24640 52020 24650
rect 52090 24640 52170 24650
rect 51870 24560 51880 24640
rect 52020 24560 52030 24640
rect 52170 24560 52180 24640
rect 51790 24460 51870 24470
rect 51940 24460 52020 24470
rect 52090 24460 52170 24470
rect 51870 24380 51880 24460
rect 52020 24380 52030 24460
rect 52170 24380 52180 24460
rect 51790 24280 51870 24290
rect 51940 24280 52020 24290
rect 52090 24280 52170 24290
rect 51870 24200 51880 24280
rect 52020 24200 52030 24280
rect 52170 24200 52180 24280
rect 51790 24100 51870 24110
rect 51940 24100 52020 24110
rect 52090 24100 52170 24110
rect 51870 24020 51880 24100
rect 52020 24020 52030 24100
rect 52170 24020 52180 24100
rect 51790 23920 51870 23930
rect 51940 23920 52020 23930
rect 52090 23920 52170 23930
rect 51870 23840 51880 23920
rect 52020 23840 52030 23920
rect 52170 23840 52180 23920
rect 51790 23740 51870 23750
rect 51940 23740 52020 23750
rect 52090 23740 52170 23750
rect 51870 23660 51880 23740
rect 52020 23660 52030 23740
rect 52170 23660 52180 23740
rect 51790 23560 51870 23570
rect 51940 23560 52020 23570
rect 52090 23560 52170 23570
rect 51870 23480 51880 23560
rect 52020 23480 52030 23560
rect 52170 23480 52180 23560
rect 51790 23380 51870 23390
rect 51940 23380 52020 23390
rect 52090 23380 52170 23390
rect 51870 23300 51880 23380
rect 52020 23300 52030 23380
rect 52170 23300 52180 23380
rect 51790 23200 51870 23210
rect 51940 23200 52020 23210
rect 52090 23200 52170 23210
rect 51870 23120 51880 23200
rect 52020 23120 52030 23200
rect 52170 23120 52180 23200
rect 51790 23020 51870 23030
rect 51940 23020 52020 23030
rect 52090 23020 52170 23030
rect 51870 22940 51880 23020
rect 52020 22940 52030 23020
rect 52170 22940 52180 23020
rect 51790 22840 51870 22850
rect 51940 22840 52020 22850
rect 52090 22840 52170 22850
rect 51870 22760 51880 22840
rect 52020 22760 52030 22840
rect 52170 22760 52180 22840
rect 51790 22660 51870 22670
rect 51940 22660 52020 22670
rect 52090 22660 52170 22670
rect 51870 22580 51880 22660
rect 52020 22580 52030 22660
rect 52170 22580 52180 22660
rect 51790 22480 51870 22490
rect 51940 22480 52020 22490
rect 52090 22480 52170 22490
rect 51870 22400 51880 22480
rect 52020 22400 52030 22480
rect 52170 22400 52180 22480
rect 51790 22300 51870 22310
rect 51940 22300 52020 22310
rect 52090 22300 52170 22310
rect 51870 22220 51880 22300
rect 52020 22220 52030 22300
rect 52170 22220 52180 22300
rect 51790 22120 51870 22130
rect 51940 22120 52020 22130
rect 52090 22120 52170 22130
rect 51870 22040 51880 22120
rect 52020 22040 52030 22120
rect 52170 22040 52180 22120
rect 51790 21940 51870 21950
rect 51940 21940 52020 21950
rect 52090 21940 52170 21950
rect 51870 21860 51880 21940
rect 52020 21860 52030 21940
rect 52170 21860 52180 21940
rect 51790 21760 51870 21770
rect 51940 21760 52020 21770
rect 52090 21760 52170 21770
rect 51870 21680 51880 21760
rect 52020 21680 52030 21760
rect 52170 21680 52180 21760
rect 51790 21580 51870 21590
rect 51940 21580 52020 21590
rect 52090 21580 52170 21590
rect 51870 21500 51880 21580
rect 52020 21500 52030 21580
rect 52170 21500 52180 21580
rect 51790 21400 51870 21410
rect 51940 21400 52020 21410
rect 52090 21400 52170 21410
rect 51870 21320 51880 21400
rect 52020 21320 52030 21400
rect 52170 21320 52180 21400
rect 51790 21220 51870 21230
rect 51940 21220 52020 21230
rect 52090 21220 52170 21230
rect 51870 21140 51880 21220
rect 52020 21140 52030 21220
rect 52170 21140 52180 21220
rect 51790 21040 51870 21050
rect 51940 21040 52020 21050
rect 52090 21040 52170 21050
rect 51870 20960 51880 21040
rect 52020 20960 52030 21040
rect 52170 20960 52180 21040
rect 51790 20860 51870 20870
rect 51940 20860 52020 20870
rect 52090 20860 52170 20870
rect 51870 20780 51880 20860
rect 52020 20780 52030 20860
rect 52170 20780 52180 20860
rect 51790 20680 51870 20690
rect 51940 20680 52020 20690
rect 52090 20680 52170 20690
rect 51870 20600 51880 20680
rect 52020 20600 52030 20680
rect 52170 20600 52180 20680
rect 51790 20500 51870 20510
rect 51940 20500 52020 20510
rect 52090 20500 52170 20510
rect 51870 20420 51880 20500
rect 52020 20420 52030 20500
rect 52170 20420 52180 20500
rect 51790 20320 51870 20330
rect 51940 20320 52020 20330
rect 52090 20320 52170 20330
rect 51870 20240 51880 20320
rect 52020 20240 52030 20320
rect 52170 20240 52180 20320
rect 51790 20140 51870 20150
rect 51940 20140 52020 20150
rect 52090 20140 52170 20150
rect 51870 20060 51880 20140
rect 52020 20060 52030 20140
rect 52170 20060 52180 20140
rect 51790 19960 51870 19970
rect 51940 19960 52020 19970
rect 52090 19960 52170 19970
rect 51870 19880 51880 19960
rect 52020 19880 52030 19960
rect 52170 19880 52180 19960
rect 52310 19800 52320 25800
rect 52430 25720 52510 25730
rect 52730 25720 52810 25730
rect 52510 25640 52520 25720
rect 52810 25640 52820 25720
rect 52430 25540 52510 25550
rect 52730 25540 52810 25550
rect 52510 25460 52520 25540
rect 52810 25460 52820 25540
rect 52430 25360 52510 25370
rect 52730 25360 52810 25370
rect 52510 25280 52520 25360
rect 52810 25280 52820 25360
rect 52430 25180 52510 25190
rect 52730 25180 52810 25190
rect 52510 25100 52520 25180
rect 52810 25100 52820 25180
rect 52430 25000 52510 25010
rect 52730 25000 52810 25010
rect 52510 24920 52520 25000
rect 52810 24920 52820 25000
rect 52430 24820 52510 24830
rect 52730 24820 52810 24830
rect 52510 24740 52520 24820
rect 52810 24740 52820 24820
rect 52430 24640 52510 24650
rect 52730 24640 52810 24650
rect 52510 24560 52520 24640
rect 52810 24560 52820 24640
rect 52430 24460 52510 24470
rect 52730 24460 52810 24470
rect 52510 24380 52520 24460
rect 52810 24380 52820 24460
rect 52430 24280 52510 24290
rect 52730 24280 52810 24290
rect 52510 24200 52520 24280
rect 52810 24200 52820 24280
rect 52430 24100 52510 24110
rect 52730 24100 52810 24110
rect 52510 24020 52520 24100
rect 52810 24020 52820 24100
rect 52430 23920 52510 23930
rect 52730 23920 52810 23930
rect 52510 23840 52520 23920
rect 52810 23840 52820 23920
rect 52430 23740 52510 23750
rect 52730 23740 52810 23750
rect 52510 23660 52520 23740
rect 52810 23660 52820 23740
rect 52430 23560 52510 23570
rect 52730 23560 52810 23570
rect 52510 23480 52520 23560
rect 52810 23480 52820 23560
rect 52430 23380 52510 23390
rect 52730 23380 52810 23390
rect 52510 23300 52520 23380
rect 52810 23300 52820 23380
rect 52430 23200 52510 23210
rect 52730 23200 52810 23210
rect 52510 23120 52520 23200
rect 52810 23120 52820 23200
rect 52430 23020 52510 23030
rect 52730 23020 52810 23030
rect 52510 22940 52520 23020
rect 52810 22940 52820 23020
rect 52430 22840 52510 22850
rect 52730 22840 52810 22850
rect 52510 22760 52520 22840
rect 52810 22760 52820 22840
rect 52430 22660 52510 22670
rect 52730 22660 52810 22670
rect 52510 22580 52520 22660
rect 52810 22580 52820 22660
rect 52430 22480 52510 22490
rect 52730 22480 52810 22490
rect 52510 22400 52520 22480
rect 52810 22400 52820 22480
rect 52430 22300 52510 22310
rect 52730 22300 52810 22310
rect 52510 22220 52520 22300
rect 52810 22220 52820 22300
rect 52430 22120 52510 22130
rect 52730 22120 52810 22130
rect 52510 22040 52520 22120
rect 52810 22040 52820 22120
rect 52430 21940 52510 21950
rect 52730 21940 52810 21950
rect 52510 21860 52520 21940
rect 52810 21860 52820 21940
rect 52430 21760 52510 21770
rect 52730 21760 52810 21770
rect 52510 21680 52520 21760
rect 52810 21680 52820 21760
rect 52430 21580 52510 21590
rect 52730 21580 52810 21590
rect 52510 21500 52520 21580
rect 52810 21500 52820 21580
rect 52430 21400 52510 21410
rect 52730 21400 52810 21410
rect 52510 21320 52520 21400
rect 52810 21320 52820 21400
rect 52430 21220 52510 21230
rect 52730 21220 52810 21230
rect 52510 21140 52520 21220
rect 52810 21140 52820 21220
rect 52430 21040 52510 21050
rect 52730 21040 52810 21050
rect 52510 20960 52520 21040
rect 52810 20960 52820 21040
rect 52430 20860 52510 20870
rect 52730 20860 52810 20870
rect 52510 20780 52520 20860
rect 52810 20780 52820 20860
rect 52430 20680 52510 20690
rect 52730 20680 52810 20690
rect 52510 20600 52520 20680
rect 52810 20600 52820 20680
rect 52430 20500 52510 20510
rect 52730 20500 52810 20510
rect 52510 20420 52520 20500
rect 52810 20420 52820 20500
rect 52430 20320 52510 20330
rect 52730 20320 52810 20330
rect 52510 20240 52520 20320
rect 52810 20240 52820 20320
rect 52430 20140 52510 20150
rect 52730 20140 52810 20150
rect 52510 20060 52520 20140
rect 52810 20060 52820 20140
rect 52430 19960 52510 19970
rect 52730 19960 52810 19970
rect 52510 19880 52520 19960
rect 52810 19880 52820 19960
rect 52990 19800 53000 25800
rect 53050 25720 53130 25730
rect 53200 25720 53280 25730
rect 53350 25720 53430 25730
rect 53130 25640 53140 25720
rect 53280 25640 53290 25720
rect 53430 25640 53440 25720
rect 53050 25540 53130 25550
rect 53200 25540 53280 25550
rect 53350 25540 53430 25550
rect 53130 25460 53140 25540
rect 53280 25460 53290 25540
rect 53430 25460 53440 25540
rect 53050 25360 53130 25370
rect 53200 25360 53280 25370
rect 53350 25360 53430 25370
rect 53130 25280 53140 25360
rect 53280 25280 53290 25360
rect 53430 25280 53440 25360
rect 53050 25180 53130 25190
rect 53200 25180 53280 25190
rect 53350 25180 53430 25190
rect 53130 25100 53140 25180
rect 53280 25100 53290 25180
rect 53430 25100 53440 25180
rect 53050 25000 53130 25010
rect 53200 25000 53280 25010
rect 53350 25000 53430 25010
rect 53130 24920 53140 25000
rect 53280 24920 53290 25000
rect 53430 24920 53440 25000
rect 53050 24820 53130 24830
rect 53200 24820 53280 24830
rect 53350 24820 53430 24830
rect 53130 24740 53140 24820
rect 53280 24740 53290 24820
rect 53430 24740 53440 24820
rect 53050 24640 53130 24650
rect 53200 24640 53280 24650
rect 53350 24640 53430 24650
rect 53130 24560 53140 24640
rect 53280 24560 53290 24640
rect 53430 24560 53440 24640
rect 53050 24460 53130 24470
rect 53200 24460 53280 24470
rect 53350 24460 53430 24470
rect 53130 24380 53140 24460
rect 53280 24380 53290 24460
rect 53430 24380 53440 24460
rect 53050 24280 53130 24290
rect 53200 24280 53280 24290
rect 53350 24280 53430 24290
rect 53130 24200 53140 24280
rect 53280 24200 53290 24280
rect 53430 24200 53440 24280
rect 53050 24100 53130 24110
rect 53200 24100 53280 24110
rect 53350 24100 53430 24110
rect 53130 24020 53140 24100
rect 53280 24020 53290 24100
rect 53430 24020 53440 24100
rect 53050 23920 53130 23930
rect 53200 23920 53280 23930
rect 53350 23920 53430 23930
rect 53130 23840 53140 23920
rect 53280 23840 53290 23920
rect 53430 23840 53440 23920
rect 53050 23740 53130 23750
rect 53200 23740 53280 23750
rect 53350 23740 53430 23750
rect 53130 23660 53140 23740
rect 53280 23660 53290 23740
rect 53430 23660 53440 23740
rect 53050 23560 53130 23570
rect 53200 23560 53280 23570
rect 53350 23560 53430 23570
rect 53130 23480 53140 23560
rect 53280 23480 53290 23560
rect 53430 23480 53440 23560
rect 53050 23380 53130 23390
rect 53200 23380 53280 23390
rect 53350 23380 53430 23390
rect 53130 23300 53140 23380
rect 53280 23300 53290 23380
rect 53430 23300 53440 23380
rect 53050 23200 53130 23210
rect 53200 23200 53280 23210
rect 53350 23200 53430 23210
rect 53130 23120 53140 23200
rect 53280 23120 53290 23200
rect 53430 23120 53440 23200
rect 53050 23020 53130 23030
rect 53200 23020 53280 23030
rect 53350 23020 53430 23030
rect 53130 22940 53140 23020
rect 53280 22940 53290 23020
rect 53430 22940 53440 23020
rect 53050 22840 53130 22850
rect 53200 22840 53280 22850
rect 53350 22840 53430 22850
rect 53130 22760 53140 22840
rect 53280 22760 53290 22840
rect 53430 22760 53440 22840
rect 53050 22660 53130 22670
rect 53200 22660 53280 22670
rect 53350 22660 53430 22670
rect 53130 22580 53140 22660
rect 53280 22580 53290 22660
rect 53430 22580 53440 22660
rect 53050 22480 53130 22490
rect 53200 22480 53280 22490
rect 53350 22480 53430 22490
rect 53130 22400 53140 22480
rect 53280 22400 53290 22480
rect 53430 22400 53440 22480
rect 53050 22300 53130 22310
rect 53200 22300 53280 22310
rect 53350 22300 53430 22310
rect 53130 22220 53140 22300
rect 53280 22220 53290 22300
rect 53430 22220 53440 22300
rect 53050 22120 53130 22130
rect 53200 22120 53280 22130
rect 53350 22120 53430 22130
rect 53130 22040 53140 22120
rect 53280 22040 53290 22120
rect 53430 22040 53440 22120
rect 53050 21940 53130 21950
rect 53200 21940 53280 21950
rect 53350 21940 53430 21950
rect 53130 21860 53140 21940
rect 53280 21860 53290 21940
rect 53430 21860 53440 21940
rect 53050 21760 53130 21770
rect 53200 21760 53280 21770
rect 53350 21760 53430 21770
rect 53130 21680 53140 21760
rect 53280 21680 53290 21760
rect 53430 21680 53440 21760
rect 53050 21580 53130 21590
rect 53200 21580 53280 21590
rect 53350 21580 53430 21590
rect 53130 21500 53140 21580
rect 53280 21500 53290 21580
rect 53430 21500 53440 21580
rect 53050 21400 53130 21410
rect 53200 21400 53280 21410
rect 53350 21400 53430 21410
rect 53130 21320 53140 21400
rect 53280 21320 53290 21400
rect 53430 21320 53440 21400
rect 53050 21220 53130 21230
rect 53200 21220 53280 21230
rect 53350 21220 53430 21230
rect 53130 21140 53140 21220
rect 53280 21140 53290 21220
rect 53430 21140 53440 21220
rect 53050 21040 53130 21050
rect 53200 21040 53280 21050
rect 53350 21040 53430 21050
rect 53130 20960 53140 21040
rect 53280 20960 53290 21040
rect 53430 20960 53440 21040
rect 53050 20860 53130 20870
rect 53200 20860 53280 20870
rect 53350 20860 53430 20870
rect 53130 20780 53140 20860
rect 53280 20780 53290 20860
rect 53430 20780 53440 20860
rect 53050 20680 53130 20690
rect 53200 20680 53280 20690
rect 53350 20680 53430 20690
rect 53130 20600 53140 20680
rect 53280 20600 53290 20680
rect 53430 20600 53440 20680
rect 53050 20500 53130 20510
rect 53200 20500 53280 20510
rect 53350 20500 53430 20510
rect 53130 20420 53140 20500
rect 53280 20420 53290 20500
rect 53430 20420 53440 20500
rect 53050 20320 53130 20330
rect 53200 20320 53280 20330
rect 53350 20320 53430 20330
rect 53130 20240 53140 20320
rect 53280 20240 53290 20320
rect 53430 20240 53440 20320
rect 53050 20140 53130 20150
rect 53200 20140 53280 20150
rect 53350 20140 53430 20150
rect 53130 20060 53140 20140
rect 53280 20060 53290 20140
rect 53430 20060 53440 20140
rect 53050 19960 53130 19970
rect 53200 19960 53280 19970
rect 53350 19960 53430 19970
rect 53130 19880 53140 19960
rect 53280 19880 53290 19960
rect 53430 19880 53440 19960
rect 53570 19800 53580 25800
rect 53690 25720 53770 25730
rect 53990 25720 54070 25730
rect 53770 25640 53780 25720
rect 54070 25640 54080 25720
rect 53690 25540 53770 25550
rect 53990 25540 54070 25550
rect 53770 25460 53780 25540
rect 54070 25460 54080 25540
rect 53690 25360 53770 25370
rect 53990 25360 54070 25370
rect 53770 25280 53780 25360
rect 54070 25280 54080 25360
rect 53690 25180 53770 25190
rect 53990 25180 54070 25190
rect 53770 25100 53780 25180
rect 54070 25100 54080 25180
rect 53690 25000 53770 25010
rect 53990 25000 54070 25010
rect 53770 24920 53780 25000
rect 54070 24920 54080 25000
rect 53690 24820 53770 24830
rect 53990 24820 54070 24830
rect 53770 24740 53780 24820
rect 54070 24740 54080 24820
rect 53690 24640 53770 24650
rect 53990 24640 54070 24650
rect 53770 24560 53780 24640
rect 54070 24560 54080 24640
rect 53690 24460 53770 24470
rect 53990 24460 54070 24470
rect 53770 24380 53780 24460
rect 54070 24380 54080 24460
rect 53690 24280 53770 24290
rect 53990 24280 54070 24290
rect 53770 24200 53780 24280
rect 54070 24200 54080 24280
rect 53690 24100 53770 24110
rect 53990 24100 54070 24110
rect 53770 24020 53780 24100
rect 54070 24020 54080 24100
rect 53690 23920 53770 23930
rect 53990 23920 54070 23930
rect 53770 23840 53780 23920
rect 54070 23840 54080 23920
rect 53690 23740 53770 23750
rect 53990 23740 54070 23750
rect 53770 23660 53780 23740
rect 54070 23660 54080 23740
rect 53690 23560 53770 23570
rect 53990 23560 54070 23570
rect 53770 23480 53780 23560
rect 54070 23480 54080 23560
rect 53690 23380 53770 23390
rect 53990 23380 54070 23390
rect 53770 23300 53780 23380
rect 54070 23300 54080 23380
rect 53690 23200 53770 23210
rect 53990 23200 54070 23210
rect 53770 23120 53780 23200
rect 54070 23120 54080 23200
rect 53690 23020 53770 23030
rect 53990 23020 54070 23030
rect 53770 22940 53780 23020
rect 54070 22940 54080 23020
rect 53690 22840 53770 22850
rect 53990 22840 54070 22850
rect 53770 22760 53780 22840
rect 54070 22760 54080 22840
rect 53690 22660 53770 22670
rect 53990 22660 54070 22670
rect 53770 22580 53780 22660
rect 54070 22580 54080 22660
rect 53690 22480 53770 22490
rect 53990 22480 54070 22490
rect 53770 22400 53780 22480
rect 54070 22400 54080 22480
rect 53690 22300 53770 22310
rect 53990 22300 54070 22310
rect 53770 22220 53780 22300
rect 54070 22220 54080 22300
rect 53690 22120 53770 22130
rect 53990 22120 54070 22130
rect 53770 22040 53780 22120
rect 54070 22040 54080 22120
rect 53690 21940 53770 21950
rect 53990 21940 54070 21950
rect 53770 21860 53780 21940
rect 54070 21860 54080 21940
rect 53690 21760 53770 21770
rect 53990 21760 54070 21770
rect 53770 21680 53780 21760
rect 54070 21680 54080 21760
rect 53690 21580 53770 21590
rect 53990 21580 54070 21590
rect 53770 21500 53780 21580
rect 54070 21500 54080 21580
rect 53690 21400 53770 21410
rect 53990 21400 54070 21410
rect 53770 21320 53780 21400
rect 54070 21320 54080 21400
rect 53690 21220 53770 21230
rect 53990 21220 54070 21230
rect 53770 21140 53780 21220
rect 54070 21140 54080 21220
rect 53690 21040 53770 21050
rect 53990 21040 54070 21050
rect 53770 20960 53780 21040
rect 54070 20960 54080 21040
rect 53690 20860 53770 20870
rect 53990 20860 54070 20870
rect 53770 20780 53780 20860
rect 54070 20780 54080 20860
rect 53690 20680 53770 20690
rect 53990 20680 54070 20690
rect 53770 20600 53780 20680
rect 54070 20600 54080 20680
rect 53690 20500 53770 20510
rect 53990 20500 54070 20510
rect 53770 20420 53780 20500
rect 54070 20420 54080 20500
rect 53690 20320 53770 20330
rect 53990 20320 54070 20330
rect 53770 20240 53780 20320
rect 54070 20240 54080 20320
rect 53690 20140 53770 20150
rect 53990 20140 54070 20150
rect 53770 20060 53780 20140
rect 54070 20060 54080 20140
rect 53690 19960 53770 19970
rect 53990 19960 54070 19970
rect 53770 19880 53780 19960
rect 54070 19880 54080 19960
rect 54250 19800 54260 25800
rect 54310 25720 54390 25730
rect 54460 25720 54540 25730
rect 54610 25720 54690 25730
rect 54390 25640 54400 25720
rect 54540 25640 54550 25720
rect 54690 25640 54700 25720
rect 54310 25540 54390 25550
rect 54460 25540 54540 25550
rect 54610 25540 54690 25550
rect 54390 25460 54400 25540
rect 54540 25460 54550 25540
rect 54690 25460 54700 25540
rect 54310 25360 54390 25370
rect 54460 25360 54540 25370
rect 54610 25360 54690 25370
rect 54390 25280 54400 25360
rect 54540 25280 54550 25360
rect 54690 25280 54700 25360
rect 54310 25180 54390 25190
rect 54460 25180 54540 25190
rect 54610 25180 54690 25190
rect 54390 25100 54400 25180
rect 54540 25100 54550 25180
rect 54690 25100 54700 25180
rect 54310 25000 54390 25010
rect 54460 25000 54540 25010
rect 54610 25000 54690 25010
rect 54390 24920 54400 25000
rect 54540 24920 54550 25000
rect 54690 24920 54700 25000
rect 54310 24820 54390 24830
rect 54460 24820 54540 24830
rect 54610 24820 54690 24830
rect 54390 24740 54400 24820
rect 54540 24740 54550 24820
rect 54690 24740 54700 24820
rect 54310 24640 54390 24650
rect 54460 24640 54540 24650
rect 54610 24640 54690 24650
rect 54390 24560 54400 24640
rect 54540 24560 54550 24640
rect 54690 24560 54700 24640
rect 54310 24460 54390 24470
rect 54460 24460 54540 24470
rect 54610 24460 54690 24470
rect 54390 24380 54400 24460
rect 54540 24380 54550 24460
rect 54690 24380 54700 24460
rect 54310 24280 54390 24290
rect 54460 24280 54540 24290
rect 54610 24280 54690 24290
rect 54390 24200 54400 24280
rect 54540 24200 54550 24280
rect 54690 24200 54700 24280
rect 54310 24100 54390 24110
rect 54460 24100 54540 24110
rect 54610 24100 54690 24110
rect 54390 24020 54400 24100
rect 54540 24020 54550 24100
rect 54690 24020 54700 24100
rect 54310 23920 54390 23930
rect 54460 23920 54540 23930
rect 54610 23920 54690 23930
rect 54390 23840 54400 23920
rect 54540 23840 54550 23920
rect 54690 23840 54700 23920
rect 54310 23740 54390 23750
rect 54460 23740 54540 23750
rect 54610 23740 54690 23750
rect 54390 23660 54400 23740
rect 54540 23660 54550 23740
rect 54690 23660 54700 23740
rect 54310 23560 54390 23570
rect 54460 23560 54540 23570
rect 54610 23560 54690 23570
rect 54390 23480 54400 23560
rect 54540 23480 54550 23560
rect 54690 23480 54700 23560
rect 54310 23380 54390 23390
rect 54460 23380 54540 23390
rect 54610 23380 54690 23390
rect 54390 23300 54400 23380
rect 54540 23300 54550 23380
rect 54690 23300 54700 23380
rect 54310 23200 54390 23210
rect 54460 23200 54540 23210
rect 54610 23200 54690 23210
rect 54390 23120 54400 23200
rect 54540 23120 54550 23200
rect 54690 23120 54700 23200
rect 54310 23020 54390 23030
rect 54460 23020 54540 23030
rect 54610 23020 54690 23030
rect 54390 22940 54400 23020
rect 54540 22940 54550 23020
rect 54690 22940 54700 23020
rect 54310 22840 54390 22850
rect 54460 22840 54540 22850
rect 54610 22840 54690 22850
rect 54390 22760 54400 22840
rect 54540 22760 54550 22840
rect 54690 22760 54700 22840
rect 54310 22660 54390 22670
rect 54460 22660 54540 22670
rect 54610 22660 54690 22670
rect 54390 22580 54400 22660
rect 54540 22580 54550 22660
rect 54690 22580 54700 22660
rect 54310 22480 54390 22490
rect 54460 22480 54540 22490
rect 54610 22480 54690 22490
rect 54390 22400 54400 22480
rect 54540 22400 54550 22480
rect 54690 22400 54700 22480
rect 54310 22300 54390 22310
rect 54460 22300 54540 22310
rect 54610 22300 54690 22310
rect 54390 22220 54400 22300
rect 54540 22220 54550 22300
rect 54690 22220 54700 22300
rect 54310 22120 54390 22130
rect 54460 22120 54540 22130
rect 54610 22120 54690 22130
rect 54390 22040 54400 22120
rect 54540 22040 54550 22120
rect 54690 22040 54700 22120
rect 54310 21940 54390 21950
rect 54460 21940 54540 21950
rect 54610 21940 54690 21950
rect 54390 21860 54400 21940
rect 54540 21860 54550 21940
rect 54690 21860 54700 21940
rect 54310 21760 54390 21770
rect 54460 21760 54540 21770
rect 54610 21760 54690 21770
rect 54390 21680 54400 21760
rect 54540 21680 54550 21760
rect 54690 21680 54700 21760
rect 54310 21580 54390 21590
rect 54460 21580 54540 21590
rect 54610 21580 54690 21590
rect 54390 21500 54400 21580
rect 54540 21500 54550 21580
rect 54690 21500 54700 21580
rect 54310 21400 54390 21410
rect 54460 21400 54540 21410
rect 54610 21400 54690 21410
rect 54390 21320 54400 21400
rect 54540 21320 54550 21400
rect 54690 21320 54700 21400
rect 54310 21220 54390 21230
rect 54460 21220 54540 21230
rect 54610 21220 54690 21230
rect 54390 21140 54400 21220
rect 54540 21140 54550 21220
rect 54690 21140 54700 21220
rect 54310 21040 54390 21050
rect 54460 21040 54540 21050
rect 54610 21040 54690 21050
rect 54390 20960 54400 21040
rect 54540 20960 54550 21040
rect 54690 20960 54700 21040
rect 54310 20860 54390 20870
rect 54460 20860 54540 20870
rect 54610 20860 54690 20870
rect 54390 20780 54400 20860
rect 54540 20780 54550 20860
rect 54690 20780 54700 20860
rect 54310 20680 54390 20690
rect 54460 20680 54540 20690
rect 54610 20680 54690 20690
rect 54390 20600 54400 20680
rect 54540 20600 54550 20680
rect 54690 20600 54700 20680
rect 54310 20500 54390 20510
rect 54460 20500 54540 20510
rect 54610 20500 54690 20510
rect 54390 20420 54400 20500
rect 54540 20420 54550 20500
rect 54690 20420 54700 20500
rect 54310 20320 54390 20330
rect 54460 20320 54540 20330
rect 54610 20320 54690 20330
rect 54390 20240 54400 20320
rect 54540 20240 54550 20320
rect 54690 20240 54700 20320
rect 54310 20140 54390 20150
rect 54460 20140 54540 20150
rect 54610 20140 54690 20150
rect 54390 20060 54400 20140
rect 54540 20060 54550 20140
rect 54690 20060 54700 20140
rect 54310 19960 54390 19970
rect 54460 19960 54540 19970
rect 54610 19960 54690 19970
rect 54390 19880 54400 19960
rect 54540 19880 54550 19960
rect 54690 19880 54700 19960
rect 54830 19800 54840 25800
rect 54950 25720 55030 25730
rect 55250 25720 55330 25730
rect 55030 25640 55040 25720
rect 55330 25640 55340 25720
rect 54950 25540 55030 25550
rect 55250 25540 55330 25550
rect 55030 25460 55040 25540
rect 55330 25460 55340 25540
rect 54950 25360 55030 25370
rect 55250 25360 55330 25370
rect 55030 25280 55040 25360
rect 55330 25280 55340 25360
rect 54950 25180 55030 25190
rect 55250 25180 55330 25190
rect 55030 25100 55040 25180
rect 55330 25100 55340 25180
rect 54950 25000 55030 25010
rect 55250 25000 55330 25010
rect 55030 24920 55040 25000
rect 55330 24920 55340 25000
rect 54950 24820 55030 24830
rect 55250 24820 55330 24830
rect 55030 24740 55040 24820
rect 55330 24740 55340 24820
rect 54950 24640 55030 24650
rect 55250 24640 55330 24650
rect 55030 24560 55040 24640
rect 55330 24560 55340 24640
rect 54950 24460 55030 24470
rect 55250 24460 55330 24470
rect 55030 24380 55040 24460
rect 55330 24380 55340 24460
rect 54950 24280 55030 24290
rect 55250 24280 55330 24290
rect 55030 24200 55040 24280
rect 55330 24200 55340 24280
rect 54950 24100 55030 24110
rect 55250 24100 55330 24110
rect 55030 24020 55040 24100
rect 55330 24020 55340 24100
rect 54950 23920 55030 23930
rect 55250 23920 55330 23930
rect 55030 23840 55040 23920
rect 55330 23840 55340 23920
rect 54950 23740 55030 23750
rect 55250 23740 55330 23750
rect 55030 23660 55040 23740
rect 55330 23660 55340 23740
rect 54950 23560 55030 23570
rect 55250 23560 55330 23570
rect 55030 23480 55040 23560
rect 55330 23480 55340 23560
rect 54950 23380 55030 23390
rect 55250 23380 55330 23390
rect 55030 23300 55040 23380
rect 55330 23300 55340 23380
rect 54950 23200 55030 23210
rect 55250 23200 55330 23210
rect 55030 23120 55040 23200
rect 55330 23120 55340 23200
rect 54950 23020 55030 23030
rect 55250 23020 55330 23030
rect 55030 22940 55040 23020
rect 55330 22940 55340 23020
rect 54950 22840 55030 22850
rect 55250 22840 55330 22850
rect 55030 22760 55040 22840
rect 55330 22760 55340 22840
rect 54950 22660 55030 22670
rect 55250 22660 55330 22670
rect 55030 22580 55040 22660
rect 55330 22580 55340 22660
rect 54950 22480 55030 22490
rect 55250 22480 55330 22490
rect 55030 22400 55040 22480
rect 55330 22400 55340 22480
rect 54950 22300 55030 22310
rect 55250 22300 55330 22310
rect 55030 22220 55040 22300
rect 55330 22220 55340 22300
rect 54950 22120 55030 22130
rect 55250 22120 55330 22130
rect 55030 22040 55040 22120
rect 55330 22040 55340 22120
rect 54950 21940 55030 21950
rect 55250 21940 55330 21950
rect 55030 21860 55040 21940
rect 55330 21860 55340 21940
rect 54950 21760 55030 21770
rect 55250 21760 55330 21770
rect 55030 21680 55040 21760
rect 55330 21680 55340 21760
rect 54950 21580 55030 21590
rect 55250 21580 55330 21590
rect 55030 21500 55040 21580
rect 55330 21500 55340 21580
rect 54950 21400 55030 21410
rect 55250 21400 55330 21410
rect 55030 21320 55040 21400
rect 55330 21320 55340 21400
rect 54950 21220 55030 21230
rect 55250 21220 55330 21230
rect 55030 21140 55040 21220
rect 55330 21140 55340 21220
rect 54950 21040 55030 21050
rect 55250 21040 55330 21050
rect 55030 20960 55040 21040
rect 55330 20960 55340 21040
rect 54950 20860 55030 20870
rect 55250 20860 55330 20870
rect 55030 20780 55040 20860
rect 55330 20780 55340 20860
rect 54950 20680 55030 20690
rect 55250 20680 55330 20690
rect 55030 20600 55040 20680
rect 55330 20600 55340 20680
rect 54950 20500 55030 20510
rect 55250 20500 55330 20510
rect 55030 20420 55040 20500
rect 55330 20420 55340 20500
rect 54950 20320 55030 20330
rect 55250 20320 55330 20330
rect 55030 20240 55040 20320
rect 55330 20240 55340 20320
rect 54950 20140 55030 20150
rect 55250 20140 55330 20150
rect 55030 20060 55040 20140
rect 55330 20060 55340 20140
rect 54950 19960 55030 19970
rect 55250 19960 55330 19970
rect 55030 19880 55040 19960
rect 55330 19880 55340 19960
rect 55510 19800 55520 25800
rect 55570 25720 55650 25730
rect 55720 25720 55800 25730
rect 55870 25720 55950 25730
rect 55650 25640 55660 25720
rect 55800 25640 55810 25720
rect 55950 25640 55960 25720
rect 55570 25540 55650 25550
rect 55720 25540 55800 25550
rect 55870 25540 55950 25550
rect 55650 25460 55660 25540
rect 55800 25460 55810 25540
rect 55950 25460 55960 25540
rect 55570 25360 55650 25370
rect 55720 25360 55800 25370
rect 55870 25360 55950 25370
rect 55650 25280 55660 25360
rect 55800 25280 55810 25360
rect 55950 25280 55960 25360
rect 55570 25180 55650 25190
rect 55720 25180 55800 25190
rect 55870 25180 55950 25190
rect 55650 25100 55660 25180
rect 55800 25100 55810 25180
rect 55950 25100 55960 25180
rect 55570 25000 55650 25010
rect 55720 25000 55800 25010
rect 55870 25000 55950 25010
rect 55650 24920 55660 25000
rect 55800 24920 55810 25000
rect 55950 24920 55960 25000
rect 55570 24820 55650 24830
rect 55720 24820 55800 24830
rect 55870 24820 55950 24830
rect 55650 24740 55660 24820
rect 55800 24740 55810 24820
rect 55950 24740 55960 24820
rect 55570 24640 55650 24650
rect 55720 24640 55800 24650
rect 55870 24640 55950 24650
rect 55650 24560 55660 24640
rect 55800 24560 55810 24640
rect 55950 24560 55960 24640
rect 55570 24460 55650 24470
rect 55720 24460 55800 24470
rect 55870 24460 55950 24470
rect 55650 24380 55660 24460
rect 55800 24380 55810 24460
rect 55950 24380 55960 24460
rect 55570 24280 55650 24290
rect 55720 24280 55800 24290
rect 55870 24280 55950 24290
rect 55650 24200 55660 24280
rect 55800 24200 55810 24280
rect 55950 24200 55960 24280
rect 55570 24100 55650 24110
rect 55720 24100 55800 24110
rect 55870 24100 55950 24110
rect 55650 24020 55660 24100
rect 55800 24020 55810 24100
rect 55950 24020 55960 24100
rect 55570 23920 55650 23930
rect 55720 23920 55800 23930
rect 55870 23920 55950 23930
rect 55650 23840 55660 23920
rect 55800 23840 55810 23920
rect 55950 23840 55960 23920
rect 55570 23740 55650 23750
rect 55720 23740 55800 23750
rect 55870 23740 55950 23750
rect 55650 23660 55660 23740
rect 55800 23660 55810 23740
rect 55950 23660 55960 23740
rect 55570 23560 55650 23570
rect 55720 23560 55800 23570
rect 55870 23560 55950 23570
rect 55650 23480 55660 23560
rect 55800 23480 55810 23560
rect 55950 23480 55960 23560
rect 55570 23380 55650 23390
rect 55720 23380 55800 23390
rect 55870 23380 55950 23390
rect 55650 23300 55660 23380
rect 55800 23300 55810 23380
rect 55950 23300 55960 23380
rect 55570 23200 55650 23210
rect 55720 23200 55800 23210
rect 55870 23200 55950 23210
rect 55650 23120 55660 23200
rect 55800 23120 55810 23200
rect 55950 23120 55960 23200
rect 55570 23020 55650 23030
rect 55720 23020 55800 23030
rect 55870 23020 55950 23030
rect 55650 22940 55660 23020
rect 55800 22940 55810 23020
rect 55950 22940 55960 23020
rect 55570 22840 55650 22850
rect 55720 22840 55800 22850
rect 55870 22840 55950 22850
rect 55650 22760 55660 22840
rect 55800 22760 55810 22840
rect 55950 22760 55960 22840
rect 55570 22660 55650 22670
rect 55720 22660 55800 22670
rect 55870 22660 55950 22670
rect 55650 22580 55660 22660
rect 55800 22580 55810 22660
rect 55950 22580 55960 22660
rect 55570 22480 55650 22490
rect 55720 22480 55800 22490
rect 55870 22480 55950 22490
rect 55650 22400 55660 22480
rect 55800 22400 55810 22480
rect 55950 22400 55960 22480
rect 55570 22300 55650 22310
rect 55720 22300 55800 22310
rect 55870 22300 55950 22310
rect 55650 22220 55660 22300
rect 55800 22220 55810 22300
rect 55950 22220 55960 22300
rect 55570 22120 55650 22130
rect 55720 22120 55800 22130
rect 55870 22120 55950 22130
rect 55650 22040 55660 22120
rect 55800 22040 55810 22120
rect 55950 22040 55960 22120
rect 55570 21940 55650 21950
rect 55720 21940 55800 21950
rect 55870 21940 55950 21950
rect 55650 21860 55660 21940
rect 55800 21860 55810 21940
rect 55950 21860 55960 21940
rect 55570 21760 55650 21770
rect 55720 21760 55800 21770
rect 55870 21760 55950 21770
rect 55650 21680 55660 21760
rect 55800 21680 55810 21760
rect 55950 21680 55960 21760
rect 55570 21580 55650 21590
rect 55720 21580 55800 21590
rect 55870 21580 55950 21590
rect 55650 21500 55660 21580
rect 55800 21500 55810 21580
rect 55950 21500 55960 21580
rect 55570 21400 55650 21410
rect 55720 21400 55800 21410
rect 55870 21400 55950 21410
rect 55650 21320 55660 21400
rect 55800 21320 55810 21400
rect 55950 21320 55960 21400
rect 55570 21220 55650 21230
rect 55720 21220 55800 21230
rect 55870 21220 55950 21230
rect 55650 21140 55660 21220
rect 55800 21140 55810 21220
rect 55950 21140 55960 21220
rect 55570 21040 55650 21050
rect 55720 21040 55800 21050
rect 55870 21040 55950 21050
rect 55650 20960 55660 21040
rect 55800 20960 55810 21040
rect 55950 20960 55960 21040
rect 55570 20860 55650 20870
rect 55720 20860 55800 20870
rect 55870 20860 55950 20870
rect 55650 20780 55660 20860
rect 55800 20780 55810 20860
rect 55950 20780 55960 20860
rect 55570 20680 55650 20690
rect 55720 20680 55800 20690
rect 55870 20680 55950 20690
rect 55650 20600 55660 20680
rect 55800 20600 55810 20680
rect 55950 20600 55960 20680
rect 55570 20500 55650 20510
rect 55720 20500 55800 20510
rect 55870 20500 55950 20510
rect 55650 20420 55660 20500
rect 55800 20420 55810 20500
rect 55950 20420 55960 20500
rect 55570 20320 55650 20330
rect 55720 20320 55800 20330
rect 55870 20320 55950 20330
rect 55650 20240 55660 20320
rect 55800 20240 55810 20320
rect 55950 20240 55960 20320
rect 55570 20140 55650 20150
rect 55720 20140 55800 20150
rect 55870 20140 55950 20150
rect 55650 20060 55660 20140
rect 55800 20060 55810 20140
rect 55950 20060 55960 20140
rect 55570 19960 55650 19970
rect 55720 19960 55800 19970
rect 55870 19960 55950 19970
rect 55650 19880 55660 19960
rect 55800 19880 55810 19960
rect 55950 19880 55960 19960
rect 56090 19800 56100 25800
rect 56210 25720 56290 25730
rect 56510 25720 56590 25730
rect 56290 25640 56300 25720
rect 56590 25640 56600 25720
rect 56210 25540 56290 25550
rect 56510 25540 56590 25550
rect 56290 25460 56300 25540
rect 56590 25460 56600 25540
rect 56210 25360 56290 25370
rect 56510 25360 56590 25370
rect 56290 25280 56300 25360
rect 56590 25280 56600 25360
rect 56210 25180 56290 25190
rect 56510 25180 56590 25190
rect 56290 25100 56300 25180
rect 56590 25100 56600 25180
rect 56210 25000 56290 25010
rect 56510 25000 56590 25010
rect 56290 24920 56300 25000
rect 56590 24920 56600 25000
rect 56210 24820 56290 24830
rect 56510 24820 56590 24830
rect 56290 24740 56300 24820
rect 56590 24740 56600 24820
rect 56210 24640 56290 24650
rect 56510 24640 56590 24650
rect 56290 24560 56300 24640
rect 56590 24560 56600 24640
rect 56210 24460 56290 24470
rect 56510 24460 56590 24470
rect 56290 24380 56300 24460
rect 56590 24380 56600 24460
rect 56210 24280 56290 24290
rect 56510 24280 56590 24290
rect 56290 24200 56300 24280
rect 56590 24200 56600 24280
rect 56210 24100 56290 24110
rect 56510 24100 56590 24110
rect 56290 24020 56300 24100
rect 56590 24020 56600 24100
rect 56210 23920 56290 23930
rect 56510 23920 56590 23930
rect 56290 23840 56300 23920
rect 56590 23840 56600 23920
rect 56210 23740 56290 23750
rect 56510 23740 56590 23750
rect 56290 23660 56300 23740
rect 56590 23660 56600 23740
rect 56210 23560 56290 23570
rect 56510 23560 56590 23570
rect 56290 23480 56300 23560
rect 56590 23480 56600 23560
rect 56210 23380 56290 23390
rect 56510 23380 56590 23390
rect 56290 23300 56300 23380
rect 56590 23300 56600 23380
rect 56210 23200 56290 23210
rect 56510 23200 56590 23210
rect 56290 23120 56300 23200
rect 56590 23120 56600 23200
rect 56210 23020 56290 23030
rect 56510 23020 56590 23030
rect 56290 22940 56300 23020
rect 56590 22940 56600 23020
rect 56210 22840 56290 22850
rect 56510 22840 56590 22850
rect 56290 22760 56300 22840
rect 56590 22760 56600 22840
rect 56210 22660 56290 22670
rect 56510 22660 56590 22670
rect 56290 22580 56300 22660
rect 56590 22580 56600 22660
rect 56210 22480 56290 22490
rect 56510 22480 56590 22490
rect 56290 22400 56300 22480
rect 56590 22400 56600 22480
rect 56210 22300 56290 22310
rect 56510 22300 56590 22310
rect 56290 22220 56300 22300
rect 56590 22220 56600 22300
rect 56210 22120 56290 22130
rect 56510 22120 56590 22130
rect 56290 22040 56300 22120
rect 56590 22040 56600 22120
rect 56210 21940 56290 21950
rect 56510 21940 56590 21950
rect 56290 21860 56300 21940
rect 56590 21860 56600 21940
rect 56210 21760 56290 21770
rect 56510 21760 56590 21770
rect 56290 21680 56300 21760
rect 56590 21680 56600 21760
rect 56210 21580 56290 21590
rect 56510 21580 56590 21590
rect 56290 21500 56300 21580
rect 56590 21500 56600 21580
rect 56210 21400 56290 21410
rect 56510 21400 56590 21410
rect 56290 21320 56300 21400
rect 56590 21320 56600 21400
rect 56210 21220 56290 21230
rect 56510 21220 56590 21230
rect 56290 21140 56300 21220
rect 56590 21140 56600 21220
rect 56210 21040 56290 21050
rect 56510 21040 56590 21050
rect 56290 20960 56300 21040
rect 56590 20960 56600 21040
rect 56210 20860 56290 20870
rect 56510 20860 56590 20870
rect 56290 20780 56300 20860
rect 56590 20780 56600 20860
rect 56210 20680 56290 20690
rect 56510 20680 56590 20690
rect 56290 20600 56300 20680
rect 56590 20600 56600 20680
rect 56210 20500 56290 20510
rect 56510 20500 56590 20510
rect 56290 20420 56300 20500
rect 56590 20420 56600 20500
rect 56210 20320 56290 20330
rect 56510 20320 56590 20330
rect 56290 20240 56300 20320
rect 56590 20240 56600 20320
rect 56210 20140 56290 20150
rect 56510 20140 56590 20150
rect 56290 20060 56300 20140
rect 56590 20060 56600 20140
rect 56210 19960 56290 19970
rect 56510 19960 56590 19970
rect 56290 19880 56300 19960
rect 56590 19880 56600 19960
rect 56770 19800 56780 25800
rect 56830 25720 56910 25730
rect 56980 25720 57060 25730
rect 57130 25720 57210 25730
rect 56910 25640 56920 25720
rect 57060 25640 57070 25720
rect 57210 25640 57220 25720
rect 56830 25540 56910 25550
rect 56980 25540 57060 25550
rect 57130 25540 57210 25550
rect 56910 25460 56920 25540
rect 57060 25460 57070 25540
rect 57210 25460 57220 25540
rect 56830 25360 56910 25370
rect 56980 25360 57060 25370
rect 57130 25360 57210 25370
rect 56910 25280 56920 25360
rect 57060 25280 57070 25360
rect 57210 25280 57220 25360
rect 56830 25180 56910 25190
rect 56980 25180 57060 25190
rect 57130 25180 57210 25190
rect 56910 25100 56920 25180
rect 57060 25100 57070 25180
rect 57210 25100 57220 25180
rect 56830 25000 56910 25010
rect 56980 25000 57060 25010
rect 57130 25000 57210 25010
rect 56910 24920 56920 25000
rect 57060 24920 57070 25000
rect 57210 24920 57220 25000
rect 56830 24820 56910 24830
rect 56980 24820 57060 24830
rect 57130 24820 57210 24830
rect 56910 24740 56920 24820
rect 57060 24740 57070 24820
rect 57210 24740 57220 24820
rect 56830 24640 56910 24650
rect 56980 24640 57060 24650
rect 57130 24640 57210 24650
rect 56910 24560 56920 24640
rect 57060 24560 57070 24640
rect 57210 24560 57220 24640
rect 56830 24460 56910 24470
rect 56980 24460 57060 24470
rect 57130 24460 57210 24470
rect 56910 24380 56920 24460
rect 57060 24380 57070 24460
rect 57210 24380 57220 24460
rect 56830 24280 56910 24290
rect 56980 24280 57060 24290
rect 57130 24280 57210 24290
rect 56910 24200 56920 24280
rect 57060 24200 57070 24280
rect 57210 24200 57220 24280
rect 56830 24100 56910 24110
rect 56980 24100 57060 24110
rect 57130 24100 57210 24110
rect 56910 24020 56920 24100
rect 57060 24020 57070 24100
rect 57210 24020 57220 24100
rect 56830 23920 56910 23930
rect 56980 23920 57060 23930
rect 57130 23920 57210 23930
rect 56910 23840 56920 23920
rect 57060 23840 57070 23920
rect 57210 23840 57220 23920
rect 56830 23740 56910 23750
rect 56980 23740 57060 23750
rect 57130 23740 57210 23750
rect 56910 23660 56920 23740
rect 57060 23660 57070 23740
rect 57210 23660 57220 23740
rect 56830 23560 56910 23570
rect 56980 23560 57060 23570
rect 57130 23560 57210 23570
rect 56910 23480 56920 23560
rect 57060 23480 57070 23560
rect 57210 23480 57220 23560
rect 56830 23380 56910 23390
rect 56980 23380 57060 23390
rect 57130 23380 57210 23390
rect 56910 23300 56920 23380
rect 57060 23300 57070 23380
rect 57210 23300 57220 23380
rect 56830 23200 56910 23210
rect 56980 23200 57060 23210
rect 57130 23200 57210 23210
rect 56910 23120 56920 23200
rect 57060 23120 57070 23200
rect 57210 23120 57220 23200
rect 56830 23020 56910 23030
rect 56980 23020 57060 23030
rect 57130 23020 57210 23030
rect 56910 22940 56920 23020
rect 57060 22940 57070 23020
rect 57210 22940 57220 23020
rect 56830 22840 56910 22850
rect 56980 22840 57060 22850
rect 57130 22840 57210 22850
rect 56910 22760 56920 22840
rect 57060 22760 57070 22840
rect 57210 22760 57220 22840
rect 56830 22660 56910 22670
rect 56980 22660 57060 22670
rect 57130 22660 57210 22670
rect 56910 22580 56920 22660
rect 57060 22580 57070 22660
rect 57210 22580 57220 22660
rect 56830 22480 56910 22490
rect 56980 22480 57060 22490
rect 57130 22480 57210 22490
rect 56910 22400 56920 22480
rect 57060 22400 57070 22480
rect 57210 22400 57220 22480
rect 56830 22300 56910 22310
rect 56980 22300 57060 22310
rect 57130 22300 57210 22310
rect 56910 22220 56920 22300
rect 57060 22220 57070 22300
rect 57210 22220 57220 22300
rect 56830 22120 56910 22130
rect 56980 22120 57060 22130
rect 57130 22120 57210 22130
rect 56910 22040 56920 22120
rect 57060 22040 57070 22120
rect 57210 22040 57220 22120
rect 56830 21940 56910 21950
rect 56980 21940 57060 21950
rect 57130 21940 57210 21950
rect 56910 21860 56920 21940
rect 57060 21860 57070 21940
rect 57210 21860 57220 21940
rect 56830 21760 56910 21770
rect 56980 21760 57060 21770
rect 57130 21760 57210 21770
rect 56910 21680 56920 21760
rect 57060 21680 57070 21760
rect 57210 21680 57220 21760
rect 56830 21580 56910 21590
rect 56980 21580 57060 21590
rect 57130 21580 57210 21590
rect 56910 21500 56920 21580
rect 57060 21500 57070 21580
rect 57210 21500 57220 21580
rect 56830 21400 56910 21410
rect 56980 21400 57060 21410
rect 57130 21400 57210 21410
rect 56910 21320 56920 21400
rect 57060 21320 57070 21400
rect 57210 21320 57220 21400
rect 56830 21220 56910 21230
rect 56980 21220 57060 21230
rect 57130 21220 57210 21230
rect 56910 21140 56920 21220
rect 57060 21140 57070 21220
rect 57210 21140 57220 21220
rect 56830 21040 56910 21050
rect 56980 21040 57060 21050
rect 57130 21040 57210 21050
rect 56910 20960 56920 21040
rect 57060 20960 57070 21040
rect 57210 20960 57220 21040
rect 56830 20860 56910 20870
rect 56980 20860 57060 20870
rect 57130 20860 57210 20870
rect 56910 20780 56920 20860
rect 57060 20780 57070 20860
rect 57210 20780 57220 20860
rect 56830 20680 56910 20690
rect 56980 20680 57060 20690
rect 57130 20680 57210 20690
rect 56910 20600 56920 20680
rect 57060 20600 57070 20680
rect 57210 20600 57220 20680
rect 56830 20500 56910 20510
rect 56980 20500 57060 20510
rect 57130 20500 57210 20510
rect 56910 20420 56920 20500
rect 57060 20420 57070 20500
rect 57210 20420 57220 20500
rect 56830 20320 56910 20330
rect 56980 20320 57060 20330
rect 57130 20320 57210 20330
rect 56910 20240 56920 20320
rect 57060 20240 57070 20320
rect 57210 20240 57220 20320
rect 56830 20140 56910 20150
rect 56980 20140 57060 20150
rect 57130 20140 57210 20150
rect 56910 20060 56920 20140
rect 57060 20060 57070 20140
rect 57210 20060 57220 20140
rect 56830 19960 56910 19970
rect 56980 19960 57060 19970
rect 57130 19960 57210 19970
rect 56910 19880 56920 19960
rect 57060 19880 57070 19960
rect 57210 19880 57220 19960
rect 57350 19800 57360 25800
rect 57470 25720 57550 25730
rect 57770 25720 57850 25730
rect 57550 25640 57560 25720
rect 57850 25640 57860 25720
rect 57470 25540 57550 25550
rect 57770 25540 57850 25550
rect 57550 25460 57560 25540
rect 57850 25460 57860 25540
rect 57470 25360 57550 25370
rect 57770 25360 57850 25370
rect 57550 25280 57560 25360
rect 57850 25280 57860 25360
rect 57470 25180 57550 25190
rect 57770 25180 57850 25190
rect 57550 25100 57560 25180
rect 57850 25100 57860 25180
rect 57470 25000 57550 25010
rect 57770 25000 57850 25010
rect 57550 24920 57560 25000
rect 57850 24920 57860 25000
rect 57470 24820 57550 24830
rect 57770 24820 57850 24830
rect 57550 24740 57560 24820
rect 57850 24740 57860 24820
rect 57470 24640 57550 24650
rect 57770 24640 57850 24650
rect 57550 24560 57560 24640
rect 57850 24560 57860 24640
rect 57470 24460 57550 24470
rect 57770 24460 57850 24470
rect 57550 24380 57560 24460
rect 57850 24380 57860 24460
rect 57470 24280 57550 24290
rect 57770 24280 57850 24290
rect 57550 24200 57560 24280
rect 57850 24200 57860 24280
rect 57470 24100 57550 24110
rect 57770 24100 57850 24110
rect 57550 24020 57560 24100
rect 57850 24020 57860 24100
rect 57470 23920 57550 23930
rect 57770 23920 57850 23930
rect 57550 23840 57560 23920
rect 57850 23840 57860 23920
rect 57470 23740 57550 23750
rect 57770 23740 57850 23750
rect 57550 23660 57560 23740
rect 57850 23660 57860 23740
rect 57470 23560 57550 23570
rect 57770 23560 57850 23570
rect 57550 23480 57560 23560
rect 57850 23480 57860 23560
rect 57470 23380 57550 23390
rect 57770 23380 57850 23390
rect 57550 23300 57560 23380
rect 57850 23300 57860 23380
rect 57470 23200 57550 23210
rect 57770 23200 57850 23210
rect 57550 23120 57560 23200
rect 57850 23120 57860 23200
rect 57470 23020 57550 23030
rect 57770 23020 57850 23030
rect 57550 22940 57560 23020
rect 57850 22940 57860 23020
rect 57470 22840 57550 22850
rect 57770 22840 57850 22850
rect 57550 22760 57560 22840
rect 57850 22760 57860 22840
rect 57470 22660 57550 22670
rect 57770 22660 57850 22670
rect 57550 22580 57560 22660
rect 57850 22580 57860 22660
rect 57470 22480 57550 22490
rect 57770 22480 57850 22490
rect 57550 22400 57560 22480
rect 57850 22400 57860 22480
rect 57470 22300 57550 22310
rect 57770 22300 57850 22310
rect 57550 22220 57560 22300
rect 57850 22220 57860 22300
rect 57470 22120 57550 22130
rect 57770 22120 57850 22130
rect 57550 22040 57560 22120
rect 57850 22040 57860 22120
rect 57470 21940 57550 21950
rect 57770 21940 57850 21950
rect 57550 21860 57560 21940
rect 57850 21860 57860 21940
rect 57470 21760 57550 21770
rect 57770 21760 57850 21770
rect 57550 21680 57560 21760
rect 57850 21680 57860 21760
rect 57470 21580 57550 21590
rect 57770 21580 57850 21590
rect 57550 21500 57560 21580
rect 57850 21500 57860 21580
rect 57470 21400 57550 21410
rect 57770 21400 57850 21410
rect 57550 21320 57560 21400
rect 57850 21320 57860 21400
rect 57470 21220 57550 21230
rect 57770 21220 57850 21230
rect 57550 21140 57560 21220
rect 57850 21140 57860 21220
rect 57470 21040 57550 21050
rect 57770 21040 57850 21050
rect 57550 20960 57560 21040
rect 57850 20960 57860 21040
rect 57470 20860 57550 20870
rect 57770 20860 57850 20870
rect 57550 20780 57560 20860
rect 57850 20780 57860 20860
rect 57470 20680 57550 20690
rect 57770 20680 57850 20690
rect 57550 20600 57560 20680
rect 57850 20600 57860 20680
rect 57470 20500 57550 20510
rect 57770 20500 57850 20510
rect 57550 20420 57560 20500
rect 57850 20420 57860 20500
rect 57470 20320 57550 20330
rect 57770 20320 57850 20330
rect 57550 20240 57560 20320
rect 57850 20240 57860 20320
rect 57470 20140 57550 20150
rect 57770 20140 57850 20150
rect 57550 20060 57560 20140
rect 57850 20060 57860 20140
rect 57470 19960 57550 19970
rect 57770 19960 57850 19970
rect 57550 19880 57560 19960
rect 57850 19880 57860 19960
rect 58030 19800 58040 25800
rect 58090 25720 58170 25730
rect 58240 25720 58320 25730
rect 58390 25720 58470 25730
rect 58170 25640 58180 25720
rect 58320 25640 58330 25720
rect 58470 25640 58480 25720
rect 58090 25540 58170 25550
rect 58240 25540 58320 25550
rect 58390 25540 58470 25550
rect 58170 25460 58180 25540
rect 58320 25460 58330 25540
rect 58470 25460 58480 25540
rect 58090 25360 58170 25370
rect 58240 25360 58320 25370
rect 58390 25360 58470 25370
rect 58170 25280 58180 25360
rect 58320 25280 58330 25360
rect 58470 25280 58480 25360
rect 58090 25180 58170 25190
rect 58240 25180 58320 25190
rect 58390 25180 58470 25190
rect 58170 25100 58180 25180
rect 58320 25100 58330 25180
rect 58470 25100 58480 25180
rect 58090 25000 58170 25010
rect 58240 25000 58320 25010
rect 58390 25000 58470 25010
rect 58170 24920 58180 25000
rect 58320 24920 58330 25000
rect 58470 24920 58480 25000
rect 58090 24820 58170 24830
rect 58240 24820 58320 24830
rect 58390 24820 58470 24830
rect 58170 24740 58180 24820
rect 58320 24740 58330 24820
rect 58470 24740 58480 24820
rect 58090 24640 58170 24650
rect 58240 24640 58320 24650
rect 58390 24640 58470 24650
rect 58170 24560 58180 24640
rect 58320 24560 58330 24640
rect 58470 24560 58480 24640
rect 58090 24460 58170 24470
rect 58240 24460 58320 24470
rect 58390 24460 58470 24470
rect 58170 24380 58180 24460
rect 58320 24380 58330 24460
rect 58470 24380 58480 24460
rect 58090 24280 58170 24290
rect 58240 24280 58320 24290
rect 58390 24280 58470 24290
rect 58170 24200 58180 24280
rect 58320 24200 58330 24280
rect 58470 24200 58480 24280
rect 58090 24100 58170 24110
rect 58240 24100 58320 24110
rect 58390 24100 58470 24110
rect 58170 24020 58180 24100
rect 58320 24020 58330 24100
rect 58470 24020 58480 24100
rect 58090 23920 58170 23930
rect 58240 23920 58320 23930
rect 58390 23920 58470 23930
rect 58170 23840 58180 23920
rect 58320 23840 58330 23920
rect 58470 23840 58480 23920
rect 58090 23740 58170 23750
rect 58240 23740 58320 23750
rect 58390 23740 58470 23750
rect 58170 23660 58180 23740
rect 58320 23660 58330 23740
rect 58470 23660 58480 23740
rect 58090 23560 58170 23570
rect 58240 23560 58320 23570
rect 58390 23560 58470 23570
rect 58170 23480 58180 23560
rect 58320 23480 58330 23560
rect 58470 23480 58480 23560
rect 58090 23380 58170 23390
rect 58240 23380 58320 23390
rect 58390 23380 58470 23390
rect 58170 23300 58180 23380
rect 58320 23300 58330 23380
rect 58470 23300 58480 23380
rect 58090 23200 58170 23210
rect 58240 23200 58320 23210
rect 58390 23200 58470 23210
rect 58170 23120 58180 23200
rect 58320 23120 58330 23200
rect 58470 23120 58480 23200
rect 58090 23020 58170 23030
rect 58240 23020 58320 23030
rect 58390 23020 58470 23030
rect 58170 22940 58180 23020
rect 58320 22940 58330 23020
rect 58470 22940 58480 23020
rect 58090 22840 58170 22850
rect 58240 22840 58320 22850
rect 58390 22840 58470 22850
rect 58170 22760 58180 22840
rect 58320 22760 58330 22840
rect 58470 22760 58480 22840
rect 58090 22660 58170 22670
rect 58240 22660 58320 22670
rect 58390 22660 58470 22670
rect 58170 22580 58180 22660
rect 58320 22580 58330 22660
rect 58470 22580 58480 22660
rect 58090 22480 58170 22490
rect 58240 22480 58320 22490
rect 58390 22480 58470 22490
rect 58170 22400 58180 22480
rect 58320 22400 58330 22480
rect 58470 22400 58480 22480
rect 58090 22300 58170 22310
rect 58240 22300 58320 22310
rect 58390 22300 58470 22310
rect 58170 22220 58180 22300
rect 58320 22220 58330 22300
rect 58470 22220 58480 22300
rect 58090 22120 58170 22130
rect 58240 22120 58320 22130
rect 58390 22120 58470 22130
rect 58170 22040 58180 22120
rect 58320 22040 58330 22120
rect 58470 22040 58480 22120
rect 58090 21940 58170 21950
rect 58240 21940 58320 21950
rect 58390 21940 58470 21950
rect 58170 21860 58180 21940
rect 58320 21860 58330 21940
rect 58470 21860 58480 21940
rect 58090 21760 58170 21770
rect 58240 21760 58320 21770
rect 58390 21760 58470 21770
rect 58170 21680 58180 21760
rect 58320 21680 58330 21760
rect 58470 21680 58480 21760
rect 58090 21580 58170 21590
rect 58240 21580 58320 21590
rect 58390 21580 58470 21590
rect 58170 21500 58180 21580
rect 58320 21500 58330 21580
rect 58470 21500 58480 21580
rect 58090 21400 58170 21410
rect 58240 21400 58320 21410
rect 58390 21400 58470 21410
rect 58170 21320 58180 21400
rect 58320 21320 58330 21400
rect 58470 21320 58480 21400
rect 58090 21220 58170 21230
rect 58240 21220 58320 21230
rect 58390 21220 58470 21230
rect 58170 21140 58180 21220
rect 58320 21140 58330 21220
rect 58470 21140 58480 21220
rect 58090 21040 58170 21050
rect 58240 21040 58320 21050
rect 58390 21040 58470 21050
rect 58170 20960 58180 21040
rect 58320 20960 58330 21040
rect 58470 20960 58480 21040
rect 58090 20860 58170 20870
rect 58240 20860 58320 20870
rect 58390 20860 58470 20870
rect 58170 20780 58180 20860
rect 58320 20780 58330 20860
rect 58470 20780 58480 20860
rect 58090 20680 58170 20690
rect 58240 20680 58320 20690
rect 58390 20680 58470 20690
rect 58170 20600 58180 20680
rect 58320 20600 58330 20680
rect 58470 20600 58480 20680
rect 58090 20500 58170 20510
rect 58240 20500 58320 20510
rect 58390 20500 58470 20510
rect 58170 20420 58180 20500
rect 58320 20420 58330 20500
rect 58470 20420 58480 20500
rect 58090 20320 58170 20330
rect 58240 20320 58320 20330
rect 58390 20320 58470 20330
rect 58170 20240 58180 20320
rect 58320 20240 58330 20320
rect 58470 20240 58480 20320
rect 58090 20140 58170 20150
rect 58240 20140 58320 20150
rect 58390 20140 58470 20150
rect 58170 20060 58180 20140
rect 58320 20060 58330 20140
rect 58470 20060 58480 20140
rect 58090 19960 58170 19970
rect 58240 19960 58320 19970
rect 58390 19960 58470 19970
rect 58170 19880 58180 19960
rect 58320 19880 58330 19960
rect 58470 19880 58480 19960
rect 58610 19800 58620 25800
rect 58730 25720 58810 25730
rect 59030 25720 59110 25730
rect 58810 25640 58820 25720
rect 59110 25640 59120 25720
rect 58730 25540 58810 25550
rect 59030 25540 59110 25550
rect 58810 25460 58820 25540
rect 59110 25460 59120 25540
rect 58730 25360 58810 25370
rect 59030 25360 59110 25370
rect 58810 25280 58820 25360
rect 59110 25280 59120 25360
rect 58730 25180 58810 25190
rect 59030 25180 59110 25190
rect 58810 25100 58820 25180
rect 59110 25100 59120 25180
rect 58730 25000 58810 25010
rect 59030 25000 59110 25010
rect 58810 24920 58820 25000
rect 59110 24920 59120 25000
rect 58730 24820 58810 24830
rect 59030 24820 59110 24830
rect 58810 24740 58820 24820
rect 59110 24740 59120 24820
rect 58730 24640 58810 24650
rect 59030 24640 59110 24650
rect 58810 24560 58820 24640
rect 59110 24560 59120 24640
rect 58730 24460 58810 24470
rect 59030 24460 59110 24470
rect 58810 24380 58820 24460
rect 59110 24380 59120 24460
rect 58730 24280 58810 24290
rect 59030 24280 59110 24290
rect 58810 24200 58820 24280
rect 59110 24200 59120 24280
rect 58730 24100 58810 24110
rect 59030 24100 59110 24110
rect 58810 24020 58820 24100
rect 59110 24020 59120 24100
rect 58730 23920 58810 23930
rect 59030 23920 59110 23930
rect 58810 23840 58820 23920
rect 59110 23840 59120 23920
rect 58730 23740 58810 23750
rect 59030 23740 59110 23750
rect 58810 23660 58820 23740
rect 59110 23660 59120 23740
rect 58730 23560 58810 23570
rect 59030 23560 59110 23570
rect 58810 23480 58820 23560
rect 59110 23480 59120 23560
rect 58730 23380 58810 23390
rect 59030 23380 59110 23390
rect 58810 23300 58820 23380
rect 59110 23300 59120 23380
rect 58730 23200 58810 23210
rect 59030 23200 59110 23210
rect 58810 23120 58820 23200
rect 59110 23120 59120 23200
rect 58730 23020 58810 23030
rect 59030 23020 59110 23030
rect 58810 22940 58820 23020
rect 59110 22940 59120 23020
rect 58730 22840 58810 22850
rect 59030 22840 59110 22850
rect 58810 22760 58820 22840
rect 59110 22760 59120 22840
rect 58730 22660 58810 22670
rect 59030 22660 59110 22670
rect 58810 22580 58820 22660
rect 59110 22580 59120 22660
rect 58730 22480 58810 22490
rect 59030 22480 59110 22490
rect 58810 22400 58820 22480
rect 59110 22400 59120 22480
rect 58730 22300 58810 22310
rect 59030 22300 59110 22310
rect 58810 22220 58820 22300
rect 59110 22220 59120 22300
rect 58730 22120 58810 22130
rect 59030 22120 59110 22130
rect 58810 22040 58820 22120
rect 59110 22040 59120 22120
rect 58730 21940 58810 21950
rect 59030 21940 59110 21950
rect 58810 21860 58820 21940
rect 59110 21860 59120 21940
rect 58730 21760 58810 21770
rect 59030 21760 59110 21770
rect 58810 21680 58820 21760
rect 59110 21680 59120 21760
rect 58730 21580 58810 21590
rect 59030 21580 59110 21590
rect 58810 21500 58820 21580
rect 59110 21500 59120 21580
rect 58730 21400 58810 21410
rect 59030 21400 59110 21410
rect 58810 21320 58820 21400
rect 59110 21320 59120 21400
rect 58730 21220 58810 21230
rect 59030 21220 59110 21230
rect 58810 21140 58820 21220
rect 59110 21140 59120 21220
rect 58730 21040 58810 21050
rect 59030 21040 59110 21050
rect 58810 20960 58820 21040
rect 59110 20960 59120 21040
rect 58730 20860 58810 20870
rect 59030 20860 59110 20870
rect 58810 20780 58820 20860
rect 59110 20780 59120 20860
rect 58730 20680 58810 20690
rect 59030 20680 59110 20690
rect 58810 20600 58820 20680
rect 59110 20600 59120 20680
rect 58730 20500 58810 20510
rect 59030 20500 59110 20510
rect 58810 20420 58820 20500
rect 59110 20420 59120 20500
rect 58730 20320 58810 20330
rect 59030 20320 59110 20330
rect 58810 20240 58820 20320
rect 59110 20240 59120 20320
rect 58730 20140 58810 20150
rect 59030 20140 59110 20150
rect 58810 20060 58820 20140
rect 59110 20060 59120 20140
rect 58730 19960 58810 19970
rect 59030 19960 59110 19970
rect 58810 19880 58820 19960
rect 59110 19880 59120 19960
rect 59290 19800 59300 25800
rect 60610 25770 60690 25780
rect 60930 25770 61010 25780
rect 61350 25770 61430 25780
rect 61670 25770 61750 25780
rect 74110 25770 74190 25780
rect 74430 25770 74510 25780
rect 74850 25770 74930 25780
rect 75170 25770 75250 25780
rect 87610 25770 87690 25780
rect 87930 25770 88010 25780
rect 88350 25770 88430 25780
rect 88670 25770 88750 25780
rect 101110 25770 101190 25780
rect 101430 25770 101510 25780
rect 101850 25770 101930 25780
rect 102170 25770 102250 25780
rect 114610 25770 114690 25780
rect 114930 25770 115010 25780
rect 115350 25770 115430 25780
rect 115670 25770 115750 25780
rect 128110 25770 128190 25780
rect 128430 25770 128510 25780
rect 128850 25770 128930 25780
rect 129170 25770 129250 25780
rect 59350 25720 59430 25730
rect 59500 25720 59580 25730
rect 59650 25720 59730 25730
rect 60060 25720 60140 25730
rect 60210 25720 60290 25730
rect 60360 25720 60440 25730
rect 59430 25640 59440 25720
rect 59580 25640 59590 25720
rect 59730 25640 59740 25720
rect 60140 25640 60150 25720
rect 60290 25640 60300 25720
rect 60440 25640 60450 25720
rect 60690 25690 60700 25770
rect 61010 25690 61020 25770
rect 61430 25690 61440 25770
rect 61750 25690 61760 25770
rect 62060 25720 62140 25730
rect 62210 25720 62290 25730
rect 73560 25720 73640 25730
rect 73710 25720 73790 25730
rect 73860 25720 73940 25730
rect 62140 25640 62150 25720
rect 62290 25640 62300 25720
rect 73640 25640 73650 25720
rect 73790 25640 73800 25720
rect 73940 25640 73950 25720
rect 74190 25690 74200 25770
rect 74510 25690 74520 25770
rect 74930 25690 74940 25770
rect 75250 25690 75260 25770
rect 75560 25720 75640 25730
rect 75710 25720 75790 25730
rect 87060 25720 87140 25730
rect 87210 25720 87290 25730
rect 87360 25720 87440 25730
rect 75640 25640 75650 25720
rect 75790 25640 75800 25720
rect 87140 25640 87150 25720
rect 87290 25640 87300 25720
rect 87440 25640 87450 25720
rect 87690 25690 87700 25770
rect 88010 25690 88020 25770
rect 88430 25690 88440 25770
rect 88750 25690 88760 25770
rect 89060 25720 89140 25730
rect 89210 25720 89290 25730
rect 100560 25720 100640 25730
rect 100710 25720 100790 25730
rect 100860 25720 100940 25730
rect 89140 25640 89150 25720
rect 89290 25640 89300 25720
rect 100640 25640 100650 25720
rect 100790 25640 100800 25720
rect 100940 25640 100950 25720
rect 101190 25690 101200 25770
rect 101510 25690 101520 25770
rect 101930 25690 101940 25770
rect 102250 25690 102260 25770
rect 102560 25720 102640 25730
rect 102710 25720 102790 25730
rect 114060 25720 114140 25730
rect 114210 25720 114290 25730
rect 114360 25720 114440 25730
rect 102640 25640 102650 25720
rect 102790 25640 102800 25720
rect 114140 25640 114150 25720
rect 114290 25640 114300 25720
rect 114440 25640 114450 25720
rect 114690 25690 114700 25770
rect 115010 25690 115020 25770
rect 115430 25690 115440 25770
rect 115750 25690 115760 25770
rect 116060 25720 116140 25730
rect 116210 25720 116290 25730
rect 127560 25720 127640 25730
rect 127710 25720 127790 25730
rect 127860 25720 127940 25730
rect 116140 25640 116150 25720
rect 116290 25640 116300 25720
rect 127640 25640 127650 25720
rect 127790 25640 127800 25720
rect 127940 25640 127950 25720
rect 128190 25690 128200 25770
rect 128510 25690 128520 25770
rect 128930 25690 128940 25770
rect 129250 25690 129260 25770
rect 129560 25720 129640 25730
rect 129710 25720 129790 25730
rect 141060 25720 141140 25730
rect 141210 25720 141290 25730
rect 141360 25720 141440 25730
rect 129640 25640 129650 25720
rect 129790 25640 129800 25720
rect 141140 25640 141150 25720
rect 141290 25640 141300 25720
rect 141440 25640 141450 25720
rect 60770 25610 60850 25620
rect 61090 25610 61170 25620
rect 61510 25610 61590 25620
rect 61830 25610 61910 25620
rect 74270 25610 74350 25620
rect 74590 25610 74670 25620
rect 75010 25610 75090 25620
rect 75330 25610 75410 25620
rect 87770 25610 87850 25620
rect 88090 25610 88170 25620
rect 88510 25610 88590 25620
rect 88830 25610 88910 25620
rect 101270 25610 101350 25620
rect 101590 25610 101670 25620
rect 102010 25610 102090 25620
rect 102330 25610 102410 25620
rect 114770 25610 114850 25620
rect 115090 25610 115170 25620
rect 115510 25610 115590 25620
rect 115830 25610 115910 25620
rect 128270 25610 128350 25620
rect 128590 25610 128670 25620
rect 129010 25610 129090 25620
rect 129330 25610 129410 25620
rect 59350 25540 59430 25550
rect 59500 25540 59580 25550
rect 59650 25540 59730 25550
rect 60060 25540 60140 25550
rect 60210 25540 60290 25550
rect 60360 25540 60440 25550
rect 59430 25460 59440 25540
rect 59580 25460 59590 25540
rect 59730 25460 59740 25540
rect 60140 25460 60150 25540
rect 60290 25460 60300 25540
rect 60440 25460 60450 25540
rect 60850 25530 60860 25610
rect 61170 25530 61180 25610
rect 61590 25530 61600 25610
rect 61910 25530 61920 25610
rect 62060 25540 62140 25550
rect 62210 25540 62290 25550
rect 73560 25540 73640 25550
rect 73710 25540 73790 25550
rect 73860 25540 73940 25550
rect 62140 25460 62150 25540
rect 62290 25460 62300 25540
rect 73640 25460 73650 25540
rect 73790 25460 73800 25540
rect 73940 25460 73950 25540
rect 74350 25530 74360 25610
rect 74670 25530 74680 25610
rect 75090 25530 75100 25610
rect 75410 25530 75420 25610
rect 75560 25540 75640 25550
rect 75710 25540 75790 25550
rect 87060 25540 87140 25550
rect 87210 25540 87290 25550
rect 87360 25540 87440 25550
rect 75640 25460 75650 25540
rect 75790 25460 75800 25540
rect 87140 25460 87150 25540
rect 87290 25460 87300 25540
rect 87440 25460 87450 25540
rect 87850 25530 87860 25610
rect 88170 25530 88180 25610
rect 88590 25530 88600 25610
rect 88910 25530 88920 25610
rect 89060 25540 89140 25550
rect 89210 25540 89290 25550
rect 100560 25540 100640 25550
rect 100710 25540 100790 25550
rect 100860 25540 100940 25550
rect 89140 25460 89150 25540
rect 89290 25460 89300 25540
rect 100640 25460 100650 25540
rect 100790 25460 100800 25540
rect 100940 25460 100950 25540
rect 101350 25530 101360 25610
rect 101670 25530 101680 25610
rect 102090 25530 102100 25610
rect 102410 25530 102420 25610
rect 102560 25540 102640 25550
rect 102710 25540 102790 25550
rect 114060 25540 114140 25550
rect 114210 25540 114290 25550
rect 114360 25540 114440 25550
rect 102640 25460 102650 25540
rect 102790 25460 102800 25540
rect 114140 25460 114150 25540
rect 114290 25460 114300 25540
rect 114440 25460 114450 25540
rect 114850 25530 114860 25610
rect 115170 25530 115180 25610
rect 115590 25530 115600 25610
rect 115910 25530 115920 25610
rect 116060 25540 116140 25550
rect 116210 25540 116290 25550
rect 127560 25540 127640 25550
rect 127710 25540 127790 25550
rect 127860 25540 127940 25550
rect 116140 25460 116150 25540
rect 116290 25460 116300 25540
rect 127640 25460 127650 25540
rect 127790 25460 127800 25540
rect 127940 25460 127950 25540
rect 128350 25530 128360 25610
rect 128670 25530 128680 25610
rect 129090 25530 129100 25610
rect 129410 25530 129420 25610
rect 129560 25540 129640 25550
rect 129710 25540 129790 25550
rect 141060 25540 141140 25550
rect 141210 25540 141290 25550
rect 141360 25540 141440 25550
rect 129640 25460 129650 25540
rect 129790 25460 129800 25540
rect 141140 25460 141150 25540
rect 141290 25460 141300 25540
rect 141440 25460 141450 25540
rect 60610 25450 60690 25460
rect 60930 25450 61010 25460
rect 61350 25450 61430 25460
rect 61670 25450 61750 25460
rect 74110 25450 74190 25460
rect 74430 25450 74510 25460
rect 74850 25450 74930 25460
rect 75170 25450 75250 25460
rect 87610 25450 87690 25460
rect 87930 25450 88010 25460
rect 88350 25450 88430 25460
rect 88670 25450 88750 25460
rect 101110 25450 101190 25460
rect 101430 25450 101510 25460
rect 101850 25450 101930 25460
rect 102170 25450 102250 25460
rect 114610 25450 114690 25460
rect 114930 25450 115010 25460
rect 115350 25450 115430 25460
rect 115670 25450 115750 25460
rect 128110 25450 128190 25460
rect 128430 25450 128510 25460
rect 128850 25450 128930 25460
rect 129170 25450 129250 25460
rect 60690 25370 60700 25450
rect 61010 25370 61020 25450
rect 61430 25370 61440 25450
rect 61750 25370 61760 25450
rect 74190 25370 74200 25450
rect 74510 25370 74520 25450
rect 74930 25370 74940 25450
rect 75250 25370 75260 25450
rect 87690 25370 87700 25450
rect 88010 25370 88020 25450
rect 88430 25370 88440 25450
rect 88750 25370 88760 25450
rect 101190 25370 101200 25450
rect 101510 25370 101520 25450
rect 101930 25370 101940 25450
rect 102250 25370 102260 25450
rect 114690 25370 114700 25450
rect 115010 25370 115020 25450
rect 115430 25370 115440 25450
rect 115750 25370 115760 25450
rect 128190 25370 128200 25450
rect 128510 25370 128520 25450
rect 128930 25370 128940 25450
rect 129250 25370 129260 25450
rect 59350 25360 59430 25370
rect 59500 25360 59580 25370
rect 59650 25360 59730 25370
rect 60060 25360 60140 25370
rect 60210 25360 60290 25370
rect 60360 25360 60440 25370
rect 62060 25360 62140 25370
rect 62210 25360 62290 25370
rect 73560 25360 73640 25370
rect 73710 25360 73790 25370
rect 73860 25360 73940 25370
rect 75560 25360 75640 25370
rect 75710 25360 75790 25370
rect 87060 25360 87140 25370
rect 87210 25360 87290 25370
rect 87360 25360 87440 25370
rect 89060 25360 89140 25370
rect 89210 25360 89290 25370
rect 100560 25360 100640 25370
rect 100710 25360 100790 25370
rect 100860 25360 100940 25370
rect 102560 25360 102640 25370
rect 102710 25360 102790 25370
rect 114060 25360 114140 25370
rect 114210 25360 114290 25370
rect 114360 25360 114440 25370
rect 116060 25360 116140 25370
rect 116210 25360 116290 25370
rect 127560 25360 127640 25370
rect 127710 25360 127790 25370
rect 127860 25360 127940 25370
rect 129560 25360 129640 25370
rect 129710 25360 129790 25370
rect 141060 25360 141140 25370
rect 141210 25360 141290 25370
rect 141360 25360 141440 25370
rect 59430 25280 59440 25360
rect 59580 25280 59590 25360
rect 59730 25280 59740 25360
rect 60140 25280 60150 25360
rect 60290 25280 60300 25360
rect 60440 25280 60450 25360
rect 60770 25290 60850 25300
rect 61090 25290 61170 25300
rect 61510 25290 61590 25300
rect 61830 25290 61910 25300
rect 60850 25210 60860 25290
rect 61170 25210 61180 25290
rect 61590 25210 61600 25290
rect 61910 25210 61920 25290
rect 62140 25280 62150 25360
rect 62290 25280 62300 25360
rect 73640 25280 73650 25360
rect 73790 25280 73800 25360
rect 73940 25280 73950 25360
rect 74270 25290 74350 25300
rect 74590 25290 74670 25300
rect 75010 25290 75090 25300
rect 75330 25290 75410 25300
rect 74350 25210 74360 25290
rect 74670 25210 74680 25290
rect 75090 25210 75100 25290
rect 75410 25210 75420 25290
rect 75640 25280 75650 25360
rect 75790 25280 75800 25360
rect 87140 25280 87150 25360
rect 87290 25280 87300 25360
rect 87440 25280 87450 25360
rect 87770 25290 87850 25300
rect 88090 25290 88170 25300
rect 88510 25290 88590 25300
rect 88830 25290 88910 25300
rect 87850 25210 87860 25290
rect 88170 25210 88180 25290
rect 88590 25210 88600 25290
rect 88910 25210 88920 25290
rect 89140 25280 89150 25360
rect 89290 25280 89300 25360
rect 100640 25280 100650 25360
rect 100790 25280 100800 25360
rect 100940 25280 100950 25360
rect 101270 25290 101350 25300
rect 101590 25290 101670 25300
rect 102010 25290 102090 25300
rect 102330 25290 102410 25300
rect 101350 25210 101360 25290
rect 101670 25210 101680 25290
rect 102090 25210 102100 25290
rect 102410 25210 102420 25290
rect 102640 25280 102650 25360
rect 102790 25280 102800 25360
rect 114140 25280 114150 25360
rect 114290 25280 114300 25360
rect 114440 25280 114450 25360
rect 114770 25290 114850 25300
rect 115090 25290 115170 25300
rect 115510 25290 115590 25300
rect 115830 25290 115910 25300
rect 114850 25210 114860 25290
rect 115170 25210 115180 25290
rect 115590 25210 115600 25290
rect 115910 25210 115920 25290
rect 116140 25280 116150 25360
rect 116290 25280 116300 25360
rect 127640 25280 127650 25360
rect 127790 25280 127800 25360
rect 127940 25280 127950 25360
rect 128270 25290 128350 25300
rect 128590 25290 128670 25300
rect 129010 25290 129090 25300
rect 129330 25290 129410 25300
rect 128350 25210 128360 25290
rect 128670 25210 128680 25290
rect 129090 25210 129100 25290
rect 129410 25210 129420 25290
rect 129640 25280 129650 25360
rect 129790 25280 129800 25360
rect 141140 25280 141150 25360
rect 141290 25280 141300 25360
rect 141440 25280 141450 25360
rect 59350 25180 59430 25190
rect 59500 25180 59580 25190
rect 59650 25180 59730 25190
rect 60060 25180 60140 25190
rect 60210 25180 60290 25190
rect 60360 25180 60440 25190
rect 62060 25180 62140 25190
rect 62210 25180 62290 25190
rect 73560 25180 73640 25190
rect 73710 25180 73790 25190
rect 73860 25180 73940 25190
rect 75560 25180 75640 25190
rect 75710 25180 75790 25190
rect 87060 25180 87140 25190
rect 87210 25180 87290 25190
rect 87360 25180 87440 25190
rect 89060 25180 89140 25190
rect 89210 25180 89290 25190
rect 100560 25180 100640 25190
rect 100710 25180 100790 25190
rect 100860 25180 100940 25190
rect 102560 25180 102640 25190
rect 102710 25180 102790 25190
rect 114060 25180 114140 25190
rect 114210 25180 114290 25190
rect 114360 25180 114440 25190
rect 116060 25180 116140 25190
rect 116210 25180 116290 25190
rect 127560 25180 127640 25190
rect 127710 25180 127790 25190
rect 127860 25180 127940 25190
rect 129560 25180 129640 25190
rect 129710 25180 129790 25190
rect 141060 25180 141140 25190
rect 141210 25180 141290 25190
rect 141360 25180 141440 25190
rect 59430 25100 59440 25180
rect 59580 25100 59590 25180
rect 59730 25100 59740 25180
rect 60140 25100 60150 25180
rect 60290 25100 60300 25180
rect 60440 25100 60450 25180
rect 60610 25130 60690 25140
rect 60930 25130 61010 25140
rect 61350 25130 61430 25140
rect 61670 25130 61750 25140
rect 60690 25050 60700 25130
rect 61010 25050 61020 25130
rect 61430 25050 61440 25130
rect 61750 25050 61760 25130
rect 62140 25100 62150 25180
rect 62290 25100 62300 25180
rect 73640 25100 73650 25180
rect 73790 25100 73800 25180
rect 73940 25100 73950 25180
rect 74110 25130 74190 25140
rect 74430 25130 74510 25140
rect 74850 25130 74930 25140
rect 75170 25130 75250 25140
rect 74190 25050 74200 25130
rect 74510 25050 74520 25130
rect 74930 25050 74940 25130
rect 75250 25050 75260 25130
rect 75640 25100 75650 25180
rect 75790 25100 75800 25180
rect 87140 25100 87150 25180
rect 87290 25100 87300 25180
rect 87440 25100 87450 25180
rect 87610 25130 87690 25140
rect 87930 25130 88010 25140
rect 88350 25130 88430 25140
rect 88670 25130 88750 25140
rect 87690 25050 87700 25130
rect 88010 25050 88020 25130
rect 88430 25050 88440 25130
rect 88750 25050 88760 25130
rect 89140 25100 89150 25180
rect 89290 25100 89300 25180
rect 100640 25100 100650 25180
rect 100790 25100 100800 25180
rect 100940 25100 100950 25180
rect 101110 25130 101190 25140
rect 101430 25130 101510 25140
rect 101850 25130 101930 25140
rect 102170 25130 102250 25140
rect 101190 25050 101200 25130
rect 101510 25050 101520 25130
rect 101930 25050 101940 25130
rect 102250 25050 102260 25130
rect 102640 25100 102650 25180
rect 102790 25100 102800 25180
rect 114140 25100 114150 25180
rect 114290 25100 114300 25180
rect 114440 25100 114450 25180
rect 114610 25130 114690 25140
rect 114930 25130 115010 25140
rect 115350 25130 115430 25140
rect 115670 25130 115750 25140
rect 114690 25050 114700 25130
rect 115010 25050 115020 25130
rect 115430 25050 115440 25130
rect 115750 25050 115760 25130
rect 116140 25100 116150 25180
rect 116290 25100 116300 25180
rect 127640 25100 127650 25180
rect 127790 25100 127800 25180
rect 127940 25100 127950 25180
rect 128110 25130 128190 25140
rect 128430 25130 128510 25140
rect 128850 25130 128930 25140
rect 129170 25130 129250 25140
rect 128190 25050 128200 25130
rect 128510 25050 128520 25130
rect 128930 25050 128940 25130
rect 129250 25050 129260 25130
rect 129640 25100 129650 25180
rect 129790 25100 129800 25180
rect 141140 25100 141150 25180
rect 141290 25100 141300 25180
rect 141440 25100 141450 25180
rect 59350 25000 59430 25010
rect 59500 25000 59580 25010
rect 59650 25000 59730 25010
rect 60060 25000 60140 25010
rect 60210 25000 60290 25010
rect 60360 25000 60440 25010
rect 62060 25000 62140 25010
rect 62210 25000 62290 25010
rect 73560 25000 73640 25010
rect 73710 25000 73790 25010
rect 73860 25000 73940 25010
rect 75560 25000 75640 25010
rect 75710 25000 75790 25010
rect 87060 25000 87140 25010
rect 87210 25000 87290 25010
rect 87360 25000 87440 25010
rect 89060 25000 89140 25010
rect 89210 25000 89290 25010
rect 100560 25000 100640 25010
rect 100710 25000 100790 25010
rect 100860 25000 100940 25010
rect 102560 25000 102640 25010
rect 102710 25000 102790 25010
rect 114060 25000 114140 25010
rect 114210 25000 114290 25010
rect 114360 25000 114440 25010
rect 116060 25000 116140 25010
rect 116210 25000 116290 25010
rect 127560 25000 127640 25010
rect 127710 25000 127790 25010
rect 127860 25000 127940 25010
rect 129560 25000 129640 25010
rect 129710 25000 129790 25010
rect 141060 25000 141140 25010
rect 141210 25000 141290 25010
rect 141360 25000 141440 25010
rect 59430 24920 59440 25000
rect 59580 24920 59590 25000
rect 59730 24920 59740 25000
rect 60140 24920 60150 25000
rect 60290 24920 60300 25000
rect 60440 24920 60450 25000
rect 60770 24970 60850 24980
rect 61090 24970 61170 24980
rect 61510 24970 61590 24980
rect 61830 24970 61910 24980
rect 60850 24890 60860 24970
rect 61170 24890 61180 24970
rect 61590 24890 61600 24970
rect 61910 24890 61920 24970
rect 62140 24920 62150 25000
rect 62290 24920 62300 25000
rect 73640 24920 73650 25000
rect 73790 24920 73800 25000
rect 73940 24920 73950 25000
rect 74270 24970 74350 24980
rect 74590 24970 74670 24980
rect 75010 24970 75090 24980
rect 75330 24970 75410 24980
rect 74350 24890 74360 24970
rect 74670 24890 74680 24970
rect 75090 24890 75100 24970
rect 75410 24890 75420 24970
rect 75640 24920 75650 25000
rect 75790 24920 75800 25000
rect 87140 24920 87150 25000
rect 87290 24920 87300 25000
rect 87440 24920 87450 25000
rect 87770 24970 87850 24980
rect 88090 24970 88170 24980
rect 88510 24970 88590 24980
rect 88830 24970 88910 24980
rect 87850 24890 87860 24970
rect 88170 24890 88180 24970
rect 88590 24890 88600 24970
rect 88910 24890 88920 24970
rect 89140 24920 89150 25000
rect 89290 24920 89300 25000
rect 100640 24920 100650 25000
rect 100790 24920 100800 25000
rect 100940 24920 100950 25000
rect 101270 24970 101350 24980
rect 101590 24970 101670 24980
rect 102010 24970 102090 24980
rect 102330 24970 102410 24980
rect 101350 24890 101360 24970
rect 101670 24890 101680 24970
rect 102090 24890 102100 24970
rect 102410 24890 102420 24970
rect 102640 24920 102650 25000
rect 102790 24920 102800 25000
rect 114140 24920 114150 25000
rect 114290 24920 114300 25000
rect 114440 24920 114450 25000
rect 114770 24970 114850 24980
rect 115090 24970 115170 24980
rect 115510 24970 115590 24980
rect 115830 24970 115910 24980
rect 114850 24890 114860 24970
rect 115170 24890 115180 24970
rect 115590 24890 115600 24970
rect 115910 24890 115920 24970
rect 116140 24920 116150 25000
rect 116290 24920 116300 25000
rect 127640 24920 127650 25000
rect 127790 24920 127800 25000
rect 127940 24920 127950 25000
rect 128270 24970 128350 24980
rect 128590 24970 128670 24980
rect 129010 24970 129090 24980
rect 129330 24970 129410 24980
rect 128350 24890 128360 24970
rect 128670 24890 128680 24970
rect 129090 24890 129100 24970
rect 129410 24890 129420 24970
rect 129640 24920 129650 25000
rect 129790 24920 129800 25000
rect 141140 24920 141150 25000
rect 141290 24920 141300 25000
rect 141440 24920 141450 25000
rect 59350 24820 59430 24830
rect 59500 24820 59580 24830
rect 59650 24820 59730 24830
rect 60060 24820 60140 24830
rect 60210 24820 60290 24830
rect 60360 24820 60440 24830
rect 62060 24820 62140 24830
rect 62210 24820 62290 24830
rect 73560 24820 73640 24830
rect 73710 24820 73790 24830
rect 73860 24820 73940 24830
rect 75560 24820 75640 24830
rect 75710 24820 75790 24830
rect 87060 24820 87140 24830
rect 87210 24820 87290 24830
rect 87360 24820 87440 24830
rect 89060 24820 89140 24830
rect 89210 24820 89290 24830
rect 100560 24820 100640 24830
rect 100710 24820 100790 24830
rect 100860 24820 100940 24830
rect 102560 24820 102640 24830
rect 102710 24820 102790 24830
rect 114060 24820 114140 24830
rect 114210 24820 114290 24830
rect 114360 24820 114440 24830
rect 116060 24820 116140 24830
rect 116210 24820 116290 24830
rect 127560 24820 127640 24830
rect 127710 24820 127790 24830
rect 127860 24820 127940 24830
rect 129560 24820 129640 24830
rect 129710 24820 129790 24830
rect 141060 24820 141140 24830
rect 141210 24820 141290 24830
rect 141360 24820 141440 24830
rect 59430 24740 59440 24820
rect 59580 24740 59590 24820
rect 59730 24740 59740 24820
rect 60140 24740 60150 24820
rect 60290 24740 60300 24820
rect 60440 24740 60450 24820
rect 60610 24810 60690 24820
rect 60930 24810 61010 24820
rect 61350 24810 61430 24820
rect 61670 24810 61750 24820
rect 60690 24730 60700 24810
rect 61010 24730 61020 24810
rect 61430 24730 61440 24810
rect 61750 24730 61760 24810
rect 62140 24740 62150 24820
rect 62290 24740 62300 24820
rect 73640 24740 73650 24820
rect 73790 24740 73800 24820
rect 73940 24740 73950 24820
rect 74110 24810 74190 24820
rect 74430 24810 74510 24820
rect 74850 24810 74930 24820
rect 75170 24810 75250 24820
rect 74190 24730 74200 24810
rect 74510 24730 74520 24810
rect 74930 24730 74940 24810
rect 75250 24730 75260 24810
rect 75640 24740 75650 24820
rect 75790 24740 75800 24820
rect 87140 24740 87150 24820
rect 87290 24740 87300 24820
rect 87440 24740 87450 24820
rect 87610 24810 87690 24820
rect 87930 24810 88010 24820
rect 88350 24810 88430 24820
rect 88670 24810 88750 24820
rect 87690 24730 87700 24810
rect 88010 24730 88020 24810
rect 88430 24730 88440 24810
rect 88750 24730 88760 24810
rect 89140 24740 89150 24820
rect 89290 24740 89300 24820
rect 100640 24740 100650 24820
rect 100790 24740 100800 24820
rect 100940 24740 100950 24820
rect 101110 24810 101190 24820
rect 101430 24810 101510 24820
rect 101850 24810 101930 24820
rect 102170 24810 102250 24820
rect 101190 24730 101200 24810
rect 101510 24730 101520 24810
rect 101930 24730 101940 24810
rect 102250 24730 102260 24810
rect 102640 24740 102650 24820
rect 102790 24740 102800 24820
rect 114140 24740 114150 24820
rect 114290 24740 114300 24820
rect 114440 24740 114450 24820
rect 114610 24810 114690 24820
rect 114930 24810 115010 24820
rect 115350 24810 115430 24820
rect 115670 24810 115750 24820
rect 114690 24730 114700 24810
rect 115010 24730 115020 24810
rect 115430 24730 115440 24810
rect 115750 24730 115760 24810
rect 116140 24740 116150 24820
rect 116290 24740 116300 24820
rect 127640 24740 127650 24820
rect 127790 24740 127800 24820
rect 127940 24740 127950 24820
rect 128110 24810 128190 24820
rect 128430 24810 128510 24820
rect 128850 24810 128930 24820
rect 129170 24810 129250 24820
rect 128190 24730 128200 24810
rect 128510 24730 128520 24810
rect 128930 24730 128940 24810
rect 129250 24730 129260 24810
rect 129640 24740 129650 24820
rect 129790 24740 129800 24820
rect 141140 24740 141150 24820
rect 141290 24740 141300 24820
rect 141440 24740 141450 24820
rect 60770 24650 60850 24660
rect 61090 24650 61170 24660
rect 61510 24650 61590 24660
rect 61830 24650 61910 24660
rect 74270 24650 74350 24660
rect 74590 24650 74670 24660
rect 75010 24650 75090 24660
rect 75330 24650 75410 24660
rect 87770 24650 87850 24660
rect 88090 24650 88170 24660
rect 88510 24650 88590 24660
rect 88830 24650 88910 24660
rect 101270 24650 101350 24660
rect 101590 24650 101670 24660
rect 102010 24650 102090 24660
rect 102330 24650 102410 24660
rect 114770 24650 114850 24660
rect 115090 24650 115170 24660
rect 115510 24650 115590 24660
rect 115830 24650 115910 24660
rect 128270 24650 128350 24660
rect 128590 24650 128670 24660
rect 129010 24650 129090 24660
rect 129330 24650 129410 24660
rect 59350 24640 59430 24650
rect 59500 24640 59580 24650
rect 59650 24640 59730 24650
rect 60060 24640 60140 24650
rect 60210 24640 60290 24650
rect 60360 24640 60440 24650
rect 59430 24560 59440 24640
rect 59580 24560 59590 24640
rect 59730 24560 59740 24640
rect 60140 24560 60150 24640
rect 60290 24560 60300 24640
rect 60440 24560 60450 24640
rect 60850 24570 60860 24650
rect 61170 24570 61180 24650
rect 61590 24570 61600 24650
rect 61910 24570 61920 24650
rect 62060 24640 62140 24650
rect 62210 24640 62290 24650
rect 73560 24640 73640 24650
rect 73710 24640 73790 24650
rect 73860 24640 73940 24650
rect 62140 24560 62150 24640
rect 62290 24560 62300 24640
rect 73640 24560 73650 24640
rect 73790 24560 73800 24640
rect 73940 24560 73950 24640
rect 74350 24570 74360 24650
rect 74670 24570 74680 24650
rect 75090 24570 75100 24650
rect 75410 24570 75420 24650
rect 75560 24640 75640 24650
rect 75710 24640 75790 24650
rect 87060 24640 87140 24650
rect 87210 24640 87290 24650
rect 87360 24640 87440 24650
rect 75640 24560 75650 24640
rect 75790 24560 75800 24640
rect 87140 24560 87150 24640
rect 87290 24560 87300 24640
rect 87440 24560 87450 24640
rect 87850 24570 87860 24650
rect 88170 24570 88180 24650
rect 88590 24570 88600 24650
rect 88910 24570 88920 24650
rect 89060 24640 89140 24650
rect 89210 24640 89290 24650
rect 100560 24640 100640 24650
rect 100710 24640 100790 24650
rect 100860 24640 100940 24650
rect 89140 24560 89150 24640
rect 89290 24560 89300 24640
rect 100640 24560 100650 24640
rect 100790 24560 100800 24640
rect 100940 24560 100950 24640
rect 101350 24570 101360 24650
rect 101670 24570 101680 24650
rect 102090 24570 102100 24650
rect 102410 24570 102420 24650
rect 102560 24640 102640 24650
rect 102710 24640 102790 24650
rect 114060 24640 114140 24650
rect 114210 24640 114290 24650
rect 114360 24640 114440 24650
rect 102640 24560 102650 24640
rect 102790 24560 102800 24640
rect 114140 24560 114150 24640
rect 114290 24560 114300 24640
rect 114440 24560 114450 24640
rect 114850 24570 114860 24650
rect 115170 24570 115180 24650
rect 115590 24570 115600 24650
rect 115910 24570 115920 24650
rect 116060 24640 116140 24650
rect 116210 24640 116290 24650
rect 127560 24640 127640 24650
rect 127710 24640 127790 24650
rect 127860 24640 127940 24650
rect 116140 24560 116150 24640
rect 116290 24560 116300 24640
rect 127640 24560 127650 24640
rect 127790 24560 127800 24640
rect 127940 24560 127950 24640
rect 128350 24570 128360 24650
rect 128670 24570 128680 24650
rect 129090 24570 129100 24650
rect 129410 24570 129420 24650
rect 129560 24640 129640 24650
rect 129710 24640 129790 24650
rect 141060 24640 141140 24650
rect 141210 24640 141290 24650
rect 141360 24640 141440 24650
rect 129640 24560 129650 24640
rect 129790 24560 129800 24640
rect 141140 24560 141150 24640
rect 141290 24560 141300 24640
rect 141440 24560 141450 24640
rect 60610 24490 60690 24500
rect 60930 24490 61010 24500
rect 61350 24490 61430 24500
rect 61670 24490 61750 24500
rect 74110 24490 74190 24500
rect 74430 24490 74510 24500
rect 74850 24490 74930 24500
rect 75170 24490 75250 24500
rect 87610 24490 87690 24500
rect 87930 24490 88010 24500
rect 88350 24490 88430 24500
rect 88670 24490 88750 24500
rect 101110 24490 101190 24500
rect 101430 24490 101510 24500
rect 101850 24490 101930 24500
rect 102170 24490 102250 24500
rect 114610 24490 114690 24500
rect 114930 24490 115010 24500
rect 115350 24490 115430 24500
rect 115670 24490 115750 24500
rect 128110 24490 128190 24500
rect 128430 24490 128510 24500
rect 128850 24490 128930 24500
rect 129170 24490 129250 24500
rect 59350 24460 59430 24470
rect 59500 24460 59580 24470
rect 59650 24460 59730 24470
rect 60060 24460 60140 24470
rect 60210 24460 60290 24470
rect 60360 24460 60440 24470
rect 59430 24380 59440 24460
rect 59580 24380 59590 24460
rect 59730 24380 59740 24460
rect 60140 24380 60150 24460
rect 60290 24380 60300 24460
rect 60440 24380 60450 24460
rect 60690 24410 60700 24490
rect 61010 24410 61020 24490
rect 61430 24410 61440 24490
rect 61750 24410 61760 24490
rect 62060 24460 62140 24470
rect 62210 24460 62290 24470
rect 73560 24460 73640 24470
rect 73710 24460 73790 24470
rect 73860 24460 73940 24470
rect 62140 24380 62150 24460
rect 62290 24380 62300 24460
rect 73640 24380 73650 24460
rect 73790 24380 73800 24460
rect 73940 24380 73950 24460
rect 74190 24410 74200 24490
rect 74510 24410 74520 24490
rect 74930 24410 74940 24490
rect 75250 24410 75260 24490
rect 75560 24460 75640 24470
rect 75710 24460 75790 24470
rect 87060 24460 87140 24470
rect 87210 24460 87290 24470
rect 87360 24460 87440 24470
rect 75640 24380 75650 24460
rect 75790 24380 75800 24460
rect 87140 24380 87150 24460
rect 87290 24380 87300 24460
rect 87440 24380 87450 24460
rect 87690 24410 87700 24490
rect 88010 24410 88020 24490
rect 88430 24410 88440 24490
rect 88750 24410 88760 24490
rect 89060 24460 89140 24470
rect 89210 24460 89290 24470
rect 100560 24460 100640 24470
rect 100710 24460 100790 24470
rect 100860 24460 100940 24470
rect 89140 24380 89150 24460
rect 89290 24380 89300 24460
rect 100640 24380 100650 24460
rect 100790 24380 100800 24460
rect 100940 24380 100950 24460
rect 101190 24410 101200 24490
rect 101510 24410 101520 24490
rect 101930 24410 101940 24490
rect 102250 24410 102260 24490
rect 102560 24460 102640 24470
rect 102710 24460 102790 24470
rect 114060 24460 114140 24470
rect 114210 24460 114290 24470
rect 114360 24460 114440 24470
rect 102640 24380 102650 24460
rect 102790 24380 102800 24460
rect 114140 24380 114150 24460
rect 114290 24380 114300 24460
rect 114440 24380 114450 24460
rect 114690 24410 114700 24490
rect 115010 24410 115020 24490
rect 115430 24410 115440 24490
rect 115750 24410 115760 24490
rect 116060 24460 116140 24470
rect 116210 24460 116290 24470
rect 127560 24460 127640 24470
rect 127710 24460 127790 24470
rect 127860 24460 127940 24470
rect 116140 24380 116150 24460
rect 116290 24380 116300 24460
rect 127640 24380 127650 24460
rect 127790 24380 127800 24460
rect 127940 24380 127950 24460
rect 128190 24410 128200 24490
rect 128510 24410 128520 24490
rect 128930 24410 128940 24490
rect 129250 24410 129260 24490
rect 129560 24460 129640 24470
rect 129710 24460 129790 24470
rect 141060 24460 141140 24470
rect 141210 24460 141290 24470
rect 141360 24460 141440 24470
rect 129640 24380 129650 24460
rect 129790 24380 129800 24460
rect 141140 24380 141150 24460
rect 141290 24380 141300 24460
rect 141440 24380 141450 24460
rect 60770 24330 60850 24340
rect 61090 24330 61170 24340
rect 61510 24330 61590 24340
rect 61830 24330 61910 24340
rect 74270 24330 74350 24340
rect 74590 24330 74670 24340
rect 75010 24330 75090 24340
rect 75330 24330 75410 24340
rect 87770 24330 87850 24340
rect 88090 24330 88170 24340
rect 88510 24330 88590 24340
rect 88830 24330 88910 24340
rect 101270 24330 101350 24340
rect 101590 24330 101670 24340
rect 102010 24330 102090 24340
rect 102330 24330 102410 24340
rect 114770 24330 114850 24340
rect 115090 24330 115170 24340
rect 115510 24330 115590 24340
rect 115830 24330 115910 24340
rect 128270 24330 128350 24340
rect 128590 24330 128670 24340
rect 129010 24330 129090 24340
rect 129330 24330 129410 24340
rect 59350 24280 59430 24290
rect 59500 24280 59580 24290
rect 59650 24280 59730 24290
rect 60060 24280 60140 24290
rect 60210 24280 60290 24290
rect 60360 24280 60440 24290
rect 59430 24200 59440 24280
rect 59580 24200 59590 24280
rect 59730 24200 59740 24280
rect 60140 24200 60150 24280
rect 60290 24200 60300 24280
rect 60440 24200 60450 24280
rect 60850 24250 60860 24330
rect 61170 24250 61180 24330
rect 61590 24250 61600 24330
rect 61910 24250 61920 24330
rect 62060 24280 62140 24290
rect 62210 24280 62290 24290
rect 73560 24280 73640 24290
rect 73710 24280 73790 24290
rect 73860 24280 73940 24290
rect 62140 24200 62150 24280
rect 62290 24200 62300 24280
rect 73640 24200 73650 24280
rect 73790 24200 73800 24280
rect 73940 24200 73950 24280
rect 74350 24250 74360 24330
rect 74670 24250 74680 24330
rect 75090 24250 75100 24330
rect 75410 24250 75420 24330
rect 75560 24280 75640 24290
rect 75710 24280 75790 24290
rect 87060 24280 87140 24290
rect 87210 24280 87290 24290
rect 87360 24280 87440 24290
rect 75640 24200 75650 24280
rect 75790 24200 75800 24280
rect 87140 24200 87150 24280
rect 87290 24200 87300 24280
rect 87440 24200 87450 24280
rect 87850 24250 87860 24330
rect 88170 24250 88180 24330
rect 88590 24250 88600 24330
rect 88910 24250 88920 24330
rect 89060 24280 89140 24290
rect 89210 24280 89290 24290
rect 100560 24280 100640 24290
rect 100710 24280 100790 24290
rect 100860 24280 100940 24290
rect 89140 24200 89150 24280
rect 89290 24200 89300 24280
rect 100640 24200 100650 24280
rect 100790 24200 100800 24280
rect 100940 24200 100950 24280
rect 101350 24250 101360 24330
rect 101670 24250 101680 24330
rect 102090 24250 102100 24330
rect 102410 24250 102420 24330
rect 102560 24280 102640 24290
rect 102710 24280 102790 24290
rect 114060 24280 114140 24290
rect 114210 24280 114290 24290
rect 114360 24280 114440 24290
rect 102640 24200 102650 24280
rect 102790 24200 102800 24280
rect 114140 24200 114150 24280
rect 114290 24200 114300 24280
rect 114440 24200 114450 24280
rect 114850 24250 114860 24330
rect 115170 24250 115180 24330
rect 115590 24250 115600 24330
rect 115910 24250 115920 24330
rect 116060 24280 116140 24290
rect 116210 24280 116290 24290
rect 127560 24280 127640 24290
rect 127710 24280 127790 24290
rect 127860 24280 127940 24290
rect 116140 24200 116150 24280
rect 116290 24200 116300 24280
rect 127640 24200 127650 24280
rect 127790 24200 127800 24280
rect 127940 24200 127950 24280
rect 128350 24250 128360 24330
rect 128670 24250 128680 24330
rect 129090 24250 129100 24330
rect 129410 24250 129420 24330
rect 129560 24280 129640 24290
rect 129710 24280 129790 24290
rect 141060 24280 141140 24290
rect 141210 24280 141290 24290
rect 141360 24280 141440 24290
rect 129640 24200 129650 24280
rect 129790 24200 129800 24280
rect 141140 24200 141150 24280
rect 141290 24200 141300 24280
rect 141440 24200 141450 24280
rect 60610 24170 60690 24180
rect 60930 24170 61010 24180
rect 61350 24170 61430 24180
rect 61670 24170 61750 24180
rect 74110 24170 74190 24180
rect 74430 24170 74510 24180
rect 74850 24170 74930 24180
rect 75170 24170 75250 24180
rect 87610 24170 87690 24180
rect 87930 24170 88010 24180
rect 88350 24170 88430 24180
rect 88670 24170 88750 24180
rect 101110 24170 101190 24180
rect 101430 24170 101510 24180
rect 101850 24170 101930 24180
rect 102170 24170 102250 24180
rect 114610 24170 114690 24180
rect 114930 24170 115010 24180
rect 115350 24170 115430 24180
rect 115670 24170 115750 24180
rect 128110 24170 128190 24180
rect 128430 24170 128510 24180
rect 128850 24170 128930 24180
rect 129170 24170 129250 24180
rect 59350 24100 59430 24110
rect 59500 24100 59580 24110
rect 59650 24100 59730 24110
rect 60060 24100 60140 24110
rect 60210 24100 60290 24110
rect 60360 24100 60440 24110
rect 59430 24020 59440 24100
rect 59580 24020 59590 24100
rect 59730 24020 59740 24100
rect 60140 24020 60150 24100
rect 60290 24020 60300 24100
rect 60440 24020 60450 24100
rect 60690 24090 60700 24170
rect 61010 24090 61020 24170
rect 61430 24090 61440 24170
rect 61750 24090 61760 24170
rect 62060 24100 62140 24110
rect 62210 24100 62290 24110
rect 73560 24100 73640 24110
rect 73710 24100 73790 24110
rect 73860 24100 73940 24110
rect 62140 24020 62150 24100
rect 62290 24020 62300 24100
rect 73640 24020 73650 24100
rect 73790 24020 73800 24100
rect 73940 24020 73950 24100
rect 74190 24090 74200 24170
rect 74510 24090 74520 24170
rect 74930 24090 74940 24170
rect 75250 24090 75260 24170
rect 75560 24100 75640 24110
rect 75710 24100 75790 24110
rect 87060 24100 87140 24110
rect 87210 24100 87290 24110
rect 87360 24100 87440 24110
rect 75640 24020 75650 24100
rect 75790 24020 75800 24100
rect 87140 24020 87150 24100
rect 87290 24020 87300 24100
rect 87440 24020 87450 24100
rect 87690 24090 87700 24170
rect 88010 24090 88020 24170
rect 88430 24090 88440 24170
rect 88750 24090 88760 24170
rect 89060 24100 89140 24110
rect 89210 24100 89290 24110
rect 100560 24100 100640 24110
rect 100710 24100 100790 24110
rect 100860 24100 100940 24110
rect 89140 24020 89150 24100
rect 89290 24020 89300 24100
rect 100640 24020 100650 24100
rect 100790 24020 100800 24100
rect 100940 24020 100950 24100
rect 101190 24090 101200 24170
rect 101510 24090 101520 24170
rect 101930 24090 101940 24170
rect 102250 24090 102260 24170
rect 102560 24100 102640 24110
rect 102710 24100 102790 24110
rect 114060 24100 114140 24110
rect 114210 24100 114290 24110
rect 114360 24100 114440 24110
rect 102640 24020 102650 24100
rect 102790 24020 102800 24100
rect 114140 24020 114150 24100
rect 114290 24020 114300 24100
rect 114440 24020 114450 24100
rect 114690 24090 114700 24170
rect 115010 24090 115020 24170
rect 115430 24090 115440 24170
rect 115750 24090 115760 24170
rect 116060 24100 116140 24110
rect 116210 24100 116290 24110
rect 127560 24100 127640 24110
rect 127710 24100 127790 24110
rect 127860 24100 127940 24110
rect 116140 24020 116150 24100
rect 116290 24020 116300 24100
rect 127640 24020 127650 24100
rect 127790 24020 127800 24100
rect 127940 24020 127950 24100
rect 128190 24090 128200 24170
rect 128510 24090 128520 24170
rect 128930 24090 128940 24170
rect 129250 24090 129260 24170
rect 129560 24100 129640 24110
rect 129710 24100 129790 24110
rect 141060 24100 141140 24110
rect 141210 24100 141290 24110
rect 141360 24100 141440 24110
rect 129640 24020 129650 24100
rect 129790 24020 129800 24100
rect 141140 24020 141150 24100
rect 141290 24020 141300 24100
rect 141440 24020 141450 24100
rect 60770 24010 60850 24020
rect 61090 24010 61170 24020
rect 61510 24010 61590 24020
rect 61830 24010 61910 24020
rect 74270 24010 74350 24020
rect 74590 24010 74670 24020
rect 75010 24010 75090 24020
rect 75330 24010 75410 24020
rect 87770 24010 87850 24020
rect 88090 24010 88170 24020
rect 88510 24010 88590 24020
rect 88830 24010 88910 24020
rect 101270 24010 101350 24020
rect 101590 24010 101670 24020
rect 102010 24010 102090 24020
rect 102330 24010 102410 24020
rect 114770 24010 114850 24020
rect 115090 24010 115170 24020
rect 115510 24010 115590 24020
rect 115830 24010 115910 24020
rect 128270 24010 128350 24020
rect 128590 24010 128670 24020
rect 129010 24010 129090 24020
rect 129330 24010 129410 24020
rect 60850 23930 60860 24010
rect 61170 23930 61180 24010
rect 61590 23930 61600 24010
rect 61910 23930 61920 24010
rect 74350 23930 74360 24010
rect 74670 23930 74680 24010
rect 75090 23930 75100 24010
rect 75410 23930 75420 24010
rect 87850 23930 87860 24010
rect 88170 23930 88180 24010
rect 88590 23930 88600 24010
rect 88910 23930 88920 24010
rect 101350 23930 101360 24010
rect 101670 23930 101680 24010
rect 102090 23930 102100 24010
rect 102410 23930 102420 24010
rect 114850 23930 114860 24010
rect 115170 23930 115180 24010
rect 115590 23930 115600 24010
rect 115910 23930 115920 24010
rect 128350 23930 128360 24010
rect 128670 23930 128680 24010
rect 129090 23930 129100 24010
rect 129410 23930 129420 24010
rect 59350 23920 59430 23930
rect 59500 23920 59580 23930
rect 59650 23920 59730 23930
rect 60060 23920 60140 23930
rect 60210 23920 60290 23930
rect 60360 23920 60440 23930
rect 62060 23920 62140 23930
rect 62210 23920 62290 23930
rect 73560 23920 73640 23930
rect 73710 23920 73790 23930
rect 73860 23920 73940 23930
rect 75560 23920 75640 23930
rect 75710 23920 75790 23930
rect 87060 23920 87140 23930
rect 87210 23920 87290 23930
rect 87360 23920 87440 23930
rect 89060 23920 89140 23930
rect 89210 23920 89290 23930
rect 100560 23920 100640 23930
rect 100710 23920 100790 23930
rect 100860 23920 100940 23930
rect 102560 23920 102640 23930
rect 102710 23920 102790 23930
rect 114060 23920 114140 23930
rect 114210 23920 114290 23930
rect 114360 23920 114440 23930
rect 116060 23920 116140 23930
rect 116210 23920 116290 23930
rect 127560 23920 127640 23930
rect 127710 23920 127790 23930
rect 127860 23920 127940 23930
rect 129560 23920 129640 23930
rect 129710 23920 129790 23930
rect 141060 23920 141140 23930
rect 141210 23920 141290 23930
rect 141360 23920 141440 23930
rect 59430 23840 59440 23920
rect 59580 23840 59590 23920
rect 59730 23840 59740 23920
rect 60140 23840 60150 23920
rect 60290 23840 60300 23920
rect 60440 23840 60450 23920
rect 60610 23850 60690 23860
rect 60930 23850 61010 23860
rect 61350 23850 61430 23860
rect 61670 23850 61750 23860
rect 60690 23770 60700 23850
rect 61010 23770 61020 23850
rect 61430 23770 61440 23850
rect 61750 23770 61760 23850
rect 62140 23840 62150 23920
rect 62290 23840 62300 23920
rect 73640 23840 73650 23920
rect 73790 23840 73800 23920
rect 73940 23840 73950 23920
rect 74110 23850 74190 23860
rect 74430 23850 74510 23860
rect 74850 23850 74930 23860
rect 75170 23850 75250 23860
rect 74190 23770 74200 23850
rect 74510 23770 74520 23850
rect 74930 23770 74940 23850
rect 75250 23770 75260 23850
rect 75640 23840 75650 23920
rect 75790 23840 75800 23920
rect 87140 23840 87150 23920
rect 87290 23840 87300 23920
rect 87440 23840 87450 23920
rect 87610 23850 87690 23860
rect 87930 23850 88010 23860
rect 88350 23850 88430 23860
rect 88670 23850 88750 23860
rect 87690 23770 87700 23850
rect 88010 23770 88020 23850
rect 88430 23770 88440 23850
rect 88750 23770 88760 23850
rect 89140 23840 89150 23920
rect 89290 23840 89300 23920
rect 100640 23840 100650 23920
rect 100790 23840 100800 23920
rect 100940 23840 100950 23920
rect 101110 23850 101190 23860
rect 101430 23850 101510 23860
rect 101850 23850 101930 23860
rect 102170 23850 102250 23860
rect 101190 23770 101200 23850
rect 101510 23770 101520 23850
rect 101930 23770 101940 23850
rect 102250 23770 102260 23850
rect 102640 23840 102650 23920
rect 102790 23840 102800 23920
rect 114140 23840 114150 23920
rect 114290 23840 114300 23920
rect 114440 23840 114450 23920
rect 114610 23850 114690 23860
rect 114930 23850 115010 23860
rect 115350 23850 115430 23860
rect 115670 23850 115750 23860
rect 114690 23770 114700 23850
rect 115010 23770 115020 23850
rect 115430 23770 115440 23850
rect 115750 23770 115760 23850
rect 116140 23840 116150 23920
rect 116290 23840 116300 23920
rect 127640 23840 127650 23920
rect 127790 23840 127800 23920
rect 127940 23840 127950 23920
rect 128110 23850 128190 23860
rect 128430 23850 128510 23860
rect 128850 23850 128930 23860
rect 129170 23850 129250 23860
rect 128190 23770 128200 23850
rect 128510 23770 128520 23850
rect 128930 23770 128940 23850
rect 129250 23770 129260 23850
rect 129640 23840 129650 23920
rect 129790 23840 129800 23920
rect 141140 23840 141150 23920
rect 141290 23840 141300 23920
rect 141440 23840 141450 23920
rect 59350 23740 59430 23750
rect 59500 23740 59580 23750
rect 59650 23740 59730 23750
rect 60060 23740 60140 23750
rect 60210 23740 60290 23750
rect 60360 23740 60440 23750
rect 62060 23740 62140 23750
rect 62210 23740 62290 23750
rect 73560 23740 73640 23750
rect 73710 23740 73790 23750
rect 73860 23740 73940 23750
rect 75560 23740 75640 23750
rect 75710 23740 75790 23750
rect 87060 23740 87140 23750
rect 87210 23740 87290 23750
rect 87360 23740 87440 23750
rect 89060 23740 89140 23750
rect 89210 23740 89290 23750
rect 100560 23740 100640 23750
rect 100710 23740 100790 23750
rect 100860 23740 100940 23750
rect 102560 23740 102640 23750
rect 102710 23740 102790 23750
rect 114060 23740 114140 23750
rect 114210 23740 114290 23750
rect 114360 23740 114440 23750
rect 116060 23740 116140 23750
rect 116210 23740 116290 23750
rect 127560 23740 127640 23750
rect 127710 23740 127790 23750
rect 127860 23740 127940 23750
rect 129560 23740 129640 23750
rect 129710 23740 129790 23750
rect 141060 23740 141140 23750
rect 141210 23740 141290 23750
rect 141360 23740 141440 23750
rect 59430 23660 59440 23740
rect 59580 23660 59590 23740
rect 59730 23660 59740 23740
rect 60140 23660 60150 23740
rect 60290 23660 60300 23740
rect 60440 23660 60450 23740
rect 60770 23690 60850 23700
rect 61090 23690 61170 23700
rect 61510 23690 61590 23700
rect 61830 23690 61910 23700
rect 60850 23610 60860 23690
rect 61170 23610 61180 23690
rect 61590 23610 61600 23690
rect 61910 23610 61920 23690
rect 62140 23660 62150 23740
rect 62290 23660 62300 23740
rect 73640 23660 73650 23740
rect 73790 23660 73800 23740
rect 73940 23660 73950 23740
rect 74270 23690 74350 23700
rect 74590 23690 74670 23700
rect 75010 23690 75090 23700
rect 75330 23690 75410 23700
rect 74350 23610 74360 23690
rect 74670 23610 74680 23690
rect 75090 23610 75100 23690
rect 75410 23610 75420 23690
rect 75640 23660 75650 23740
rect 75790 23660 75800 23740
rect 87140 23660 87150 23740
rect 87290 23660 87300 23740
rect 87440 23660 87450 23740
rect 87770 23690 87850 23700
rect 88090 23690 88170 23700
rect 88510 23690 88590 23700
rect 88830 23690 88910 23700
rect 87850 23610 87860 23690
rect 88170 23610 88180 23690
rect 88590 23610 88600 23690
rect 88910 23610 88920 23690
rect 89140 23660 89150 23740
rect 89290 23660 89300 23740
rect 100640 23660 100650 23740
rect 100790 23660 100800 23740
rect 100940 23660 100950 23740
rect 101270 23690 101350 23700
rect 101590 23690 101670 23700
rect 102010 23690 102090 23700
rect 102330 23690 102410 23700
rect 101350 23610 101360 23690
rect 101670 23610 101680 23690
rect 102090 23610 102100 23690
rect 102410 23610 102420 23690
rect 102640 23660 102650 23740
rect 102790 23660 102800 23740
rect 114140 23660 114150 23740
rect 114290 23660 114300 23740
rect 114440 23660 114450 23740
rect 114770 23690 114850 23700
rect 115090 23690 115170 23700
rect 115510 23690 115590 23700
rect 115830 23690 115910 23700
rect 114850 23610 114860 23690
rect 115170 23610 115180 23690
rect 115590 23610 115600 23690
rect 115910 23610 115920 23690
rect 116140 23660 116150 23740
rect 116290 23660 116300 23740
rect 127640 23660 127650 23740
rect 127790 23660 127800 23740
rect 127940 23660 127950 23740
rect 128270 23690 128350 23700
rect 128590 23690 128670 23700
rect 129010 23690 129090 23700
rect 129330 23690 129410 23700
rect 128350 23610 128360 23690
rect 128670 23610 128680 23690
rect 129090 23610 129100 23690
rect 129410 23610 129420 23690
rect 129640 23660 129650 23740
rect 129790 23660 129800 23740
rect 141140 23660 141150 23740
rect 141290 23660 141300 23740
rect 141440 23660 141450 23740
rect 59350 23560 59430 23570
rect 59500 23560 59580 23570
rect 59650 23560 59730 23570
rect 60060 23560 60140 23570
rect 60210 23560 60290 23570
rect 60360 23560 60440 23570
rect 62060 23560 62140 23570
rect 62210 23560 62290 23570
rect 73560 23560 73640 23570
rect 73710 23560 73790 23570
rect 73860 23560 73940 23570
rect 75560 23560 75640 23570
rect 75710 23560 75790 23570
rect 87060 23560 87140 23570
rect 87210 23560 87290 23570
rect 87360 23560 87440 23570
rect 89060 23560 89140 23570
rect 89210 23560 89290 23570
rect 100560 23560 100640 23570
rect 100710 23560 100790 23570
rect 100860 23560 100940 23570
rect 102560 23560 102640 23570
rect 102710 23560 102790 23570
rect 114060 23560 114140 23570
rect 114210 23560 114290 23570
rect 114360 23560 114440 23570
rect 116060 23560 116140 23570
rect 116210 23560 116290 23570
rect 127560 23560 127640 23570
rect 127710 23560 127790 23570
rect 127860 23560 127940 23570
rect 129560 23560 129640 23570
rect 129710 23560 129790 23570
rect 141060 23560 141140 23570
rect 141210 23560 141290 23570
rect 141360 23560 141440 23570
rect 59430 23480 59440 23560
rect 59580 23480 59590 23560
rect 59730 23480 59740 23560
rect 60140 23480 60150 23560
rect 60290 23480 60300 23560
rect 60440 23480 60450 23560
rect 60610 23530 60690 23540
rect 60930 23530 61010 23540
rect 61350 23530 61430 23540
rect 61670 23530 61750 23540
rect 60690 23450 60700 23530
rect 61010 23450 61020 23530
rect 61430 23450 61440 23530
rect 61750 23450 61760 23530
rect 62140 23480 62150 23560
rect 62290 23480 62300 23560
rect 73640 23480 73650 23560
rect 73790 23480 73800 23560
rect 73940 23480 73950 23560
rect 74110 23530 74190 23540
rect 74430 23530 74510 23540
rect 74850 23530 74930 23540
rect 75170 23530 75250 23540
rect 74190 23450 74200 23530
rect 74510 23450 74520 23530
rect 74930 23450 74940 23530
rect 75250 23450 75260 23530
rect 75640 23480 75650 23560
rect 75790 23480 75800 23560
rect 87140 23480 87150 23560
rect 87290 23480 87300 23560
rect 87440 23480 87450 23560
rect 87610 23530 87690 23540
rect 87930 23530 88010 23540
rect 88350 23530 88430 23540
rect 88670 23530 88750 23540
rect 87690 23450 87700 23530
rect 88010 23450 88020 23530
rect 88430 23450 88440 23530
rect 88750 23450 88760 23530
rect 89140 23480 89150 23560
rect 89290 23480 89300 23560
rect 100640 23480 100650 23560
rect 100790 23480 100800 23560
rect 100940 23480 100950 23560
rect 101110 23530 101190 23540
rect 101430 23530 101510 23540
rect 101850 23530 101930 23540
rect 102170 23530 102250 23540
rect 101190 23450 101200 23530
rect 101510 23450 101520 23530
rect 101930 23450 101940 23530
rect 102250 23450 102260 23530
rect 102640 23480 102650 23560
rect 102790 23480 102800 23560
rect 114140 23480 114150 23560
rect 114290 23480 114300 23560
rect 114440 23480 114450 23560
rect 114610 23530 114690 23540
rect 114930 23530 115010 23540
rect 115350 23530 115430 23540
rect 115670 23530 115750 23540
rect 114690 23450 114700 23530
rect 115010 23450 115020 23530
rect 115430 23450 115440 23530
rect 115750 23450 115760 23530
rect 116140 23480 116150 23560
rect 116290 23480 116300 23560
rect 127640 23480 127650 23560
rect 127790 23480 127800 23560
rect 127940 23480 127950 23560
rect 128110 23530 128190 23540
rect 128430 23530 128510 23540
rect 128850 23530 128930 23540
rect 129170 23530 129250 23540
rect 128190 23450 128200 23530
rect 128510 23450 128520 23530
rect 128930 23450 128940 23530
rect 129250 23450 129260 23530
rect 129640 23480 129650 23560
rect 129790 23480 129800 23560
rect 141140 23480 141150 23560
rect 141290 23480 141300 23560
rect 141440 23480 141450 23560
rect 59350 23380 59430 23390
rect 59500 23380 59580 23390
rect 59650 23380 59730 23390
rect 60060 23380 60140 23390
rect 60210 23380 60290 23390
rect 60360 23380 60440 23390
rect 62060 23380 62140 23390
rect 62210 23380 62290 23390
rect 73560 23380 73640 23390
rect 73710 23380 73790 23390
rect 73860 23380 73940 23390
rect 75560 23380 75640 23390
rect 75710 23380 75790 23390
rect 87060 23380 87140 23390
rect 87210 23380 87290 23390
rect 87360 23380 87440 23390
rect 89060 23380 89140 23390
rect 89210 23380 89290 23390
rect 100560 23380 100640 23390
rect 100710 23380 100790 23390
rect 100860 23380 100940 23390
rect 102560 23380 102640 23390
rect 102710 23380 102790 23390
rect 114060 23380 114140 23390
rect 114210 23380 114290 23390
rect 114360 23380 114440 23390
rect 116060 23380 116140 23390
rect 116210 23380 116290 23390
rect 127560 23380 127640 23390
rect 127710 23380 127790 23390
rect 127860 23380 127940 23390
rect 129560 23380 129640 23390
rect 129710 23380 129790 23390
rect 141060 23380 141140 23390
rect 141210 23380 141290 23390
rect 141360 23380 141440 23390
rect 59430 23300 59440 23380
rect 59580 23300 59590 23380
rect 59730 23300 59740 23380
rect 60140 23300 60150 23380
rect 60290 23300 60300 23380
rect 60440 23300 60450 23380
rect 60770 23370 60850 23380
rect 61090 23370 61170 23380
rect 61510 23370 61590 23380
rect 61830 23370 61910 23380
rect 60850 23290 60860 23370
rect 61170 23290 61180 23370
rect 61590 23290 61600 23370
rect 61910 23290 61920 23370
rect 62140 23300 62150 23380
rect 62290 23300 62300 23380
rect 73640 23300 73650 23380
rect 73790 23300 73800 23380
rect 73940 23300 73950 23380
rect 74270 23370 74350 23380
rect 74590 23370 74670 23380
rect 75010 23370 75090 23380
rect 75330 23370 75410 23380
rect 74350 23290 74360 23370
rect 74670 23290 74680 23370
rect 75090 23290 75100 23370
rect 75410 23290 75420 23370
rect 75640 23300 75650 23380
rect 75790 23300 75800 23380
rect 87140 23300 87150 23380
rect 87290 23300 87300 23380
rect 87440 23300 87450 23380
rect 87770 23370 87850 23380
rect 88090 23370 88170 23380
rect 88510 23370 88590 23380
rect 88830 23370 88910 23380
rect 87850 23290 87860 23370
rect 88170 23290 88180 23370
rect 88590 23290 88600 23370
rect 88910 23290 88920 23370
rect 89140 23300 89150 23380
rect 89290 23300 89300 23380
rect 100640 23300 100650 23380
rect 100790 23300 100800 23380
rect 100940 23300 100950 23380
rect 101270 23370 101350 23380
rect 101590 23370 101670 23380
rect 102010 23370 102090 23380
rect 102330 23370 102410 23380
rect 101350 23290 101360 23370
rect 101670 23290 101680 23370
rect 102090 23290 102100 23370
rect 102410 23290 102420 23370
rect 102640 23300 102650 23380
rect 102790 23300 102800 23380
rect 114140 23300 114150 23380
rect 114290 23300 114300 23380
rect 114440 23300 114450 23380
rect 114770 23370 114850 23380
rect 115090 23370 115170 23380
rect 115510 23370 115590 23380
rect 115830 23370 115910 23380
rect 114850 23290 114860 23370
rect 115170 23290 115180 23370
rect 115590 23290 115600 23370
rect 115910 23290 115920 23370
rect 116140 23300 116150 23380
rect 116290 23300 116300 23380
rect 127640 23300 127650 23380
rect 127790 23300 127800 23380
rect 127940 23300 127950 23380
rect 128270 23370 128350 23380
rect 128590 23370 128670 23380
rect 129010 23370 129090 23380
rect 129330 23370 129410 23380
rect 128350 23290 128360 23370
rect 128670 23290 128680 23370
rect 129090 23290 129100 23370
rect 129410 23290 129420 23370
rect 129640 23300 129650 23380
rect 129790 23300 129800 23380
rect 141140 23300 141150 23380
rect 141290 23300 141300 23380
rect 141440 23300 141450 23380
rect 60610 23210 60690 23220
rect 60930 23210 61010 23220
rect 61350 23210 61430 23220
rect 61670 23210 61750 23220
rect 74110 23210 74190 23220
rect 74430 23210 74510 23220
rect 74850 23210 74930 23220
rect 75170 23210 75250 23220
rect 87610 23210 87690 23220
rect 87930 23210 88010 23220
rect 88350 23210 88430 23220
rect 88670 23210 88750 23220
rect 101110 23210 101190 23220
rect 101430 23210 101510 23220
rect 101850 23210 101930 23220
rect 102170 23210 102250 23220
rect 114610 23210 114690 23220
rect 114930 23210 115010 23220
rect 115350 23210 115430 23220
rect 115670 23210 115750 23220
rect 128110 23210 128190 23220
rect 128430 23210 128510 23220
rect 128850 23210 128930 23220
rect 129170 23210 129250 23220
rect 59350 23200 59430 23210
rect 59500 23200 59580 23210
rect 59650 23200 59730 23210
rect 60060 23200 60140 23210
rect 60210 23200 60290 23210
rect 60360 23200 60440 23210
rect 59430 23120 59440 23200
rect 59580 23120 59590 23200
rect 59730 23120 59740 23200
rect 60140 23120 60150 23200
rect 60290 23120 60300 23200
rect 60440 23120 60450 23200
rect 60690 23130 60700 23210
rect 61010 23130 61020 23210
rect 61430 23130 61440 23210
rect 61750 23130 61760 23210
rect 62060 23200 62140 23210
rect 62210 23200 62290 23210
rect 73560 23200 73640 23210
rect 73710 23200 73790 23210
rect 73860 23200 73940 23210
rect 62140 23120 62150 23200
rect 62290 23120 62300 23200
rect 73640 23120 73650 23200
rect 73790 23120 73800 23200
rect 73940 23120 73950 23200
rect 74190 23130 74200 23210
rect 74510 23130 74520 23210
rect 74930 23130 74940 23210
rect 75250 23130 75260 23210
rect 75560 23200 75640 23210
rect 75710 23200 75790 23210
rect 87060 23200 87140 23210
rect 87210 23200 87290 23210
rect 87360 23200 87440 23210
rect 75640 23120 75650 23200
rect 75790 23120 75800 23200
rect 87140 23120 87150 23200
rect 87290 23120 87300 23200
rect 87440 23120 87450 23200
rect 87690 23130 87700 23210
rect 88010 23130 88020 23210
rect 88430 23130 88440 23210
rect 88750 23130 88760 23210
rect 89060 23200 89140 23210
rect 89210 23200 89290 23210
rect 100560 23200 100640 23210
rect 100710 23200 100790 23210
rect 100860 23200 100940 23210
rect 89140 23120 89150 23200
rect 89290 23120 89300 23200
rect 100640 23120 100650 23200
rect 100790 23120 100800 23200
rect 100940 23120 100950 23200
rect 101190 23130 101200 23210
rect 101510 23130 101520 23210
rect 101930 23130 101940 23210
rect 102250 23130 102260 23210
rect 102560 23200 102640 23210
rect 102710 23200 102790 23210
rect 114060 23200 114140 23210
rect 114210 23200 114290 23210
rect 114360 23200 114440 23210
rect 102640 23120 102650 23200
rect 102790 23120 102800 23200
rect 114140 23120 114150 23200
rect 114290 23120 114300 23200
rect 114440 23120 114450 23200
rect 114690 23130 114700 23210
rect 115010 23130 115020 23210
rect 115430 23130 115440 23210
rect 115750 23130 115760 23210
rect 116060 23200 116140 23210
rect 116210 23200 116290 23210
rect 127560 23200 127640 23210
rect 127710 23200 127790 23210
rect 127860 23200 127940 23210
rect 116140 23120 116150 23200
rect 116290 23120 116300 23200
rect 127640 23120 127650 23200
rect 127790 23120 127800 23200
rect 127940 23120 127950 23200
rect 128190 23130 128200 23210
rect 128510 23130 128520 23210
rect 128930 23130 128940 23210
rect 129250 23130 129260 23210
rect 129560 23200 129640 23210
rect 129710 23200 129790 23210
rect 141060 23200 141140 23210
rect 141210 23200 141290 23210
rect 141360 23200 141440 23210
rect 129640 23120 129650 23200
rect 129790 23120 129800 23200
rect 141140 23120 141150 23200
rect 141290 23120 141300 23200
rect 141440 23120 141450 23200
rect 60770 23050 60850 23060
rect 61090 23050 61170 23060
rect 61510 23050 61590 23060
rect 61830 23050 61910 23060
rect 74270 23050 74350 23060
rect 74590 23050 74670 23060
rect 75010 23050 75090 23060
rect 75330 23050 75410 23060
rect 87770 23050 87850 23060
rect 88090 23050 88170 23060
rect 88510 23050 88590 23060
rect 88830 23050 88910 23060
rect 101270 23050 101350 23060
rect 101590 23050 101670 23060
rect 102010 23050 102090 23060
rect 102330 23050 102410 23060
rect 114770 23050 114850 23060
rect 115090 23050 115170 23060
rect 115510 23050 115590 23060
rect 115830 23050 115910 23060
rect 128270 23050 128350 23060
rect 128590 23050 128670 23060
rect 129010 23050 129090 23060
rect 129330 23050 129410 23060
rect 59350 23020 59430 23030
rect 59500 23020 59580 23030
rect 59650 23020 59730 23030
rect 60060 23020 60140 23030
rect 60210 23020 60290 23030
rect 60360 23020 60440 23030
rect 59430 22940 59440 23020
rect 59580 22940 59590 23020
rect 59730 22940 59740 23020
rect 60140 22940 60150 23020
rect 60290 22940 60300 23020
rect 60440 22940 60450 23020
rect 60850 22970 60860 23050
rect 61170 22970 61180 23050
rect 61590 22970 61600 23050
rect 61910 22970 61920 23050
rect 62060 23020 62140 23030
rect 62210 23020 62290 23030
rect 73560 23020 73640 23030
rect 73710 23020 73790 23030
rect 73860 23020 73940 23030
rect 62140 22940 62150 23020
rect 62290 22940 62300 23020
rect 73640 22940 73650 23020
rect 73790 22940 73800 23020
rect 73940 22940 73950 23020
rect 74350 22970 74360 23050
rect 74670 22970 74680 23050
rect 75090 22970 75100 23050
rect 75410 22970 75420 23050
rect 75560 23020 75640 23030
rect 75710 23020 75790 23030
rect 87060 23020 87140 23030
rect 87210 23020 87290 23030
rect 87360 23020 87440 23030
rect 75640 22940 75650 23020
rect 75790 22940 75800 23020
rect 87140 22940 87150 23020
rect 87290 22940 87300 23020
rect 87440 22940 87450 23020
rect 87850 22970 87860 23050
rect 88170 22970 88180 23050
rect 88590 22970 88600 23050
rect 88910 22970 88920 23050
rect 89060 23020 89140 23030
rect 89210 23020 89290 23030
rect 100560 23020 100640 23030
rect 100710 23020 100790 23030
rect 100860 23020 100940 23030
rect 89140 22940 89150 23020
rect 89290 22940 89300 23020
rect 100640 22940 100650 23020
rect 100790 22940 100800 23020
rect 100940 22940 100950 23020
rect 101350 22970 101360 23050
rect 101670 22970 101680 23050
rect 102090 22970 102100 23050
rect 102410 22970 102420 23050
rect 102560 23020 102640 23030
rect 102710 23020 102790 23030
rect 114060 23020 114140 23030
rect 114210 23020 114290 23030
rect 114360 23020 114440 23030
rect 102640 22940 102650 23020
rect 102790 22940 102800 23020
rect 114140 22940 114150 23020
rect 114290 22940 114300 23020
rect 114440 22940 114450 23020
rect 114850 22970 114860 23050
rect 115170 22970 115180 23050
rect 115590 22970 115600 23050
rect 115910 22970 115920 23050
rect 116060 23020 116140 23030
rect 116210 23020 116290 23030
rect 127560 23020 127640 23030
rect 127710 23020 127790 23030
rect 127860 23020 127940 23030
rect 116140 22940 116150 23020
rect 116290 22940 116300 23020
rect 127640 22940 127650 23020
rect 127790 22940 127800 23020
rect 127940 22940 127950 23020
rect 128350 22970 128360 23050
rect 128670 22970 128680 23050
rect 129090 22970 129100 23050
rect 129410 22970 129420 23050
rect 129560 23020 129640 23030
rect 129710 23020 129790 23030
rect 141060 23020 141140 23030
rect 141210 23020 141290 23030
rect 141360 23020 141440 23030
rect 129640 22940 129650 23020
rect 129790 22940 129800 23020
rect 141140 22940 141150 23020
rect 141290 22940 141300 23020
rect 141440 22940 141450 23020
rect 60610 22890 60690 22900
rect 60930 22890 61010 22900
rect 61350 22890 61430 22900
rect 61670 22890 61750 22900
rect 74110 22890 74190 22900
rect 74430 22890 74510 22900
rect 74850 22890 74930 22900
rect 75170 22890 75250 22900
rect 87610 22890 87690 22900
rect 87930 22890 88010 22900
rect 88350 22890 88430 22900
rect 88670 22890 88750 22900
rect 101110 22890 101190 22900
rect 101430 22890 101510 22900
rect 101850 22890 101930 22900
rect 102170 22890 102250 22900
rect 114610 22890 114690 22900
rect 114930 22890 115010 22900
rect 115350 22890 115430 22900
rect 115670 22890 115750 22900
rect 128110 22890 128190 22900
rect 128430 22890 128510 22900
rect 128850 22890 128930 22900
rect 129170 22890 129250 22900
rect 59350 22840 59430 22850
rect 59500 22840 59580 22850
rect 59650 22840 59730 22850
rect 60060 22840 60140 22850
rect 60210 22840 60290 22850
rect 60360 22840 60440 22850
rect 59430 22760 59440 22840
rect 59580 22760 59590 22840
rect 59730 22760 59740 22840
rect 60140 22760 60150 22840
rect 60290 22760 60300 22840
rect 60440 22760 60450 22840
rect 60690 22810 60700 22890
rect 61010 22810 61020 22890
rect 61430 22810 61440 22890
rect 61750 22810 61760 22890
rect 62060 22840 62140 22850
rect 62210 22840 62290 22850
rect 73560 22840 73640 22850
rect 73710 22840 73790 22850
rect 73860 22840 73940 22850
rect 62140 22760 62150 22840
rect 62290 22760 62300 22840
rect 73640 22760 73650 22840
rect 73790 22760 73800 22840
rect 73940 22760 73950 22840
rect 74190 22810 74200 22890
rect 74510 22810 74520 22890
rect 74930 22810 74940 22890
rect 75250 22810 75260 22890
rect 75560 22840 75640 22850
rect 75710 22840 75790 22850
rect 87060 22840 87140 22850
rect 87210 22840 87290 22850
rect 87360 22840 87440 22850
rect 75640 22760 75650 22840
rect 75790 22760 75800 22840
rect 87140 22760 87150 22840
rect 87290 22760 87300 22840
rect 87440 22760 87450 22840
rect 87690 22810 87700 22890
rect 88010 22810 88020 22890
rect 88430 22810 88440 22890
rect 88750 22810 88760 22890
rect 89060 22840 89140 22850
rect 89210 22840 89290 22850
rect 100560 22840 100640 22850
rect 100710 22840 100790 22850
rect 100860 22840 100940 22850
rect 89140 22760 89150 22840
rect 89290 22760 89300 22840
rect 100640 22760 100650 22840
rect 100790 22760 100800 22840
rect 100940 22760 100950 22840
rect 101190 22810 101200 22890
rect 101510 22810 101520 22890
rect 101930 22810 101940 22890
rect 102250 22810 102260 22890
rect 102560 22840 102640 22850
rect 102710 22840 102790 22850
rect 114060 22840 114140 22850
rect 114210 22840 114290 22850
rect 114360 22840 114440 22850
rect 102640 22760 102650 22840
rect 102790 22760 102800 22840
rect 114140 22760 114150 22840
rect 114290 22760 114300 22840
rect 114440 22760 114450 22840
rect 114690 22810 114700 22890
rect 115010 22810 115020 22890
rect 115430 22810 115440 22890
rect 115750 22810 115760 22890
rect 116060 22840 116140 22850
rect 116210 22840 116290 22850
rect 127560 22840 127640 22850
rect 127710 22840 127790 22850
rect 127860 22840 127940 22850
rect 116140 22760 116150 22840
rect 116290 22760 116300 22840
rect 127640 22760 127650 22840
rect 127790 22760 127800 22840
rect 127940 22760 127950 22840
rect 128190 22810 128200 22890
rect 128510 22810 128520 22890
rect 128930 22810 128940 22890
rect 129250 22810 129260 22890
rect 129560 22840 129640 22850
rect 129710 22840 129790 22850
rect 141060 22840 141140 22850
rect 141210 22840 141290 22850
rect 141360 22840 141440 22850
rect 129640 22760 129650 22840
rect 129790 22760 129800 22840
rect 141140 22760 141150 22840
rect 141290 22760 141300 22840
rect 141440 22760 141450 22840
rect 60770 22730 60850 22740
rect 61090 22730 61170 22740
rect 61510 22730 61590 22740
rect 61830 22730 61910 22740
rect 74270 22730 74350 22740
rect 74590 22730 74670 22740
rect 75010 22730 75090 22740
rect 75330 22730 75410 22740
rect 87770 22730 87850 22740
rect 88090 22730 88170 22740
rect 88510 22730 88590 22740
rect 88830 22730 88910 22740
rect 101270 22730 101350 22740
rect 101590 22730 101670 22740
rect 102010 22730 102090 22740
rect 102330 22730 102410 22740
rect 114770 22730 114850 22740
rect 115090 22730 115170 22740
rect 115510 22730 115590 22740
rect 115830 22730 115910 22740
rect 128270 22730 128350 22740
rect 128590 22730 128670 22740
rect 129010 22730 129090 22740
rect 129330 22730 129410 22740
rect 59350 22660 59430 22670
rect 59500 22660 59580 22670
rect 59650 22660 59730 22670
rect 60060 22660 60140 22670
rect 60210 22660 60290 22670
rect 60360 22660 60440 22670
rect 59430 22580 59440 22660
rect 59580 22580 59590 22660
rect 59730 22580 59740 22660
rect 60140 22580 60150 22660
rect 60290 22580 60300 22660
rect 60440 22580 60450 22660
rect 60850 22650 60860 22730
rect 61170 22650 61180 22730
rect 61590 22650 61600 22730
rect 61910 22650 61920 22730
rect 62060 22660 62140 22670
rect 62210 22660 62290 22670
rect 73560 22660 73640 22670
rect 73710 22660 73790 22670
rect 73860 22660 73940 22670
rect 62140 22580 62150 22660
rect 62290 22580 62300 22660
rect 73640 22580 73650 22660
rect 73790 22580 73800 22660
rect 73940 22580 73950 22660
rect 74350 22650 74360 22730
rect 74670 22650 74680 22730
rect 75090 22650 75100 22730
rect 75410 22650 75420 22730
rect 75560 22660 75640 22670
rect 75710 22660 75790 22670
rect 87060 22660 87140 22670
rect 87210 22660 87290 22670
rect 87360 22660 87440 22670
rect 75640 22580 75650 22660
rect 75790 22580 75800 22660
rect 87140 22580 87150 22660
rect 87290 22580 87300 22660
rect 87440 22580 87450 22660
rect 87850 22650 87860 22730
rect 88170 22650 88180 22730
rect 88590 22650 88600 22730
rect 88910 22650 88920 22730
rect 89060 22660 89140 22670
rect 89210 22660 89290 22670
rect 100560 22660 100640 22670
rect 100710 22660 100790 22670
rect 100860 22660 100940 22670
rect 89140 22580 89150 22660
rect 89290 22580 89300 22660
rect 100640 22580 100650 22660
rect 100790 22580 100800 22660
rect 100940 22580 100950 22660
rect 101350 22650 101360 22730
rect 101670 22650 101680 22730
rect 102090 22650 102100 22730
rect 102410 22650 102420 22730
rect 102560 22660 102640 22670
rect 102710 22660 102790 22670
rect 114060 22660 114140 22670
rect 114210 22660 114290 22670
rect 114360 22660 114440 22670
rect 102640 22580 102650 22660
rect 102790 22580 102800 22660
rect 114140 22580 114150 22660
rect 114290 22580 114300 22660
rect 114440 22580 114450 22660
rect 114850 22650 114860 22730
rect 115170 22650 115180 22730
rect 115590 22650 115600 22730
rect 115910 22650 115920 22730
rect 116060 22660 116140 22670
rect 116210 22660 116290 22670
rect 127560 22660 127640 22670
rect 127710 22660 127790 22670
rect 127860 22660 127940 22670
rect 116140 22580 116150 22660
rect 116290 22580 116300 22660
rect 127640 22580 127650 22660
rect 127790 22580 127800 22660
rect 127940 22580 127950 22660
rect 128350 22650 128360 22730
rect 128670 22650 128680 22730
rect 129090 22650 129100 22730
rect 129410 22650 129420 22730
rect 129560 22660 129640 22670
rect 129710 22660 129790 22670
rect 141060 22660 141140 22670
rect 141210 22660 141290 22670
rect 141360 22660 141440 22670
rect 129640 22580 129650 22660
rect 129790 22580 129800 22660
rect 141140 22580 141150 22660
rect 141290 22580 141300 22660
rect 141440 22580 141450 22660
rect 60610 22570 60690 22580
rect 60930 22570 61010 22580
rect 61350 22570 61430 22580
rect 61670 22570 61750 22580
rect 74110 22570 74190 22580
rect 74430 22570 74510 22580
rect 74850 22570 74930 22580
rect 75170 22570 75250 22580
rect 87610 22570 87690 22580
rect 87930 22570 88010 22580
rect 88350 22570 88430 22580
rect 88670 22570 88750 22580
rect 101110 22570 101190 22580
rect 101430 22570 101510 22580
rect 101850 22570 101930 22580
rect 102170 22570 102250 22580
rect 114610 22570 114690 22580
rect 114930 22570 115010 22580
rect 115350 22570 115430 22580
rect 115670 22570 115750 22580
rect 128110 22570 128190 22580
rect 128430 22570 128510 22580
rect 128850 22570 128930 22580
rect 129170 22570 129250 22580
rect 60690 22490 60700 22570
rect 61010 22490 61020 22570
rect 61430 22490 61440 22570
rect 61750 22490 61760 22570
rect 74190 22490 74200 22570
rect 74510 22490 74520 22570
rect 74930 22490 74940 22570
rect 75250 22490 75260 22570
rect 87690 22490 87700 22570
rect 88010 22490 88020 22570
rect 88430 22490 88440 22570
rect 88750 22490 88760 22570
rect 101190 22490 101200 22570
rect 101510 22490 101520 22570
rect 101930 22490 101940 22570
rect 102250 22490 102260 22570
rect 114690 22490 114700 22570
rect 115010 22490 115020 22570
rect 115430 22490 115440 22570
rect 115750 22490 115760 22570
rect 128190 22490 128200 22570
rect 128510 22490 128520 22570
rect 128930 22490 128940 22570
rect 129250 22490 129260 22570
rect 59350 22480 59430 22490
rect 59500 22480 59580 22490
rect 59650 22480 59730 22490
rect 60060 22480 60140 22490
rect 60210 22480 60290 22490
rect 60360 22480 60440 22490
rect 62060 22480 62140 22490
rect 62210 22480 62290 22490
rect 73560 22480 73640 22490
rect 73710 22480 73790 22490
rect 73860 22480 73940 22490
rect 75560 22480 75640 22490
rect 75710 22480 75790 22490
rect 87060 22480 87140 22490
rect 87210 22480 87290 22490
rect 87360 22480 87440 22490
rect 89060 22480 89140 22490
rect 89210 22480 89290 22490
rect 100560 22480 100640 22490
rect 100710 22480 100790 22490
rect 100860 22480 100940 22490
rect 102560 22480 102640 22490
rect 102710 22480 102790 22490
rect 114060 22480 114140 22490
rect 114210 22480 114290 22490
rect 114360 22480 114440 22490
rect 116060 22480 116140 22490
rect 116210 22480 116290 22490
rect 127560 22480 127640 22490
rect 127710 22480 127790 22490
rect 127860 22480 127940 22490
rect 129560 22480 129640 22490
rect 129710 22480 129790 22490
rect 141060 22480 141140 22490
rect 141210 22480 141290 22490
rect 141360 22480 141440 22490
rect 59430 22400 59440 22480
rect 59580 22400 59590 22480
rect 59730 22400 59740 22480
rect 60140 22400 60150 22480
rect 60290 22400 60300 22480
rect 60440 22400 60450 22480
rect 60770 22410 60850 22420
rect 61090 22410 61170 22420
rect 61510 22410 61590 22420
rect 61830 22410 61910 22420
rect 60850 22330 60860 22410
rect 61170 22330 61180 22410
rect 61590 22330 61600 22410
rect 61910 22330 61920 22410
rect 62140 22400 62150 22480
rect 62290 22400 62300 22480
rect 73640 22400 73650 22480
rect 73790 22400 73800 22480
rect 73940 22400 73950 22480
rect 74270 22410 74350 22420
rect 74590 22410 74670 22420
rect 75010 22410 75090 22420
rect 75330 22410 75410 22420
rect 74350 22330 74360 22410
rect 74670 22330 74680 22410
rect 75090 22330 75100 22410
rect 75410 22330 75420 22410
rect 75640 22400 75650 22480
rect 75790 22400 75800 22480
rect 87140 22400 87150 22480
rect 87290 22400 87300 22480
rect 87440 22400 87450 22480
rect 87770 22410 87850 22420
rect 88090 22410 88170 22420
rect 88510 22410 88590 22420
rect 88830 22410 88910 22420
rect 87850 22330 87860 22410
rect 88170 22330 88180 22410
rect 88590 22330 88600 22410
rect 88910 22330 88920 22410
rect 89140 22400 89150 22480
rect 89290 22400 89300 22480
rect 100640 22400 100650 22480
rect 100790 22400 100800 22480
rect 100940 22400 100950 22480
rect 101270 22410 101350 22420
rect 101590 22410 101670 22420
rect 102010 22410 102090 22420
rect 102330 22410 102410 22420
rect 101350 22330 101360 22410
rect 101670 22330 101680 22410
rect 102090 22330 102100 22410
rect 102410 22330 102420 22410
rect 102640 22400 102650 22480
rect 102790 22400 102800 22480
rect 114140 22400 114150 22480
rect 114290 22400 114300 22480
rect 114440 22400 114450 22480
rect 114770 22410 114850 22420
rect 115090 22410 115170 22420
rect 115510 22410 115590 22420
rect 115830 22410 115910 22420
rect 114850 22330 114860 22410
rect 115170 22330 115180 22410
rect 115590 22330 115600 22410
rect 115910 22330 115920 22410
rect 116140 22400 116150 22480
rect 116290 22400 116300 22480
rect 127640 22400 127650 22480
rect 127790 22400 127800 22480
rect 127940 22400 127950 22480
rect 128270 22410 128350 22420
rect 128590 22410 128670 22420
rect 129010 22410 129090 22420
rect 129330 22410 129410 22420
rect 128350 22330 128360 22410
rect 128670 22330 128680 22410
rect 129090 22330 129100 22410
rect 129410 22330 129420 22410
rect 129640 22400 129650 22480
rect 129790 22400 129800 22480
rect 141140 22400 141150 22480
rect 141290 22400 141300 22480
rect 141440 22400 141450 22480
rect 59350 22300 59430 22310
rect 59500 22300 59580 22310
rect 59650 22300 59730 22310
rect 60060 22300 60140 22310
rect 60210 22300 60290 22310
rect 60360 22300 60440 22310
rect 62060 22300 62140 22310
rect 62210 22300 62290 22310
rect 73560 22300 73640 22310
rect 73710 22300 73790 22310
rect 73860 22300 73940 22310
rect 75560 22300 75640 22310
rect 75710 22300 75790 22310
rect 87060 22300 87140 22310
rect 87210 22300 87290 22310
rect 87360 22300 87440 22310
rect 89060 22300 89140 22310
rect 89210 22300 89290 22310
rect 100560 22300 100640 22310
rect 100710 22300 100790 22310
rect 100860 22300 100940 22310
rect 102560 22300 102640 22310
rect 102710 22300 102790 22310
rect 114060 22300 114140 22310
rect 114210 22300 114290 22310
rect 114360 22300 114440 22310
rect 116060 22300 116140 22310
rect 116210 22300 116290 22310
rect 127560 22300 127640 22310
rect 127710 22300 127790 22310
rect 127860 22300 127940 22310
rect 129560 22300 129640 22310
rect 129710 22300 129790 22310
rect 141060 22300 141140 22310
rect 141210 22300 141290 22310
rect 141360 22300 141440 22310
rect 59430 22220 59440 22300
rect 59580 22220 59590 22300
rect 59730 22220 59740 22300
rect 60140 22220 60150 22300
rect 60290 22220 60300 22300
rect 60440 22220 60450 22300
rect 60610 22250 60690 22260
rect 60930 22250 61010 22260
rect 61350 22250 61430 22260
rect 61670 22250 61750 22260
rect 60690 22170 60700 22250
rect 61010 22170 61020 22250
rect 61430 22170 61440 22250
rect 61750 22170 61760 22250
rect 62140 22220 62150 22300
rect 62290 22220 62300 22300
rect 73640 22220 73650 22300
rect 73790 22220 73800 22300
rect 73940 22220 73950 22300
rect 74110 22250 74190 22260
rect 74430 22250 74510 22260
rect 74850 22250 74930 22260
rect 75170 22250 75250 22260
rect 74190 22170 74200 22250
rect 74510 22170 74520 22250
rect 74930 22170 74940 22250
rect 75250 22170 75260 22250
rect 75640 22220 75650 22300
rect 75790 22220 75800 22300
rect 87140 22220 87150 22300
rect 87290 22220 87300 22300
rect 87440 22220 87450 22300
rect 87610 22250 87690 22260
rect 87930 22250 88010 22260
rect 88350 22250 88430 22260
rect 88670 22250 88750 22260
rect 87690 22170 87700 22250
rect 88010 22170 88020 22250
rect 88430 22170 88440 22250
rect 88750 22170 88760 22250
rect 89140 22220 89150 22300
rect 89290 22220 89300 22300
rect 100640 22220 100650 22300
rect 100790 22220 100800 22300
rect 100940 22220 100950 22300
rect 101110 22250 101190 22260
rect 101430 22250 101510 22260
rect 101850 22250 101930 22260
rect 102170 22250 102250 22260
rect 101190 22170 101200 22250
rect 101510 22170 101520 22250
rect 101930 22170 101940 22250
rect 102250 22170 102260 22250
rect 102640 22220 102650 22300
rect 102790 22220 102800 22300
rect 114140 22220 114150 22300
rect 114290 22220 114300 22300
rect 114440 22220 114450 22300
rect 114610 22250 114690 22260
rect 114930 22250 115010 22260
rect 115350 22250 115430 22260
rect 115670 22250 115750 22260
rect 114690 22170 114700 22250
rect 115010 22170 115020 22250
rect 115430 22170 115440 22250
rect 115750 22170 115760 22250
rect 116140 22220 116150 22300
rect 116290 22220 116300 22300
rect 127640 22220 127650 22300
rect 127790 22220 127800 22300
rect 127940 22220 127950 22300
rect 128110 22250 128190 22260
rect 128430 22250 128510 22260
rect 128850 22250 128930 22260
rect 129170 22250 129250 22260
rect 128190 22170 128200 22250
rect 128510 22170 128520 22250
rect 128930 22170 128940 22250
rect 129250 22170 129260 22250
rect 129640 22220 129650 22300
rect 129790 22220 129800 22300
rect 141140 22220 141150 22300
rect 141290 22220 141300 22300
rect 141440 22220 141450 22300
rect 59350 22120 59430 22130
rect 59500 22120 59580 22130
rect 59650 22120 59730 22130
rect 60060 22120 60140 22130
rect 60210 22120 60290 22130
rect 60360 22120 60440 22130
rect 62060 22120 62140 22130
rect 62210 22120 62290 22130
rect 73560 22120 73640 22130
rect 73710 22120 73790 22130
rect 73860 22120 73940 22130
rect 75560 22120 75640 22130
rect 75710 22120 75790 22130
rect 87060 22120 87140 22130
rect 87210 22120 87290 22130
rect 87360 22120 87440 22130
rect 89060 22120 89140 22130
rect 89210 22120 89290 22130
rect 100560 22120 100640 22130
rect 100710 22120 100790 22130
rect 100860 22120 100940 22130
rect 102560 22120 102640 22130
rect 102710 22120 102790 22130
rect 114060 22120 114140 22130
rect 114210 22120 114290 22130
rect 114360 22120 114440 22130
rect 116060 22120 116140 22130
rect 116210 22120 116290 22130
rect 127560 22120 127640 22130
rect 127710 22120 127790 22130
rect 127860 22120 127940 22130
rect 129560 22120 129640 22130
rect 129710 22120 129790 22130
rect 141060 22120 141140 22130
rect 141210 22120 141290 22130
rect 141360 22120 141440 22130
rect 59430 22040 59440 22120
rect 59580 22040 59590 22120
rect 59730 22040 59740 22120
rect 60140 22040 60150 22120
rect 60290 22040 60300 22120
rect 60440 22040 60450 22120
rect 60770 22090 60850 22100
rect 61090 22090 61170 22100
rect 61510 22090 61590 22100
rect 61830 22090 61910 22100
rect 60850 22010 60860 22090
rect 61170 22010 61180 22090
rect 61590 22010 61600 22090
rect 61910 22010 61920 22090
rect 62140 22040 62150 22120
rect 62290 22040 62300 22120
rect 73640 22040 73650 22120
rect 73790 22040 73800 22120
rect 73940 22040 73950 22120
rect 74270 22090 74350 22100
rect 74590 22090 74670 22100
rect 75010 22090 75090 22100
rect 75330 22090 75410 22100
rect 74350 22010 74360 22090
rect 74670 22010 74680 22090
rect 75090 22010 75100 22090
rect 75410 22010 75420 22090
rect 75640 22040 75650 22120
rect 75790 22040 75800 22120
rect 87140 22040 87150 22120
rect 87290 22040 87300 22120
rect 87440 22040 87450 22120
rect 87770 22090 87850 22100
rect 88090 22090 88170 22100
rect 88510 22090 88590 22100
rect 88830 22090 88910 22100
rect 87850 22010 87860 22090
rect 88170 22010 88180 22090
rect 88590 22010 88600 22090
rect 88910 22010 88920 22090
rect 89140 22040 89150 22120
rect 89290 22040 89300 22120
rect 100640 22040 100650 22120
rect 100790 22040 100800 22120
rect 100940 22040 100950 22120
rect 101270 22090 101350 22100
rect 101590 22090 101670 22100
rect 102010 22090 102090 22100
rect 102330 22090 102410 22100
rect 101350 22010 101360 22090
rect 101670 22010 101680 22090
rect 102090 22010 102100 22090
rect 102410 22010 102420 22090
rect 102640 22040 102650 22120
rect 102790 22040 102800 22120
rect 114140 22040 114150 22120
rect 114290 22040 114300 22120
rect 114440 22040 114450 22120
rect 114770 22090 114850 22100
rect 115090 22090 115170 22100
rect 115510 22090 115590 22100
rect 115830 22090 115910 22100
rect 114850 22010 114860 22090
rect 115170 22010 115180 22090
rect 115590 22010 115600 22090
rect 115910 22010 115920 22090
rect 116140 22040 116150 22120
rect 116290 22040 116300 22120
rect 127640 22040 127650 22120
rect 127790 22040 127800 22120
rect 127940 22040 127950 22120
rect 128270 22090 128350 22100
rect 128590 22090 128670 22100
rect 129010 22090 129090 22100
rect 129330 22090 129410 22100
rect 128350 22010 128360 22090
rect 128670 22010 128680 22090
rect 129090 22010 129100 22090
rect 129410 22010 129420 22090
rect 129640 22040 129650 22120
rect 129790 22040 129800 22120
rect 141140 22040 141150 22120
rect 141290 22040 141300 22120
rect 141440 22040 141450 22120
rect 59350 21940 59430 21950
rect 59500 21940 59580 21950
rect 59650 21940 59730 21950
rect 60060 21940 60140 21950
rect 60210 21940 60290 21950
rect 60360 21940 60440 21950
rect 62060 21940 62140 21950
rect 62210 21940 62290 21950
rect 73560 21940 73640 21950
rect 73710 21940 73790 21950
rect 73860 21940 73940 21950
rect 75560 21940 75640 21950
rect 75710 21940 75790 21950
rect 87060 21940 87140 21950
rect 87210 21940 87290 21950
rect 87360 21940 87440 21950
rect 89060 21940 89140 21950
rect 89210 21940 89290 21950
rect 100560 21940 100640 21950
rect 100710 21940 100790 21950
rect 100860 21940 100940 21950
rect 102560 21940 102640 21950
rect 102710 21940 102790 21950
rect 114060 21940 114140 21950
rect 114210 21940 114290 21950
rect 114360 21940 114440 21950
rect 116060 21940 116140 21950
rect 116210 21940 116290 21950
rect 127560 21940 127640 21950
rect 127710 21940 127790 21950
rect 127860 21940 127940 21950
rect 129560 21940 129640 21950
rect 129710 21940 129790 21950
rect 141060 21940 141140 21950
rect 141210 21940 141290 21950
rect 141360 21940 141440 21950
rect 59430 21860 59440 21940
rect 59580 21860 59590 21940
rect 59730 21860 59740 21940
rect 60140 21860 60150 21940
rect 60290 21860 60300 21940
rect 60440 21860 60450 21940
rect 60610 21930 60690 21940
rect 60930 21930 61010 21940
rect 61350 21930 61430 21940
rect 61670 21930 61750 21940
rect 60690 21850 60700 21930
rect 61010 21850 61020 21930
rect 61430 21850 61440 21930
rect 61750 21850 61760 21930
rect 62140 21860 62150 21940
rect 62290 21860 62300 21940
rect 73640 21860 73650 21940
rect 73790 21860 73800 21940
rect 73940 21860 73950 21940
rect 74110 21930 74190 21940
rect 74430 21930 74510 21940
rect 74850 21930 74930 21940
rect 75170 21930 75250 21940
rect 74190 21850 74200 21930
rect 74510 21850 74520 21930
rect 74930 21850 74940 21930
rect 75250 21850 75260 21930
rect 75640 21860 75650 21940
rect 75790 21860 75800 21940
rect 87140 21860 87150 21940
rect 87290 21860 87300 21940
rect 87440 21860 87450 21940
rect 87610 21930 87690 21940
rect 87930 21930 88010 21940
rect 88350 21930 88430 21940
rect 88670 21930 88750 21940
rect 87690 21850 87700 21930
rect 88010 21850 88020 21930
rect 88430 21850 88440 21930
rect 88750 21850 88760 21930
rect 89140 21860 89150 21940
rect 89290 21860 89300 21940
rect 100640 21860 100650 21940
rect 100790 21860 100800 21940
rect 100940 21860 100950 21940
rect 101110 21930 101190 21940
rect 101430 21930 101510 21940
rect 101850 21930 101930 21940
rect 102170 21930 102250 21940
rect 101190 21850 101200 21930
rect 101510 21850 101520 21930
rect 101930 21850 101940 21930
rect 102250 21850 102260 21930
rect 102640 21860 102650 21940
rect 102790 21860 102800 21940
rect 114140 21860 114150 21940
rect 114290 21860 114300 21940
rect 114440 21860 114450 21940
rect 114610 21930 114690 21940
rect 114930 21930 115010 21940
rect 115350 21930 115430 21940
rect 115670 21930 115750 21940
rect 114690 21850 114700 21930
rect 115010 21850 115020 21930
rect 115430 21850 115440 21930
rect 115750 21850 115760 21930
rect 116140 21860 116150 21940
rect 116290 21860 116300 21940
rect 127640 21860 127650 21940
rect 127790 21860 127800 21940
rect 127940 21860 127950 21940
rect 128110 21930 128190 21940
rect 128430 21930 128510 21940
rect 128850 21930 128930 21940
rect 129170 21930 129250 21940
rect 128190 21850 128200 21930
rect 128510 21850 128520 21930
rect 128930 21850 128940 21930
rect 129250 21850 129260 21930
rect 129640 21860 129650 21940
rect 129790 21860 129800 21940
rect 141140 21860 141150 21940
rect 141290 21860 141300 21940
rect 141440 21860 141450 21940
rect 60770 21770 60850 21780
rect 61090 21770 61170 21780
rect 61510 21770 61590 21780
rect 61830 21770 61910 21780
rect 74270 21770 74350 21780
rect 74590 21770 74670 21780
rect 75010 21770 75090 21780
rect 75330 21770 75410 21780
rect 87770 21770 87850 21780
rect 88090 21770 88170 21780
rect 88510 21770 88590 21780
rect 88830 21770 88910 21780
rect 101270 21770 101350 21780
rect 101590 21770 101670 21780
rect 102010 21770 102090 21780
rect 102330 21770 102410 21780
rect 114770 21770 114850 21780
rect 115090 21770 115170 21780
rect 115510 21770 115590 21780
rect 115830 21770 115910 21780
rect 128270 21770 128350 21780
rect 128590 21770 128670 21780
rect 129010 21770 129090 21780
rect 129330 21770 129410 21780
rect 59350 21760 59430 21770
rect 59500 21760 59580 21770
rect 59650 21760 59730 21770
rect 60060 21760 60140 21770
rect 60210 21760 60290 21770
rect 60360 21760 60440 21770
rect 59430 21680 59440 21760
rect 59580 21680 59590 21760
rect 59730 21680 59740 21760
rect 60140 21680 60150 21760
rect 60290 21680 60300 21760
rect 60440 21680 60450 21760
rect 60850 21690 60860 21770
rect 61170 21690 61180 21770
rect 61590 21690 61600 21770
rect 61910 21690 61920 21770
rect 62060 21760 62140 21770
rect 62210 21760 62290 21770
rect 73560 21760 73640 21770
rect 73710 21760 73790 21770
rect 73860 21760 73940 21770
rect 62140 21680 62150 21760
rect 62290 21680 62300 21760
rect 73640 21680 73650 21760
rect 73790 21680 73800 21760
rect 73940 21680 73950 21760
rect 74350 21690 74360 21770
rect 74670 21690 74680 21770
rect 75090 21690 75100 21770
rect 75410 21690 75420 21770
rect 75560 21760 75640 21770
rect 75710 21760 75790 21770
rect 87060 21760 87140 21770
rect 87210 21760 87290 21770
rect 87360 21760 87440 21770
rect 75640 21680 75650 21760
rect 75790 21680 75800 21760
rect 87140 21680 87150 21760
rect 87290 21680 87300 21760
rect 87440 21680 87450 21760
rect 87850 21690 87860 21770
rect 88170 21690 88180 21770
rect 88590 21690 88600 21770
rect 88910 21690 88920 21770
rect 89060 21760 89140 21770
rect 89210 21760 89290 21770
rect 100560 21760 100640 21770
rect 100710 21760 100790 21770
rect 100860 21760 100940 21770
rect 89140 21680 89150 21760
rect 89290 21680 89300 21760
rect 100640 21680 100650 21760
rect 100790 21680 100800 21760
rect 100940 21680 100950 21760
rect 101350 21690 101360 21770
rect 101670 21690 101680 21770
rect 102090 21690 102100 21770
rect 102410 21690 102420 21770
rect 102560 21760 102640 21770
rect 102710 21760 102790 21770
rect 114060 21760 114140 21770
rect 114210 21760 114290 21770
rect 114360 21760 114440 21770
rect 102640 21680 102650 21760
rect 102790 21680 102800 21760
rect 114140 21680 114150 21760
rect 114290 21680 114300 21760
rect 114440 21680 114450 21760
rect 114850 21690 114860 21770
rect 115170 21690 115180 21770
rect 115590 21690 115600 21770
rect 115910 21690 115920 21770
rect 116060 21760 116140 21770
rect 116210 21760 116290 21770
rect 127560 21760 127640 21770
rect 127710 21760 127790 21770
rect 127860 21760 127940 21770
rect 116140 21680 116150 21760
rect 116290 21680 116300 21760
rect 127640 21680 127650 21760
rect 127790 21680 127800 21760
rect 127940 21680 127950 21760
rect 128350 21690 128360 21770
rect 128670 21690 128680 21770
rect 129090 21690 129100 21770
rect 129410 21690 129420 21770
rect 129560 21760 129640 21770
rect 129710 21760 129790 21770
rect 141060 21760 141140 21770
rect 141210 21760 141290 21770
rect 141360 21760 141440 21770
rect 129640 21680 129650 21760
rect 129790 21680 129800 21760
rect 141140 21680 141150 21760
rect 141290 21680 141300 21760
rect 141440 21680 141450 21760
rect 60610 21610 60690 21620
rect 60930 21610 61010 21620
rect 61350 21610 61430 21620
rect 61670 21610 61750 21620
rect 74110 21610 74190 21620
rect 74430 21610 74510 21620
rect 74850 21610 74930 21620
rect 75170 21610 75250 21620
rect 87610 21610 87690 21620
rect 87930 21610 88010 21620
rect 88350 21610 88430 21620
rect 88670 21610 88750 21620
rect 101110 21610 101190 21620
rect 101430 21610 101510 21620
rect 101850 21610 101930 21620
rect 102170 21610 102250 21620
rect 114610 21610 114690 21620
rect 114930 21610 115010 21620
rect 115350 21610 115430 21620
rect 115670 21610 115750 21620
rect 128110 21610 128190 21620
rect 128430 21610 128510 21620
rect 128850 21610 128930 21620
rect 129170 21610 129250 21620
rect 59350 21580 59430 21590
rect 59500 21580 59580 21590
rect 59650 21580 59730 21590
rect 60060 21580 60140 21590
rect 60210 21580 60290 21590
rect 60360 21580 60440 21590
rect 59430 21500 59440 21580
rect 59580 21500 59590 21580
rect 59730 21500 59740 21580
rect 60140 21500 60150 21580
rect 60290 21500 60300 21580
rect 60440 21500 60450 21580
rect 60690 21530 60700 21610
rect 61010 21530 61020 21610
rect 61430 21530 61440 21610
rect 61750 21530 61760 21610
rect 62060 21580 62140 21590
rect 62210 21580 62290 21590
rect 73560 21580 73640 21590
rect 73710 21580 73790 21590
rect 73860 21580 73940 21590
rect 62140 21500 62150 21580
rect 62290 21500 62300 21580
rect 73640 21500 73650 21580
rect 73790 21500 73800 21580
rect 73940 21500 73950 21580
rect 74190 21530 74200 21610
rect 74510 21530 74520 21610
rect 74930 21530 74940 21610
rect 75250 21530 75260 21610
rect 75560 21580 75640 21590
rect 75710 21580 75790 21590
rect 87060 21580 87140 21590
rect 87210 21580 87290 21590
rect 87360 21580 87440 21590
rect 75640 21500 75650 21580
rect 75790 21500 75800 21580
rect 87140 21500 87150 21580
rect 87290 21500 87300 21580
rect 87440 21500 87450 21580
rect 87690 21530 87700 21610
rect 88010 21530 88020 21610
rect 88430 21530 88440 21610
rect 88750 21530 88760 21610
rect 89060 21580 89140 21590
rect 89210 21580 89290 21590
rect 100560 21580 100640 21590
rect 100710 21580 100790 21590
rect 100860 21580 100940 21590
rect 89140 21500 89150 21580
rect 89290 21500 89300 21580
rect 100640 21500 100650 21580
rect 100790 21500 100800 21580
rect 100940 21500 100950 21580
rect 101190 21530 101200 21610
rect 101510 21530 101520 21610
rect 101930 21530 101940 21610
rect 102250 21530 102260 21610
rect 102560 21580 102640 21590
rect 102710 21580 102790 21590
rect 114060 21580 114140 21590
rect 114210 21580 114290 21590
rect 114360 21580 114440 21590
rect 102640 21500 102650 21580
rect 102790 21500 102800 21580
rect 114140 21500 114150 21580
rect 114290 21500 114300 21580
rect 114440 21500 114450 21580
rect 114690 21530 114700 21610
rect 115010 21530 115020 21610
rect 115430 21530 115440 21610
rect 115750 21530 115760 21610
rect 116060 21580 116140 21590
rect 116210 21580 116290 21590
rect 127560 21580 127640 21590
rect 127710 21580 127790 21590
rect 127860 21580 127940 21590
rect 116140 21500 116150 21580
rect 116290 21500 116300 21580
rect 127640 21500 127650 21580
rect 127790 21500 127800 21580
rect 127940 21500 127950 21580
rect 128190 21530 128200 21610
rect 128510 21530 128520 21610
rect 128930 21530 128940 21610
rect 129250 21530 129260 21610
rect 129560 21580 129640 21590
rect 129710 21580 129790 21590
rect 141060 21580 141140 21590
rect 141210 21580 141290 21590
rect 141360 21580 141440 21590
rect 129640 21500 129650 21580
rect 129790 21500 129800 21580
rect 141140 21500 141150 21580
rect 141290 21500 141300 21580
rect 141440 21500 141450 21580
rect 60770 21450 60850 21460
rect 61090 21450 61170 21460
rect 61510 21450 61590 21460
rect 61830 21450 61910 21460
rect 74270 21450 74350 21460
rect 74590 21450 74670 21460
rect 75010 21450 75090 21460
rect 75330 21450 75410 21460
rect 87770 21450 87850 21460
rect 88090 21450 88170 21460
rect 88510 21450 88590 21460
rect 88830 21450 88910 21460
rect 101270 21450 101350 21460
rect 101590 21450 101670 21460
rect 102010 21450 102090 21460
rect 102330 21450 102410 21460
rect 114770 21450 114850 21460
rect 115090 21450 115170 21460
rect 115510 21450 115590 21460
rect 115830 21450 115910 21460
rect 128270 21450 128350 21460
rect 128590 21450 128670 21460
rect 129010 21450 129090 21460
rect 129330 21450 129410 21460
rect 59350 21400 59430 21410
rect 59500 21400 59580 21410
rect 59650 21400 59730 21410
rect 60060 21400 60140 21410
rect 60210 21400 60290 21410
rect 60360 21400 60440 21410
rect 59430 21320 59440 21400
rect 59580 21320 59590 21400
rect 59730 21320 59740 21400
rect 60140 21320 60150 21400
rect 60290 21320 60300 21400
rect 60440 21320 60450 21400
rect 60850 21370 60860 21450
rect 61170 21370 61180 21450
rect 61590 21370 61600 21450
rect 61910 21370 61920 21450
rect 62060 21400 62140 21410
rect 62210 21400 62290 21410
rect 73560 21400 73640 21410
rect 73710 21400 73790 21410
rect 73860 21400 73940 21410
rect 62140 21320 62150 21400
rect 62290 21320 62300 21400
rect 73640 21320 73650 21400
rect 73790 21320 73800 21400
rect 73940 21320 73950 21400
rect 74350 21370 74360 21450
rect 74670 21370 74680 21450
rect 75090 21370 75100 21450
rect 75410 21370 75420 21450
rect 75560 21400 75640 21410
rect 75710 21400 75790 21410
rect 87060 21400 87140 21410
rect 87210 21400 87290 21410
rect 87360 21400 87440 21410
rect 75640 21320 75650 21400
rect 75790 21320 75800 21400
rect 87140 21320 87150 21400
rect 87290 21320 87300 21400
rect 87440 21320 87450 21400
rect 87850 21370 87860 21450
rect 88170 21370 88180 21450
rect 88590 21370 88600 21450
rect 88910 21370 88920 21450
rect 89060 21400 89140 21410
rect 89210 21400 89290 21410
rect 100560 21400 100640 21410
rect 100710 21400 100790 21410
rect 100860 21400 100940 21410
rect 89140 21320 89150 21400
rect 89290 21320 89300 21400
rect 100640 21320 100650 21400
rect 100790 21320 100800 21400
rect 100940 21320 100950 21400
rect 101350 21370 101360 21450
rect 101670 21370 101680 21450
rect 102090 21370 102100 21450
rect 102410 21370 102420 21450
rect 102560 21400 102640 21410
rect 102710 21400 102790 21410
rect 114060 21400 114140 21410
rect 114210 21400 114290 21410
rect 114360 21400 114440 21410
rect 102640 21320 102650 21400
rect 102790 21320 102800 21400
rect 114140 21320 114150 21400
rect 114290 21320 114300 21400
rect 114440 21320 114450 21400
rect 114850 21370 114860 21450
rect 115170 21370 115180 21450
rect 115590 21370 115600 21450
rect 115910 21370 115920 21450
rect 116060 21400 116140 21410
rect 116210 21400 116290 21410
rect 127560 21400 127640 21410
rect 127710 21400 127790 21410
rect 127860 21400 127940 21410
rect 116140 21320 116150 21400
rect 116290 21320 116300 21400
rect 127640 21320 127650 21400
rect 127790 21320 127800 21400
rect 127940 21320 127950 21400
rect 128350 21370 128360 21450
rect 128670 21370 128680 21450
rect 129090 21370 129100 21450
rect 129410 21370 129420 21450
rect 129560 21400 129640 21410
rect 129710 21400 129790 21410
rect 141060 21400 141140 21410
rect 141210 21400 141290 21410
rect 141360 21400 141440 21410
rect 129640 21320 129650 21400
rect 129790 21320 129800 21400
rect 141140 21320 141150 21400
rect 141290 21320 141300 21400
rect 141440 21320 141450 21400
rect 60610 21290 60690 21300
rect 60930 21290 61010 21300
rect 61350 21290 61430 21300
rect 61670 21290 61750 21300
rect 74110 21290 74190 21300
rect 74430 21290 74510 21300
rect 74850 21290 74930 21300
rect 75170 21290 75250 21300
rect 87610 21290 87690 21300
rect 87930 21290 88010 21300
rect 88350 21290 88430 21300
rect 88670 21290 88750 21300
rect 101110 21290 101190 21300
rect 101430 21290 101510 21300
rect 101850 21290 101930 21300
rect 102170 21290 102250 21300
rect 114610 21290 114690 21300
rect 114930 21290 115010 21300
rect 115350 21290 115430 21300
rect 115670 21290 115750 21300
rect 128110 21290 128190 21300
rect 128430 21290 128510 21300
rect 128850 21290 128930 21300
rect 129170 21290 129250 21300
rect 59350 21220 59430 21230
rect 59500 21220 59580 21230
rect 59650 21220 59730 21230
rect 60060 21220 60140 21230
rect 60210 21220 60290 21230
rect 60360 21220 60440 21230
rect 59430 21140 59440 21220
rect 59580 21140 59590 21220
rect 59730 21140 59740 21220
rect 60140 21140 60150 21220
rect 60290 21140 60300 21220
rect 60440 21140 60450 21220
rect 60690 21210 60700 21290
rect 61010 21210 61020 21290
rect 61430 21210 61440 21290
rect 61750 21210 61760 21290
rect 62060 21220 62140 21230
rect 62210 21220 62290 21230
rect 73560 21220 73640 21230
rect 73710 21220 73790 21230
rect 73860 21220 73940 21230
rect 62140 21140 62150 21220
rect 62290 21140 62300 21220
rect 73640 21140 73650 21220
rect 73790 21140 73800 21220
rect 73940 21140 73950 21220
rect 74190 21210 74200 21290
rect 74510 21210 74520 21290
rect 74930 21210 74940 21290
rect 75250 21210 75260 21290
rect 75560 21220 75640 21230
rect 75710 21220 75790 21230
rect 87060 21220 87140 21230
rect 87210 21220 87290 21230
rect 87360 21220 87440 21230
rect 75640 21140 75650 21220
rect 75790 21140 75800 21220
rect 87140 21140 87150 21220
rect 87290 21140 87300 21220
rect 87440 21140 87450 21220
rect 87690 21210 87700 21290
rect 88010 21210 88020 21290
rect 88430 21210 88440 21290
rect 88750 21210 88760 21290
rect 89060 21220 89140 21230
rect 89210 21220 89290 21230
rect 100560 21220 100640 21230
rect 100710 21220 100790 21230
rect 100860 21220 100940 21230
rect 89140 21140 89150 21220
rect 89290 21140 89300 21220
rect 100640 21140 100650 21220
rect 100790 21140 100800 21220
rect 100940 21140 100950 21220
rect 101190 21210 101200 21290
rect 101510 21210 101520 21290
rect 101930 21210 101940 21290
rect 102250 21210 102260 21290
rect 102560 21220 102640 21230
rect 102710 21220 102790 21230
rect 114060 21220 114140 21230
rect 114210 21220 114290 21230
rect 114360 21220 114440 21230
rect 102640 21140 102650 21220
rect 102790 21140 102800 21220
rect 114140 21140 114150 21220
rect 114290 21140 114300 21220
rect 114440 21140 114450 21220
rect 114690 21210 114700 21290
rect 115010 21210 115020 21290
rect 115430 21210 115440 21290
rect 115750 21210 115760 21290
rect 116060 21220 116140 21230
rect 116210 21220 116290 21230
rect 127560 21220 127640 21230
rect 127710 21220 127790 21230
rect 127860 21220 127940 21230
rect 116140 21140 116150 21220
rect 116290 21140 116300 21220
rect 127640 21140 127650 21220
rect 127790 21140 127800 21220
rect 127940 21140 127950 21220
rect 128190 21210 128200 21290
rect 128510 21210 128520 21290
rect 128930 21210 128940 21290
rect 129250 21210 129260 21290
rect 129560 21220 129640 21230
rect 129710 21220 129790 21230
rect 141060 21220 141140 21230
rect 141210 21220 141290 21230
rect 141360 21220 141440 21230
rect 129640 21140 129650 21220
rect 129790 21140 129800 21220
rect 141140 21140 141150 21220
rect 141290 21140 141300 21220
rect 141440 21140 141450 21220
rect 60770 21130 60850 21140
rect 61090 21130 61170 21140
rect 61510 21130 61590 21140
rect 61830 21130 61910 21140
rect 74270 21130 74350 21140
rect 74590 21130 74670 21140
rect 75010 21130 75090 21140
rect 75330 21130 75410 21140
rect 87770 21130 87850 21140
rect 88090 21130 88170 21140
rect 88510 21130 88590 21140
rect 88830 21130 88910 21140
rect 101270 21130 101350 21140
rect 101590 21130 101670 21140
rect 102010 21130 102090 21140
rect 102330 21130 102410 21140
rect 114770 21130 114850 21140
rect 115090 21130 115170 21140
rect 115510 21130 115590 21140
rect 115830 21130 115910 21140
rect 128270 21130 128350 21140
rect 128590 21130 128670 21140
rect 129010 21130 129090 21140
rect 129330 21130 129410 21140
rect 60850 21050 60860 21130
rect 61170 21050 61180 21130
rect 61590 21050 61600 21130
rect 61910 21050 61920 21130
rect 74350 21050 74360 21130
rect 74670 21050 74680 21130
rect 75090 21050 75100 21130
rect 75410 21050 75420 21130
rect 87850 21050 87860 21130
rect 88170 21050 88180 21130
rect 88590 21050 88600 21130
rect 88910 21050 88920 21130
rect 101350 21050 101360 21130
rect 101670 21050 101680 21130
rect 102090 21050 102100 21130
rect 102410 21050 102420 21130
rect 114850 21050 114860 21130
rect 115170 21050 115180 21130
rect 115590 21050 115600 21130
rect 115910 21050 115920 21130
rect 128350 21050 128360 21130
rect 128670 21050 128680 21130
rect 129090 21050 129100 21130
rect 129410 21050 129420 21130
rect 59350 21040 59430 21050
rect 59500 21040 59580 21050
rect 59650 21040 59730 21050
rect 60060 21040 60140 21050
rect 60210 21040 60290 21050
rect 60360 21040 60440 21050
rect 62060 21040 62140 21050
rect 62210 21040 62290 21050
rect 73560 21040 73640 21050
rect 73710 21040 73790 21050
rect 73860 21040 73940 21050
rect 75560 21040 75640 21050
rect 75710 21040 75790 21050
rect 87060 21040 87140 21050
rect 87210 21040 87290 21050
rect 87360 21040 87440 21050
rect 89060 21040 89140 21050
rect 89210 21040 89290 21050
rect 100560 21040 100640 21050
rect 100710 21040 100790 21050
rect 100860 21040 100940 21050
rect 102560 21040 102640 21050
rect 102710 21040 102790 21050
rect 114060 21040 114140 21050
rect 114210 21040 114290 21050
rect 114360 21040 114440 21050
rect 116060 21040 116140 21050
rect 116210 21040 116290 21050
rect 127560 21040 127640 21050
rect 127710 21040 127790 21050
rect 127860 21040 127940 21050
rect 129560 21040 129640 21050
rect 129710 21040 129790 21050
rect 141060 21040 141140 21050
rect 141210 21040 141290 21050
rect 141360 21040 141440 21050
rect 59430 20960 59440 21040
rect 59580 20960 59590 21040
rect 59730 20960 59740 21040
rect 60140 20960 60150 21040
rect 60290 20960 60300 21040
rect 60440 20960 60450 21040
rect 60610 20970 60690 20980
rect 60930 20970 61010 20980
rect 61350 20970 61430 20980
rect 61670 20970 61750 20980
rect 60690 20890 60700 20970
rect 61010 20890 61020 20970
rect 61430 20890 61440 20970
rect 61750 20890 61760 20970
rect 62140 20960 62150 21040
rect 62290 20960 62300 21040
rect 73640 20960 73650 21040
rect 73790 20960 73800 21040
rect 73940 20960 73950 21040
rect 74110 20970 74190 20980
rect 74430 20970 74510 20980
rect 74850 20970 74930 20980
rect 75170 20970 75250 20980
rect 74190 20890 74200 20970
rect 74510 20890 74520 20970
rect 74930 20890 74940 20970
rect 75250 20890 75260 20970
rect 75640 20960 75650 21040
rect 75790 20960 75800 21040
rect 87140 20960 87150 21040
rect 87290 20960 87300 21040
rect 87440 20960 87450 21040
rect 87610 20970 87690 20980
rect 87930 20970 88010 20980
rect 88350 20970 88430 20980
rect 88670 20970 88750 20980
rect 87690 20890 87700 20970
rect 88010 20890 88020 20970
rect 88430 20890 88440 20970
rect 88750 20890 88760 20970
rect 89140 20960 89150 21040
rect 89290 20960 89300 21040
rect 100640 20960 100650 21040
rect 100790 20960 100800 21040
rect 100940 20960 100950 21040
rect 101110 20970 101190 20980
rect 101430 20970 101510 20980
rect 101850 20970 101930 20980
rect 102170 20970 102250 20980
rect 101190 20890 101200 20970
rect 101510 20890 101520 20970
rect 101930 20890 101940 20970
rect 102250 20890 102260 20970
rect 102640 20960 102650 21040
rect 102790 20960 102800 21040
rect 114140 20960 114150 21040
rect 114290 20960 114300 21040
rect 114440 20960 114450 21040
rect 114610 20970 114690 20980
rect 114930 20970 115010 20980
rect 115350 20970 115430 20980
rect 115670 20970 115750 20980
rect 114690 20890 114700 20970
rect 115010 20890 115020 20970
rect 115430 20890 115440 20970
rect 115750 20890 115760 20970
rect 116140 20960 116150 21040
rect 116290 20960 116300 21040
rect 127640 20960 127650 21040
rect 127790 20960 127800 21040
rect 127940 20960 127950 21040
rect 128110 20970 128190 20980
rect 128430 20970 128510 20980
rect 128850 20970 128930 20980
rect 129170 20970 129250 20980
rect 128190 20890 128200 20970
rect 128510 20890 128520 20970
rect 128930 20890 128940 20970
rect 129250 20890 129260 20970
rect 129640 20960 129650 21040
rect 129790 20960 129800 21040
rect 141140 20960 141150 21040
rect 141290 20960 141300 21040
rect 141440 20960 141450 21040
rect 59350 20860 59430 20870
rect 59500 20860 59580 20870
rect 59650 20860 59730 20870
rect 60060 20860 60140 20870
rect 60210 20860 60290 20870
rect 60360 20860 60440 20870
rect 62060 20860 62140 20870
rect 62210 20860 62290 20870
rect 73560 20860 73640 20870
rect 73710 20860 73790 20870
rect 73860 20860 73940 20870
rect 75560 20860 75640 20870
rect 75710 20860 75790 20870
rect 87060 20860 87140 20870
rect 87210 20860 87290 20870
rect 87360 20860 87440 20870
rect 89060 20860 89140 20870
rect 89210 20860 89290 20870
rect 100560 20860 100640 20870
rect 100710 20860 100790 20870
rect 100860 20860 100940 20870
rect 102560 20860 102640 20870
rect 102710 20860 102790 20870
rect 114060 20860 114140 20870
rect 114210 20860 114290 20870
rect 114360 20860 114440 20870
rect 116060 20860 116140 20870
rect 116210 20860 116290 20870
rect 127560 20860 127640 20870
rect 127710 20860 127790 20870
rect 127860 20860 127940 20870
rect 129560 20860 129640 20870
rect 129710 20860 129790 20870
rect 141060 20860 141140 20870
rect 141210 20860 141290 20870
rect 141360 20860 141440 20870
rect 59430 20780 59440 20860
rect 59580 20780 59590 20860
rect 59730 20780 59740 20860
rect 60140 20780 60150 20860
rect 60290 20780 60300 20860
rect 60440 20780 60450 20860
rect 60770 20810 60850 20820
rect 61090 20810 61170 20820
rect 61510 20810 61590 20820
rect 61830 20810 61910 20820
rect 60850 20730 60860 20810
rect 61170 20730 61180 20810
rect 61590 20730 61600 20810
rect 61910 20730 61920 20810
rect 62140 20780 62150 20860
rect 62290 20780 62300 20860
rect 73640 20780 73650 20860
rect 73790 20780 73800 20860
rect 73940 20780 73950 20860
rect 74270 20810 74350 20820
rect 74590 20810 74670 20820
rect 75010 20810 75090 20820
rect 75330 20810 75410 20820
rect 74350 20730 74360 20810
rect 74670 20730 74680 20810
rect 75090 20730 75100 20810
rect 75410 20730 75420 20810
rect 75640 20780 75650 20860
rect 75790 20780 75800 20860
rect 87140 20780 87150 20860
rect 87290 20780 87300 20860
rect 87440 20780 87450 20860
rect 87770 20810 87850 20820
rect 88090 20810 88170 20820
rect 88510 20810 88590 20820
rect 88830 20810 88910 20820
rect 87850 20730 87860 20810
rect 88170 20730 88180 20810
rect 88590 20730 88600 20810
rect 88910 20730 88920 20810
rect 89140 20780 89150 20860
rect 89290 20780 89300 20860
rect 100640 20780 100650 20860
rect 100790 20780 100800 20860
rect 100940 20780 100950 20860
rect 101270 20810 101350 20820
rect 101590 20810 101670 20820
rect 102010 20810 102090 20820
rect 102330 20810 102410 20820
rect 101350 20730 101360 20810
rect 101670 20730 101680 20810
rect 102090 20730 102100 20810
rect 102410 20730 102420 20810
rect 102640 20780 102650 20860
rect 102790 20780 102800 20860
rect 114140 20780 114150 20860
rect 114290 20780 114300 20860
rect 114440 20780 114450 20860
rect 114770 20810 114850 20820
rect 115090 20810 115170 20820
rect 115510 20810 115590 20820
rect 115830 20810 115910 20820
rect 114850 20730 114860 20810
rect 115170 20730 115180 20810
rect 115590 20730 115600 20810
rect 115910 20730 115920 20810
rect 116140 20780 116150 20860
rect 116290 20780 116300 20860
rect 127640 20780 127650 20860
rect 127790 20780 127800 20860
rect 127940 20780 127950 20860
rect 128270 20810 128350 20820
rect 128590 20810 128670 20820
rect 129010 20810 129090 20820
rect 129330 20810 129410 20820
rect 128350 20730 128360 20810
rect 128670 20730 128680 20810
rect 129090 20730 129100 20810
rect 129410 20730 129420 20810
rect 129640 20780 129650 20860
rect 129790 20780 129800 20860
rect 141140 20780 141150 20860
rect 141290 20780 141300 20860
rect 141440 20780 141450 20860
rect 59350 20680 59430 20690
rect 59500 20680 59580 20690
rect 59650 20680 59730 20690
rect 60060 20680 60140 20690
rect 60210 20680 60290 20690
rect 60360 20680 60440 20690
rect 62060 20680 62140 20690
rect 62210 20680 62290 20690
rect 73560 20680 73640 20690
rect 73710 20680 73790 20690
rect 73860 20680 73940 20690
rect 75560 20680 75640 20690
rect 75710 20680 75790 20690
rect 87060 20680 87140 20690
rect 87210 20680 87290 20690
rect 87360 20680 87440 20690
rect 89060 20680 89140 20690
rect 89210 20680 89290 20690
rect 100560 20680 100640 20690
rect 100710 20680 100790 20690
rect 100860 20680 100940 20690
rect 102560 20680 102640 20690
rect 102710 20680 102790 20690
rect 114060 20680 114140 20690
rect 114210 20680 114290 20690
rect 114360 20680 114440 20690
rect 116060 20680 116140 20690
rect 116210 20680 116290 20690
rect 127560 20680 127640 20690
rect 127710 20680 127790 20690
rect 127860 20680 127940 20690
rect 129560 20680 129640 20690
rect 129710 20680 129790 20690
rect 141060 20680 141140 20690
rect 141210 20680 141290 20690
rect 141360 20680 141440 20690
rect 59430 20600 59440 20680
rect 59580 20600 59590 20680
rect 59730 20600 59740 20680
rect 60140 20600 60150 20680
rect 60290 20600 60300 20680
rect 60440 20600 60450 20680
rect 60610 20650 60690 20660
rect 60930 20650 61010 20660
rect 61350 20650 61430 20660
rect 61670 20650 61750 20660
rect 60690 20570 60700 20650
rect 61010 20570 61020 20650
rect 61430 20570 61440 20650
rect 61750 20570 61760 20650
rect 62140 20600 62150 20680
rect 62290 20600 62300 20680
rect 73640 20600 73650 20680
rect 73790 20600 73800 20680
rect 73940 20600 73950 20680
rect 74110 20650 74190 20660
rect 74430 20650 74510 20660
rect 74850 20650 74930 20660
rect 75170 20650 75250 20660
rect 74190 20570 74200 20650
rect 74510 20570 74520 20650
rect 74930 20570 74940 20650
rect 75250 20570 75260 20650
rect 75640 20600 75650 20680
rect 75790 20600 75800 20680
rect 87140 20600 87150 20680
rect 87290 20600 87300 20680
rect 87440 20600 87450 20680
rect 87610 20650 87690 20660
rect 87930 20650 88010 20660
rect 88350 20650 88430 20660
rect 88670 20650 88750 20660
rect 87690 20570 87700 20650
rect 88010 20570 88020 20650
rect 88430 20570 88440 20650
rect 88750 20570 88760 20650
rect 89140 20600 89150 20680
rect 89290 20600 89300 20680
rect 100640 20600 100650 20680
rect 100790 20600 100800 20680
rect 100940 20600 100950 20680
rect 101110 20650 101190 20660
rect 101430 20650 101510 20660
rect 101850 20650 101930 20660
rect 102170 20650 102250 20660
rect 101190 20570 101200 20650
rect 101510 20570 101520 20650
rect 101930 20570 101940 20650
rect 102250 20570 102260 20650
rect 102640 20600 102650 20680
rect 102790 20600 102800 20680
rect 114140 20600 114150 20680
rect 114290 20600 114300 20680
rect 114440 20600 114450 20680
rect 114610 20650 114690 20660
rect 114930 20650 115010 20660
rect 115350 20650 115430 20660
rect 115670 20650 115750 20660
rect 114690 20570 114700 20650
rect 115010 20570 115020 20650
rect 115430 20570 115440 20650
rect 115750 20570 115760 20650
rect 116140 20600 116150 20680
rect 116290 20600 116300 20680
rect 127640 20600 127650 20680
rect 127790 20600 127800 20680
rect 127940 20600 127950 20680
rect 128110 20650 128190 20660
rect 128430 20650 128510 20660
rect 128850 20650 128930 20660
rect 129170 20650 129250 20660
rect 128190 20570 128200 20650
rect 128510 20570 128520 20650
rect 128930 20570 128940 20650
rect 129250 20570 129260 20650
rect 129640 20600 129650 20680
rect 129790 20600 129800 20680
rect 141140 20600 141150 20680
rect 141290 20600 141300 20680
rect 141440 20600 141450 20680
rect 59350 20500 59430 20510
rect 59500 20500 59580 20510
rect 59650 20500 59730 20510
rect 60060 20500 60140 20510
rect 60210 20500 60290 20510
rect 60360 20500 60440 20510
rect 62060 20500 62140 20510
rect 62210 20500 62290 20510
rect 73560 20500 73640 20510
rect 73710 20500 73790 20510
rect 73860 20500 73940 20510
rect 75560 20500 75640 20510
rect 75710 20500 75790 20510
rect 87060 20500 87140 20510
rect 87210 20500 87290 20510
rect 87360 20500 87440 20510
rect 89060 20500 89140 20510
rect 89210 20500 89290 20510
rect 100560 20500 100640 20510
rect 100710 20500 100790 20510
rect 100860 20500 100940 20510
rect 102560 20500 102640 20510
rect 102710 20500 102790 20510
rect 114060 20500 114140 20510
rect 114210 20500 114290 20510
rect 114360 20500 114440 20510
rect 116060 20500 116140 20510
rect 116210 20500 116290 20510
rect 127560 20500 127640 20510
rect 127710 20500 127790 20510
rect 127860 20500 127940 20510
rect 129560 20500 129640 20510
rect 129710 20500 129790 20510
rect 141060 20500 141140 20510
rect 141210 20500 141290 20510
rect 141360 20500 141440 20510
rect 59430 20420 59440 20500
rect 59580 20420 59590 20500
rect 59730 20420 59740 20500
rect 60140 20420 60150 20500
rect 60290 20420 60300 20500
rect 60440 20420 60450 20500
rect 60770 20490 60850 20500
rect 61090 20490 61170 20500
rect 61510 20490 61590 20500
rect 61830 20490 61910 20500
rect 60850 20410 60860 20490
rect 61170 20410 61180 20490
rect 61590 20410 61600 20490
rect 61910 20410 61920 20490
rect 62140 20420 62150 20500
rect 62290 20420 62300 20500
rect 73640 20420 73650 20500
rect 73790 20420 73800 20500
rect 73940 20420 73950 20500
rect 74270 20490 74350 20500
rect 74590 20490 74670 20500
rect 75010 20490 75090 20500
rect 75330 20490 75410 20500
rect 74350 20410 74360 20490
rect 74670 20410 74680 20490
rect 75090 20410 75100 20490
rect 75410 20410 75420 20490
rect 75640 20420 75650 20500
rect 75790 20420 75800 20500
rect 87140 20420 87150 20500
rect 87290 20420 87300 20500
rect 87440 20420 87450 20500
rect 87770 20490 87850 20500
rect 88090 20490 88170 20500
rect 88510 20490 88590 20500
rect 88830 20490 88910 20500
rect 87850 20410 87860 20490
rect 88170 20410 88180 20490
rect 88590 20410 88600 20490
rect 88910 20410 88920 20490
rect 89140 20420 89150 20500
rect 89290 20420 89300 20500
rect 100640 20420 100650 20500
rect 100790 20420 100800 20500
rect 100940 20420 100950 20500
rect 101270 20490 101350 20500
rect 101590 20490 101670 20500
rect 102010 20490 102090 20500
rect 102330 20490 102410 20500
rect 101350 20410 101360 20490
rect 101670 20410 101680 20490
rect 102090 20410 102100 20490
rect 102410 20410 102420 20490
rect 102640 20420 102650 20500
rect 102790 20420 102800 20500
rect 114140 20420 114150 20500
rect 114290 20420 114300 20500
rect 114440 20420 114450 20500
rect 114770 20490 114850 20500
rect 115090 20490 115170 20500
rect 115510 20490 115590 20500
rect 115830 20490 115910 20500
rect 114850 20410 114860 20490
rect 115170 20410 115180 20490
rect 115590 20410 115600 20490
rect 115910 20410 115920 20490
rect 116140 20420 116150 20500
rect 116290 20420 116300 20500
rect 127640 20420 127650 20500
rect 127790 20420 127800 20500
rect 127940 20420 127950 20500
rect 128270 20490 128350 20500
rect 128590 20490 128670 20500
rect 129010 20490 129090 20500
rect 129330 20490 129410 20500
rect 128350 20410 128360 20490
rect 128670 20410 128680 20490
rect 129090 20410 129100 20490
rect 129410 20410 129420 20490
rect 129640 20420 129650 20500
rect 129790 20420 129800 20500
rect 141140 20420 141150 20500
rect 141290 20420 141300 20500
rect 141440 20420 141450 20500
rect 60610 20330 60690 20340
rect 60930 20330 61010 20340
rect 61350 20330 61430 20340
rect 61670 20330 61750 20340
rect 74110 20330 74190 20340
rect 74430 20330 74510 20340
rect 74850 20330 74930 20340
rect 75170 20330 75250 20340
rect 87610 20330 87690 20340
rect 87930 20330 88010 20340
rect 88350 20330 88430 20340
rect 88670 20330 88750 20340
rect 101110 20330 101190 20340
rect 101430 20330 101510 20340
rect 101850 20330 101930 20340
rect 102170 20330 102250 20340
rect 114610 20330 114690 20340
rect 114930 20330 115010 20340
rect 115350 20330 115430 20340
rect 115670 20330 115750 20340
rect 128110 20330 128190 20340
rect 128430 20330 128510 20340
rect 128850 20330 128930 20340
rect 129170 20330 129250 20340
rect 59350 20320 59430 20330
rect 59500 20320 59580 20330
rect 59650 20320 59730 20330
rect 60060 20320 60140 20330
rect 60210 20320 60290 20330
rect 60360 20320 60440 20330
rect 59430 20240 59440 20320
rect 59580 20240 59590 20320
rect 59730 20240 59740 20320
rect 60140 20240 60150 20320
rect 60290 20240 60300 20320
rect 60440 20240 60450 20320
rect 60690 20250 60700 20330
rect 61010 20250 61020 20330
rect 61430 20250 61440 20330
rect 61750 20250 61760 20330
rect 62060 20320 62140 20330
rect 62210 20320 62290 20330
rect 73560 20320 73640 20330
rect 73710 20320 73790 20330
rect 73860 20320 73940 20330
rect 62140 20240 62150 20320
rect 62290 20240 62300 20320
rect 73640 20240 73650 20320
rect 73790 20240 73800 20320
rect 73940 20240 73950 20320
rect 74190 20250 74200 20330
rect 74510 20250 74520 20330
rect 74930 20250 74940 20330
rect 75250 20250 75260 20330
rect 75560 20320 75640 20330
rect 75710 20320 75790 20330
rect 87060 20320 87140 20330
rect 87210 20320 87290 20330
rect 87360 20320 87440 20330
rect 75640 20240 75650 20320
rect 75790 20240 75800 20320
rect 87140 20240 87150 20320
rect 87290 20240 87300 20320
rect 87440 20240 87450 20320
rect 87690 20250 87700 20330
rect 88010 20250 88020 20330
rect 88430 20250 88440 20330
rect 88750 20250 88760 20330
rect 89060 20320 89140 20330
rect 89210 20320 89290 20330
rect 100560 20320 100640 20330
rect 100710 20320 100790 20330
rect 100860 20320 100940 20330
rect 89140 20240 89150 20320
rect 89290 20240 89300 20320
rect 100640 20240 100650 20320
rect 100790 20240 100800 20320
rect 100940 20240 100950 20320
rect 101190 20250 101200 20330
rect 101510 20250 101520 20330
rect 101930 20250 101940 20330
rect 102250 20250 102260 20330
rect 102560 20320 102640 20330
rect 102710 20320 102790 20330
rect 114060 20320 114140 20330
rect 114210 20320 114290 20330
rect 114360 20320 114440 20330
rect 102640 20240 102650 20320
rect 102790 20240 102800 20320
rect 114140 20240 114150 20320
rect 114290 20240 114300 20320
rect 114440 20240 114450 20320
rect 114690 20250 114700 20330
rect 115010 20250 115020 20330
rect 115430 20250 115440 20330
rect 115750 20250 115760 20330
rect 116060 20320 116140 20330
rect 116210 20320 116290 20330
rect 127560 20320 127640 20330
rect 127710 20320 127790 20330
rect 127860 20320 127940 20330
rect 116140 20240 116150 20320
rect 116290 20240 116300 20320
rect 127640 20240 127650 20320
rect 127790 20240 127800 20320
rect 127940 20240 127950 20320
rect 128190 20250 128200 20330
rect 128510 20250 128520 20330
rect 128930 20250 128940 20330
rect 129250 20250 129260 20330
rect 129560 20320 129640 20330
rect 129710 20320 129790 20330
rect 141060 20320 141140 20330
rect 141210 20320 141290 20330
rect 141360 20320 141440 20330
rect 129640 20240 129650 20320
rect 129790 20240 129800 20320
rect 141140 20240 141150 20320
rect 141290 20240 141300 20320
rect 141440 20240 141450 20320
rect 60770 20170 60850 20180
rect 61090 20170 61170 20180
rect 61510 20170 61590 20180
rect 61830 20170 61910 20180
rect 74270 20170 74350 20180
rect 74590 20170 74670 20180
rect 75010 20170 75090 20180
rect 75330 20170 75410 20180
rect 87770 20170 87850 20180
rect 88090 20170 88170 20180
rect 88510 20170 88590 20180
rect 88830 20170 88910 20180
rect 101270 20170 101350 20180
rect 101590 20170 101670 20180
rect 102010 20170 102090 20180
rect 102330 20170 102410 20180
rect 114770 20170 114850 20180
rect 115090 20170 115170 20180
rect 115510 20170 115590 20180
rect 115830 20170 115910 20180
rect 128270 20170 128350 20180
rect 128590 20170 128670 20180
rect 129010 20170 129090 20180
rect 129330 20170 129410 20180
rect 59350 20140 59430 20150
rect 59500 20140 59580 20150
rect 59650 20140 59730 20150
rect 60060 20140 60140 20150
rect 60210 20140 60290 20150
rect 60360 20140 60440 20150
rect 59430 20060 59440 20140
rect 59580 20060 59590 20140
rect 59730 20060 59740 20140
rect 60140 20060 60150 20140
rect 60290 20060 60300 20140
rect 60440 20060 60450 20140
rect 60850 20090 60860 20170
rect 61170 20090 61180 20170
rect 61590 20090 61600 20170
rect 61910 20090 61920 20170
rect 62060 20140 62140 20150
rect 62210 20140 62290 20150
rect 73560 20140 73640 20150
rect 73710 20140 73790 20150
rect 73860 20140 73940 20150
rect 62140 20060 62150 20140
rect 62290 20060 62300 20140
rect 73640 20060 73650 20140
rect 73790 20060 73800 20140
rect 73940 20060 73950 20140
rect 74350 20090 74360 20170
rect 74670 20090 74680 20170
rect 75090 20090 75100 20170
rect 75410 20090 75420 20170
rect 75560 20140 75640 20150
rect 75710 20140 75790 20150
rect 87060 20140 87140 20150
rect 87210 20140 87290 20150
rect 87360 20140 87440 20150
rect 75640 20060 75650 20140
rect 75790 20060 75800 20140
rect 87140 20060 87150 20140
rect 87290 20060 87300 20140
rect 87440 20060 87450 20140
rect 87850 20090 87860 20170
rect 88170 20090 88180 20170
rect 88590 20090 88600 20170
rect 88910 20090 88920 20170
rect 89060 20140 89140 20150
rect 89210 20140 89290 20150
rect 100560 20140 100640 20150
rect 100710 20140 100790 20150
rect 100860 20140 100940 20150
rect 89140 20060 89150 20140
rect 89290 20060 89300 20140
rect 100640 20060 100650 20140
rect 100790 20060 100800 20140
rect 100940 20060 100950 20140
rect 101350 20090 101360 20170
rect 101670 20090 101680 20170
rect 102090 20090 102100 20170
rect 102410 20090 102420 20170
rect 102560 20140 102640 20150
rect 102710 20140 102790 20150
rect 114060 20140 114140 20150
rect 114210 20140 114290 20150
rect 114360 20140 114440 20150
rect 102640 20060 102650 20140
rect 102790 20060 102800 20140
rect 114140 20060 114150 20140
rect 114290 20060 114300 20140
rect 114440 20060 114450 20140
rect 114850 20090 114860 20170
rect 115170 20090 115180 20170
rect 115590 20090 115600 20170
rect 115910 20090 115920 20170
rect 116060 20140 116140 20150
rect 116210 20140 116290 20150
rect 127560 20140 127640 20150
rect 127710 20140 127790 20150
rect 127860 20140 127940 20150
rect 116140 20060 116150 20140
rect 116290 20060 116300 20140
rect 127640 20060 127650 20140
rect 127790 20060 127800 20140
rect 127940 20060 127950 20140
rect 128350 20090 128360 20170
rect 128670 20090 128680 20170
rect 129090 20090 129100 20170
rect 129410 20090 129420 20170
rect 129560 20140 129640 20150
rect 129710 20140 129790 20150
rect 141060 20140 141140 20150
rect 141210 20140 141290 20150
rect 141360 20140 141440 20150
rect 129640 20060 129650 20140
rect 129790 20060 129800 20140
rect 141140 20060 141150 20140
rect 141290 20060 141300 20140
rect 141440 20060 141450 20140
rect 60610 20010 60690 20020
rect 60930 20010 61010 20020
rect 61350 20010 61430 20020
rect 61670 20010 61750 20020
rect 74110 20010 74190 20020
rect 74430 20010 74510 20020
rect 74850 20010 74930 20020
rect 75170 20010 75250 20020
rect 87610 20010 87690 20020
rect 87930 20010 88010 20020
rect 88350 20010 88430 20020
rect 88670 20010 88750 20020
rect 101110 20010 101190 20020
rect 101430 20010 101510 20020
rect 101850 20010 101930 20020
rect 102170 20010 102250 20020
rect 114610 20010 114690 20020
rect 114930 20010 115010 20020
rect 115350 20010 115430 20020
rect 115670 20010 115750 20020
rect 128110 20010 128190 20020
rect 128430 20010 128510 20020
rect 128850 20010 128930 20020
rect 129170 20010 129250 20020
rect 59350 19960 59430 19970
rect 59500 19960 59580 19970
rect 59650 19960 59730 19970
rect 60060 19960 60140 19970
rect 60210 19960 60290 19970
rect 60360 19960 60440 19970
rect 59430 19880 59440 19960
rect 59580 19880 59590 19960
rect 59730 19880 59740 19960
rect 60140 19880 60150 19960
rect 60290 19880 60300 19960
rect 60440 19880 60450 19960
rect 60690 19930 60700 20010
rect 61010 19930 61020 20010
rect 61430 19930 61440 20010
rect 61750 19930 61760 20010
rect 62060 19960 62140 19970
rect 62210 19960 62290 19970
rect 73560 19960 73640 19970
rect 73710 19960 73790 19970
rect 73860 19960 73940 19970
rect 62140 19880 62150 19960
rect 62290 19880 62300 19960
rect 73640 19880 73650 19960
rect 73790 19880 73800 19960
rect 73940 19880 73950 19960
rect 74190 19930 74200 20010
rect 74510 19930 74520 20010
rect 74930 19930 74940 20010
rect 75250 19930 75260 20010
rect 75560 19960 75640 19970
rect 75710 19960 75790 19970
rect 87060 19960 87140 19970
rect 87210 19960 87290 19970
rect 87360 19960 87440 19970
rect 75640 19880 75650 19960
rect 75790 19880 75800 19960
rect 87140 19880 87150 19960
rect 87290 19880 87300 19960
rect 87440 19880 87450 19960
rect 87690 19930 87700 20010
rect 88010 19930 88020 20010
rect 88430 19930 88440 20010
rect 88750 19930 88760 20010
rect 89060 19960 89140 19970
rect 89210 19960 89290 19970
rect 100560 19960 100640 19970
rect 100710 19960 100790 19970
rect 100860 19960 100940 19970
rect 89140 19880 89150 19960
rect 89290 19880 89300 19960
rect 100640 19880 100650 19960
rect 100790 19880 100800 19960
rect 100940 19880 100950 19960
rect 101190 19930 101200 20010
rect 101510 19930 101520 20010
rect 101930 19930 101940 20010
rect 102250 19930 102260 20010
rect 102560 19960 102640 19970
rect 102710 19960 102790 19970
rect 114060 19960 114140 19970
rect 114210 19960 114290 19970
rect 114360 19960 114440 19970
rect 102640 19880 102650 19960
rect 102790 19880 102800 19960
rect 114140 19880 114150 19960
rect 114290 19880 114300 19960
rect 114440 19880 114450 19960
rect 114690 19930 114700 20010
rect 115010 19930 115020 20010
rect 115430 19930 115440 20010
rect 115750 19930 115760 20010
rect 116060 19960 116140 19970
rect 116210 19960 116290 19970
rect 127560 19960 127640 19970
rect 127710 19960 127790 19970
rect 127860 19960 127940 19970
rect 116140 19880 116150 19960
rect 116290 19880 116300 19960
rect 127640 19880 127650 19960
rect 127790 19880 127800 19960
rect 127940 19880 127950 19960
rect 128190 19930 128200 20010
rect 128510 19930 128520 20010
rect 128930 19930 128940 20010
rect 129250 19930 129260 20010
rect 129560 19960 129640 19970
rect 129710 19960 129790 19970
rect 141060 19960 141140 19970
rect 141210 19960 141290 19970
rect 141360 19960 141440 19970
rect 129640 19880 129650 19960
rect 129790 19880 129800 19960
rect 141140 19880 141150 19960
rect 141290 19880 141300 19960
rect 141440 19880 141450 19960
rect 60770 19850 60850 19860
rect 61090 19850 61170 19860
rect 61510 19850 61590 19860
rect 61830 19850 61910 19860
rect 74270 19850 74350 19860
rect 74590 19850 74670 19860
rect 75010 19850 75090 19860
rect 75330 19850 75410 19860
rect 87770 19850 87850 19860
rect 88090 19850 88170 19860
rect 88510 19850 88590 19860
rect 88830 19850 88910 19860
rect 101270 19850 101350 19860
rect 101590 19850 101670 19860
rect 102010 19850 102090 19860
rect 102330 19850 102410 19860
rect 114770 19850 114850 19860
rect 115090 19850 115170 19860
rect 115510 19850 115590 19860
rect 115830 19850 115910 19860
rect 128270 19850 128350 19860
rect 128590 19850 128670 19860
rect 129010 19850 129090 19860
rect 129330 19850 129410 19860
rect 48500 19780 48640 19790
rect 48710 19780 48790 19790
rect 60060 19780 60140 19790
rect 60210 19780 60290 19790
rect 60360 19780 60440 19790
rect 44065 19690 44145 19700
rect 44385 19690 44465 19700
rect 44705 19690 44785 19700
rect 45025 19690 45105 19700
rect 45345 19690 45425 19700
rect 45665 19690 45745 19700
rect 45985 19690 46065 19700
rect 46305 19690 46385 19700
rect 46625 19690 46705 19700
rect 46945 19690 47025 19700
rect 47265 19690 47345 19700
rect 47585 19690 47665 19700
rect 47905 19690 47985 19700
rect 48225 19690 48305 19700
rect 42950 19620 42980 19630
rect 43220 19620 43300 19630
rect 42980 19540 42990 19620
rect 43300 19540 43310 19620
rect 44145 19610 44155 19690
rect 44465 19610 44475 19690
rect 44785 19610 44795 19690
rect 45105 19610 45115 19690
rect 45425 19610 45435 19690
rect 45745 19610 45755 19690
rect 46065 19610 46075 19690
rect 46385 19610 46395 19690
rect 46705 19610 46715 19690
rect 47025 19610 47035 19690
rect 47345 19610 47355 19690
rect 47665 19610 47675 19690
rect 47985 19610 47995 19690
rect 48305 19610 48315 19690
rect 48500 19610 48605 19780
rect 48640 19700 48650 19780
rect 48790 19700 48800 19780
rect 60140 19700 60150 19780
rect 60290 19700 60300 19780
rect 60440 19700 60450 19780
rect 60850 19770 60860 19850
rect 61170 19770 61180 19850
rect 61590 19770 61600 19850
rect 61910 19770 61920 19850
rect 62060 19780 62140 19790
rect 62210 19780 62290 19790
rect 73560 19780 73640 19790
rect 73710 19780 73790 19790
rect 73860 19780 73940 19790
rect 62140 19700 62150 19780
rect 62290 19700 62300 19780
rect 73640 19700 73650 19780
rect 73790 19700 73800 19780
rect 73940 19700 73950 19780
rect 74350 19770 74360 19850
rect 74670 19770 74680 19850
rect 75090 19770 75100 19850
rect 75410 19770 75420 19850
rect 75560 19780 75640 19790
rect 75710 19780 75790 19790
rect 87060 19780 87140 19790
rect 87210 19780 87290 19790
rect 87360 19780 87440 19790
rect 75640 19700 75650 19780
rect 75790 19700 75800 19780
rect 87140 19700 87150 19780
rect 87290 19700 87300 19780
rect 87440 19700 87450 19780
rect 87850 19770 87860 19850
rect 88170 19770 88180 19850
rect 88590 19770 88600 19850
rect 88910 19770 88920 19850
rect 89060 19780 89140 19790
rect 89210 19780 89290 19790
rect 100560 19780 100640 19790
rect 100710 19780 100790 19790
rect 100860 19780 100940 19790
rect 89140 19700 89150 19780
rect 89290 19700 89300 19780
rect 100640 19700 100650 19780
rect 100790 19700 100800 19780
rect 100940 19700 100950 19780
rect 101350 19770 101360 19850
rect 101670 19770 101680 19850
rect 102090 19770 102100 19850
rect 102410 19770 102420 19850
rect 102560 19780 102640 19790
rect 102710 19780 102790 19790
rect 114060 19780 114140 19790
rect 114210 19780 114290 19790
rect 114360 19780 114440 19790
rect 102640 19700 102650 19780
rect 102790 19700 102800 19780
rect 114140 19700 114150 19780
rect 114290 19700 114300 19780
rect 114440 19700 114450 19780
rect 114850 19770 114860 19850
rect 115170 19770 115180 19850
rect 115590 19770 115600 19850
rect 115910 19770 115920 19850
rect 116060 19780 116140 19790
rect 116210 19780 116290 19790
rect 127560 19780 127640 19790
rect 127710 19780 127790 19790
rect 127860 19780 127940 19790
rect 116140 19700 116150 19780
rect 116290 19700 116300 19780
rect 127640 19700 127650 19780
rect 127790 19700 127800 19780
rect 127940 19700 127950 19780
rect 128350 19770 128360 19850
rect 128670 19770 128680 19850
rect 129090 19770 129100 19850
rect 129410 19770 129420 19850
rect 129560 19780 129640 19790
rect 129710 19780 129790 19790
rect 141060 19780 141140 19790
rect 141210 19780 141290 19790
rect 141360 19780 141440 19790
rect 129640 19700 129650 19780
rect 129790 19700 129800 19780
rect 141140 19700 141150 19780
rect 141290 19700 141300 19780
rect 141440 19700 141450 19780
rect 60610 19690 60690 19700
rect 60930 19690 61010 19700
rect 61350 19690 61430 19700
rect 61670 19690 61750 19700
rect 74110 19690 74190 19700
rect 74430 19690 74510 19700
rect 74850 19690 74930 19700
rect 75170 19690 75250 19700
rect 87610 19690 87690 19700
rect 87930 19690 88010 19700
rect 88350 19690 88430 19700
rect 88670 19690 88750 19700
rect 101110 19690 101190 19700
rect 101430 19690 101510 19700
rect 101850 19690 101930 19700
rect 102170 19690 102250 19700
rect 114610 19690 114690 19700
rect 114930 19690 115010 19700
rect 115350 19690 115430 19700
rect 115670 19690 115750 19700
rect 128110 19690 128190 19700
rect 128430 19690 128510 19700
rect 128850 19690 128930 19700
rect 129170 19690 129250 19700
rect 60690 19610 60700 19690
rect 61010 19610 61020 19690
rect 61430 19610 61440 19690
rect 61750 19610 61760 19690
rect 74190 19610 74200 19690
rect 74510 19610 74520 19690
rect 74930 19610 74940 19690
rect 75250 19610 75260 19690
rect 87690 19610 87700 19690
rect 88010 19610 88020 19690
rect 88430 19610 88440 19690
rect 88750 19610 88760 19690
rect 101190 19610 101200 19690
rect 101510 19610 101520 19690
rect 101930 19610 101940 19690
rect 102250 19610 102260 19690
rect 114690 19610 114700 19690
rect 115010 19610 115020 19690
rect 115430 19610 115440 19690
rect 115750 19610 115760 19690
rect 128190 19610 128200 19690
rect 128510 19610 128520 19690
rect 128930 19610 128940 19690
rect 129250 19610 129260 19690
rect 48500 19600 48640 19610
rect 48710 19600 48790 19610
rect 60060 19600 60140 19610
rect 60210 19600 60290 19610
rect 60360 19600 60440 19610
rect 62060 19600 62140 19610
rect 62210 19600 62290 19610
rect 73560 19600 73640 19610
rect 73710 19600 73790 19610
rect 73860 19600 73940 19610
rect 75560 19600 75640 19610
rect 75710 19600 75790 19610
rect 87060 19600 87140 19610
rect 87210 19600 87290 19610
rect 87360 19600 87440 19610
rect 89060 19600 89140 19610
rect 89210 19600 89290 19610
rect 100560 19600 100640 19610
rect 100710 19600 100790 19610
rect 100860 19600 100940 19610
rect 102560 19600 102640 19610
rect 102710 19600 102790 19610
rect 114060 19600 114140 19610
rect 114210 19600 114290 19610
rect 114360 19600 114440 19610
rect 116060 19600 116140 19610
rect 116210 19600 116290 19610
rect 127560 19600 127640 19610
rect 127710 19600 127790 19610
rect 127860 19600 127940 19610
rect 129560 19600 129640 19610
rect 129710 19600 129790 19610
rect 141060 19600 141140 19610
rect 141210 19600 141290 19610
rect 141360 19600 141440 19610
rect 43905 19530 43985 19540
rect 44225 19530 44305 19540
rect 44545 19530 44625 19540
rect 44865 19530 44945 19540
rect 45185 19530 45265 19540
rect 45505 19530 45585 19540
rect 45825 19530 45905 19540
rect 46145 19530 46225 19540
rect 46465 19530 46545 19540
rect 46785 19530 46865 19540
rect 47105 19530 47185 19540
rect 47425 19530 47505 19540
rect 47745 19530 47825 19540
rect 48065 19530 48145 19540
rect 43060 19460 43140 19470
rect 43380 19460 43460 19470
rect 43140 19380 43150 19460
rect 43460 19380 43470 19460
rect 43985 19450 43995 19530
rect 44305 19450 44315 19530
rect 44625 19450 44635 19530
rect 44945 19450 44955 19530
rect 45265 19450 45275 19530
rect 45585 19450 45595 19530
rect 45905 19450 45915 19530
rect 46225 19450 46235 19530
rect 46545 19450 46555 19530
rect 46865 19450 46875 19530
rect 47185 19450 47195 19530
rect 47505 19450 47515 19530
rect 47825 19450 47835 19530
rect 48145 19450 48155 19530
rect 48500 19430 48605 19600
rect 48640 19520 48650 19600
rect 48790 19520 48800 19600
rect 60140 19520 60150 19600
rect 60290 19520 60300 19600
rect 60440 19520 60450 19600
rect 60770 19530 60850 19540
rect 61090 19530 61170 19540
rect 61510 19530 61590 19540
rect 61830 19530 61910 19540
rect 60850 19450 60860 19530
rect 61170 19450 61180 19530
rect 61590 19450 61600 19530
rect 61910 19450 61920 19530
rect 62140 19520 62150 19600
rect 62290 19520 62300 19600
rect 73640 19520 73650 19600
rect 73790 19520 73800 19600
rect 73940 19520 73950 19600
rect 74270 19530 74350 19540
rect 74590 19530 74670 19540
rect 75010 19530 75090 19540
rect 75330 19530 75410 19540
rect 74350 19450 74360 19530
rect 74670 19450 74680 19530
rect 75090 19450 75100 19530
rect 75410 19450 75420 19530
rect 75640 19520 75650 19600
rect 75790 19520 75800 19600
rect 87140 19520 87150 19600
rect 87290 19520 87300 19600
rect 87440 19520 87450 19600
rect 87770 19530 87850 19540
rect 88090 19530 88170 19540
rect 88510 19530 88590 19540
rect 88830 19530 88910 19540
rect 87850 19450 87860 19530
rect 88170 19450 88180 19530
rect 88590 19450 88600 19530
rect 88910 19450 88920 19530
rect 89140 19520 89150 19600
rect 89290 19520 89300 19600
rect 100640 19520 100650 19600
rect 100790 19520 100800 19600
rect 100940 19520 100950 19600
rect 101270 19530 101350 19540
rect 101590 19530 101670 19540
rect 102010 19530 102090 19540
rect 102330 19530 102410 19540
rect 101350 19450 101360 19530
rect 101670 19450 101680 19530
rect 102090 19450 102100 19530
rect 102410 19450 102420 19530
rect 102640 19520 102650 19600
rect 102790 19520 102800 19600
rect 114140 19520 114150 19600
rect 114290 19520 114300 19600
rect 114440 19520 114450 19600
rect 114770 19530 114850 19540
rect 115090 19530 115170 19540
rect 115510 19530 115590 19540
rect 115830 19530 115910 19540
rect 114850 19450 114860 19530
rect 115170 19450 115180 19530
rect 115590 19450 115600 19530
rect 115910 19450 115920 19530
rect 116140 19520 116150 19600
rect 116290 19520 116300 19600
rect 127640 19520 127650 19600
rect 127790 19520 127800 19600
rect 127940 19520 127950 19600
rect 128270 19530 128350 19540
rect 128590 19530 128670 19540
rect 129010 19530 129090 19540
rect 129330 19530 129410 19540
rect 128350 19450 128360 19530
rect 128670 19450 128680 19530
rect 129090 19450 129100 19530
rect 129410 19450 129420 19530
rect 129640 19520 129650 19600
rect 129790 19520 129800 19600
rect 141140 19520 141150 19600
rect 141290 19520 141300 19600
rect 141440 19520 141450 19600
rect 48500 19420 48640 19430
rect 48710 19420 48790 19430
rect 60060 19420 60140 19430
rect 60210 19420 60290 19430
rect 60360 19420 60440 19430
rect 62060 19420 62140 19430
rect 62210 19420 62290 19430
rect 73560 19420 73640 19430
rect 73710 19420 73790 19430
rect 73860 19420 73940 19430
rect 75560 19420 75640 19430
rect 75710 19420 75790 19430
rect 87060 19420 87140 19430
rect 87210 19420 87290 19430
rect 87360 19420 87440 19430
rect 89060 19420 89140 19430
rect 89210 19420 89290 19430
rect 100560 19420 100640 19430
rect 100710 19420 100790 19430
rect 100860 19420 100940 19430
rect 102560 19420 102640 19430
rect 102710 19420 102790 19430
rect 114060 19420 114140 19430
rect 114210 19420 114290 19430
rect 114360 19420 114440 19430
rect 116060 19420 116140 19430
rect 116210 19420 116290 19430
rect 127560 19420 127640 19430
rect 127710 19420 127790 19430
rect 127860 19420 127940 19430
rect 129560 19420 129640 19430
rect 129710 19420 129790 19430
rect 141060 19420 141140 19430
rect 141210 19420 141290 19430
rect 141360 19420 141440 19430
rect 44065 19370 44145 19380
rect 44385 19370 44465 19380
rect 44705 19370 44785 19380
rect 45025 19370 45105 19380
rect 45345 19370 45425 19380
rect 45665 19370 45745 19380
rect 45985 19370 46065 19380
rect 46305 19370 46385 19380
rect 46625 19370 46705 19380
rect 46945 19370 47025 19380
rect 47265 19370 47345 19380
rect 47585 19370 47665 19380
rect 47905 19370 47985 19380
rect 48225 19370 48305 19380
rect 42950 19300 42980 19310
rect 43220 19300 43300 19310
rect 42980 19220 42990 19300
rect 43300 19220 43310 19300
rect 44145 19290 44155 19370
rect 44465 19290 44475 19370
rect 44785 19290 44795 19370
rect 45105 19290 45115 19370
rect 45425 19290 45435 19370
rect 45745 19290 45755 19370
rect 46065 19290 46075 19370
rect 46385 19290 46395 19370
rect 46705 19290 46715 19370
rect 47025 19290 47035 19370
rect 47345 19290 47355 19370
rect 47665 19290 47675 19370
rect 47985 19290 47995 19370
rect 48305 19290 48315 19370
rect 48500 19250 48605 19420
rect 48640 19340 48650 19420
rect 48790 19340 48800 19420
rect 60140 19340 60150 19420
rect 60290 19340 60300 19420
rect 60440 19340 60450 19420
rect 60610 19370 60690 19380
rect 60930 19370 61010 19380
rect 61350 19370 61430 19380
rect 61670 19370 61750 19380
rect 49180 19280 49210 19310
rect 49300 19280 49330 19310
rect 49420 19280 49450 19310
rect 49540 19280 49570 19310
rect 49660 19280 49690 19310
rect 49780 19280 49810 19310
rect 49900 19280 49930 19310
rect 50020 19280 50050 19310
rect 50140 19280 50170 19310
rect 50260 19280 50290 19310
rect 50380 19280 50410 19310
rect 50500 19280 50530 19310
rect 50620 19280 50650 19310
rect 50740 19280 50770 19310
rect 50860 19280 50890 19310
rect 50980 19280 51010 19310
rect 51100 19280 51130 19310
rect 51220 19280 51250 19310
rect 51340 19280 51370 19310
rect 51460 19280 51490 19310
rect 51580 19280 51610 19310
rect 51700 19280 51730 19310
rect 51820 19280 51850 19310
rect 51940 19280 51970 19310
rect 52060 19280 52090 19310
rect 52180 19280 52210 19310
rect 52300 19280 52330 19310
rect 52420 19280 52450 19310
rect 52540 19280 52570 19310
rect 52660 19280 52690 19310
rect 52780 19280 52810 19310
rect 52900 19280 52930 19310
rect 53020 19280 53050 19310
rect 53140 19280 53170 19310
rect 53260 19280 53290 19310
rect 53380 19280 53410 19310
rect 53500 19280 53530 19310
rect 53620 19280 53650 19310
rect 53740 19280 53770 19310
rect 53860 19280 53890 19310
rect 53980 19280 54010 19310
rect 54100 19280 54130 19310
rect 54220 19280 54250 19310
rect 54340 19280 54370 19310
rect 54460 19280 54490 19310
rect 54580 19280 54610 19310
rect 54700 19280 54730 19310
rect 54820 19280 54850 19310
rect 54940 19280 54970 19310
rect 55060 19280 55090 19310
rect 55180 19280 55210 19310
rect 55300 19280 55330 19310
rect 55420 19280 55450 19310
rect 55540 19280 55570 19310
rect 55660 19280 55690 19310
rect 55780 19280 55810 19310
rect 55900 19280 55930 19310
rect 56020 19280 56050 19310
rect 56140 19280 56170 19310
rect 56260 19280 56290 19310
rect 56380 19280 56410 19310
rect 56500 19280 56530 19310
rect 56620 19280 56650 19310
rect 56740 19280 56770 19310
rect 56860 19280 56890 19310
rect 56980 19280 57010 19310
rect 57100 19280 57130 19310
rect 57220 19280 57250 19310
rect 57340 19280 57370 19310
rect 57460 19280 57490 19310
rect 57580 19280 57610 19310
rect 57700 19280 57730 19310
rect 57820 19280 57850 19310
rect 57940 19280 57970 19310
rect 58060 19280 58090 19310
rect 58180 19280 58210 19310
rect 58300 19280 58330 19310
rect 58420 19280 58450 19310
rect 58540 19280 58570 19310
rect 58660 19280 58690 19310
rect 58780 19280 58810 19310
rect 58900 19280 58930 19310
rect 59020 19280 59050 19310
rect 59140 19280 59170 19310
rect 59260 19280 59290 19310
rect 59380 19280 59410 19310
rect 59500 19280 59530 19310
rect 59620 19280 59650 19310
rect 59740 19280 59770 19310
rect 60690 19290 60700 19370
rect 61010 19290 61020 19370
rect 61430 19290 61440 19370
rect 61750 19290 61760 19370
rect 62140 19340 62150 19420
rect 62290 19340 62300 19420
rect 73640 19340 73650 19420
rect 73790 19340 73800 19420
rect 73940 19340 73950 19420
rect 74110 19370 74190 19380
rect 74430 19370 74510 19380
rect 74850 19370 74930 19380
rect 75170 19370 75250 19380
rect 62680 19280 62710 19310
rect 73245 19280 73270 19310
rect 74190 19290 74200 19370
rect 74510 19290 74520 19370
rect 74930 19290 74940 19370
rect 75250 19290 75260 19370
rect 75640 19340 75650 19420
rect 75790 19340 75800 19420
rect 87140 19340 87150 19420
rect 87290 19340 87300 19420
rect 87440 19340 87450 19420
rect 87610 19370 87690 19380
rect 87930 19370 88010 19380
rect 88350 19370 88430 19380
rect 88670 19370 88750 19380
rect 76180 19280 76210 19310
rect 86745 19280 86770 19310
rect 87690 19290 87700 19370
rect 88010 19290 88020 19370
rect 88430 19290 88440 19370
rect 88750 19290 88760 19370
rect 89140 19340 89150 19420
rect 89290 19340 89300 19420
rect 100640 19340 100650 19420
rect 100790 19340 100800 19420
rect 100940 19340 100950 19420
rect 101110 19370 101190 19380
rect 101430 19370 101510 19380
rect 101850 19370 101930 19380
rect 102170 19370 102250 19380
rect 89680 19280 89710 19310
rect 100245 19280 100270 19310
rect 101190 19290 101200 19370
rect 101510 19290 101520 19370
rect 101930 19290 101940 19370
rect 102250 19290 102260 19370
rect 102640 19340 102650 19420
rect 102790 19340 102800 19420
rect 114140 19340 114150 19420
rect 114290 19340 114300 19420
rect 114440 19340 114450 19420
rect 114610 19370 114690 19380
rect 114930 19370 115010 19380
rect 115350 19370 115430 19380
rect 115670 19370 115750 19380
rect 103180 19280 103210 19310
rect 113745 19280 113770 19310
rect 114690 19290 114700 19370
rect 115010 19290 115020 19370
rect 115430 19290 115440 19370
rect 115750 19290 115760 19370
rect 116140 19340 116150 19420
rect 116290 19340 116300 19420
rect 127640 19340 127650 19420
rect 127790 19340 127800 19420
rect 127940 19340 127950 19420
rect 128110 19370 128190 19380
rect 128430 19370 128510 19380
rect 128850 19370 128930 19380
rect 129170 19370 129250 19380
rect 116680 19280 116710 19310
rect 127245 19280 127270 19310
rect 128190 19290 128200 19370
rect 128510 19290 128520 19370
rect 128930 19290 128940 19370
rect 129250 19290 129260 19370
rect 129640 19340 129650 19420
rect 129790 19340 129800 19420
rect 141140 19340 141150 19420
rect 141290 19340 141300 19420
rect 141440 19340 141450 19420
rect 130180 19280 130210 19310
rect 49060 19250 49120 19280
rect 49180 19250 49240 19280
rect 49300 19250 49360 19280
rect 49420 19250 49480 19280
rect 49540 19250 49600 19280
rect 49660 19250 49720 19280
rect 49780 19250 49840 19280
rect 49900 19250 49960 19280
rect 50020 19250 50080 19280
rect 50140 19250 50200 19280
rect 50260 19250 50320 19280
rect 50380 19250 50440 19280
rect 50500 19250 50560 19280
rect 50620 19250 50680 19280
rect 50740 19250 50800 19280
rect 50860 19250 50920 19280
rect 50980 19250 51040 19280
rect 51100 19250 51160 19280
rect 51220 19250 51280 19280
rect 51340 19250 51400 19280
rect 51460 19250 51520 19280
rect 51580 19250 51640 19280
rect 51700 19250 51760 19280
rect 51820 19250 51880 19280
rect 51940 19250 52000 19280
rect 52060 19250 52120 19280
rect 52180 19250 52240 19280
rect 52300 19250 52360 19280
rect 52420 19250 52480 19280
rect 52540 19250 52600 19280
rect 52660 19250 52720 19280
rect 52780 19250 52840 19280
rect 52900 19250 52960 19280
rect 53020 19250 53080 19280
rect 53140 19250 53200 19280
rect 53260 19250 53320 19280
rect 53380 19250 53440 19280
rect 53500 19250 53560 19280
rect 53620 19250 53680 19280
rect 53740 19250 53800 19280
rect 53860 19250 53920 19280
rect 53980 19250 54040 19280
rect 54100 19250 54160 19280
rect 54220 19250 54280 19280
rect 54340 19250 54400 19280
rect 54460 19250 54520 19280
rect 54580 19250 54640 19280
rect 54700 19250 54760 19280
rect 54820 19250 54880 19280
rect 54940 19250 55000 19280
rect 55060 19250 55120 19280
rect 55180 19250 55240 19280
rect 55300 19250 55360 19280
rect 55420 19250 55480 19280
rect 55540 19250 55600 19280
rect 55660 19250 55720 19280
rect 55780 19250 55840 19280
rect 55900 19250 55960 19280
rect 56020 19250 56080 19280
rect 56140 19250 56200 19280
rect 56260 19250 56320 19280
rect 56380 19250 56440 19280
rect 56500 19250 56560 19280
rect 56620 19250 56680 19280
rect 56740 19250 56800 19280
rect 56860 19250 56920 19280
rect 56980 19250 57040 19280
rect 57100 19250 57160 19280
rect 57220 19250 57280 19280
rect 57340 19250 57400 19280
rect 57460 19250 57520 19280
rect 57580 19250 57640 19280
rect 57700 19250 57760 19280
rect 57820 19250 57880 19280
rect 57940 19250 58000 19280
rect 58060 19250 58120 19280
rect 58180 19250 58240 19280
rect 58300 19250 58360 19280
rect 58420 19250 58480 19280
rect 58540 19250 58600 19280
rect 58660 19250 58720 19280
rect 58780 19250 58840 19280
rect 58900 19250 58960 19280
rect 59020 19250 59080 19280
rect 59140 19250 59200 19280
rect 59260 19250 59320 19280
rect 59380 19250 59440 19280
rect 59500 19250 59560 19280
rect 59620 19250 59680 19280
rect 59740 19250 59800 19280
rect 62560 19250 62620 19280
rect 62680 19250 62740 19280
rect 73245 19250 73300 19280
rect 76060 19250 76120 19280
rect 76180 19250 76240 19280
rect 86745 19250 86800 19280
rect 89560 19250 89620 19280
rect 89680 19250 89740 19280
rect 100245 19250 100300 19280
rect 103060 19250 103120 19280
rect 103180 19250 103240 19280
rect 113745 19250 113800 19280
rect 116560 19250 116620 19280
rect 116680 19250 116740 19280
rect 127245 19250 127300 19280
rect 130060 19250 130120 19280
rect 130180 19250 130240 19280
rect 48500 19240 48640 19250
rect 48710 19240 48790 19250
rect 60060 19240 60140 19250
rect 60210 19240 60290 19250
rect 60360 19240 60440 19250
rect 62060 19240 62140 19250
rect 62210 19240 62290 19250
rect 73560 19240 73640 19250
rect 73710 19240 73790 19250
rect 73860 19240 73940 19250
rect 75560 19240 75640 19250
rect 75710 19240 75790 19250
rect 87060 19240 87140 19250
rect 87210 19240 87290 19250
rect 87360 19240 87440 19250
rect 89060 19240 89140 19250
rect 89210 19240 89290 19250
rect 100560 19240 100640 19250
rect 100710 19240 100790 19250
rect 100860 19240 100940 19250
rect 102560 19240 102640 19250
rect 102710 19240 102790 19250
rect 114060 19240 114140 19250
rect 114210 19240 114290 19250
rect 114360 19240 114440 19250
rect 116060 19240 116140 19250
rect 116210 19240 116290 19250
rect 127560 19240 127640 19250
rect 127710 19240 127790 19250
rect 127860 19240 127940 19250
rect 129560 19240 129640 19250
rect 129710 19240 129790 19250
rect 141060 19240 141140 19250
rect 141210 19240 141290 19250
rect 141360 19240 141440 19250
rect 43905 19210 43985 19220
rect 44225 19210 44305 19220
rect 44545 19210 44625 19220
rect 44865 19210 44945 19220
rect 45185 19210 45265 19220
rect 45505 19210 45585 19220
rect 45825 19210 45905 19220
rect 46145 19210 46225 19220
rect 46465 19210 46545 19220
rect 46785 19210 46865 19220
rect 47105 19210 47185 19220
rect 47425 19210 47505 19220
rect 47745 19210 47825 19220
rect 48065 19210 48145 19220
rect 43060 19140 43140 19150
rect 43380 19140 43460 19150
rect 43140 19060 43150 19140
rect 43460 19060 43470 19140
rect 43985 19130 43995 19210
rect 44305 19130 44315 19210
rect 44625 19130 44635 19210
rect 44945 19130 44955 19210
rect 45265 19130 45275 19210
rect 45585 19130 45595 19210
rect 45905 19130 45915 19210
rect 46225 19130 46235 19210
rect 46545 19130 46555 19210
rect 46865 19130 46875 19210
rect 47185 19130 47195 19210
rect 47505 19130 47515 19210
rect 47825 19130 47835 19210
rect 48145 19130 48155 19210
rect 48500 19070 48605 19240
rect 48640 19160 48650 19240
rect 48790 19160 48800 19240
rect 49180 19160 49210 19190
rect 49300 19160 49330 19190
rect 49420 19160 49450 19190
rect 49540 19160 49570 19190
rect 49660 19160 49690 19190
rect 49780 19160 49810 19190
rect 49900 19160 49930 19190
rect 50020 19160 50050 19190
rect 50140 19160 50170 19190
rect 50260 19160 50290 19190
rect 50380 19160 50410 19190
rect 50500 19160 50530 19190
rect 50620 19160 50650 19190
rect 50740 19160 50770 19190
rect 50860 19160 50890 19190
rect 50980 19160 51010 19190
rect 51100 19160 51130 19190
rect 51220 19160 51250 19190
rect 51340 19160 51370 19190
rect 51460 19160 51490 19190
rect 51580 19160 51610 19190
rect 51700 19160 51730 19190
rect 51820 19160 51850 19190
rect 51940 19160 51970 19190
rect 52060 19160 52090 19190
rect 52180 19160 52210 19190
rect 52300 19160 52330 19190
rect 52420 19160 52450 19190
rect 52540 19160 52570 19190
rect 52660 19160 52690 19190
rect 52780 19160 52810 19190
rect 52900 19160 52930 19190
rect 53020 19160 53050 19190
rect 53140 19160 53170 19190
rect 53260 19160 53290 19190
rect 53380 19160 53410 19190
rect 53500 19160 53530 19190
rect 53620 19160 53650 19190
rect 53740 19160 53770 19190
rect 53860 19160 53890 19190
rect 53980 19160 54010 19190
rect 54100 19160 54130 19190
rect 54220 19160 54250 19190
rect 54340 19160 54370 19190
rect 54460 19160 54490 19190
rect 54580 19160 54610 19190
rect 54700 19160 54730 19190
rect 54820 19160 54850 19190
rect 54940 19160 54970 19190
rect 55060 19160 55090 19190
rect 55180 19160 55210 19190
rect 55300 19160 55330 19190
rect 55420 19160 55450 19190
rect 55540 19160 55570 19190
rect 55660 19160 55690 19190
rect 55780 19160 55810 19190
rect 55900 19160 55930 19190
rect 56020 19160 56050 19190
rect 56140 19160 56170 19190
rect 56260 19160 56290 19190
rect 56380 19160 56410 19190
rect 56500 19160 56530 19190
rect 56620 19160 56650 19190
rect 56740 19160 56770 19190
rect 56860 19160 56890 19190
rect 56980 19160 57010 19190
rect 57100 19160 57130 19190
rect 57220 19160 57250 19190
rect 57340 19160 57370 19190
rect 57460 19160 57490 19190
rect 57580 19160 57610 19190
rect 57700 19160 57730 19190
rect 57820 19160 57850 19190
rect 57940 19160 57970 19190
rect 58060 19160 58090 19190
rect 58180 19160 58210 19190
rect 58300 19160 58330 19190
rect 58420 19160 58450 19190
rect 58540 19160 58570 19190
rect 58660 19160 58690 19190
rect 58780 19160 58810 19190
rect 58900 19160 58930 19190
rect 59020 19160 59050 19190
rect 59140 19160 59170 19190
rect 59260 19160 59290 19190
rect 59380 19160 59410 19190
rect 59500 19160 59530 19190
rect 59620 19160 59650 19190
rect 59740 19160 59770 19190
rect 60140 19160 60150 19240
rect 60290 19160 60300 19240
rect 60440 19160 60450 19240
rect 60770 19210 60850 19220
rect 61090 19210 61170 19220
rect 61510 19210 61590 19220
rect 61830 19210 61910 19220
rect 49060 19130 49120 19160
rect 49180 19130 49240 19160
rect 49300 19130 49360 19160
rect 49420 19130 49480 19160
rect 49540 19130 49600 19160
rect 49660 19130 49720 19160
rect 49780 19130 49840 19160
rect 49900 19130 49960 19160
rect 50020 19130 50080 19160
rect 50140 19130 50200 19160
rect 50260 19130 50320 19160
rect 50380 19130 50440 19160
rect 50500 19130 50560 19160
rect 50620 19130 50680 19160
rect 50740 19130 50800 19160
rect 50860 19130 50920 19160
rect 50980 19130 51040 19160
rect 51100 19130 51160 19160
rect 51220 19130 51280 19160
rect 51340 19130 51400 19160
rect 51460 19130 51520 19160
rect 51580 19130 51640 19160
rect 51700 19130 51760 19160
rect 51820 19130 51880 19160
rect 51940 19130 52000 19160
rect 52060 19130 52120 19160
rect 52180 19130 52240 19160
rect 52300 19130 52360 19160
rect 52420 19130 52480 19160
rect 52540 19130 52600 19160
rect 52660 19130 52720 19160
rect 52780 19130 52840 19160
rect 52900 19130 52960 19160
rect 53020 19130 53080 19160
rect 53140 19130 53200 19160
rect 53260 19130 53320 19160
rect 53380 19130 53440 19160
rect 53500 19130 53560 19160
rect 53620 19130 53680 19160
rect 53740 19130 53800 19160
rect 53860 19130 53920 19160
rect 53980 19130 54040 19160
rect 54100 19130 54160 19160
rect 54220 19130 54280 19160
rect 54340 19130 54400 19160
rect 54460 19130 54520 19160
rect 54580 19130 54640 19160
rect 54700 19130 54760 19160
rect 54820 19130 54880 19160
rect 54940 19130 55000 19160
rect 55060 19130 55120 19160
rect 55180 19130 55240 19160
rect 55300 19130 55360 19160
rect 55420 19130 55480 19160
rect 55540 19130 55600 19160
rect 55660 19130 55720 19160
rect 55780 19130 55840 19160
rect 55900 19130 55960 19160
rect 56020 19130 56080 19160
rect 56140 19130 56200 19160
rect 56260 19130 56320 19160
rect 56380 19130 56440 19160
rect 56500 19130 56560 19160
rect 56620 19130 56680 19160
rect 56740 19130 56800 19160
rect 56860 19130 56920 19160
rect 56980 19130 57040 19160
rect 57100 19130 57160 19160
rect 57220 19130 57280 19160
rect 57340 19130 57400 19160
rect 57460 19130 57520 19160
rect 57580 19130 57640 19160
rect 57700 19130 57760 19160
rect 57820 19130 57880 19160
rect 57940 19130 58000 19160
rect 58060 19130 58120 19160
rect 58180 19130 58240 19160
rect 58300 19130 58360 19160
rect 58420 19130 58480 19160
rect 58540 19130 58600 19160
rect 58660 19130 58720 19160
rect 58780 19130 58840 19160
rect 58900 19130 58960 19160
rect 59020 19130 59080 19160
rect 59140 19130 59200 19160
rect 59260 19130 59320 19160
rect 59380 19130 59440 19160
rect 59500 19130 59560 19160
rect 59620 19130 59680 19160
rect 59740 19130 59800 19160
rect 60850 19130 60860 19210
rect 61170 19130 61180 19210
rect 61590 19130 61600 19210
rect 61910 19130 61920 19210
rect 62140 19160 62150 19240
rect 62290 19160 62300 19240
rect 62680 19160 62710 19190
rect 73245 19160 73270 19190
rect 73640 19160 73650 19240
rect 73790 19160 73800 19240
rect 73940 19160 73950 19240
rect 74270 19210 74350 19220
rect 74590 19210 74670 19220
rect 75010 19210 75090 19220
rect 75330 19210 75410 19220
rect 62560 19130 62620 19160
rect 62680 19130 62740 19160
rect 73245 19130 73300 19160
rect 74350 19130 74360 19210
rect 74670 19130 74680 19210
rect 75090 19130 75100 19210
rect 75410 19130 75420 19210
rect 75640 19160 75650 19240
rect 75790 19160 75800 19240
rect 76180 19160 76210 19190
rect 86745 19160 86770 19190
rect 87140 19160 87150 19240
rect 87290 19160 87300 19240
rect 87440 19160 87450 19240
rect 87770 19210 87850 19220
rect 88090 19210 88170 19220
rect 88510 19210 88590 19220
rect 88830 19210 88910 19220
rect 76060 19130 76120 19160
rect 76180 19130 76240 19160
rect 86745 19130 86800 19160
rect 87850 19130 87860 19210
rect 88170 19130 88180 19210
rect 88590 19130 88600 19210
rect 88910 19130 88920 19210
rect 89140 19160 89150 19240
rect 89290 19160 89300 19240
rect 89680 19160 89710 19190
rect 100245 19160 100270 19190
rect 100640 19160 100650 19240
rect 100790 19160 100800 19240
rect 100940 19160 100950 19240
rect 101270 19210 101350 19220
rect 101590 19210 101670 19220
rect 102010 19210 102090 19220
rect 102330 19210 102410 19220
rect 89560 19130 89620 19160
rect 89680 19130 89740 19160
rect 100245 19130 100300 19160
rect 101350 19130 101360 19210
rect 101670 19130 101680 19210
rect 102090 19130 102100 19210
rect 102410 19130 102420 19210
rect 102640 19160 102650 19240
rect 102790 19160 102800 19240
rect 103180 19160 103210 19190
rect 113745 19160 113770 19190
rect 114140 19160 114150 19240
rect 114290 19160 114300 19240
rect 114440 19160 114450 19240
rect 114770 19210 114850 19220
rect 115090 19210 115170 19220
rect 115510 19210 115590 19220
rect 115830 19210 115910 19220
rect 103060 19130 103120 19160
rect 103180 19130 103240 19160
rect 113745 19130 113800 19160
rect 114850 19130 114860 19210
rect 115170 19130 115180 19210
rect 115590 19130 115600 19210
rect 115910 19130 115920 19210
rect 116140 19160 116150 19240
rect 116290 19160 116300 19240
rect 116680 19160 116710 19190
rect 127245 19160 127270 19190
rect 127640 19160 127650 19240
rect 127790 19160 127800 19240
rect 127940 19160 127950 19240
rect 128270 19210 128350 19220
rect 128590 19210 128670 19220
rect 129010 19210 129090 19220
rect 129330 19210 129410 19220
rect 116560 19130 116620 19160
rect 116680 19130 116740 19160
rect 127245 19130 127300 19160
rect 128350 19130 128360 19210
rect 128670 19130 128680 19210
rect 129090 19130 129100 19210
rect 129410 19130 129420 19210
rect 129640 19160 129650 19240
rect 129790 19160 129800 19240
rect 130180 19160 130210 19190
rect 141140 19160 141150 19240
rect 141290 19160 141300 19240
rect 141440 19160 141450 19240
rect 130060 19130 130120 19160
rect 130180 19130 130240 19160
rect 48500 19060 48640 19070
rect 48710 19060 48790 19070
rect 44065 19050 44145 19060
rect 44385 19050 44465 19060
rect 44705 19050 44785 19060
rect 45025 19050 45105 19060
rect 45345 19050 45425 19060
rect 45665 19050 45745 19060
rect 45985 19050 46065 19060
rect 46305 19050 46385 19060
rect 46625 19050 46705 19060
rect 46945 19050 47025 19060
rect 47265 19050 47345 19060
rect 47585 19050 47665 19060
rect 47905 19050 47985 19060
rect 48225 19050 48305 19060
rect 44145 18970 44155 19050
rect 44465 18970 44475 19050
rect 44785 18970 44795 19050
rect 45105 18970 45115 19050
rect 45425 18970 45435 19050
rect 45745 18970 45755 19050
rect 46065 18970 46075 19050
rect 46385 18970 46395 19050
rect 46705 18970 46715 19050
rect 47025 18970 47035 19050
rect 47345 18970 47355 19050
rect 47665 18970 47675 19050
rect 47985 18970 47995 19050
rect 48305 18970 48315 19050
rect 48500 18900 48605 19060
rect 48640 18980 48650 19060
rect 48790 18980 48800 19060
rect 49180 19010 49210 19070
rect 49300 19010 49330 19070
rect 49420 19010 49450 19070
rect 49540 19010 49570 19070
rect 49660 19010 49690 19070
rect 49780 19010 49810 19070
rect 49900 19010 49930 19070
rect 50020 19010 50050 19070
rect 50140 19010 50170 19070
rect 50260 19010 50290 19070
rect 50380 19010 50410 19070
rect 50500 19010 50530 19070
rect 50620 19010 50650 19070
rect 50740 19010 50770 19070
rect 50860 19010 50890 19070
rect 50980 19010 51010 19070
rect 51100 19010 51130 19070
rect 51220 19010 51250 19070
rect 51340 19010 51370 19070
rect 51460 19010 51490 19070
rect 51580 19010 51610 19070
rect 51700 19010 51730 19070
rect 51820 19010 51850 19070
rect 51940 19010 51970 19070
rect 52060 19010 52090 19070
rect 52180 19010 52210 19070
rect 52300 19010 52330 19070
rect 52420 19010 52450 19070
rect 52540 19010 52570 19070
rect 52660 19010 52690 19070
rect 52780 19010 52810 19070
rect 52900 19010 52930 19070
rect 53020 19010 53050 19070
rect 53140 19010 53170 19070
rect 53260 19010 53290 19070
rect 53380 19010 53410 19070
rect 53500 19010 53530 19070
rect 53620 19010 53650 19070
rect 53740 19010 53770 19070
rect 53860 19010 53890 19070
rect 53980 19010 54010 19070
rect 54100 19010 54130 19070
rect 54220 19010 54250 19070
rect 54340 19010 54370 19070
rect 54460 19010 54490 19070
rect 54580 19010 54610 19070
rect 54700 19010 54730 19070
rect 54820 19010 54850 19070
rect 54940 19010 54970 19070
rect 55060 19010 55090 19070
rect 55180 19010 55210 19070
rect 55300 19010 55330 19070
rect 55420 19010 55450 19070
rect 55540 19010 55570 19070
rect 55660 19010 55690 19070
rect 55780 19010 55810 19070
rect 55900 19010 55930 19070
rect 56020 19010 56050 19070
rect 56140 19010 56170 19070
rect 56260 19010 56290 19070
rect 56380 19010 56410 19070
rect 56500 19010 56530 19070
rect 56620 19010 56650 19070
rect 56740 19010 56770 19070
rect 56860 19010 56890 19070
rect 56980 19010 57010 19070
rect 57100 19010 57130 19070
rect 57220 19010 57250 19070
rect 57340 19010 57370 19070
rect 57460 19010 57490 19070
rect 57580 19010 57610 19070
rect 57700 19010 57730 19070
rect 57820 19010 57850 19070
rect 57940 19010 57970 19070
rect 58060 19010 58090 19070
rect 58180 19010 58210 19070
rect 58300 19010 58330 19070
rect 58420 19010 58450 19070
rect 58540 19010 58570 19070
rect 58660 19010 58690 19070
rect 58780 19010 58810 19070
rect 58900 19010 58930 19070
rect 59020 19010 59050 19070
rect 59140 19010 59170 19070
rect 59260 19010 59290 19070
rect 59380 19010 59410 19070
rect 59500 19010 59530 19070
rect 59620 19010 59650 19070
rect 59740 19010 59770 19070
rect 60060 19060 60140 19070
rect 60210 19060 60290 19070
rect 60360 19060 60440 19070
rect 62060 19060 62140 19070
rect 62210 19060 62290 19070
rect 60140 18980 60150 19060
rect 60290 18980 60300 19060
rect 60440 18980 60450 19060
rect 60610 19050 60690 19060
rect 60930 19050 61010 19060
rect 61350 19050 61430 19060
rect 61670 19050 61750 19060
rect 60690 18970 60700 19050
rect 61010 18970 61020 19050
rect 61430 18970 61440 19050
rect 61750 18970 61760 19050
rect 62140 18980 62150 19060
rect 62290 18980 62300 19060
rect 62680 19010 62710 19070
rect 73245 19010 73270 19070
rect 73560 19060 73640 19070
rect 73710 19060 73790 19070
rect 73860 19060 73940 19070
rect 75560 19060 75640 19070
rect 75710 19060 75790 19070
rect 73640 18980 73650 19060
rect 73790 18980 73800 19060
rect 73940 18980 73950 19060
rect 74110 19050 74190 19060
rect 74430 19050 74510 19060
rect 74850 19050 74930 19060
rect 75170 19050 75250 19060
rect 74190 18970 74200 19050
rect 74510 18970 74520 19050
rect 74930 18970 74940 19050
rect 75250 18970 75260 19050
rect 75640 18980 75650 19060
rect 75790 18980 75800 19060
rect 76180 19010 76210 19070
rect 86745 19010 86770 19070
rect 87060 19060 87140 19070
rect 87210 19060 87290 19070
rect 87360 19060 87440 19070
rect 89060 19060 89140 19070
rect 89210 19060 89290 19070
rect 87140 18980 87150 19060
rect 87290 18980 87300 19060
rect 87440 18980 87450 19060
rect 87610 19050 87690 19060
rect 87930 19050 88010 19060
rect 88350 19050 88430 19060
rect 88670 19050 88750 19060
rect 87690 18970 87700 19050
rect 88010 18970 88020 19050
rect 88430 18970 88440 19050
rect 88750 18970 88760 19050
rect 89140 18980 89150 19060
rect 89290 18980 89300 19060
rect 89680 19010 89710 19070
rect 100245 19010 100270 19070
rect 100560 19060 100640 19070
rect 100710 19060 100790 19070
rect 100860 19060 100940 19070
rect 102560 19060 102640 19070
rect 102710 19060 102790 19070
rect 100640 18980 100650 19060
rect 100790 18980 100800 19060
rect 100940 18980 100950 19060
rect 101110 19050 101190 19060
rect 101430 19050 101510 19060
rect 101850 19050 101930 19060
rect 102170 19050 102250 19060
rect 101190 18970 101200 19050
rect 101510 18970 101520 19050
rect 101930 18970 101940 19050
rect 102250 18970 102260 19050
rect 102640 18980 102650 19060
rect 102790 18980 102800 19060
rect 103180 19010 103210 19070
rect 113745 19010 113770 19070
rect 114060 19060 114140 19070
rect 114210 19060 114290 19070
rect 114360 19060 114440 19070
rect 116060 19060 116140 19070
rect 116210 19060 116290 19070
rect 114140 18980 114150 19060
rect 114290 18980 114300 19060
rect 114440 18980 114450 19060
rect 114610 19050 114690 19060
rect 114930 19050 115010 19060
rect 115350 19050 115430 19060
rect 115670 19050 115750 19060
rect 114690 18970 114700 19050
rect 115010 18970 115020 19050
rect 115430 18970 115440 19050
rect 115750 18970 115760 19050
rect 116140 18980 116150 19060
rect 116290 18980 116300 19060
rect 116680 19010 116710 19070
rect 127245 19010 127270 19070
rect 127560 19060 127640 19070
rect 127710 19060 127790 19070
rect 127860 19060 127940 19070
rect 129560 19060 129640 19070
rect 129710 19060 129790 19070
rect 127640 18980 127650 19060
rect 127790 18980 127800 19060
rect 127940 18980 127950 19060
rect 128110 19050 128190 19060
rect 128430 19050 128510 19060
rect 128850 19050 128930 19060
rect 129170 19050 129250 19060
rect 128190 18970 128200 19050
rect 128510 18970 128520 19050
rect 128930 18970 128940 19050
rect 129250 18970 129260 19050
rect 129640 18980 129650 19060
rect 129790 18980 129800 19060
rect 130180 19010 130210 19070
rect 141060 19060 141140 19070
rect 141210 19060 141290 19070
rect 141360 19060 141440 19070
rect 141140 18980 141150 19060
rect 141290 18980 141300 19060
rect 141440 18980 141450 19060
rect 141565 18900 141620 26700
rect 146540 26500 146620 26510
rect 146860 26500 146940 26510
rect 146620 26420 146630 26500
rect 146940 26420 146950 26500
rect 141945 26410 142025 26420
rect 145200 26410 145225 26420
rect 145465 26410 145545 26420
rect 145785 26410 145865 26420
rect 146105 26410 146185 26420
rect 142025 26330 142035 26410
rect 145225 26330 145235 26410
rect 145545 26330 145555 26410
rect 145865 26330 145875 26410
rect 146185 26330 146195 26410
rect 146700 26340 146780 26350
rect 147020 26340 147100 26350
rect 146780 26260 146790 26340
rect 141785 26250 141865 26260
rect 142105 26250 142185 26260
rect 145305 26250 145385 26260
rect 145625 26250 145705 26260
rect 145945 26250 146025 26260
rect 141865 26170 141875 26250
rect 142185 26170 142195 26250
rect 145385 26170 145395 26250
rect 145705 26170 145715 26250
rect 146025 26170 146035 26250
rect 146540 26180 146620 26190
rect 146860 26180 146940 26190
rect 146620 26100 146630 26180
rect 146940 26100 146950 26180
rect 141945 26090 142025 26100
rect 145200 26090 145225 26100
rect 145465 26090 145545 26100
rect 145785 26090 145865 26100
rect 146105 26090 146185 26100
rect 142025 26010 142035 26090
rect 145225 26010 145235 26090
rect 145545 26010 145555 26090
rect 145865 26010 145875 26090
rect 146185 26010 146195 26090
rect 146700 26020 146780 26030
rect 147020 26020 147100 26030
rect 146780 25940 146790 26020
rect 141785 25930 141865 25940
rect 142105 25930 142185 25940
rect 145305 25930 145385 25940
rect 145625 25930 145705 25940
rect 145945 25930 146025 25940
rect 141865 25850 141875 25930
rect 142185 25850 142195 25930
rect 145385 25850 145395 25930
rect 145705 25850 145715 25930
rect 146025 25850 146035 25930
rect 146540 25860 146620 25870
rect 146860 25860 146940 25870
rect 146620 25780 146630 25860
rect 146940 25780 146950 25860
rect 141945 25770 142025 25780
rect 145200 25770 145225 25780
rect 145465 25770 145545 25780
rect 145785 25770 145865 25780
rect 146105 25770 146185 25780
rect 142025 25690 142035 25770
rect 145225 25690 145235 25770
rect 145545 25690 145555 25770
rect 145865 25690 145875 25770
rect 146185 25690 146195 25770
rect 146700 25700 146780 25710
rect 147020 25700 147100 25710
rect 146780 25620 146790 25700
rect 141785 25610 141865 25620
rect 142105 25610 142185 25620
rect 145305 25610 145385 25620
rect 145625 25610 145705 25620
rect 145945 25610 146025 25620
rect 141865 25530 141875 25610
rect 142185 25530 142195 25610
rect 145385 25530 145395 25610
rect 145705 25530 145715 25610
rect 146025 25530 146035 25610
rect 146540 25540 146620 25550
rect 146860 25540 146940 25550
rect 146620 25460 146630 25540
rect 146940 25460 146950 25540
rect 141945 25450 142025 25460
rect 145200 25450 145225 25460
rect 145465 25450 145545 25460
rect 145785 25450 145865 25460
rect 146105 25450 146185 25460
rect 142025 25370 142035 25450
rect 145225 25370 145235 25450
rect 145545 25370 145555 25450
rect 145865 25370 145875 25450
rect 146185 25370 146195 25450
rect 146700 25380 146780 25390
rect 147020 25380 147100 25390
rect 146780 25300 146790 25380
rect 141785 25290 141865 25300
rect 142105 25290 142185 25300
rect 145305 25290 145385 25300
rect 145625 25290 145705 25300
rect 145945 25290 146025 25300
rect 141865 25210 141875 25290
rect 142185 25210 142195 25290
rect 145385 25210 145395 25290
rect 145705 25210 145715 25290
rect 146025 25210 146035 25290
rect 146540 25220 146620 25230
rect 146860 25220 146940 25230
rect 146620 25140 146630 25220
rect 146940 25140 146950 25220
rect 141945 25130 142025 25140
rect 145200 25130 145225 25140
rect 145465 25130 145545 25140
rect 145785 25130 145865 25140
rect 146105 25130 146185 25140
rect 142025 25050 142035 25130
rect 145225 25050 145235 25130
rect 145545 25050 145555 25130
rect 145865 25050 145875 25130
rect 146185 25050 146195 25130
rect 146700 25060 146780 25070
rect 147020 25060 147100 25070
rect 146780 24980 146790 25060
rect 141785 24970 141865 24980
rect 142105 24970 142185 24980
rect 145305 24970 145385 24980
rect 145625 24970 145705 24980
rect 145945 24970 146025 24980
rect 141865 24890 141875 24970
rect 142185 24890 142195 24970
rect 145385 24890 145395 24970
rect 145705 24890 145715 24970
rect 146025 24890 146035 24970
rect 146540 24900 146620 24910
rect 146860 24900 146940 24910
rect 146620 24820 146630 24900
rect 146940 24820 146950 24900
rect 141945 24810 142025 24820
rect 145200 24810 145225 24820
rect 145465 24810 145545 24820
rect 145785 24810 145865 24820
rect 146105 24810 146185 24820
rect 142025 24730 142035 24810
rect 145225 24730 145235 24810
rect 145545 24730 145555 24810
rect 145865 24730 145875 24810
rect 146185 24730 146195 24810
rect 146700 24740 146780 24750
rect 147020 24740 147100 24750
rect 146780 24660 146790 24740
rect 141785 24650 141865 24660
rect 142105 24650 142185 24660
rect 145305 24650 145385 24660
rect 145625 24650 145705 24660
rect 145945 24650 146025 24660
rect 141865 24570 141875 24650
rect 142185 24570 142195 24650
rect 145385 24570 145395 24650
rect 145705 24570 145715 24650
rect 146025 24570 146035 24650
rect 146540 24580 146620 24590
rect 146860 24580 146940 24590
rect 146620 24500 146630 24580
rect 146940 24500 146950 24580
rect 141945 24490 142025 24500
rect 145200 24490 145225 24500
rect 145465 24490 145545 24500
rect 145785 24490 145865 24500
rect 146105 24490 146185 24500
rect 142025 24410 142035 24490
rect 145225 24410 145235 24490
rect 145545 24410 145555 24490
rect 145865 24410 145875 24490
rect 146185 24410 146195 24490
rect 146700 24420 146780 24430
rect 147020 24420 147100 24430
rect 146780 24340 146790 24420
rect 141785 24330 141865 24340
rect 142105 24330 142185 24340
rect 145305 24330 145385 24340
rect 145625 24330 145705 24340
rect 145945 24330 146025 24340
rect 141865 24250 141875 24330
rect 142185 24250 142195 24330
rect 145385 24250 145395 24330
rect 145705 24250 145715 24330
rect 146025 24250 146035 24330
rect 146540 24260 146620 24270
rect 146860 24260 146940 24270
rect 146620 24180 146630 24260
rect 146940 24180 146950 24260
rect 141945 24170 142025 24180
rect 145200 24170 145225 24180
rect 145465 24170 145545 24180
rect 145785 24170 145865 24180
rect 146105 24170 146185 24180
rect 142025 24090 142035 24170
rect 145225 24090 145235 24170
rect 145545 24090 145555 24170
rect 145865 24090 145875 24170
rect 146185 24090 146195 24170
rect 146700 24100 146780 24110
rect 147020 24100 147100 24110
rect 146780 24020 146790 24100
rect 141785 24010 141865 24020
rect 142105 24010 142185 24020
rect 145305 24010 145385 24020
rect 145625 24010 145705 24020
rect 145945 24010 146025 24020
rect 141865 23930 141875 24010
rect 142185 23930 142195 24010
rect 145385 23930 145395 24010
rect 145705 23930 145715 24010
rect 146025 23930 146035 24010
rect 146540 23940 146620 23950
rect 146860 23940 146940 23950
rect 146620 23860 146630 23940
rect 146940 23860 146950 23940
rect 141945 23850 142025 23860
rect 145200 23850 145225 23860
rect 145465 23850 145545 23860
rect 145785 23850 145865 23860
rect 146105 23850 146185 23860
rect 142025 23770 142035 23850
rect 145225 23770 145235 23850
rect 145545 23770 145555 23850
rect 145865 23770 145875 23850
rect 146185 23770 146195 23850
rect 146700 23780 146780 23790
rect 147020 23780 147100 23790
rect 146780 23700 146790 23780
rect 141785 23690 141865 23700
rect 142105 23690 142185 23700
rect 145305 23690 145385 23700
rect 145625 23690 145705 23700
rect 145945 23690 146025 23700
rect 141865 23610 141875 23690
rect 142185 23610 142195 23690
rect 145385 23610 145395 23690
rect 145705 23610 145715 23690
rect 146025 23610 146035 23690
rect 146540 23620 146620 23630
rect 146860 23620 146940 23630
rect 146620 23540 146630 23620
rect 146940 23540 146950 23620
rect 141945 23530 142025 23540
rect 145200 23530 145225 23540
rect 145465 23530 145545 23540
rect 145785 23530 145865 23540
rect 146105 23530 146185 23540
rect 142025 23450 142035 23530
rect 145225 23450 145235 23530
rect 145545 23450 145555 23530
rect 145865 23450 145875 23530
rect 146185 23450 146195 23530
rect 146700 23460 146780 23470
rect 147020 23460 147100 23470
rect 146780 23380 146790 23460
rect 141785 23370 141865 23380
rect 142105 23370 142185 23380
rect 145305 23370 145385 23380
rect 145625 23370 145705 23380
rect 145945 23370 146025 23380
rect 141865 23290 141875 23370
rect 142185 23290 142195 23370
rect 145385 23290 145395 23370
rect 145705 23290 145715 23370
rect 146025 23290 146035 23370
rect 146540 23300 146620 23310
rect 146860 23300 146940 23310
rect 146620 23220 146630 23300
rect 146940 23220 146950 23300
rect 141945 23210 142025 23220
rect 145200 23210 145225 23220
rect 145465 23210 145545 23220
rect 145785 23210 145865 23220
rect 146105 23210 146185 23220
rect 142025 23130 142035 23210
rect 145225 23130 145235 23210
rect 145545 23130 145555 23210
rect 145865 23130 145875 23210
rect 146185 23130 146195 23210
rect 146700 23140 146780 23150
rect 147020 23140 147100 23150
rect 146780 23060 146790 23140
rect 141785 23050 141865 23060
rect 142105 23050 142185 23060
rect 145305 23050 145385 23060
rect 145625 23050 145705 23060
rect 145945 23050 146025 23060
rect 141865 22970 141875 23050
rect 142185 22970 142195 23050
rect 145385 22970 145395 23050
rect 145705 22970 145715 23050
rect 146025 22970 146035 23050
rect 146540 22980 146620 22990
rect 146860 22980 146940 22990
rect 146620 22900 146630 22980
rect 146940 22900 146950 22980
rect 141945 22890 142025 22900
rect 145200 22890 145225 22900
rect 145465 22890 145545 22900
rect 145785 22890 145865 22900
rect 146105 22890 146185 22900
rect 142025 22810 142035 22890
rect 145225 22810 145235 22890
rect 145545 22810 145555 22890
rect 145865 22810 145875 22890
rect 146185 22810 146195 22890
rect 146700 22820 146780 22830
rect 147020 22820 147100 22830
rect 146780 22740 146790 22820
rect 141785 22730 141865 22740
rect 142105 22730 142185 22740
rect 145305 22730 145385 22740
rect 145625 22730 145705 22740
rect 145945 22730 146025 22740
rect 141865 22650 141875 22730
rect 142185 22650 142195 22730
rect 145385 22650 145395 22730
rect 145705 22650 145715 22730
rect 146025 22650 146035 22730
rect 146540 22660 146620 22670
rect 146860 22660 146940 22670
rect 146620 22580 146630 22660
rect 146940 22580 146950 22660
rect 141945 22570 142025 22580
rect 145200 22570 145225 22580
rect 145465 22570 145545 22580
rect 145785 22570 145865 22580
rect 146105 22570 146185 22580
rect 142025 22490 142035 22570
rect 145225 22490 145235 22570
rect 145545 22490 145555 22570
rect 145865 22490 145875 22570
rect 146185 22490 146195 22570
rect 146700 22500 146780 22510
rect 147020 22500 147100 22510
rect 146780 22420 146790 22500
rect 141785 22410 141865 22420
rect 142105 22410 142185 22420
rect 145305 22410 145385 22420
rect 145625 22410 145705 22420
rect 145945 22410 146025 22420
rect 141865 22330 141875 22410
rect 142185 22330 142195 22410
rect 145385 22330 145395 22410
rect 145705 22330 145715 22410
rect 146025 22330 146035 22410
rect 146540 22340 146620 22350
rect 146860 22340 146940 22350
rect 146620 22260 146630 22340
rect 146940 22260 146950 22340
rect 141945 22250 142025 22260
rect 145200 22250 145225 22260
rect 145465 22250 145545 22260
rect 145785 22250 145865 22260
rect 146105 22250 146185 22260
rect 142025 22170 142035 22250
rect 145225 22170 145235 22250
rect 145545 22170 145555 22250
rect 145865 22170 145875 22250
rect 146185 22170 146195 22250
rect 146700 22180 146780 22190
rect 147020 22180 147100 22190
rect 146780 22100 146790 22180
rect 141785 22090 141865 22100
rect 142105 22090 142185 22100
rect 145305 22090 145385 22100
rect 145625 22090 145705 22100
rect 145945 22090 146025 22100
rect 141865 22010 141875 22090
rect 142185 22010 142195 22090
rect 145385 22010 145395 22090
rect 145705 22010 145715 22090
rect 146025 22010 146035 22090
rect 146540 22020 146620 22030
rect 146860 22020 146940 22030
rect 146620 21940 146630 22020
rect 146940 21940 146950 22020
rect 141945 21930 142025 21940
rect 145200 21930 145225 21940
rect 145465 21930 145545 21940
rect 145785 21930 145865 21940
rect 146105 21930 146185 21940
rect 142025 21850 142035 21930
rect 145225 21850 145235 21930
rect 145545 21850 145555 21930
rect 145865 21850 145875 21930
rect 146185 21850 146195 21930
rect 146700 21860 146780 21870
rect 147020 21860 147100 21870
rect 146780 21780 146790 21860
rect 141785 21770 141865 21780
rect 142105 21770 142185 21780
rect 145305 21770 145385 21780
rect 145625 21770 145705 21780
rect 145945 21770 146025 21780
rect 141865 21690 141875 21770
rect 142185 21690 142195 21770
rect 145385 21690 145395 21770
rect 145705 21690 145715 21770
rect 146025 21690 146035 21770
rect 146540 21700 146620 21710
rect 146860 21700 146940 21710
rect 146620 21620 146630 21700
rect 146940 21620 146950 21700
rect 141945 21610 142025 21620
rect 145200 21610 145225 21620
rect 145465 21610 145545 21620
rect 145785 21610 145865 21620
rect 146105 21610 146185 21620
rect 142025 21530 142035 21610
rect 145225 21530 145235 21610
rect 145545 21530 145555 21610
rect 145865 21530 145875 21610
rect 146185 21530 146195 21610
rect 146700 21540 146780 21550
rect 147020 21540 147100 21550
rect 146780 21460 146790 21540
rect 141785 21450 141865 21460
rect 142105 21450 142185 21460
rect 145305 21450 145385 21460
rect 145625 21450 145705 21460
rect 145945 21450 146025 21460
rect 141865 21370 141875 21450
rect 142185 21370 142195 21450
rect 145385 21370 145395 21450
rect 145705 21370 145715 21450
rect 146025 21370 146035 21450
rect 146540 21380 146620 21390
rect 146860 21380 146940 21390
rect 146620 21300 146630 21380
rect 146940 21300 146950 21380
rect 141945 21290 142025 21300
rect 145200 21290 145225 21300
rect 145465 21290 145545 21300
rect 145785 21290 145865 21300
rect 146105 21290 146185 21300
rect 142025 21210 142035 21290
rect 145225 21210 145235 21290
rect 145545 21210 145555 21290
rect 145865 21210 145875 21290
rect 146185 21210 146195 21290
rect 146700 21220 146780 21230
rect 147020 21220 147100 21230
rect 146780 21140 146790 21220
rect 141785 21130 141865 21140
rect 142105 21130 142185 21140
rect 145305 21130 145385 21140
rect 145625 21130 145705 21140
rect 145945 21130 146025 21140
rect 141865 21050 141875 21130
rect 142185 21050 142195 21130
rect 145385 21050 145395 21130
rect 145705 21050 145715 21130
rect 146025 21050 146035 21130
rect 146540 21060 146620 21070
rect 146860 21060 146940 21070
rect 146620 20980 146630 21060
rect 146940 20980 146950 21060
rect 141945 20970 142025 20980
rect 145200 20970 145225 20980
rect 145465 20970 145545 20980
rect 145785 20970 145865 20980
rect 146105 20970 146185 20980
rect 142025 20890 142035 20970
rect 145225 20890 145235 20970
rect 145545 20890 145555 20970
rect 145865 20890 145875 20970
rect 146185 20890 146195 20970
rect 146700 20900 146780 20910
rect 147020 20900 147100 20910
rect 146780 20820 146790 20900
rect 141785 20810 141865 20820
rect 142105 20810 142185 20820
rect 145305 20810 145385 20820
rect 145625 20810 145705 20820
rect 145945 20810 146025 20820
rect 141865 20730 141875 20810
rect 142185 20730 142195 20810
rect 145385 20730 145395 20810
rect 145705 20730 145715 20810
rect 146025 20730 146035 20810
rect 146540 20740 146620 20750
rect 146860 20740 146940 20750
rect 146620 20660 146630 20740
rect 146940 20660 146950 20740
rect 141945 20650 142025 20660
rect 145200 20650 145225 20660
rect 145465 20650 145545 20660
rect 145785 20650 145865 20660
rect 146105 20650 146185 20660
rect 142025 20570 142035 20650
rect 145225 20570 145235 20650
rect 145545 20570 145555 20650
rect 145865 20570 145875 20650
rect 146185 20570 146195 20650
rect 146700 20580 146780 20590
rect 147020 20580 147100 20590
rect 146780 20500 146790 20580
rect 141785 20490 141865 20500
rect 142105 20490 142185 20500
rect 145305 20490 145385 20500
rect 145625 20490 145705 20500
rect 145945 20490 146025 20500
rect 141865 20410 141875 20490
rect 142185 20410 142195 20490
rect 145385 20410 145395 20490
rect 145705 20410 145715 20490
rect 146025 20410 146035 20490
rect 146540 20420 146620 20430
rect 146860 20420 146940 20430
rect 146620 20340 146630 20420
rect 146940 20340 146950 20420
rect 141945 20330 142025 20340
rect 145200 20330 145225 20340
rect 145465 20330 145545 20340
rect 145785 20330 145865 20340
rect 146105 20330 146185 20340
rect 142025 20250 142035 20330
rect 145225 20250 145235 20330
rect 145545 20250 145555 20330
rect 145865 20250 145875 20330
rect 146185 20250 146195 20330
rect 146700 20260 146780 20270
rect 147020 20260 147100 20270
rect 146780 20180 146790 20260
rect 141785 20170 141865 20180
rect 142105 20170 142185 20180
rect 145305 20170 145385 20180
rect 145625 20170 145705 20180
rect 145945 20170 146025 20180
rect 141865 20090 141875 20170
rect 142185 20090 142195 20170
rect 145385 20090 145395 20170
rect 145705 20090 145715 20170
rect 146025 20090 146035 20170
rect 146540 20100 146620 20110
rect 146860 20100 146940 20110
rect 146620 20020 146630 20100
rect 146940 20020 146950 20100
rect 141945 20010 142025 20020
rect 145200 20010 145225 20020
rect 145465 20010 145545 20020
rect 145785 20010 145865 20020
rect 146105 20010 146185 20020
rect 142025 19930 142035 20010
rect 145225 19930 145235 20010
rect 145545 19930 145555 20010
rect 145865 19930 145875 20010
rect 146185 19930 146195 20010
rect 146700 19940 146780 19950
rect 147020 19940 147100 19950
rect 146780 19860 146790 19940
rect 141785 19850 141865 19860
rect 142105 19850 142185 19860
rect 145305 19850 145385 19860
rect 145625 19850 145705 19860
rect 145945 19850 146025 19860
rect 141865 19770 141875 19850
rect 142185 19770 142195 19850
rect 145385 19770 145395 19850
rect 145705 19770 145715 19850
rect 146025 19770 146035 19850
rect 146540 19780 146620 19790
rect 146860 19780 146940 19790
rect 146620 19700 146630 19780
rect 146940 19700 146950 19780
rect 141945 19690 142025 19700
rect 145200 19690 145225 19700
rect 145465 19690 145545 19700
rect 145785 19690 145865 19700
rect 146105 19690 146185 19700
rect 142025 19610 142035 19690
rect 145225 19610 145235 19690
rect 145545 19610 145555 19690
rect 145865 19610 145875 19690
rect 146185 19610 146195 19690
rect 146700 19620 146780 19630
rect 147020 19620 147100 19630
rect 146780 19540 146790 19620
rect 141785 19530 141865 19540
rect 142105 19530 142185 19540
rect 145305 19530 145385 19540
rect 145625 19530 145705 19540
rect 145945 19530 146025 19540
rect 141865 19450 141875 19530
rect 142185 19450 142195 19530
rect 145385 19450 145395 19530
rect 145705 19450 145715 19530
rect 146025 19450 146035 19530
rect 146540 19460 146620 19470
rect 146860 19460 146940 19470
rect 146620 19380 146630 19460
rect 146940 19380 146950 19460
rect 141945 19370 142025 19380
rect 145200 19370 145225 19380
rect 145465 19370 145545 19380
rect 145785 19370 145865 19380
rect 146105 19370 146185 19380
rect 142025 19290 142035 19370
rect 145225 19290 145235 19370
rect 145545 19290 145555 19370
rect 145865 19290 145875 19370
rect 146185 19290 146195 19370
rect 146700 19300 146780 19310
rect 147020 19300 147100 19310
rect 146780 19220 146790 19300
rect 141785 19210 141865 19220
rect 142105 19210 142185 19220
rect 145305 19210 145385 19220
rect 145625 19210 145705 19220
rect 145945 19210 146025 19220
rect 141865 19130 141875 19210
rect 142185 19130 142195 19210
rect 145385 19130 145395 19210
rect 145705 19130 145715 19210
rect 146025 19130 146035 19210
rect 146540 19140 146620 19150
rect 146860 19140 146940 19150
rect 146620 19060 146630 19140
rect 146940 19060 146950 19140
rect 141945 19050 142025 19060
rect 145200 19050 145225 19060
rect 145465 19050 145545 19060
rect 145785 19050 145865 19060
rect 146105 19050 146185 19060
rect 142025 18970 142035 19050
rect 145225 18970 145235 19050
rect 145545 18970 145555 19050
rect 145865 18970 145875 19050
rect 146185 18970 146195 19050
<< metal1 >>
rect 103800 143060 104500 144200
rect 106100 143700 144145 144500
rect 143245 140000 144145 143700
rect 143650 114035 143860 114460
rect 143650 113320 144075 113530
rect 145400 87120 145650 103000
rect 145395 86800 145910 87120
rect 45955 75940 46235 76360
rect 143690 59375 143900 59815
rect 143740 57040 144260 57255
rect 145400 56820 145650 86800
rect 143740 56440 144260 56655
rect 98400 46240 99600 46475
rect 98400 45900 98700 46240
rect 60120 45600 98700 45900
rect 99000 45600 106555 45900
rect 99000 45300 99300 45600
rect 73620 45000 99300 45300
rect 73300 44135 73620 45000
<< m2contact >>
rect 106100 144500 113245 146000
rect 143440 115960 143860 116260
rect 145400 103000 145940 103320
rect 45655 78080 46530 84930
rect 145400 56440 145650 56820
rect 99600 46240 100050 46475
rect 59800 45445 60120 45900
rect 106555 45600 106945 45900
rect 73300 45000 73620 45300
<< metal2 >>
rect 49000 145510 49320 145940
rect 62500 144205 62820 145940
rect 76000 142900 76320 145940
rect 76000 142100 79780 142900
rect 79235 140900 79780 142100
rect 89500 141350 89820 145940
rect 101700 140800 102440 142970
rect 103800 140800 104500 143060
rect 116500 141800 116820 145940
rect 130000 143100 130320 145940
rect 130000 142400 135745 143100
rect 116500 141100 133045 141800
rect 135300 141000 135745 142400
rect 44060 129880 45500 130200
rect 44060 116380 44900 116700
rect 44500 105415 44900 116380
rect 45100 106015 45500 129880
rect 144900 130000 145940 130320
rect 143650 113530 143860 114035
rect 44900 105040 45720 105160
rect 44500 103200 44900 104185
rect 44060 102880 44900 103200
rect 45500 103840 45996 103960
rect 45100 102500 45500 103585
rect 44500 102100 45500 102500
rect 44500 89699 44900 102100
rect 44060 89379 44900 89699
rect 42300 78080 45655 84930
rect 44500 75940 45955 76360
rect 44500 62700 44900 75940
rect 44060 62380 44900 62700
rect 144400 59585 144650 116360
rect 143900 59375 144650 59585
rect 144900 57255 145150 130000
rect 144260 57040 145150 57255
rect 144260 56440 145400 56655
rect 44060 48880 45100 49200
rect 59800 44060 60120 45445
rect 67540 45000 67645 46265
rect 94240 45600 94505 46345
rect 94840 46200 94945 46365
rect 106840 45900 106945 46350
rect 107440 45300 107545 46285
rect 73300 44135 73620 45000
rect 99600 45000 107545 45300
rect 99600 44400 99900 45000
rect 108640 44400 108745 46465
rect 86800 44100 99900 44400
rect 100300 44100 108745 44400
rect 113800 44060 114120 44535
rect 127300 44060 127620 45200
rect 140800 44060 141120 45775
<< m3contact >>
rect 49000 144700 50845 145510
rect 62500 143400 64455 144205
rect 77850 140900 78750 141350
rect 88400 140900 89820 141350
rect 101700 142970 102440 144200
rect 103800 143060 104500 144200
rect 144400 116360 144650 116820
rect 143440 115540 143860 115960
rect 143650 114035 143860 114460
rect 143650 113320 144075 113530
rect 45100 105640 45500 106015
rect 44500 105040 44900 105415
rect 44500 104185 44900 104560
rect 45100 103585 45500 103960
rect 45955 75940 46360 76360
rect 143690 59375 143900 59815
rect 145440 116500 145940 116820
rect 145650 100300 145940 100905
rect 145395 86800 145940 87120
rect 145360 73300 145940 73620
rect 145545 59800 145940 60120
rect 143740 57040 144260 57255
rect 143740 56440 144260 56655
rect 45100 48880 45500 49415
rect 94840 45900 95325 46200
rect 94240 45300 94725 45600
rect 67540 44700 68070 45000
rect 140800 45775 141120 46200
rect 127300 45200 127620 45600
rect 113800 44535 114120 45000
<< metal3 >>
rect 50845 144700 104500 145500
rect 103800 144200 104500 144700
rect 64455 143400 101700 144200
rect 78750 140900 88400 141350
rect 144650 116500 145440 116820
rect 144105 113740 145900 113950
rect 144075 113320 145400 113530
rect 143695 112240 144900 112360
rect 143840 111640 144400 111760
rect 45500 105640 46315 105760
rect 44900 105040 46590 105160
rect 44900 104440 46785 104560
rect 45500 103840 46530 103960
rect 45100 101440 47970 101561
rect 45100 49415 45500 101440
rect 143690 59815 143900 60460
rect 144150 60120 144400 111640
rect 144650 73620 144900 112240
rect 145150 87120 145400 113320
rect 145650 100905 145900 113740
rect 145150 86800 145395 87120
rect 144650 73300 145360 73620
rect 144150 59800 145545 60120
rect 95325 45900 140800 46200
rect 94725 45300 127300 45600
rect 68070 44700 113800 45000
use PIC  CIN0_2 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN1_6
timestamp 1537935238
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN2_5
timestamp 1537935238
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN3_11
timestamp 1537935238
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  CIN4_15
timestamp 1537935238
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  CIN5_16
timestamp 1537935238
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  CIN6_17
timestamp 1537935238
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  CLK_4
timestamp 1537935238
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1718295485
transform 1 0 46600 0 1 46600
box -945 -360 97560 94545
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1709081121
transform 0 -1 171100 -1 0 75646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_1
timestamp 1709081121
transform 0 -1 171100 -1 0 62146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_2
timestamp 1709081121
transform 0 -1 171100 -1 0 102646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_3
timestamp 1709081121
transform 0 -1 171100 -1 0 89146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_4
timestamp 1709081121
transform 0 -1 171100 -1 0 129646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_5
timestamp 1709081121
transform 0 -1 171100 -1 0 116146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_6
timestamp 1709081121
transform 1 0 73845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_7
timestamp 1709081121
transform 1 0 60345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_8
timestamp 1709081121
transform 1 0 100845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_9
timestamp 1709081121
transform 1 0 87345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_10
timestamp 1709081121
transform 1 0 127845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_11
timestamp 1709081121
transform 1 0 114345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_12
timestamp 1709081121
transform 0 1 18900 -1 0 75655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_13
timestamp 1709081121
transform 0 1 18900 -1 0 62155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_14
timestamp 1709081121
transform 0 1 18900 -1 0 102655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_15
timestamp 1709081121
transform 0 1 18900 -1 0 89155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_16
timestamp 1709081121
transform 1 0 73845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_17
timestamp 1709081121
transform 0 1 18900 -1 0 116155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_18
timestamp 1709081121
transform 0 1 18900 -1 0 129655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_19
timestamp 1709081121
transform 1 0 60345 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_20
timestamp 1709081121
transform 1 0 100845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_21
timestamp 1709081121
transform 1 0 87345 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_22
timestamp 1709081121
transform 1 0 127845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_23
timestamp 1709081121
transform 1 0 114345 0 -1 171099
box 0 0 1810 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 43675 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 141375 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 43675 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 18900 -1 0 48685
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 18900 -1 0 146205
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 171100 -1 0 146325
box -35 0 5035 25060
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PVDD  PVDD_10 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 0 1 18900 -1 0 87500
box 0 -9150 12000 25300
use PVSS  PVSS_22 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 102500 0 -1 171100
box 0 -9150 12000 25300
use PIC  RDY_3
timestamp 1537935238
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  VLD_14 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use PIC  XIN0_12
timestamp 1537935238
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN1_9
timestamp 1537935238
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN2_27
timestamp 1537935238
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  XIN3_13
timestamp 1537935238
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use POB8  XOUT0_24
timestamp 1537935238
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT1_23
timestamp 1537935238
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT2_21
timestamp 1537935238
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT3_20
timestamp 1537935238
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  YIN0_1
timestamp 1537935238
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN1_0
timestamp 1537935238
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN2_7
timestamp 1537935238
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PIC  YIN3_8
timestamp 1537935238
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB8  YOUT0_19
timestamp 1537935238
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  YOUT1_18
timestamp 1537935238
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB8  YOUT2_25
timestamp 1537935238
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT3_26
timestamp 1537935238
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
<< end >>
