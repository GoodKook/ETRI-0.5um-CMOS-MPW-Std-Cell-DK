magic
tech scmos
magscale 1 30
timestamp 1537935238
<< checkpaint >>
rect -700 -9750 12700 25951
<< metal2 >>
rect 255 25160 575 25300
rect 1720 25160 2040 25300
rect 11300 25160 11620 25300
use CMD_TR  CMD_TR_0
timestamp 1537935238
transform 1 0 7620 0 1 23990
box 50 -175 1270 890
use DOUBLE_GUARD  DOUBLE_GUARD_0
timestamp 1537935238
transform 1 0 0 0 1 8300
box -100 -100 12095 2500
use GUARD  GUARD_0
timestamp 1537935238
transform 1 0 0 0 1 21100
box -100 -100 12095 3960
use INV2  INV2_0
timestamp 1537935238
transform 1 0 9570 0 1 21570
box -10 -210 2130 3230
use INV  INV_0
timestamp 1537935238
transform 1 0 8690 0 1 21570
box -10 -210 930 3070
use LTSLOGIC  LTSLOGIC_0
timestamp 1537935238
transform 1 0 300 0 1 21100
box 0 -300 5590 4200
use METAL_RING  METAL_RING_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 0 0 12000 25060
use NDRV  NDRV_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 0 0 12000 7800
use PAD_80  PAD_80_0
timestamp 1537935238
transform 1 0 6000 0 1 -4900
box -4250 -4250 4250 4900
use PAD_METAL_PBCT4  PAD_METAL_PBCT4_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 0 0 12000 25300
use PDRV  PDRV_0
timestamp 1537935238
transform 1 0 0 0 1 11300
box -100 -100 12100 7900
use SINGLE_GUARD  SINGLE_GUARD_0
timestamp 1537935238
transform 1 0 0 0 1 19600
box 0 0 12000 1000
<< labels >>
flabel space 6000 -4900 6000 -4900 0 FreeSans 5000 0 0 0 PAD
flabel m3p s 0 15090 0 15090 0 FreeSans 5000 0 0 0 VDD
flabel m3p s 0 21695 0 21695 0 FreeSans 5000 0 0 0 VDD
flabel m3p s 0 23940 0 23940 0 FreeSans 5000 0 0 0 VSS
flabel m3p s 0 3760 0 3760 0 FreeSans 5000 0 0 0 VSS
flabel m2p s 11460 25300 11460 25300 0 FreeSans 2000 0 0 0 Y
flabel m2p s 1895 25300 1895 25300 0 FreeSans 2000 0 0 0 A
flabel m2p s 405 25300 405 25300 0 FreeSans 2000 0 0 0 OE
<< end >>
