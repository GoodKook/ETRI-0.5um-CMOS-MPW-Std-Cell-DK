magic
tech scmos
magscale 1 6
timestamp 1725338759
<< checkpaint >>
rect -66 350 206 402
rect -92 346 232 350
rect -92 -90 286 346
<< nwell >>
rect 0 0 176 260
<< ptransistor >>
rect 65 30 75 230
<< pdiffusion >>
rect 62 30 65 230
rect 75 30 78 230
<< ndcontact >>
rect 134 30 166 226
<< pdcontact >>
rect 28 30 62 230
rect 78 30 112 230
<< polysilicon >>
rect 65 230 75 250
rect 65 20 75 30
<< polycontact >>
rect 54 250 86 282
<< metal1 >>
rect 52 282 88 284
rect 52 250 54 282
rect 86 250 88 282
rect 52 248 88 250
rect 26 230 62 232
rect 26 30 28 230
rect 26 28 62 30
rect 78 230 114 232
rect 112 30 114 230
rect 78 28 114 30
rect 132 226 168 228
rect 132 30 134 226
rect 166 30 168 226
rect 132 28 168 30
<< end >>
