magic
tech scmos
magscale 1 2
timestamp 1727443468
<< checkpaint >>
rect 1133 2416 1227 2521
<< error_s >>
rect 4 5464 5536 5476
rect 4 5204 5536 5216
rect 4 4944 5536 4956
rect 4 4684 5536 4696
rect 4 4424 5536 4436
rect 4 4164 5536 4176
rect 4 3904 5536 3916
rect 4 3644 5536 3656
rect 4 3384 5536 3396
rect 4 3124 5536 3136
rect 4 2864 5536 2876
rect 4 2604 5536 2616
rect 4 2344 5536 2356
rect 4 2084 5536 2096
rect 4 1824 5536 1836
rect 4 1564 5536 1576
rect 4 1304 5536 1316
rect 4 1044 5536 1056
rect 4 784 5536 796
rect 4 524 5536 536
rect 4 264 5536 276
rect 4 4 5536 16
<< nwell >>
rect 664 4076 690 4084
<< metal1 >>
rect -63 5218 -3 5478
rect 5510 5462 5603 5478
rect 647 5403 660 5407
rect 647 5397 673 5403
rect 4767 5397 4813 5403
rect 647 5393 660 5397
rect 47 5373 53 5387
rect 447 5377 513 5383
rect 1567 5377 1613 5383
rect 1827 5377 1873 5383
rect 2167 5373 2173 5387
rect 2287 5373 2293 5387
rect 2667 5383 2680 5387
rect 2667 5377 2693 5383
rect 2667 5373 2680 5377
rect 2907 5377 2953 5383
rect 3047 5377 3093 5383
rect 3147 5373 3153 5387
rect 3247 5377 3313 5383
rect 3760 5383 3773 5387
rect 3747 5377 3773 5383
rect 3760 5373 3773 5377
rect 3867 5377 3953 5383
rect 4307 5377 4373 5383
rect 4647 5377 4693 5383
rect 4980 5383 4993 5387
rect 4967 5377 4993 5383
rect 4980 5373 4993 5377
rect 5107 5377 5193 5383
rect 487 5357 553 5363
rect 621 5357 653 5363
rect 4413 5367 4427 5373
rect 4207 5357 4253 5363
rect 4527 5353 4533 5367
rect 367 5333 373 5347
rect 827 5343 840 5347
rect 827 5337 853 5343
rect 827 5333 840 5337
rect 1747 5337 1793 5343
rect 1947 5333 1953 5347
rect 3187 5343 3200 5347
rect 3187 5337 3213 5343
rect 3187 5333 3200 5337
rect 1307 5317 1373 5323
rect 1707 5317 1753 5323
rect 2467 5313 2472 5327
rect 2507 5317 2553 5323
rect 2807 5323 2820 5327
rect 2807 5317 2833 5323
rect 2807 5313 2820 5317
rect 3627 5313 3633 5327
rect 3927 5317 3973 5323
rect 4300 5323 4313 5327
rect 4287 5317 4313 5323
rect 4300 5313 4313 5317
rect 5280 5323 5293 5327
rect 5267 5317 5293 5323
rect 5280 5313 5293 5317
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 1327 5097 1373 5103
rect 1627 5097 1673 5103
rect 2047 5103 2060 5107
rect 2047 5097 2073 5103
rect 2047 5093 2060 5097
rect 2187 5093 2193 5107
rect 2307 5103 2320 5107
rect 2307 5097 2333 5103
rect 2307 5093 2320 5097
rect 2667 5093 2673 5107
rect 3007 5093 3013 5107
rect 3247 5093 3253 5107
rect 3580 5103 3593 5107
rect 3567 5097 3593 5103
rect 3580 5093 3593 5097
rect 187 5073 193 5087
rect 1047 5077 1113 5083
rect 2447 5073 2453 5087
rect 2727 5077 2793 5083
rect 3900 5083 3913 5087
rect 3887 5077 3913 5083
rect 3900 5073 3913 5077
rect 4061 5077 4093 5083
rect 727 5057 773 5063
rect 3047 5066 3063 5067
rect 3047 5053 3053 5066
rect 3687 5060 3723 5063
rect 3687 5057 3727 5060
rect 4227 5057 4273 5063
rect 287 5033 292 5047
rect 317 5040 393 5043
rect 313 5037 393 5040
rect 153 5027 167 5033
rect 313 5027 327 5037
rect 1080 5043 1093 5047
rect 1067 5037 1093 5043
rect 1080 5033 1093 5037
rect 1347 5037 1433 5043
rect 1547 5033 1553 5047
rect 1787 5043 1800 5047
rect 1787 5037 1813 5043
rect 1787 5033 1800 5037
rect 2007 5033 2013 5047
rect 2267 5037 2313 5043
rect 3713 5047 3727 5057
rect 4340 5063 4353 5067
rect 4327 5057 4353 5063
rect 4340 5053 4353 5057
rect 4540 5063 4553 5067
rect 4527 5057 4553 5063
rect 4540 5053 4553 5057
rect 2517 5037 2553 5043
rect 2517 5003 2523 5037
rect 3167 5037 3233 5043
rect 3347 5043 3360 5047
rect 3347 5037 3373 5043
rect 3347 5033 3360 5037
rect 4027 5037 4073 5043
rect 4787 5037 4853 5043
rect 4947 5033 4953 5047
rect 5367 5033 5372 5047
rect 5407 5043 5420 5047
rect 5407 5037 5433 5043
rect 5407 5033 5420 5037
rect 4427 5017 4493 5023
rect 2487 4997 2523 5003
rect 5543 4958 5603 5462
rect 5510 4942 5603 4958
rect 967 4883 980 4887
rect 967 4873 983 4883
rect 633 4867 647 4873
rect 147 4857 213 4863
rect 267 4857 313 4863
rect 567 4857 633 4863
rect 687 4857 733 4863
rect 867 4853 873 4867
rect 187 4813 193 4827
rect 587 4823 600 4827
rect 587 4817 613 4823
rect 587 4813 600 4817
rect 977 4826 983 4873
rect 4327 4877 4393 4883
rect 1107 4857 1153 4863
rect 1197 4857 1233 4863
rect 1667 4853 1673 4867
rect 1787 4857 1852 4863
rect 1887 4853 1893 4867
rect 2107 4857 2173 4863
rect 2647 4857 2693 4863
rect 2747 4857 2793 4863
rect 2893 4863 2907 4873
rect 2893 4860 2933 4863
rect 2897 4857 2933 4860
rect 3167 4853 3173 4867
rect 3267 4853 3273 4867
rect 3807 4853 3813 4867
rect 4220 4863 4233 4867
rect 4207 4857 4233 4863
rect 4220 4854 4233 4857
rect 4477 4857 4533 4863
rect 4220 4853 4240 4854
rect 2307 4833 2313 4847
rect 2847 4833 2853 4847
rect 3973 4843 3987 4853
rect 3927 4840 3987 4843
rect 3927 4837 3983 4840
rect 4477 4843 4483 4857
rect 4427 4837 4483 4843
rect 5307 4837 5353 4843
rect 4667 4817 4713 4823
rect 467 4803 480 4807
rect 467 4797 493 4803
rect 467 4793 480 4797
rect 1367 4793 1373 4807
rect 2100 4803 2113 4807
rect 2087 4797 2113 4803
rect 2100 4793 2113 4797
rect 2407 4803 2420 4807
rect 2407 4797 2433 4803
rect 2407 4793 2420 4797
rect 2547 4803 2560 4807
rect 2547 4797 2573 4803
rect 2547 4793 2560 4797
rect 5267 4793 5273 4807
rect 5427 4793 5433 4807
rect 1437 4777 1473 4783
rect 1827 4717 1853 4723
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 2727 4617 2753 4623
rect 2847 4597 2883 4603
rect 2313 4587 2327 4593
rect 1027 4573 1033 4587
rect 1147 4583 1160 4587
rect 1537 4586 1553 4587
rect 1147 4577 1173 4583
rect 1147 4573 1160 4577
rect 267 4553 273 4567
rect 673 4563 687 4573
rect 1547 4573 1553 4586
rect 2267 4573 2273 4587
rect 673 4560 713 4563
rect 677 4557 713 4560
rect 1707 4553 1713 4567
rect 2187 4537 2233 4543
rect 2307 4533 2313 4547
rect 2877 4543 2883 4597
rect 3007 4593 3013 4607
rect 2927 4573 2933 4587
rect 4467 4573 4473 4587
rect 4607 4573 4613 4587
rect 4747 4573 4753 4587
rect 4867 4577 4913 4583
rect 3867 4557 3913 4563
rect 4047 4557 4073 4563
rect 4087 4553 4093 4567
rect 2877 4537 2913 4543
rect 3037 4540 3073 4543
rect 3033 4537 3073 4540
rect 3033 4527 3047 4537
rect 3767 4537 3813 4543
rect 5307 4537 5373 4543
rect 247 4517 293 4523
rect 347 4513 352 4527
rect 387 4523 400 4527
rect 387 4517 413 4523
rect 467 4517 512 4523
rect 387 4513 400 4517
rect 547 4523 560 4527
rect 547 4517 573 4523
rect 547 4513 560 4517
rect 1347 4513 1353 4527
rect 2367 4513 2373 4527
rect 2687 4517 2733 4523
rect 2827 4517 2873 4523
rect 3200 4523 3213 4527
rect 3187 4517 3213 4523
rect 3200 4513 3213 4517
rect 3327 4513 3333 4527
rect 3427 4513 3433 4527
rect 3487 4517 3533 4523
rect 3557 4507 3563 4533
rect 3987 4517 4073 4523
rect 4207 4513 4213 4527
rect 1887 4497 1933 4503
rect 3807 4497 3833 4503
rect 5057 4497 5113 4503
rect 5057 4487 5063 4497
rect 5047 4477 5063 4487
rect 5047 4473 5060 4477
rect 967 4457 1013 4463
rect 5543 4438 5603 4942
rect 5510 4422 5603 4438
rect 927 4363 940 4367
rect 927 4357 953 4363
rect 927 4353 940 4357
rect 3607 4357 3653 4363
rect 5187 4357 5253 4363
rect 620 4343 633 4347
rect 487 4337 553 4343
rect 607 4337 633 4343
rect 620 4333 633 4337
rect 1247 4333 1253 4347
rect 1360 4346 1380 4347
rect 1367 4343 1380 4346
rect 1367 4337 1393 4343
rect 1367 4333 1380 4337
rect 1707 4333 1713 4347
rect 3433 4347 3447 4353
rect 2667 4337 2713 4343
rect 3747 4337 3813 4343
rect 4667 4337 4753 4343
rect 1027 4323 1040 4327
rect 1027 4317 1053 4323
rect 1027 4313 1040 4317
rect 1167 4317 1213 4323
rect 1807 4317 1853 4323
rect 2347 4313 2353 4327
rect 2547 4317 2593 4323
rect 3007 4317 3073 4323
rect 4247 4317 4293 4323
rect 5193 4323 5207 4333
rect 5167 4320 5207 4323
rect 5167 4317 5203 4320
rect 5313 4323 5327 4333
rect 5313 4320 5353 4323
rect 5317 4317 5353 4320
rect 467 4293 473 4307
rect 527 4293 533 4307
rect 687 4293 693 4307
rect 1627 4293 1633 4307
rect 2193 4303 2207 4313
rect 2193 4300 2253 4303
rect 2197 4297 2253 4300
rect 2647 4297 2693 4303
rect 3187 4297 3233 4303
rect 3393 4303 3407 4313
rect 3367 4300 3407 4303
rect 3367 4297 3403 4300
rect 4207 4293 4213 4307
rect 4427 4297 4473 4303
rect 4747 4303 4760 4307
rect 4747 4297 4773 4303
rect 4787 4297 4833 4303
rect 4747 4293 4760 4297
rect 1633 4287 1647 4293
rect 5447 4293 5453 4307
rect 67 4273 73 4287
rect 167 4283 180 4287
rect 167 4277 193 4283
rect 167 4273 180 4277
rect 1840 4286 1860 4287
rect 1840 4283 1853 4286
rect 1827 4277 1853 4283
rect 1840 4273 1853 4277
rect 1773 4267 1787 4273
rect 2167 4277 2213 4283
rect 2367 4277 2413 4283
rect 2787 4277 2833 4283
rect 3887 4273 3893 4287
rect 4927 4277 4972 4283
rect 5007 4273 5013 4287
rect 2313 4267 2327 4273
rect 327 4253 333 4267
rect 5087 4253 5093 4267
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 367 4057 413 4063
rect 2267 4063 2280 4067
rect 2267 4057 2293 4063
rect 2267 4053 2280 4057
rect 2887 4053 2893 4067
rect 3840 4063 3853 4067
rect 3827 4057 3853 4063
rect 3840 4053 3853 4057
rect 4267 4053 4273 4067
rect 4667 4057 4713 4063
rect 5367 4063 5380 4067
rect 5367 4057 5393 4063
rect 5367 4053 5380 4057
rect 1553 4043 1567 4053
rect 2693 4047 2707 4053
rect 1553 4040 1593 4043
rect 1557 4037 1593 4040
rect 3507 4033 3513 4047
rect 4887 4037 4973 4043
rect 5087 4033 5093 4047
rect 5187 4037 5233 4043
rect 100 4023 113 4027
rect 87 4017 113 4023
rect 100 4013 113 4017
rect 787 4017 833 4023
rect 2220 4023 2233 4027
rect 2207 4017 2233 4023
rect 2220 4013 2233 4017
rect 2407 4023 2420 4027
rect 2407 4017 2433 4023
rect 2407 4013 2420 4017
rect 2907 4013 2913 4027
rect 3340 4023 3353 4027
rect 3267 4017 3313 4023
rect 3327 4017 3353 4023
rect 3340 4013 3353 4017
rect 2733 4007 2747 4013
rect 3607 4017 3633 4023
rect 3687 4017 3733 4023
rect 4007 4013 4013 4027
rect 4067 4017 4113 4023
rect 487 3997 573 4003
rect 1640 4003 1653 4007
rect 1627 3997 1653 4003
rect 1640 3993 1653 3997
rect 1867 3997 1953 4003
rect 2047 4003 2060 4007
rect 2047 3997 2073 4003
rect 2047 3993 2060 3997
rect 2627 3997 2673 4003
rect 3087 3997 3153 4003
rect 3847 3997 3893 4003
rect 4387 3993 4393 4007
rect 4527 3997 4593 4003
rect 4747 3993 4753 4007
rect 3407 3973 3413 3987
rect 127 3957 173 3963
rect 5543 3918 5603 4422
rect 5510 3902 5603 3918
rect 1500 3843 1513 3847
rect 1497 3833 1513 3843
rect 4767 3833 4773 3847
rect 5127 3837 5193 3843
rect 5287 3833 5293 3847
rect 5440 3843 5453 3847
rect 5427 3837 5453 3843
rect 5440 3833 5453 3837
rect 247 3817 293 3823
rect 587 3817 653 3823
rect 787 3813 793 3827
rect 807 3813 813 3827
rect 987 3817 1033 3823
rect 1207 3817 1253 3823
rect 1367 3813 1373 3827
rect 1497 3823 1503 3833
rect 1427 3817 1503 3823
rect 1907 3823 1920 3827
rect 1907 3817 1933 3823
rect 1907 3813 1920 3817
rect 2087 3817 2153 3823
rect 2687 3813 2693 3827
rect 2760 3823 2773 3827
rect 2747 3817 2773 3823
rect 2760 3813 2773 3817
rect 2887 3817 2933 3823
rect 3307 3817 3373 3823
rect 3647 3813 3653 3827
rect 3807 3817 3873 3823
rect 4187 3817 4233 3823
rect 4427 3813 4433 3827
rect 4567 3813 4573 3827
rect 4907 3813 4913 3827
rect 947 3797 993 3803
rect 1307 3793 1313 3807
rect 1507 3803 1520 3807
rect 1507 3797 1533 3803
rect 1507 3793 1520 3797
rect 2307 3803 2320 3807
rect 2307 3797 2333 3803
rect 2307 3793 2320 3797
rect 2827 3793 2833 3807
rect 3200 3803 3213 3807
rect 3187 3797 3213 3803
rect 3200 3793 3213 3797
rect 4087 3793 4093 3807
rect 4287 3797 4333 3803
rect 4487 3803 4500 3807
rect 4487 3797 4513 3803
rect 4647 3797 4713 3803
rect 4487 3793 4500 3797
rect 1967 3773 1973 3787
rect 2240 3783 2253 3787
rect 2227 3777 2253 3783
rect 2240 3773 2253 3777
rect 3087 3773 3093 3787
rect 3627 3773 3633 3787
rect 3687 3777 3773 3783
rect 5120 3783 5133 3787
rect 5107 3777 5133 3783
rect 5120 3773 5133 3777
rect 167 3753 173 3767
rect 657 3766 673 3767
rect 667 3753 673 3766
rect 4247 3753 4253 3767
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 1007 3577 1033 3583
rect 187 3553 193 3567
rect 1400 3543 1413 3547
rect 1387 3537 1413 3543
rect 1400 3533 1413 3537
rect 2413 3547 2427 3553
rect 3907 3533 3913 3547
rect 5287 3543 5300 3547
rect 5287 3537 5313 3543
rect 5287 3533 5300 3537
rect 327 3513 333 3527
rect 760 3526 780 3527
rect 760 3523 773 3526
rect 747 3517 773 3523
rect 760 3513 773 3517
rect 2977 3517 3013 3523
rect 2693 3507 2707 3513
rect 967 3493 973 3507
rect 1967 3493 1973 3507
rect 2047 3493 2053 3507
rect 2167 3493 2173 3507
rect 2460 3503 2473 3507
rect 2447 3497 2473 3503
rect 2460 3493 2473 3497
rect 2977 3503 2983 3517
rect 2927 3497 2983 3503
rect 3173 3507 3187 3513
rect 3413 3507 3427 3513
rect 3607 3497 3653 3503
rect 3947 3503 3960 3507
rect 3947 3497 3973 3503
rect 4087 3497 4133 3503
rect 3947 3493 3960 3497
rect 4640 3503 4653 3507
rect 4447 3497 4493 3503
rect 4627 3497 4653 3503
rect 4640 3494 4653 3497
rect 4640 3493 4660 3494
rect 5167 3503 5180 3507
rect 5167 3497 5193 3503
rect 5167 3493 5180 3497
rect 5433 3487 5447 3493
rect 47 3483 60 3487
rect 47 3477 73 3483
rect 47 3473 60 3477
rect 437 3486 453 3487
rect 447 3473 453 3486
rect 687 3483 700 3487
rect 687 3477 713 3483
rect 687 3473 700 3477
rect 1067 3473 1073 3487
rect 1167 3477 1233 3483
rect 1547 3477 1593 3483
rect 1787 3477 1833 3483
rect 2507 3473 2513 3487
rect 3787 3473 3793 3487
rect 3807 3477 3833 3483
rect 4240 3483 4253 3487
rect 4227 3477 4253 3483
rect 4240 3473 4253 3477
rect 4387 3473 4393 3487
rect 4667 3477 4713 3483
rect 5027 3477 5073 3483
rect 5487 3473 5493 3487
rect 4807 3457 4853 3463
rect 5543 3398 5603 3902
rect 5510 3382 5603 3398
rect 3817 3337 3853 3343
rect 1027 3317 1113 3323
rect 3547 3317 3593 3323
rect 3817 3323 3823 3337
rect 3767 3317 3823 3323
rect 87 3297 153 3303
rect 487 3293 493 3307
rect 1567 3293 1573 3307
rect 2147 3297 2193 3303
rect 3687 3293 3693 3307
rect 4440 3303 4453 3307
rect 4427 3297 4453 3303
rect 4440 3293 4453 3297
rect 4560 3303 4573 3307
rect 4547 3297 4573 3303
rect 4560 3293 4573 3297
rect 5167 3297 5213 3303
rect 1173 3283 1187 3293
rect 1173 3280 1213 3283
rect 1177 3277 1213 3280
rect 1467 3273 1473 3287
rect 1500 3283 1513 3287
rect 1487 3277 1513 3283
rect 1500 3273 1513 3277
rect 2027 3273 2033 3287
rect 2247 3273 2253 3287
rect 133 3263 147 3273
rect 2860 3283 2873 3287
rect 2687 3277 2733 3283
rect 2847 3277 2873 3283
rect 2860 3273 2873 3277
rect 2947 3277 2993 3283
rect 3080 3283 3093 3287
rect 3067 3277 3093 3283
rect 3080 3273 3093 3277
rect 4007 3277 4053 3283
rect 4987 3283 5000 3287
rect 4987 3277 5013 3283
rect 5217 3277 5273 3283
rect 4987 3273 5000 3277
rect 133 3260 193 3263
rect 137 3257 193 3260
rect 367 3257 413 3263
rect 877 3266 893 3267
rect 887 3253 893 3266
rect 947 3257 993 3263
rect 1687 3263 1700 3267
rect 1687 3257 1713 3263
rect 1687 3253 1700 3257
rect 2087 3263 2100 3267
rect 2087 3257 2113 3263
rect 2087 3253 2100 3257
rect 3900 3263 3913 3267
rect 3887 3257 3913 3263
rect 3900 3253 3913 3257
rect 4120 3263 4133 3267
rect 4107 3257 4133 3263
rect 4120 3253 4133 3257
rect 4287 3263 4300 3267
rect 4287 3257 4313 3263
rect 4287 3254 4300 3257
rect 4280 3253 4300 3254
rect 4887 3263 4900 3267
rect 4887 3257 4913 3263
rect 4887 3253 4900 3257
rect 1287 3237 1333 3243
rect 4227 3237 4273 3243
rect 227 3223 240 3227
rect 227 3217 253 3223
rect 227 3213 240 3217
rect 2037 3220 2043 3233
rect 4607 3243 4620 3247
rect 4607 3237 4633 3243
rect 4607 3233 4620 3237
rect 2033 3207 2047 3220
rect 4687 3213 4693 3227
rect 5217 3226 5223 3277
rect 5447 3257 5493 3263
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 47 3013 53 3027
rect 547 3023 560 3027
rect 547 3017 573 3023
rect 547 3013 560 3017
rect 1247 3017 1293 3023
rect 2120 3023 2133 3027
rect 2107 3017 2133 3023
rect 2120 3013 2133 3017
rect 947 2997 993 3003
rect 1687 2993 1693 3007
rect 4347 2993 4353 3007
rect 4820 3003 4833 3007
rect 4807 2997 4833 3003
rect 4820 2993 4833 2997
rect 5167 2997 5233 3003
rect 3033 2987 3047 2993
rect 1287 2983 1300 2987
rect 1287 2977 1313 2983
rect 1287 2973 1300 2977
rect 1367 2977 1433 2983
rect 2727 2973 2733 2987
rect 3247 2983 3260 2987
rect 3247 2977 3273 2983
rect 3247 2973 3260 2977
rect 4107 2973 4113 2987
rect 4417 2986 4433 2987
rect 4427 2973 4433 2986
rect 4580 2983 4593 2987
rect 4567 2977 4593 2983
rect 4580 2973 4593 2977
rect 4720 2983 4733 2987
rect 4707 2977 4733 2983
rect 4720 2973 4733 2977
rect 5453 2967 5467 2973
rect 227 2953 233 2967
rect 307 2963 320 2967
rect 307 2957 333 2963
rect 307 2953 320 2957
rect 647 2957 733 2963
rect 1067 2963 1080 2967
rect 1067 2957 1093 2963
rect 1067 2953 1080 2957
rect 1640 2963 1653 2967
rect 1627 2957 1653 2963
rect 1640 2953 1653 2957
rect 1807 2953 1813 2967
rect 1827 2953 1832 2967
rect 1867 2957 1913 2963
rect 1967 2957 2033 2963
rect 5067 2963 5080 2967
rect 5067 2957 5093 2963
rect 5067 2953 5080 2957
rect 5507 2953 5513 2967
rect 4887 2933 4893 2947
rect 4967 2937 5013 2943
rect 5543 2878 5603 3382
rect 5510 2862 5603 2878
rect 1893 2803 1907 2813
rect 1893 2800 1933 2803
rect 1897 2797 1933 2800
rect 147 2773 153 2787
rect 407 2786 420 2787
rect 407 2773 413 2786
rect 507 2773 513 2787
rect 747 2783 760 2787
rect 747 2777 773 2783
rect 747 2773 760 2777
rect 987 2783 1000 2787
rect 987 2777 1013 2783
rect 987 2773 1000 2777
rect 1287 2777 1353 2783
rect 1687 2777 1753 2783
rect 1807 2773 1813 2787
rect 2133 2783 2147 2793
rect 3687 2797 3753 2803
rect 3920 2803 3933 2807
rect 3907 2797 3933 2803
rect 3920 2793 3933 2797
rect 2433 2787 2447 2793
rect 2067 2780 2147 2783
rect 2067 2777 2143 2780
rect 3047 2777 3093 2783
rect 3853 2783 3867 2793
rect 3827 2780 3867 2783
rect 3827 2777 3863 2780
rect 4687 2777 4753 2783
rect 5347 2773 5353 2787
rect 1207 2753 1213 2767
rect 2127 2757 2173 2763
rect 2507 2753 2513 2767
rect 2747 2757 2823 2763
rect 3007 2757 3053 2763
rect 100 2743 113 2747
rect 87 2737 113 2743
rect 100 2733 113 2737
rect 873 2743 887 2753
rect 873 2740 913 2743
rect 877 2737 913 2740
rect 473 2727 487 2733
rect 1587 2740 1623 2743
rect 1587 2737 1627 2740
rect 1613 2727 1627 2737
rect 2007 2743 2020 2747
rect 2007 2737 2033 2743
rect 2007 2733 2020 2737
rect 2817 2743 2823 2757
rect 5500 2763 5513 2767
rect 5487 2757 5513 2763
rect 5500 2753 5513 2757
rect 3373 2747 3387 2753
rect 2817 2737 2853 2743
rect 3647 2733 3653 2747
rect 3807 2733 3813 2747
rect 3867 2733 3873 2747
rect 4047 2733 4053 2747
rect 4347 2737 4393 2743
rect 4693 2743 4707 2753
rect 4693 2740 4733 2743
rect 4697 2737 4733 2740
rect 4817 2740 4873 2743
rect 4813 2737 4873 2740
rect 4813 2727 4827 2737
rect 5367 2733 5373 2747
rect 647 2713 653 2727
rect 2207 2713 2213 2727
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 5467 2517 5493 2523
rect 187 2503 200 2507
rect 187 2497 213 2503
rect 187 2493 200 2497
rect 667 2493 673 2507
rect 887 2493 893 2507
rect 1127 2503 1140 2507
rect 1127 2497 1153 2503
rect 1127 2493 1140 2497
rect 427 2473 433 2487
rect 840 2483 853 2487
rect 827 2477 853 2483
rect 840 2473 853 2477
rect 2967 2473 2973 2487
rect 3667 2473 3673 2487
rect 4287 2483 4300 2487
rect 4287 2477 4313 2483
rect 4287 2473 4300 2477
rect 5267 2473 5273 2487
rect 1687 2453 1693 2467
rect 1873 2463 1887 2473
rect 3493 2467 3507 2473
rect 4433 2467 4447 2473
rect 4993 2467 5007 2473
rect 1847 2460 1887 2463
rect 1847 2457 1883 2460
rect 2547 2453 2553 2467
rect 4887 2453 4893 2467
rect 27 2437 73 2443
rect 527 2433 533 2447
rect 1067 2433 1073 2447
rect 1567 2443 1580 2447
rect 1567 2437 1593 2443
rect 1567 2433 1580 2437
rect 2227 2437 2273 2443
rect 2827 2443 2840 2447
rect 2827 2437 2853 2443
rect 2827 2433 2840 2437
rect 3147 2433 3153 2447
rect 307 2417 353 2423
rect 1947 2413 1953 2427
rect 2967 2423 2980 2427
rect 2967 2417 2993 2423
rect 2967 2413 2980 2417
rect 3687 2413 3693 2427
rect 4360 2423 4373 2427
rect 4347 2417 4373 2423
rect 4360 2413 4373 2417
rect 5260 2423 5273 2427
rect 4467 2417 4503 2423
rect 5247 2417 5273 2423
rect 4497 2407 4503 2417
rect 5260 2413 5273 2417
rect 4497 2397 4513 2407
rect 4500 2393 4513 2397
rect 5543 2358 5603 2862
rect 5510 2342 5603 2358
rect 1767 2273 1773 2287
rect 3127 2283 3140 2287
rect 3127 2277 3153 2283
rect 3127 2273 3140 2277
rect 3207 2277 3293 2283
rect 3987 2277 4033 2283
rect 5247 2283 5260 2287
rect 5247 2277 5273 2283
rect 5247 2273 5260 2277
rect 5387 2273 5393 2287
rect 267 2253 273 2267
rect 567 2257 633 2263
rect 1607 2253 1613 2267
rect 2293 2263 2307 2273
rect 2293 2260 2333 2263
rect 2297 2257 2333 2260
rect 2987 2263 3000 2267
rect 2987 2257 3013 2263
rect 2987 2253 3000 2257
rect 4380 2263 4393 2267
rect 4367 2257 4393 2263
rect 4380 2253 4393 2257
rect 1193 2247 1207 2253
rect 47 2243 60 2247
rect 47 2237 73 2243
rect 47 2233 60 2237
rect 540 2246 560 2247
rect 540 2243 553 2246
rect 527 2237 553 2243
rect 540 2233 553 2237
rect 687 2237 733 2243
rect 907 2243 920 2247
rect 907 2237 933 2243
rect 907 2233 920 2237
rect 2427 2233 2433 2247
rect 3427 2237 3473 2243
rect 4127 2234 4133 2247
rect 4260 2243 4273 2247
rect 4247 2237 4273 2243
rect 4127 2233 4143 2234
rect 4260 2233 4273 2237
rect 187 2217 253 2223
rect 1813 2223 1827 2233
rect 2033 2227 2047 2233
rect 3313 2227 3327 2233
rect 4593 2227 4607 2233
rect 1787 2220 1827 2223
rect 1787 2217 1823 2220
rect 3927 2223 3940 2227
rect 3927 2217 3953 2223
rect 3927 2213 3940 2217
rect 5367 2213 5373 2227
rect 497 2180 503 2193
rect 493 2167 507 2180
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 3893 1987 3907 1993
rect 5393 1983 5407 1993
rect 5367 1980 5407 1983
rect 5367 1977 5403 1980
rect 2653 1967 2667 1973
rect 827 1953 833 1967
rect 887 1953 893 1967
rect 1267 1953 1273 1967
rect 493 1947 507 1953
rect 1847 1953 1853 1967
rect 2080 1963 2093 1967
rect 2067 1957 2093 1963
rect 2080 1953 2093 1957
rect 5067 1963 5080 1967
rect 5067 1957 5093 1963
rect 5067 1953 5080 1957
rect 5187 1957 5233 1963
rect 2313 1947 2327 1953
rect 287 1933 293 1947
rect 1747 1937 1793 1943
rect 1987 1943 2000 1947
rect 1987 1937 2013 1943
rect 1987 1933 2000 1937
rect 2867 1933 2873 1947
rect 3307 1943 3320 1947
rect 3307 1937 3333 1943
rect 3307 1933 3320 1937
rect 3887 1943 3900 1947
rect 3887 1937 3913 1943
rect 3887 1933 3900 1937
rect 5360 1943 5373 1947
rect 5347 1937 5373 1943
rect 5360 1934 5373 1937
rect 5360 1933 5380 1934
rect 727 1917 793 1923
rect 2660 1923 2672 1927
rect 2647 1917 2672 1923
rect 2660 1913 2672 1917
rect 2707 1917 2773 1923
rect 3007 1914 3013 1927
rect 3007 1913 3023 1914
rect 3767 1923 3780 1927
rect 3767 1917 3793 1923
rect 3767 1913 3780 1917
rect 4287 1917 4352 1923
rect 4387 1913 4393 1927
rect 4487 1913 4493 1927
rect 4907 1917 4993 1923
rect 5187 1923 5200 1927
rect 5187 1917 5213 1923
rect 5187 1913 5200 1917
rect 1940 1903 1953 1907
rect 1727 1897 1813 1903
rect 1927 1897 1953 1903
rect 1940 1893 1953 1897
rect 2047 1893 2053 1907
rect 3500 1903 3513 1907
rect 3487 1897 3513 1903
rect 3500 1893 3513 1897
rect 4027 1897 4093 1903
rect 4160 1903 4173 1907
rect 4147 1897 4173 1903
rect 4160 1893 4173 1897
rect 4760 1906 4780 1907
rect 4760 1903 4773 1906
rect 4577 1900 4653 1903
rect 4573 1897 4653 1900
rect 4747 1897 4773 1903
rect 4573 1887 4587 1897
rect 4760 1893 4773 1897
rect 5127 1893 5133 1907
rect 5543 1838 5603 2342
rect 5510 1822 5603 1838
rect 1467 1757 1553 1763
rect 1687 1757 1733 1763
rect 1927 1757 1973 1763
rect 2913 1760 2927 1773
rect 257 1737 292 1743
rect 93 1707 107 1713
rect 257 1686 263 1737
rect 327 1733 333 1747
rect 1620 1743 1633 1747
rect 1607 1737 1633 1743
rect 1620 1733 1633 1737
rect 2140 1743 2153 1747
rect 2127 1737 2153 1743
rect 2140 1733 2153 1737
rect 2917 1747 2923 1760
rect 3773 1763 3787 1773
rect 3747 1760 3787 1763
rect 3747 1757 3783 1760
rect 4387 1757 4433 1763
rect 5087 1763 5100 1767
rect 5087 1757 5113 1763
rect 5087 1753 5100 1757
rect 2787 1743 2800 1747
rect 2787 1737 2813 1743
rect 2787 1733 2800 1737
rect 3347 1737 3393 1743
rect 3907 1737 3973 1743
rect 4053 1743 4067 1753
rect 4053 1740 4093 1743
rect 4057 1737 4093 1740
rect 4540 1743 4553 1747
rect 4527 1737 4553 1743
rect 4540 1733 4553 1737
rect 5187 1743 5200 1747
rect 5187 1737 5213 1743
rect 5187 1733 5200 1737
rect 2267 1717 2313 1723
rect 4607 1717 4653 1723
rect 4807 1717 4853 1723
rect 4907 1717 4973 1723
rect 1013 1707 1027 1713
rect 1427 1693 1433 1707
rect 1527 1697 1573 1703
rect 1627 1703 1640 1707
rect 1627 1697 1653 1703
rect 1627 1693 1640 1697
rect 2177 1700 2213 1703
rect 2173 1697 2213 1700
rect 2173 1687 2187 1697
rect 2627 1697 2673 1703
rect 2927 1693 2933 1707
rect 3027 1693 3033 1707
rect 3087 1706 3103 1707
rect 3087 1693 3093 1706
rect 3327 1697 3413 1703
rect 4007 1700 4043 1703
rect 4007 1697 4047 1700
rect 4033 1687 4047 1697
rect 4207 1697 4253 1703
rect 1387 1657 1413 1663
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 1800 1463 1813 1467
rect 1787 1457 1813 1463
rect 1800 1453 1813 1457
rect 2587 1443 2600 1447
rect 2587 1437 2613 1443
rect 2587 1433 2600 1437
rect 2987 1433 2993 1447
rect 3207 1433 3213 1447
rect 3347 1443 3360 1447
rect 3347 1437 3373 1443
rect 3347 1433 3360 1437
rect 3587 1437 3633 1443
rect 3827 1443 3840 1447
rect 3827 1437 3853 1443
rect 3827 1433 3840 1437
rect 953 1427 967 1433
rect 1113 1427 1127 1433
rect 5287 1437 5333 1443
rect 5387 1437 5433 1443
rect 367 1413 373 1427
rect 907 1413 913 1427
rect 1327 1417 1393 1423
rect 2367 1423 2380 1427
rect 2367 1417 2393 1423
rect 2367 1413 2380 1417
rect 3267 1413 3273 1427
rect 4107 1413 4113 1427
rect 4807 1413 4813 1427
rect 5197 1426 5213 1427
rect 5207 1413 5213 1426
rect 1267 1397 1353 1403
rect 1647 1397 1713 1403
rect 1927 1406 1943 1407
rect 1927 1393 1933 1406
rect 2047 1393 2053 1407
rect 2547 1397 2633 1403
rect 4387 1393 4393 1407
rect 4333 1387 4347 1393
rect 267 1377 333 1383
rect 487 1377 533 1383
rect 587 1377 633 1383
rect 927 1373 933 1387
rect 1027 1377 1093 1383
rect 3407 1377 3453 1383
rect 3707 1383 3720 1387
rect 3707 1377 3733 1383
rect 3707 1373 3720 1377
rect 4587 1377 4632 1383
rect 4667 1373 4673 1387
rect 5413 1386 5427 1393
rect 5543 1318 5603 1822
rect 5510 1302 5603 1318
rect 2067 1243 2080 1247
rect 2067 1237 2093 1243
rect 2687 1237 2733 1243
rect 2067 1233 2080 1237
rect 4687 1237 4733 1243
rect 4807 1237 4853 1243
rect 1847 1217 1923 1223
rect 500 1206 520 1207
rect 233 1187 247 1193
rect 507 1203 520 1206
rect 573 1203 587 1213
rect 507 1197 533 1203
rect 573 1200 603 1203
rect 577 1197 603 1200
rect 507 1193 520 1197
rect 597 1187 603 1197
rect 1547 1203 1560 1207
rect 1547 1197 1573 1203
rect 1547 1193 1560 1197
rect 1293 1187 1307 1193
rect 597 1177 613 1187
rect 600 1173 613 1177
rect 1917 1186 1923 1217
rect 1947 1213 1953 1227
rect 2240 1223 2253 1227
rect 2227 1217 2253 1223
rect 2240 1214 2253 1217
rect 2240 1213 2260 1214
rect 2727 1217 2773 1223
rect 3507 1213 3513 1227
rect 3827 1217 3893 1223
rect 4507 1217 4553 1223
rect 4620 1223 4633 1227
rect 4607 1217 4633 1223
rect 4620 1213 4633 1217
rect 5127 1217 5193 1223
rect 2627 1203 2640 1207
rect 2877 1206 2893 1207
rect 2627 1197 2653 1203
rect 2627 1193 2640 1197
rect 2887 1193 2893 1206
rect 3287 1193 3293 1207
rect 3407 1197 3453 1203
rect 4827 1193 4833 1207
rect 5177 1197 5233 1203
rect 2273 1183 2287 1192
rect 2273 1180 2333 1183
rect 2277 1177 2333 1180
rect 4467 1173 4473 1187
rect 4940 1183 4953 1187
rect 4927 1177 4953 1183
rect 4940 1173 4953 1177
rect 5020 1183 5033 1187
rect 5007 1177 5033 1183
rect 5020 1173 5033 1177
rect 5177 1183 5183 1197
rect 5147 1177 5183 1183
rect 3427 1153 3433 1167
rect 5253 1147 5267 1153
rect 2267 1137 2313 1143
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 2633 947 2647 953
rect 4607 933 4613 947
rect 5307 943 5320 947
rect 5307 933 5323 943
rect 107 913 113 927
rect 360 923 373 927
rect 347 917 373 923
rect 360 913 373 917
rect 1007 913 1013 927
rect 1507 917 1553 923
rect 2900 923 2913 927
rect 2897 913 2913 923
rect 3427 913 3433 927
rect 4167 923 4180 927
rect 4167 917 4193 923
rect 4167 913 4180 917
rect 5317 923 5323 933
rect 5317 917 5373 923
rect 267 903 280 907
rect 267 897 293 903
rect 267 893 280 897
rect 827 897 873 903
rect 1627 893 1633 907
rect 1747 897 1813 903
rect 2247 897 2313 903
rect 2367 897 2413 903
rect 2567 897 2613 903
rect 2067 877 2113 883
rect 2507 877 2573 883
rect 267 857 313 863
rect 607 863 620 867
rect 607 857 633 863
rect 607 853 620 857
rect 907 857 973 863
rect 2897 866 2903 913
rect 4027 903 4040 907
rect 4027 897 4053 903
rect 4027 893 4040 897
rect 4647 897 4713 903
rect 5427 903 5440 907
rect 5427 897 5453 903
rect 5427 893 5440 897
rect 3147 873 3153 887
rect 3907 873 3913 887
rect 3533 863 3547 873
rect 4173 867 4187 873
rect 4727 877 4773 883
rect 4887 873 4893 887
rect 5120 886 5140 887
rect 5127 883 5140 886
rect 5127 877 5153 883
rect 5127 873 5140 877
rect 3533 860 3573 863
rect 3537 857 3573 860
rect 5247 853 5253 867
rect 5267 857 5323 863
rect 5317 843 5323 857
rect 5317 837 5353 843
rect 5543 798 5603 1302
rect 5510 782 5603 798
rect 107 717 153 723
rect 207 717 253 723
rect 2047 717 2093 723
rect 3167 713 3173 727
rect 1193 707 1207 713
rect 287 693 293 707
rect 1507 693 1513 707
rect 1620 703 1633 707
rect 1607 697 1633 703
rect 1620 693 1633 697
rect 1747 697 1793 703
rect 2187 697 2233 703
rect 3787 703 3800 707
rect 3787 700 3803 703
rect 3787 693 3807 700
rect 3827 693 3833 707
rect 4027 697 4093 703
rect 4407 693 4413 707
rect 4827 697 4873 703
rect 500 683 513 687
rect 487 677 513 683
rect 500 673 513 677
rect 567 677 613 683
rect 680 683 693 687
rect 667 677 693 683
rect 680 673 693 677
rect 767 677 833 683
rect 1147 674 1153 687
rect 1147 673 1163 674
rect 1667 683 1680 687
rect 1667 677 1693 683
rect 1667 673 1680 677
rect 3033 687 3047 693
rect 3793 687 3807 693
rect 2767 674 2773 687
rect 2757 673 2773 674
rect 3127 673 3133 687
rect 3747 673 3753 687
rect 4087 677 4133 683
rect 113 667 127 673
rect 1313 667 1327 673
rect 5213 667 5227 673
rect 1040 663 1053 667
rect 1027 657 1053 663
rect 1040 653 1053 657
rect 3327 663 3340 667
rect 3327 657 3353 663
rect 3327 653 3340 657
rect 3567 653 3573 667
rect 4937 657 4973 663
rect 3407 633 3413 647
rect 3687 643 3700 647
rect 3687 637 3713 643
rect 3687 633 3700 637
rect 4080 646 4100 647
rect 1677 603 1683 633
rect 4087 643 4100 646
rect 4087 637 4113 643
rect 4087 633 4100 637
rect 3347 613 3353 627
rect 1627 597 1683 603
rect -63 522 30 538
rect -63 18 -3 522
rect 887 423 900 427
rect 887 417 913 423
rect 887 413 900 417
rect 1387 413 1393 427
rect 1727 413 1733 427
rect 1947 423 1960 427
rect 1947 417 1973 423
rect 1947 413 1960 417
rect 2347 403 2360 407
rect 2347 397 2373 403
rect 2347 393 2360 397
rect 393 387 407 393
rect 4667 393 4673 407
rect 5080 403 5093 407
rect 5067 397 5093 403
rect 5080 393 5093 397
rect 927 373 933 387
rect 1367 377 1413 383
rect 1747 373 1753 387
rect 1967 383 1980 387
rect 1967 377 1993 383
rect 1967 373 1980 377
rect 4887 373 4893 387
rect 1080 363 1093 367
rect 1067 357 1093 363
rect 1080 353 1093 357
rect 1807 357 1873 363
rect 2813 363 2827 373
rect 2813 360 2853 363
rect 2817 357 2853 360
rect 3267 357 3353 363
rect 4147 363 4160 367
rect 4147 357 4173 363
rect 4147 353 4160 357
rect 4627 363 4640 367
rect 4627 357 4653 363
rect 4627 353 4640 357
rect 4747 357 4793 363
rect 4947 297 4973 303
rect 5543 278 5603 782
rect 5510 262 5603 278
rect 187 197 253 203
rect 387 193 393 207
rect 2107 203 2120 207
rect 2107 197 2133 203
rect 2107 193 2120 197
rect 3607 194 3613 207
rect 3597 193 3613 194
rect 4807 203 4820 207
rect 4807 197 4833 203
rect 4807 193 4820 197
rect 507 177 553 183
rect 840 183 853 187
rect 827 177 853 183
rect 840 173 853 177
rect 1400 183 1413 187
rect 1387 177 1413 183
rect 1400 173 1413 177
rect 2427 183 2440 187
rect 2427 177 2453 183
rect 2427 173 2440 177
rect 3687 177 3753 183
rect 4647 177 4693 183
rect 5320 183 5333 187
rect 5307 177 5333 183
rect 5320 173 5333 177
rect 5253 167 5267 173
rect 127 163 140 167
rect 127 157 153 163
rect 127 153 140 157
rect 347 153 353 167
rect 1180 163 1193 167
rect 1167 157 1193 163
rect 1180 153 1193 157
rect 1247 153 1253 167
rect 2900 163 2913 167
rect 2887 157 2913 163
rect 2900 153 2913 157
rect 3140 163 3153 167
rect 3127 157 3153 163
rect 3140 153 3153 157
rect 3307 153 3313 167
rect 3407 153 3413 167
rect 3847 153 3853 167
rect 4167 157 4213 163
rect 4327 163 4340 167
rect 4327 157 4353 163
rect 4327 153 4340 157
rect 5407 157 5513 163
rect 233 143 247 153
rect 5133 147 5147 153
rect 207 140 247 143
rect 207 137 243 140
rect 407 133 413 147
rect 627 137 673 143
rect 740 143 753 147
rect 727 137 753 143
rect 740 133 753 137
rect 940 143 953 147
rect 927 137 953 143
rect 940 133 953 137
rect 4867 133 4873 147
rect 4967 133 4973 147
rect 1060 123 1073 127
rect 1047 117 1073 123
rect 1060 113 1073 117
rect 4187 113 4193 127
rect -63 2 30 18
rect 5543 2 5603 262
<< m2contact >>
rect 633 5393 647 5407
rect 4813 5393 4827 5407
rect 33 5373 47 5387
rect 93 5373 107 5387
rect 333 5373 347 5387
rect 393 5373 407 5387
rect 513 5373 527 5387
rect 873 5373 887 5387
rect 913 5373 927 5387
rect 1113 5373 1127 5387
rect 1233 5373 1247 5387
rect 1513 5373 1527 5387
rect 1613 5373 1627 5387
rect 1773 5373 1787 5387
rect 1873 5373 1887 5387
rect 1913 5373 1927 5387
rect 2053 5373 2067 5387
rect 2093 5373 2107 5387
rect 2153 5373 2167 5387
rect 2227 5373 2241 5387
rect 2273 5373 2287 5387
rect 2333 5373 2347 5387
rect 2653 5373 2667 5387
rect 2733 5373 2747 5387
rect 2893 5373 2907 5387
rect 2993 5373 3007 5387
rect 3033 5373 3047 5387
rect 3093 5373 3107 5387
rect 3153 5373 3167 5387
rect 3193 5373 3207 5387
rect 3233 5373 3247 5387
rect 3353 5373 3367 5387
rect 3413 5373 3427 5387
rect 3453 5373 3467 5387
rect 3693 5373 3707 5387
rect 3773 5373 3787 5387
rect 3813 5373 3827 5387
rect 3953 5373 3967 5387
rect 4113 5373 4127 5387
rect 4153 5373 4167 5387
rect 4293 5373 4307 5387
rect 4413 5373 4427 5387
rect 4593 5373 4607 5387
rect 4693 5373 4707 5387
rect 4913 5373 4927 5387
rect 4993 5373 5007 5387
rect 5053 5373 5067 5387
rect 5193 5373 5207 5387
rect 5453 5373 5467 5387
rect 5493 5373 5507 5387
rect 193 5353 207 5367
rect 473 5353 487 5367
rect 607 5353 621 5367
rect 753 5353 767 5367
rect 1013 5353 1027 5367
rect 1153 5353 1167 5367
rect 1293 5353 1307 5367
rect 1393 5353 1407 5367
rect 1673 5353 1687 5367
rect 2433 5354 2447 5368
rect 2573 5353 2587 5367
rect 2853 5353 2867 5367
rect 3593 5353 3607 5367
rect 3993 5353 4007 5367
rect 4193 5353 4207 5367
rect 4533 5353 4547 5367
rect 4733 5353 4747 5367
rect 4833 5353 4847 5367
rect 5233 5353 5247 5367
rect 5353 5354 5367 5368
rect 73 5333 87 5347
rect 113 5333 127 5347
rect 213 5333 227 5347
rect 313 5333 327 5347
rect 353 5333 367 5347
rect 413 5333 427 5347
rect 693 5333 707 5347
rect 813 5333 827 5347
rect 893 5333 907 5347
rect 1253 5333 1267 5347
rect 1413 5333 1427 5347
rect 1493 5333 1507 5347
rect 1533 5333 1547 5347
rect 1653 5333 1667 5347
rect 1733 5333 1747 5347
rect 1833 5333 1847 5347
rect 1953 5333 1967 5347
rect 2033 5333 2047 5347
rect 2073 5333 2087 5347
rect 2153 5332 2167 5346
rect 2193 5333 2207 5347
rect 2313 5333 2327 5347
rect 2353 5333 2367 5347
rect 2413 5333 2427 5347
rect 2593 5333 2607 5347
rect 2713 5333 2727 5347
rect 2753 5333 2767 5347
rect 2873 5333 2887 5347
rect 2973 5333 2987 5347
rect 3013 5333 3027 5347
rect 3073 5333 3087 5347
rect 3113 5333 3127 5347
rect 3173 5333 3187 5347
rect 3293 5333 3307 5347
rect 3333 5333 3347 5347
rect 3433 5333 3447 5347
rect 3473 5333 3487 5347
rect 3573 5333 3587 5347
rect 3673 5333 3687 5347
rect 3713 5333 3727 5347
rect 3833 5333 3847 5347
rect 3873 5333 3887 5347
rect 4013 5333 4027 5347
rect 4093 5333 4107 5347
rect 4133 5333 4147 5347
rect 4573 5333 4587 5347
rect 4613 5333 4627 5347
rect 4773 5333 4787 5347
rect 4933 5333 4947 5347
rect 4973 5333 4987 5347
rect 5073 5333 5087 5347
rect 5113 5333 5127 5347
rect 5213 5333 5227 5347
rect 5373 5333 5387 5347
rect 5433 5333 5447 5347
rect 5473 5333 5487 5347
rect 173 5313 187 5327
rect 533 5313 547 5327
rect 573 5313 587 5327
rect 733 5313 747 5327
rect 773 5313 787 5327
rect 993 5313 1007 5327
rect 1033 5313 1047 5327
rect 1293 5312 1307 5326
rect 1753 5313 1767 5327
rect 2472 5313 2486 5327
rect 2493 5313 2507 5327
rect 2793 5313 2807 5327
rect 3633 5313 3647 5327
rect 3913 5313 3927 5327
rect 4233 5313 4247 5327
rect 4273 5313 4287 5327
rect 4313 5313 4327 5327
rect 4493 5313 4507 5327
rect 4533 5312 4547 5326
rect 4813 5313 4827 5327
rect 4853 5313 4867 5327
rect 5293 5313 5307 5327
rect 5333 5313 5347 5327
rect 233 5293 247 5307
rect 1433 5293 1447 5307
rect 1633 5293 1647 5307
rect 2393 5293 2407 5307
rect 2613 5293 2627 5307
rect 2893 5293 2907 5307
rect 3553 5293 3567 5307
rect 4033 5293 4047 5307
rect 5193 5293 5207 5307
rect 5393 5293 5407 5307
rect 493 5113 507 5127
rect 633 5113 647 5127
rect 1253 5113 1267 5127
rect 1733 5113 1747 5127
rect 2133 5113 2147 5127
rect 2253 5113 2267 5127
rect 2393 5113 2407 5127
rect 2733 5113 2747 5127
rect 3313 5113 3327 5127
rect 3493 5113 3507 5127
rect 5233 5112 5247 5126
rect 553 5093 567 5107
rect 693 5093 707 5107
rect 753 5093 767 5107
rect 793 5093 807 5107
rect 853 5093 867 5107
rect 893 5093 907 5107
rect 1373 5093 1387 5107
rect 1613 5093 1627 5107
rect 2033 5093 2047 5107
rect 2173 5093 2187 5107
rect 2293 5093 2307 5107
rect 2653 5093 2667 5107
rect 2993 5093 3007 5107
rect 3053 5093 3067 5107
rect 3233 5093 3247 5107
rect 3593 5093 3607 5107
rect 3653 5093 3667 5107
rect 3693 5093 3707 5107
rect 4193 5092 4207 5106
rect 4233 5093 4247 5107
rect 4293 5093 4307 5107
rect 4333 5093 4347 5107
rect 4493 5093 4507 5107
rect 4533 5093 4547 5107
rect 5173 5093 5187 5107
rect 53 5073 67 5087
rect 93 5073 107 5087
rect 193 5073 207 5087
rect 253 5073 267 5087
rect 293 5073 307 5087
rect 413 5073 427 5087
rect 453 5073 467 5087
rect 513 5073 527 5087
rect 653 5074 667 5088
rect 993 5072 1007 5086
rect 1033 5073 1047 5087
rect 1113 5073 1127 5087
rect 1173 5073 1187 5087
rect 1213 5073 1227 5087
rect 1273 5073 1287 5087
rect 1413 5073 1427 5087
rect 1453 5073 1467 5087
rect 1533 5074 1547 5088
rect 1573 5073 1587 5087
rect 1713 5073 1727 5087
rect 1833 5073 1847 5087
rect 1873 5073 1887 5087
rect 1933 5073 1947 5087
rect 1973 5073 1987 5087
rect 2113 5074 2127 5088
rect 2233 5074 2247 5088
rect 2373 5073 2387 5087
rect 2433 5073 2447 5087
rect 2573 5074 2587 5088
rect 2613 5073 2627 5087
rect 2713 5073 2727 5087
rect 2913 5073 2927 5087
rect 2953 5073 2967 5087
rect 3133 5073 3147 5087
rect 3173 5073 3187 5087
rect 3293 5073 3307 5087
rect 3393 5073 3407 5087
rect 3433 5073 3447 5087
rect 3513 5073 3527 5087
rect 3753 5073 3767 5087
rect 3793 5073 3807 5087
rect 3913 5073 3927 5087
rect 3953 5073 3967 5087
rect 3993 5073 4007 5087
rect 4047 5073 4061 5087
rect 4393 5073 4407 5087
rect 4633 5073 4647 5087
rect 4673 5073 4687 5087
rect 4753 5073 4767 5087
rect 4793 5073 4807 5087
rect 4873 5073 4887 5087
rect 4913 5073 4927 5087
rect 5033 5073 5047 5087
rect 5073 5073 5087 5087
rect 5213 5073 5227 5087
rect 5293 5073 5307 5087
rect 5333 5073 5347 5087
rect 5453 5073 5467 5087
rect 5493 5073 5507 5087
rect 533 5053 547 5067
rect 673 5054 687 5068
rect 713 5053 727 5067
rect 873 5053 887 5067
rect 1293 5053 1307 5067
rect 1693 5053 1707 5067
rect 2093 5053 2107 5067
rect 2213 5053 2227 5067
rect 2353 5053 2367 5067
rect 2693 5053 2707 5067
rect 3053 5052 3067 5066
rect 3273 5053 3287 5067
rect 3533 5053 3547 5067
rect 73 5033 87 5047
rect 113 5033 127 5047
rect 233 5033 247 5047
rect 292 5033 306 5047
rect 153 5013 167 5027
rect 433 5033 447 5047
rect 973 5033 987 5047
rect 1013 5033 1027 5047
rect 1053 5033 1067 5047
rect 1093 5033 1107 5047
rect 1153 5033 1167 5047
rect 1193 5033 1207 5047
rect 1333 5033 1347 5047
rect 1473 5033 1487 5047
rect 1533 5033 1547 5047
rect 1593 5033 1607 5047
rect 1773 5033 1787 5047
rect 1853 5033 1867 5047
rect 1953 5033 1967 5047
rect 2013 5033 2027 5047
rect 2253 5033 2267 5047
rect 2313 5033 2327 5047
rect 2473 5034 2487 5048
rect 4273 5053 4287 5067
rect 4353 5053 4367 5067
rect 4433 5053 4447 5067
rect 4553 5053 4567 5067
rect 5193 5052 5207 5066
rect 313 5013 327 5027
rect 2473 4993 2487 5007
rect 2593 5033 2607 5047
rect 2773 5033 2787 5047
rect 2893 5033 2907 5047
rect 2933 5033 2947 5047
rect 2973 5033 2987 5047
rect 3113 5033 3127 5047
rect 3233 5033 3247 5047
rect 3333 5033 3347 5047
rect 3413 5033 3427 5047
rect 3713 5033 3727 5047
rect 3773 5033 3787 5047
rect 3813 5033 3827 5047
rect 3853 5033 3867 5047
rect 3933 5033 3947 5047
rect 3973 5033 3987 5047
rect 4013 5033 4027 5047
rect 4073 5033 4087 5047
rect 4113 5033 4127 5047
rect 4653 5033 4667 5047
rect 4693 5033 4707 5047
rect 4733 5033 4747 5047
rect 4853 5033 4867 5047
rect 4893 5033 4907 5047
rect 4953 5033 4967 5047
rect 5013 5033 5027 5047
rect 5053 5033 5067 5047
rect 5313 5033 5327 5047
rect 5372 5033 5386 5047
rect 5393 5033 5407 5047
rect 5433 5033 5447 5047
rect 5473 5033 5487 5047
rect 4493 5013 4507 5027
rect 633 4873 647 4887
rect 953 4873 967 4887
rect 133 4854 147 4868
rect 313 4853 327 4867
rect 553 4853 567 4867
rect 733 4853 747 4867
rect 773 4853 787 4867
rect 813 4853 827 4867
rect 853 4853 867 4867
rect 93 4833 107 4847
rect 373 4833 387 4847
rect 513 4833 527 4847
rect 933 4833 947 4847
rect 113 4813 127 4827
rect 173 4813 187 4827
rect 233 4813 247 4827
rect 393 4813 407 4827
rect 533 4813 547 4827
rect 573 4813 587 4827
rect 653 4813 667 4827
rect 753 4813 767 4827
rect 793 4813 807 4827
rect 893 4813 907 4827
rect 2893 4873 2907 4887
rect 4393 4873 4407 4887
rect 1013 4853 1027 4867
rect 1093 4853 1107 4867
rect 1233 4853 1247 4867
rect 1273 4853 1287 4867
rect 1613 4853 1627 4867
rect 1673 4853 1687 4867
rect 1733 4853 1747 4867
rect 1852 4853 1866 4867
rect 1873 4853 1887 4867
rect 1933 4853 1947 4867
rect 2093 4853 2107 4867
rect 2633 4853 2647 4867
rect 2693 4853 2707 4867
rect 2793 4853 2807 4867
rect 3073 4853 3087 4867
rect 3113 4853 3127 4867
rect 3153 4853 3167 4867
rect 3173 4853 3187 4867
rect 3253 4853 3267 4867
rect 3353 4853 3367 4867
rect 3513 4853 3527 4867
rect 3613 4853 3627 4867
rect 3653 4853 3667 4867
rect 3693 4853 3707 4867
rect 3793 4853 3807 4867
rect 3973 4853 3987 4867
rect 4013 4853 4027 4867
rect 4053 4853 4067 4867
rect 4233 4854 4247 4868
rect 1053 4833 1067 4847
rect 1393 4834 1407 4848
rect 1513 4833 1527 4847
rect 2053 4833 2067 4847
rect 2233 4833 2247 4847
rect 2293 4833 2307 4847
rect 2453 4833 2467 4847
rect 2593 4834 2607 4848
rect 2833 4833 2847 4847
rect 2993 4833 3007 4847
rect 3213 4833 3227 4847
rect 3413 4833 3427 4847
rect 3453 4833 3467 4847
rect 3753 4833 3767 4847
rect 4133 4833 4147 4847
rect 4293 4833 4307 4847
rect 4573 4853 4587 4867
rect 4633 4853 4647 4867
rect 4773 4853 4787 4867
rect 4813 4853 4827 4867
rect 4953 4833 4967 4847
rect 5093 4833 5107 4847
rect 5233 4833 5247 4847
rect 5293 4833 5307 4847
rect 5453 4833 5467 4847
rect 973 4812 987 4826
rect 1133 4813 1147 4827
rect 1173 4813 1187 4827
rect 1253 4813 1267 4827
rect 1293 4813 1307 4827
rect 1413 4813 1427 4827
rect 1493 4813 1507 4827
rect 1593 4813 1607 4827
rect 1633 4813 1647 4827
rect 1753 4813 1767 4827
rect 1793 4813 1807 4827
rect 1913 4813 1927 4827
rect 1953 4813 1967 4827
rect 2033 4813 2047 4827
rect 2193 4813 2207 4827
rect 2473 4813 2487 4827
rect 2613 4813 2627 4827
rect 2713 4813 2727 4827
rect 2753 4813 2767 4827
rect 2953 4813 2967 4827
rect 3093 4813 3107 4827
rect 3133 4813 3147 4827
rect 3253 4813 3267 4827
rect 3373 4813 3387 4827
rect 3493 4813 3507 4827
rect 3633 4813 3647 4827
rect 3673 4813 3687 4827
rect 3793 4813 3807 4827
rect 4033 4813 4047 4827
rect 4073 4813 4087 4827
rect 4173 4813 4187 4827
rect 4333 4813 4347 4827
rect 4513 4813 4527 4827
rect 4553 4813 4567 4827
rect 4713 4813 4727 4827
rect 4753 4813 4767 4827
rect 4833 4813 4847 4827
rect 4973 4813 4987 4827
rect 5073 4813 5087 4827
rect 5213 4813 5227 4827
rect 5473 4812 5487 4826
rect 73 4793 87 4807
rect 353 4793 367 4807
rect 453 4793 467 4807
rect 1353 4793 1367 4807
rect 1533 4793 1547 4807
rect 2113 4793 2127 4807
rect 2293 4793 2307 4807
rect 2333 4793 2347 4807
rect 2393 4793 2407 4807
rect 2533 4793 2547 4807
rect 2833 4793 2847 4807
rect 2873 4793 2887 4807
rect 3893 4793 3907 4807
rect 3933 4793 3947 4807
rect 4393 4793 4407 4807
rect 4433 4793 4447 4807
rect 4933 4793 4947 4807
rect 5113 4793 5127 4807
rect 5273 4793 5287 4807
rect 5333 4793 5347 4807
rect 5373 4793 5387 4807
rect 5413 4793 5427 4807
rect 133 4773 147 4787
rect 413 4773 427 4787
rect 553 4773 567 4787
rect 1473 4773 1487 4787
rect 2013 4773 2027 4787
rect 2493 4773 2507 4787
rect 2633 4773 2647 4787
rect 4993 4773 5007 4787
rect 5053 4773 5067 4787
rect 5193 4773 5207 4787
rect 5493 4773 5507 4787
rect 1813 4713 1827 4727
rect 1853 4713 1867 4727
rect 2713 4613 2727 4627
rect 2753 4613 2767 4627
rect 153 4593 167 4607
rect 1093 4593 1107 4607
rect 1233 4593 1247 4607
rect 1613 4593 1627 4607
rect 2013 4593 2027 4607
rect 2313 4593 2327 4607
rect 2573 4593 2587 4607
rect 2833 4593 2847 4607
rect 73 4573 87 4587
rect 113 4573 127 4587
rect 213 4573 227 4587
rect 673 4573 687 4587
rect 893 4573 907 4587
rect 933 4573 947 4587
rect 1013 4573 1027 4587
rect 1133 4573 1147 4587
rect 173 4553 187 4567
rect 253 4553 267 4567
rect 313 4553 327 4567
rect 433 4553 447 4567
rect 473 4553 487 4567
rect 593 4553 607 4567
rect 633 4553 647 4567
rect 1533 4572 1547 4586
rect 2073 4573 2087 4587
rect 2153 4573 2167 4587
rect 2193 4573 2207 4587
rect 2253 4573 2267 4587
rect 2513 4573 2527 4587
rect 813 4553 827 4567
rect 1073 4554 1087 4568
rect 1213 4553 1227 4567
rect 1273 4553 1287 4567
rect 1313 4553 1327 4567
rect 1453 4553 1467 4567
rect 1493 4553 1507 4567
rect 1593 4553 1607 4567
rect 1713 4553 1727 4567
rect 1773 4553 1787 4567
rect 1813 4553 1827 4567
rect 1913 4553 1927 4567
rect 2033 4553 2047 4567
rect 2393 4553 2407 4567
rect 2433 4553 2447 4567
rect 2553 4554 2567 4568
rect 2653 4553 2667 4567
rect 2693 4553 2707 4567
rect 2793 4553 2807 4567
rect 2833 4553 2847 4567
rect 93 4533 107 4547
rect 193 4532 207 4546
rect 853 4533 867 4547
rect 913 4533 927 4547
rect 1053 4533 1067 4547
rect 1193 4533 1207 4547
rect 1573 4533 1587 4547
rect 1953 4533 1967 4547
rect 2053 4533 2067 4547
rect 2233 4534 2247 4548
rect 2313 4533 2327 4547
rect 2533 4533 2547 4547
rect 3013 4593 3027 4607
rect 4353 4593 4367 4607
rect 4393 4593 4407 4607
rect 4533 4593 4547 4607
rect 4673 4593 4687 4607
rect 4793 4593 4807 4607
rect 2913 4573 2927 4587
rect 3053 4573 3067 4587
rect 3093 4573 3107 4587
rect 3733 4573 3747 4587
rect 3773 4573 3787 4587
rect 4293 4573 4307 4587
rect 4473 4573 4487 4587
rect 4613 4573 4627 4587
rect 4753 4573 4767 4587
rect 4913 4573 4927 4587
rect 5353 4573 5367 4587
rect 5393 4573 5407 4587
rect 2973 4554 2987 4568
rect 3233 4554 3247 4568
rect 3453 4553 3467 4567
rect 3493 4553 3507 4567
rect 3613 4554 3627 4568
rect 3653 4553 3667 4567
rect 3913 4553 3927 4567
rect 3953 4553 3967 4567
rect 3993 4553 4007 4567
rect 4033 4553 4047 4567
rect 4073 4553 4087 4567
rect 4173 4553 4187 4567
rect 4213 4554 4227 4568
rect 4333 4553 4347 4567
rect 4413 4553 4427 4567
rect 4553 4554 4567 4568
rect 4693 4554 4707 4568
rect 4813 4553 4827 4567
rect 4953 4553 4967 4567
rect 4993 4553 5007 4567
rect 5133 4553 5147 4567
rect 5213 4553 5227 4567
rect 5253 4553 5267 4567
rect 5433 4553 5447 4567
rect 5473 4553 5487 4567
rect 2913 4533 2927 4547
rect 2953 4533 2967 4547
rect 3133 4533 3147 4547
rect 3373 4533 3387 4547
rect 3553 4533 3567 4547
rect 3813 4533 3827 4547
rect 4313 4533 4327 4547
rect 4433 4533 4447 4547
rect 4573 4533 4587 4547
rect 4713 4533 4727 4547
rect 4833 4533 4847 4547
rect 5093 4533 5107 4547
rect 5293 4533 5307 4547
rect 233 4513 247 4527
rect 352 4513 366 4527
rect 373 4513 387 4527
rect 512 4513 526 4527
rect 533 4513 547 4527
rect 613 4513 627 4527
rect 693 4513 707 4527
rect 793 4513 807 4527
rect 1293 4513 1307 4527
rect 1353 4513 1367 4527
rect 1433 4513 1447 4527
rect 1473 4513 1487 4527
rect 1673 4513 1687 4527
rect 1753 4513 1767 4527
rect 1793 4513 1807 4527
rect 1833 4513 1847 4527
rect 2353 4513 2367 4527
rect 2413 4513 2427 4527
rect 2633 4513 2647 4527
rect 2733 4513 2747 4527
rect 2773 4513 2787 4527
rect 2873 4513 2887 4527
rect 3033 4513 3047 4527
rect 3213 4513 3227 4527
rect 3253 4513 3267 4527
rect 3313 4513 3327 4527
rect 3413 4513 3427 4527
rect 3533 4513 3547 4527
rect 3593 4513 3607 4527
rect 3633 4513 3647 4527
rect 3673 4513 3687 4527
rect 3873 4513 3887 4527
rect 3933 4513 3947 4527
rect 4073 4513 4087 4527
rect 4113 4513 4127 4527
rect 4153 4513 4167 4527
rect 4213 4513 4227 4527
rect 4933 4513 4947 4527
rect 4973 4513 4987 4527
rect 5013 4513 5027 4527
rect 5193 4513 5207 4527
rect 5233 4513 5247 4527
rect 5453 4513 5467 4527
rect 5493 4513 5507 4527
rect 1873 4493 1887 4507
rect 3553 4493 3567 4507
rect 3793 4494 3807 4508
rect 3833 4493 3847 4507
rect 5033 4473 5047 4487
rect 953 4453 967 4467
rect 1013 4453 1027 4467
rect 913 4353 927 4367
rect 3433 4353 3447 4367
rect 3653 4353 3667 4367
rect 5173 4353 5187 4367
rect 433 4333 447 4347
rect 473 4333 487 4347
rect 633 4333 647 4347
rect 713 4333 727 4347
rect 813 4333 827 4347
rect 853 4332 867 4346
rect 1233 4333 1247 4347
rect 1353 4332 1367 4346
rect 1433 4333 1447 4347
rect 1533 4333 1547 4347
rect 1573 4333 1587 4347
rect 1653 4333 1667 4347
rect 1713 4333 1727 4347
rect 1913 4333 1927 4347
rect 1953 4333 1967 4347
rect 2013 4333 2027 4347
rect 2273 4334 2287 4348
rect 2433 4333 2447 4347
rect 2653 4333 2667 4347
rect 2713 4333 2727 4347
rect 3113 4333 3127 4347
rect 3153 4333 3167 4347
rect 3193 4333 3207 4347
rect 3293 4333 3307 4347
rect 3333 4333 3347 4347
rect 3473 4333 3487 4347
rect 3513 4333 3527 4347
rect 3693 4333 3707 4347
rect 3813 4333 3827 4347
rect 4053 4333 4067 4347
rect 4093 4333 4107 4347
rect 4173 4333 4187 4347
rect 4433 4333 4447 4347
rect 4493 4333 4507 4347
rect 4533 4333 4547 4347
rect 4613 4333 4627 4347
rect 4753 4333 4767 4347
rect 4793 4333 4807 4347
rect 5193 4333 5207 4347
rect 93 4313 107 4327
rect 213 4313 227 4327
rect 353 4314 367 4328
rect 933 4313 947 4327
rect 1013 4313 1027 4327
rect 1153 4313 1167 4327
rect 1213 4313 1227 4327
rect 1293 4313 1307 4327
rect 1853 4313 1867 4327
rect 2133 4314 2147 4328
rect 2193 4313 2207 4327
rect 2353 4313 2367 4327
rect 2593 4313 2607 4327
rect 2753 4313 2767 4327
rect 2893 4313 2907 4327
rect 3073 4313 3087 4327
rect 3393 4313 3407 4327
rect 3613 4313 3627 4327
rect 3853 4313 3867 4327
rect 3953 4313 3967 4327
rect 4233 4313 4247 4327
rect 4893 4313 4907 4327
rect 5033 4313 5047 4327
rect 5313 4333 5327 4347
rect 5233 4313 5247 4327
rect 5473 4313 5487 4327
rect 233 4293 247 4307
rect 333 4293 347 4307
rect 473 4293 487 4307
rect 513 4293 527 4307
rect 573 4293 587 4307
rect 673 4293 687 4307
rect 793 4293 807 4307
rect 833 4293 847 4307
rect 973 4292 987 4306
rect 1373 4293 1387 4307
rect 1413 4293 1427 4307
rect 1513 4293 1527 4307
rect 1553 4293 1567 4307
rect 1613 4293 1627 4307
rect 1673 4293 1687 4307
rect 1893 4293 1907 4307
rect 1933 4293 1947 4307
rect 2033 4293 2047 4307
rect 2113 4293 2127 4307
rect 2453 4293 2467 4307
rect 2693 4293 2707 4307
rect 2733 4293 2747 4307
rect 2913 4293 2927 4307
rect 3133 4293 3147 4307
rect 3173 4294 3187 4308
rect 3233 4293 3247 4307
rect 3273 4293 3287 4307
rect 3453 4293 3467 4307
rect 3493 4293 3507 4307
rect 3573 4293 3587 4307
rect 3673 4293 3687 4307
rect 3713 4293 3727 4307
rect 3833 4293 3847 4307
rect 4073 4293 4087 4307
rect 4113 4293 4127 4307
rect 4213 4293 4227 4307
rect 4473 4293 4487 4307
rect 4513 4293 4527 4307
rect 4553 4293 4567 4307
rect 4633 4293 4647 4307
rect 4673 4293 4687 4307
rect 4733 4293 4747 4307
rect 4833 4292 4847 4306
rect 4873 4293 4887 4307
rect 5053 4293 5067 4307
rect 5273 4293 5287 4307
rect 5433 4293 5447 4307
rect 5453 4293 5467 4307
rect 53 4273 67 4287
rect 73 4273 87 4287
rect 113 4273 127 4287
rect 153 4273 167 4287
rect 373 4273 387 4287
rect 1033 4272 1047 4286
rect 1073 4273 1087 4287
rect 1133 4273 1147 4287
rect 1173 4273 1187 4287
rect 1633 4273 1647 4287
rect 1853 4272 1867 4286
rect 2213 4273 2227 4287
rect 2413 4273 2427 4287
rect 2513 4273 2527 4287
rect 2553 4273 2567 4287
rect 2833 4273 2847 4287
rect 2873 4273 2887 4287
rect 2973 4273 2987 4287
rect 3013 4273 3027 4287
rect 3893 4273 3907 4287
rect 3933 4273 3947 4287
rect 3973 4273 3987 4287
rect 4273 4273 4287 4287
rect 4313 4273 4327 4287
rect 4972 4273 4986 4287
rect 4993 4273 5007 4287
rect 5133 4273 5147 4287
rect 5173 4273 5187 4287
rect 5333 4273 5347 4287
rect 5373 4273 5387 4287
rect 5493 4273 5507 4287
rect 253 4253 267 4267
rect 313 4253 327 4267
rect 333 4253 347 4267
rect 1773 4253 1787 4267
rect 2093 4253 2107 4267
rect 2313 4253 2327 4267
rect 2713 4253 2727 4267
rect 2933 4253 2947 4267
rect 3813 4253 3827 4267
rect 4853 4253 4867 4267
rect 5073 4253 5087 4267
rect 5093 4253 5107 4267
rect 5433 4253 5447 4267
rect 233 4073 247 4087
rect 473 4073 487 4087
rect 673 4073 687 4087
rect 1433 4073 1447 4087
rect 1653 4073 1667 4087
rect 2353 4073 2367 4087
rect 3753 4073 3767 4087
rect 4193 4073 4207 4087
rect 4593 4073 4607 4087
rect 5253 4073 5267 4087
rect 5453 4073 5467 4087
rect 53 4053 67 4067
rect 93 4053 107 4067
rect 173 4053 187 4067
rect 353 4053 367 4067
rect 733 4053 747 4067
rect 813 4053 827 4067
rect 853 4053 867 4067
rect 1493 4053 1507 4067
rect 1553 4053 1567 4067
rect 1713 4053 1727 4067
rect 1793 4054 1807 4068
rect 1833 4053 1847 4067
rect 2173 4053 2187 4067
rect 2213 4053 2227 4067
rect 2253 4053 2267 4067
rect 2413 4053 2427 4067
rect 2453 4053 2467 4067
rect 2693 4053 2707 4067
rect 2873 4053 2887 4067
rect 2933 4053 2947 4067
rect 3293 4053 3307 4067
rect 3333 4053 3347 4067
rect 3653 4053 3667 4067
rect 3693 4053 3707 4067
rect 3853 4053 3867 4067
rect 3973 4053 3987 4067
rect 4013 4053 4027 4067
rect 4093 4053 4107 4067
rect 4133 4053 4147 4067
rect 4273 4053 4287 4067
rect 4713 4053 4727 4067
rect 5313 4053 5327 4067
rect 5353 4053 5367 4067
rect 213 4033 227 4047
rect 313 4033 327 4047
rect 453 4033 467 4047
rect 553 4033 567 4047
rect 593 4033 607 4047
rect 693 4033 707 4047
rect 933 4033 947 4047
rect 973 4033 987 4047
rect 1053 4033 1067 4047
rect 1093 4033 1107 4047
rect 1213 4033 1227 4047
rect 1253 4033 1267 4047
rect 1333 4033 1347 4047
rect 1453 4033 1467 4047
rect 1673 4033 1687 4047
rect 1933 4032 1947 4046
rect 1973 4033 1987 4047
rect 2093 4033 2107 4047
rect 2333 4033 2347 4047
rect 2533 4033 2547 4047
rect 2573 4033 2587 4047
rect 2793 4033 2807 4047
rect 2833 4033 2847 4047
rect 3013 4033 3027 4047
rect 3053 4033 3067 4047
rect 3173 4033 3187 4047
rect 3393 4033 3407 4047
rect 3493 4033 3507 4047
rect 3553 4033 3567 4047
rect 3773 4033 3787 4047
rect 3913 4033 3927 4047
rect 4213 4033 4227 4047
rect 4313 4033 4327 4047
rect 4353 4033 4367 4047
rect 4453 4033 4467 4047
rect 4493 4033 4507 4047
rect 4613 4033 4627 4047
rect 4773 4033 4787 4047
rect 4813 4033 4827 4047
rect 5013 4033 5027 4047
rect 5073 4033 5087 4047
rect 5233 4033 5247 4047
rect 5273 4034 5287 4048
rect 5433 4033 5447 4047
rect 113 4013 127 4027
rect 193 4013 207 4027
rect 433 4013 447 4027
rect 713 4013 727 4027
rect 773 4013 787 4027
rect 1473 4012 1487 4026
rect 1693 4013 1707 4027
rect 1813 4013 1827 4027
rect 2133 4013 2147 4027
rect 2233 4013 2247 4027
rect 2313 4013 2327 4027
rect 2393 4013 2407 4027
rect 2893 4013 2907 4027
rect 3213 4013 3227 4027
rect 3253 4013 3267 4027
rect 3353 4013 3367 4027
rect 3433 4012 3447 4026
rect 3593 4012 3607 4026
rect 3633 4013 3647 4027
rect 3733 4013 3747 4027
rect 3793 4013 3807 4027
rect 4013 4013 4027 4027
rect 4053 4013 4067 4027
rect 4233 4013 4247 4027
rect 4633 4013 4647 4027
rect 5293 4013 5307 4027
rect 5413 4013 5427 4027
rect 333 3993 347 4007
rect 473 3993 487 4007
rect 613 3993 627 4007
rect 913 3992 927 4006
rect 953 3993 967 4007
rect 1033 3993 1047 4007
rect 1073 3993 1087 4007
rect 1113 3993 1127 4007
rect 1193 3993 1207 4007
rect 1233 3992 1247 4006
rect 1273 3993 1287 4007
rect 1353 3993 1367 4007
rect 1613 3993 1627 4007
rect 1653 3993 1667 4007
rect 1853 3993 1867 4007
rect 1993 3993 2007 4007
rect 2033 3993 2047 4007
rect 2513 3993 2527 4007
rect 2553 3993 2567 4007
rect 2613 3993 2627 4007
rect 2733 3993 2747 4007
rect 2773 3993 2787 4007
rect 2813 3992 2827 4006
rect 2993 3993 3007 4007
rect 3033 3993 3047 4007
rect 3073 3994 3087 4008
rect 3493 3993 3507 4007
rect 3533 3993 3547 4007
rect 3833 3993 3847 4007
rect 4333 3993 4347 4007
rect 4393 3993 4407 4007
rect 4473 3993 4487 4007
rect 4593 3993 4607 4007
rect 4733 3993 4747 4007
rect 4793 3993 4807 4007
rect 4893 3993 4907 4007
rect 4993 3993 5007 4007
rect 5033 3993 5047 4007
rect 5113 3993 5127 4007
rect 5153 3993 5167 4007
rect 3393 3973 3407 3987
rect 113 3953 127 3967
rect 173 3953 187 3967
rect 1513 3833 1527 3847
rect 4753 3833 4767 3847
rect 5113 3833 5127 3847
rect 5273 3833 5287 3847
rect 5453 3833 5467 3847
rect 53 3813 67 3827
rect 93 3813 107 3827
rect 233 3814 247 3828
rect 333 3813 347 3827
rect 533 3812 547 3826
rect 573 3813 587 3827
rect 653 3813 667 3827
rect 773 3813 787 3827
rect 813 3813 827 3827
rect 973 3813 987 3827
rect 1033 3813 1047 3827
rect 1253 3813 1267 3827
rect 1353 3813 1367 3827
rect 1373 3813 1387 3827
rect 1673 3813 1687 3827
rect 1713 3813 1727 3827
rect 1773 3813 1787 3827
rect 1853 3813 1867 3827
rect 1893 3813 1907 3827
rect 1933 3813 1947 3827
rect 2153 3813 2167 3827
rect 2193 3813 2207 3827
rect 2233 3813 2247 3827
rect 2433 3813 2447 3827
rect 2473 3813 2487 3827
rect 2553 3813 2567 3827
rect 2673 3813 2687 3827
rect 2773 3813 2787 3827
rect 2873 3813 2887 3827
rect 2973 3813 2987 3827
rect 3053 3813 3067 3827
rect 3253 3813 3267 3827
rect 3373 3813 3387 3827
rect 3413 3812 3427 3826
rect 3513 3813 3527 3827
rect 3553 3813 3567 3827
rect 3633 3813 3647 3827
rect 3693 3813 3707 3827
rect 3753 3813 3767 3827
rect 3873 3812 3887 3826
rect 3933 3813 3947 3827
rect 3973 3813 3987 3827
rect 4033 3813 4047 3827
rect 4133 3813 4147 3827
rect 4233 3813 4247 3827
rect 4373 3813 4387 3827
rect 4433 3813 4447 3827
rect 4573 3813 4587 3827
rect 4913 3813 4927 3827
rect 5013 3813 5027 3827
rect 5073 3813 5087 3827
rect 193 3793 207 3807
rect 433 3793 447 3807
rect 693 3793 707 3807
rect 853 3793 867 3807
rect 993 3793 1007 3807
rect 1073 3793 1087 3807
rect 1133 3793 1147 3807
rect 1313 3793 1327 3807
rect 1493 3793 1507 3807
rect 2013 3793 2027 3807
rect 2293 3793 2307 3807
rect 2613 3793 2627 3807
rect 2833 3793 2847 3807
rect 3213 3793 3227 3807
rect 4093 3793 4107 3807
rect 4333 3793 4347 3807
rect 4473 3793 4487 3807
rect 4713 3793 4727 3807
rect 4753 3793 4767 3807
rect 4833 3793 4847 3807
rect 5213 3793 5227 3807
rect 5313 3793 5327 3807
rect 5433 3793 5447 3807
rect 73 3773 87 3787
rect 113 3773 127 3787
rect 213 3773 227 3787
rect 313 3773 327 3787
rect 353 3773 367 3787
rect 553 3773 567 3787
rect 593 3773 607 3787
rect 713 3773 727 3787
rect 813 3773 827 3787
rect 1173 3772 1187 3786
rect 1393 3773 1407 3787
rect 1433 3773 1447 3787
rect 1653 3773 1667 3787
rect 1693 3773 1707 3787
rect 1753 3774 1767 3788
rect 1833 3773 1847 3787
rect 1953 3773 1967 3787
rect 1973 3773 1987 3787
rect 2053 3773 2067 3787
rect 2173 3773 2187 3787
rect 2253 3773 2267 3787
rect 2413 3773 2427 3787
rect 2453 3773 2467 3787
rect 2573 3773 2587 3787
rect 2673 3773 2687 3787
rect 2713 3773 2727 3787
rect 2913 3773 2927 3787
rect 2953 3773 2967 3787
rect 3073 3773 3087 3787
rect 3093 3773 3107 3787
rect 3273 3773 3287 3787
rect 3313 3773 3327 3787
rect 3433 3773 3447 3787
rect 3493 3773 3507 3787
rect 3533 3773 3547 3787
rect 3613 3773 3627 3787
rect 3773 3773 3787 3787
rect 3813 3773 3827 3787
rect 3913 3773 3927 3787
rect 3953 3773 3967 3787
rect 4013 3773 4027 3787
rect 4153 3773 4167 3787
rect 4193 3773 4207 3787
rect 4393 3773 4407 3787
rect 4433 3773 4447 3787
rect 4793 3773 4807 3787
rect 4873 3773 4887 3787
rect 4993 3773 5007 3787
rect 5133 3773 5147 3787
rect 5173 3773 5187 3787
rect 5273 3772 5287 3786
rect 5393 3773 5407 3787
rect 153 3753 167 3767
rect 413 3753 427 3767
rect 453 3753 467 3767
rect 653 3752 667 3766
rect 913 3753 927 3767
rect 953 3753 967 3767
rect 1273 3753 1287 3767
rect 1313 3753 1327 3767
rect 1513 3753 1527 3767
rect 1553 3753 1567 3767
rect 2313 3753 2327 3767
rect 2353 3752 2367 3766
rect 2793 3753 2807 3767
rect 2833 3753 2847 3767
rect 3153 3753 3167 3767
rect 3193 3753 3207 3767
rect 4233 3753 4247 3767
rect 4293 3753 4307 3767
rect 4613 3753 4627 3767
rect 4653 3753 4667 3767
rect 233 3733 247 3747
rect 733 3733 747 3747
rect 993 3573 1007 3587
rect 1033 3573 1047 3587
rect 173 3553 187 3567
rect 193 3553 207 3567
rect 2413 3553 2427 3567
rect 3833 3553 3847 3567
rect 5373 3553 5387 3567
rect 253 3533 267 3547
rect 953 3533 967 3547
rect 993 3533 1007 3547
rect 1333 3533 1347 3547
rect 1373 3533 1387 3547
rect 1413 3533 1427 3547
rect 1933 3533 1947 3547
rect 1973 3534 1987 3548
rect 2013 3533 2027 3547
rect 2053 3533 2067 3547
rect 2133 3533 2147 3547
rect 2173 3533 2187 3547
rect 2453 3533 2467 3547
rect 2893 3533 2907 3547
rect 2933 3533 2947 3547
rect 3633 3533 3647 3547
rect 3673 3533 3687 3547
rect 3913 3533 3927 3547
rect 3953 3533 3967 3547
rect 3993 3533 4007 3547
rect 4053 3533 4067 3547
rect 4093 3533 4107 3547
rect 4473 3533 4487 3547
rect 4513 3533 4527 3547
rect 5173 3533 5187 3547
rect 5213 3533 5227 3547
rect 5273 3533 5287 3547
rect 93 3513 107 3527
rect 133 3513 147 3527
rect 213 3514 227 3528
rect 313 3513 327 3527
rect 433 3513 447 3527
rect 473 3513 487 3527
rect 553 3513 567 3527
rect 593 3513 607 3527
rect 693 3513 707 3527
rect 733 3513 747 3527
rect 773 3512 787 3526
rect 813 3513 827 3527
rect 853 3513 867 3527
rect 1093 3513 1107 3527
rect 1133 3513 1147 3527
rect 1213 3513 1227 3527
rect 1253 3513 1267 3527
rect 1473 3513 1487 3527
rect 1513 3513 1527 3527
rect 1693 3513 1707 3527
rect 1733 3513 1747 3527
rect 1813 3513 1827 3527
rect 1853 3513 1867 3527
rect 2273 3513 2287 3527
rect 2313 3513 2327 3527
rect 2533 3513 2547 3527
rect 2573 3513 2587 3527
rect 233 3493 247 3507
rect 953 3493 967 3507
rect 1353 3493 1367 3507
rect 1633 3493 1647 3507
rect 1973 3493 1987 3507
rect 2053 3493 2067 3507
rect 2173 3493 2187 3507
rect 2473 3493 2487 3507
rect 2693 3493 2707 3507
rect 2733 3493 2747 3507
rect 3053 3513 3067 3527
rect 3753 3513 3767 3527
rect 3853 3513 3867 3527
rect 4193 3513 4207 3527
rect 4233 3513 4247 3527
rect 4353 3513 4367 3527
rect 4553 3513 4567 3527
rect 4733 3513 4747 3527
rect 4773 3514 4787 3528
rect 4873 3513 4887 3527
rect 4933 3513 4947 3527
rect 4973 3513 4987 3527
rect 5053 3513 5067 3527
rect 5093 3513 5107 3527
rect 5353 3513 5367 3527
rect 3173 3493 3187 3507
rect 3213 3493 3227 3507
rect 3413 3493 3427 3507
rect 3453 3493 3467 3507
rect 3593 3493 3607 3507
rect 3713 3494 3727 3508
rect 3873 3493 3887 3507
rect 3933 3493 3947 3507
rect 4133 3493 4147 3507
rect 4313 3493 4327 3507
rect 4433 3493 4447 3507
rect 4653 3494 4667 3508
rect 4833 3493 4847 3507
rect 5153 3493 5167 3507
rect 5333 3493 5347 3507
rect 33 3473 47 3487
rect 113 3473 127 3487
rect 353 3473 367 3487
rect 433 3472 447 3486
rect 493 3473 507 3487
rect 533 3473 547 3487
rect 573 3473 587 3487
rect 673 3473 687 3487
rect 753 3473 767 3487
rect 793 3473 807 3487
rect 833 3473 847 3487
rect 1053 3473 1067 3487
rect 1113 3473 1127 3487
rect 1153 3473 1167 3487
rect 1273 3472 1287 3486
rect 1453 3473 1467 3487
rect 1493 3473 1507 3487
rect 1533 3473 1547 3487
rect 1673 3473 1687 3487
rect 1713 3473 1727 3487
rect 1773 3473 1787 3487
rect 1873 3473 1887 3487
rect 2293 3473 2307 3487
rect 2333 3473 2347 3487
rect 2493 3473 2507 3487
rect 2513 3473 2527 3487
rect 2553 3473 2567 3487
rect 2813 3473 2827 3487
rect 3033 3473 3047 3487
rect 3073 3473 3087 3487
rect 3293 3473 3307 3487
rect 3533 3473 3547 3487
rect 3793 3473 3807 3487
rect 3833 3473 3847 3487
rect 4173 3473 4187 3487
rect 4253 3473 4267 3487
rect 4393 3473 4407 3487
rect 4573 3473 4587 3487
rect 4653 3472 4667 3486
rect 4753 3473 4767 3487
rect 4913 3473 4927 3487
rect 4953 3473 4967 3487
rect 5013 3473 5027 3487
rect 5113 3473 5127 3487
rect 5433 3473 5447 3487
rect 5493 3473 5507 3487
rect 4793 3453 4807 3467
rect 1013 3313 1027 3327
rect 3593 3313 3607 3327
rect 3853 3333 3867 3347
rect 33 3293 47 3307
rect 153 3293 167 3307
rect 213 3293 227 3307
rect 433 3293 447 3307
rect 473 3293 487 3307
rect 533 3293 547 3307
rect 773 3293 787 3307
rect 813 3293 827 3307
rect 873 3293 887 3307
rect 973 3293 987 3307
rect 1173 3293 1187 3307
rect 1553 3293 1567 3307
rect 1693 3293 1707 3307
rect 1813 3293 1827 3307
rect 2093 3293 2107 3307
rect 2193 3293 2207 3307
rect 2313 3293 2327 3307
rect 2573 3293 2587 3307
rect 2613 3293 2627 3307
rect 3153 3293 3167 3307
rect 3193 3293 3207 3307
rect 3293 3293 3307 3307
rect 3333 3293 3347 3307
rect 3393 3293 3407 3307
rect 3433 3293 3447 3307
rect 3633 3293 3647 3307
rect 3693 3293 3707 3307
rect 3853 3293 3867 3307
rect 4113 3293 4127 3307
rect 4333 3293 4347 3307
rect 4373 3293 4387 3307
rect 4453 3293 4467 3307
rect 4493 3293 4507 3307
rect 4573 3293 4587 3307
rect 4753 3293 4767 3307
rect 4793 3293 4807 3307
rect 4933 3293 4947 3307
rect 5113 3293 5127 3307
rect 5213 3293 5227 3307
rect 5473 3293 5487 3307
rect 133 3273 147 3287
rect 293 3273 307 3287
rect 653 3273 667 3287
rect 1093 3273 1107 3287
rect 1353 3273 1367 3287
rect 1453 3273 1467 3287
rect 1513 3273 1527 3287
rect 1633 3273 1647 3287
rect 1893 3273 1907 3287
rect 2033 3273 2047 3287
rect 2253 3273 2267 3287
rect 53 3254 67 3268
rect 93 3253 107 3267
rect 2393 3272 2407 3286
rect 2673 3273 2687 3287
rect 2873 3273 2887 3287
rect 2993 3273 3007 3287
rect 3093 3273 3107 3287
rect 3553 3273 3567 3287
rect 3773 3273 3787 3287
rect 4053 3273 4067 3287
rect 4193 3273 4207 3287
rect 4653 3273 4667 3287
rect 4973 3273 4987 3287
rect 273 3253 287 3267
rect 353 3253 367 3267
rect 513 3253 527 3267
rect 553 3253 567 3267
rect 673 3253 687 3267
rect 793 3253 807 3267
rect 833 3253 847 3267
rect 873 3252 887 3266
rect 933 3252 947 3266
rect 1133 3253 1147 3267
rect 1373 3253 1387 3267
rect 1593 3253 1607 3267
rect 1673 3253 1687 3267
rect 1713 3253 1727 3267
rect 1793 3253 1807 3267
rect 1913 3253 1927 3267
rect 2073 3253 2087 3267
rect 2153 3253 2167 3267
rect 2433 3253 2447 3267
rect 2593 3253 2607 3267
rect 2633 3253 2647 3267
rect 3133 3253 3147 3267
rect 3173 3253 3187 3267
rect 3273 3253 3287 3267
rect 3313 3253 3327 3267
rect 3413 3253 3427 3267
rect 3453 3253 3467 3267
rect 3513 3253 3527 3267
rect 3613 3253 3627 3267
rect 3653 3253 3667 3267
rect 3733 3253 3747 3267
rect 3913 3253 3927 3267
rect 4133 3253 4147 3267
rect 4173 3253 4187 3267
rect 4273 3254 4287 3268
rect 4393 3253 4407 3267
rect 4433 3253 4447 3267
rect 4513 3253 4527 3267
rect 4553 3253 4567 3267
rect 4673 3254 4687 3268
rect 4773 3253 4787 3267
rect 4813 3253 4827 3267
rect 4873 3253 4887 3267
rect 5133 3253 5147 3267
rect 5173 3253 5187 3267
rect 313 3233 327 3247
rect 633 3233 647 3247
rect 1193 3233 1207 3247
rect 1233 3233 1247 3247
rect 1273 3233 1287 3247
rect 1453 3233 1467 3247
rect 1493 3233 1507 3247
rect 1873 3233 1887 3247
rect 1993 3233 2007 3247
rect 2213 3233 2227 3247
rect 2253 3233 2267 3247
rect 2713 3233 2727 3247
rect 2753 3233 2767 3247
rect 2813 3233 2827 3247
rect 2853 3233 2867 3247
rect 2913 3234 2927 3248
rect 2953 3233 2967 3247
rect 3033 3233 3047 3247
rect 3073 3233 3087 3247
rect 3973 3233 3987 3247
rect 4013 3233 4027 3247
rect 213 3213 227 3227
rect 253 3213 267 3227
rect 693 3213 707 3227
rect 1393 3213 1407 3227
rect 1933 3213 1947 3227
rect 4273 3232 4287 3246
rect 4593 3233 4607 3247
rect 4993 3233 5007 3247
rect 5033 3233 5047 3247
rect 4153 3213 4167 3227
rect 4673 3213 4687 3227
rect 4693 3213 4707 3227
rect 5373 3273 5387 3287
rect 5393 3253 5407 3267
rect 5433 3253 5447 3267
rect 5253 3233 5267 3247
rect 5293 3233 5307 3247
rect 5353 3233 5367 3247
rect 5213 3212 5227 3226
rect 5413 3213 5427 3227
rect 2033 3193 2047 3207
rect 113 3033 127 3047
rect 493 3033 507 3047
rect 633 3033 647 3047
rect 2033 3033 2047 3047
rect 5313 3033 5327 3047
rect 33 3013 47 3027
rect 433 3013 447 3027
rect 533 3013 547 3027
rect 1233 3013 1247 3027
rect 1293 3013 1307 3027
rect 1333 3013 1347 3027
rect 1413 3013 1427 3027
rect 1453 3013 1467 3027
rect 2133 3013 2147 3027
rect 3253 3013 3267 3027
rect 3293 3013 3307 3027
rect 4413 3013 4427 3027
rect 4453 3013 4467 3027
rect 4533 3013 4547 3027
rect 4573 3013 4587 3027
rect 5373 3013 5387 3027
rect 93 2993 107 3007
rect 153 2993 167 3007
rect 193 2993 207 3007
rect 313 2993 327 3007
rect 353 2993 367 3007
rect 473 2993 487 3007
rect 613 2993 627 3007
rect 713 2993 727 3007
rect 753 2993 767 3007
rect 853 2993 867 3007
rect 893 2993 907 3007
rect 933 2993 947 3007
rect 1073 2993 1087 3007
rect 1113 2993 1127 3007
rect 1173 2993 1187 3007
rect 1553 2993 1567 3007
rect 1593 2993 1607 3007
rect 1673 2993 1687 3007
rect 1793 2993 1807 3007
rect 1933 2993 1947 3007
rect 1973 2993 1987 3007
rect 2053 2993 2067 3007
rect 2173 2992 2187 3006
rect 2213 2993 2227 3007
rect 2393 2993 2407 3007
rect 2673 2993 2687 3007
rect 3373 2993 3387 3007
rect 3413 2993 3427 3007
rect 3473 2993 3487 3007
rect 3613 2993 3627 3007
rect 3833 2993 3847 3007
rect 3873 2993 3887 3007
rect 4213 2993 4227 3007
rect 4253 2993 4267 3007
rect 4333 2993 4347 3007
rect 4633 2993 4647 3007
rect 4833 2993 4847 3007
rect 4873 2993 4887 3007
rect 5033 2993 5047 3007
rect 5073 2993 5087 3007
rect 5113 2993 5127 3007
rect 5153 2993 5167 3007
rect 5333 2993 5347 3007
rect 73 2973 87 2987
rect 453 2973 467 2987
rect 593 2973 607 2987
rect 1213 2973 1227 2987
rect 1273 2973 1287 2987
rect 1353 2973 1367 2987
rect 1753 2973 1767 2987
rect 2073 2973 2087 2987
rect 2353 2973 2367 2987
rect 2513 2973 2527 2987
rect 2713 2973 2727 2987
rect 2733 2973 2747 2987
rect 2873 2973 2887 2987
rect 3033 2973 3047 2987
rect 3073 2973 3087 2987
rect 3233 2973 3247 2987
rect 3653 2973 3667 2987
rect 3973 2973 3987 2987
rect 4093 2973 4107 2987
rect 4413 2972 4427 2986
rect 4593 2973 4607 2987
rect 4733 2973 4747 2987
rect 4913 2973 4927 2987
rect 4993 2973 5007 2987
rect 5353 2973 5367 2987
rect 173 2953 187 2967
rect 233 2953 247 2967
rect 293 2953 307 2967
rect 373 2953 387 2967
rect 633 2953 647 2967
rect 773 2953 787 2967
rect 833 2953 847 2967
rect 873 2953 887 2967
rect 1013 2953 1027 2967
rect 1053 2953 1067 2967
rect 1133 2953 1147 2967
rect 1533 2953 1547 2967
rect 1573 2953 1587 2967
rect 1613 2953 1627 2967
rect 1653 2953 1667 2967
rect 1713 2953 1727 2967
rect 1793 2953 1807 2967
rect 1832 2953 1846 2967
rect 1853 2953 1867 2967
rect 1953 2953 1967 2967
rect 2033 2953 2047 2967
rect 2153 2953 2167 2967
rect 2193 2953 2207 2967
rect 2273 2953 2287 2967
rect 2553 2953 2567 2967
rect 2793 2953 2807 2967
rect 2913 2953 2927 2967
rect 3153 2953 3167 2967
rect 3353 2953 3367 2967
rect 3393 2953 3407 2967
rect 3493 2953 3507 2967
rect 3733 2953 3747 2967
rect 3813 2953 3827 2967
rect 3853 2953 3867 2967
rect 4233 2953 4247 2967
rect 4273 2953 4287 2967
rect 4373 2953 4387 2967
rect 4653 2953 4667 2967
rect 4773 2953 4787 2967
rect 5053 2953 5067 2967
rect 5093 2953 5107 2967
rect 5133 2953 5147 2967
rect 5213 2953 5227 2967
rect 5453 2953 5467 2967
rect 5513 2953 5527 2967
rect 1193 2932 1207 2946
rect 4873 2933 4887 2947
rect 4953 2933 4967 2947
rect 1893 2813 1907 2827
rect 1133 2793 1147 2807
rect 1473 2793 1487 2807
rect 2133 2793 2147 2807
rect 93 2773 107 2787
rect 133 2773 147 2787
rect 193 2773 207 2787
rect 393 2773 407 2787
rect 413 2772 427 2786
rect 453 2773 467 2787
rect 513 2773 527 2787
rect 733 2773 747 2787
rect 813 2773 827 2787
rect 933 2772 947 2786
rect 973 2773 987 2787
rect 1053 2773 1067 2787
rect 1273 2773 1287 2787
rect 1393 2773 1407 2787
rect 1553 2773 1567 2787
rect 1633 2772 1647 2786
rect 1753 2773 1767 2787
rect 1793 2773 1807 2787
rect 1853 2773 1867 2787
rect 2013 2773 2027 2787
rect 2433 2793 2447 2807
rect 3753 2793 3767 2807
rect 3853 2793 3867 2807
rect 3933 2793 3947 2807
rect 2873 2773 2887 2787
rect 2913 2773 2927 2787
rect 3033 2772 3047 2786
rect 3233 2773 3247 2787
rect 3273 2773 3287 2787
rect 3493 2773 3507 2787
rect 3613 2773 3627 2787
rect 4153 2773 4167 2787
rect 4233 2774 4247 2788
rect 4273 2773 4287 2787
rect 4313 2773 4327 2787
rect 4413 2773 4427 2787
rect 4453 2773 4467 2787
rect 4673 2773 4687 2787
rect 4793 2773 4807 2787
rect 4893 2773 4907 2787
rect 4973 2773 4987 2787
rect 5013 2773 5027 2787
rect 5053 2773 5067 2787
rect 5273 2773 5287 2787
rect 5333 2773 5347 2787
rect 293 2753 307 2767
rect 553 2753 567 2767
rect 673 2753 687 2767
rect 873 2753 887 2767
rect 1113 2753 1127 2767
rect 1193 2753 1207 2767
rect 1494 2753 1508 2767
rect 1953 2753 1967 2767
rect 2113 2753 2127 2767
rect 2353 2753 2367 2767
rect 2493 2753 2507 2767
rect 2653 2753 2667 2767
rect 113 2733 127 2747
rect 173 2733 187 2747
rect 213 2733 227 2747
rect 313 2733 327 2747
rect 433 2733 447 2747
rect 693 2733 707 2747
rect 793 2733 807 2747
rect 833 2733 847 2747
rect 993 2733 1007 2747
rect 1033 2733 1047 2747
rect 1153 2733 1167 2747
rect 1333 2733 1347 2747
rect 1373 2732 1387 2746
rect 1453 2733 1467 2747
rect 1653 2733 1667 2747
rect 1693 2733 1707 2747
rect 1793 2733 1807 2747
rect 1833 2733 1847 2747
rect 1913 2733 1927 2747
rect 1993 2733 2007 2747
rect 2073 2733 2087 2747
rect 2313 2733 2327 2747
rect 3053 2753 3067 2767
rect 3133 2753 3147 2767
rect 3373 2753 3387 2767
rect 3413 2753 3427 2767
rect 3693 2753 3707 2767
rect 3913 2753 3927 2767
rect 4073 2753 4087 2767
rect 4533 2753 4547 2767
rect 4693 2753 4707 2767
rect 5193 2753 5207 2767
rect 5513 2753 5527 2767
rect 2893 2733 2907 2747
rect 3213 2733 3227 2747
rect 3253 2733 3267 2747
rect 3593 2733 3607 2747
rect 3633 2733 3647 2747
rect 3813 2733 3827 2747
rect 3853 2733 3867 2747
rect 4053 2733 4067 2747
rect 4253 2733 4267 2747
rect 4293 2733 4307 2747
rect 4333 2733 4347 2747
rect 4573 2733 4587 2747
rect 4733 2733 4747 2747
rect 4773 2733 4787 2747
rect 4993 2733 5007 2747
rect 5033 2733 5047 2747
rect 5153 2733 5167 2747
rect 5353 2733 5367 2747
rect 273 2713 287 2727
rect 473 2713 487 2727
rect 533 2713 547 2727
rect 573 2713 587 2727
rect 633 2713 647 2727
rect 1193 2713 1207 2727
rect 1233 2713 1247 2727
rect 1613 2713 1627 2727
rect 2153 2713 2167 2727
rect 2213 2713 2227 2727
rect 2713 2713 2727 2727
rect 2753 2713 2767 2727
rect 2973 2713 2987 2727
rect 3013 2713 3027 2727
rect 4813 2713 4827 2727
rect 5453 2713 5467 2727
rect 5493 2713 5507 2727
rect 333 2693 347 2707
rect 713 2693 727 2707
rect 273 2512 287 2526
rect 733 2513 747 2527
rect 953 2513 967 2527
rect 1213 2513 1227 2527
rect 5453 2513 5467 2527
rect 5493 2513 5507 2527
rect 173 2493 187 2507
rect 653 2493 667 2507
rect 873 2493 887 2507
rect 1113 2493 1127 2507
rect 93 2473 107 2487
rect 133 2473 147 2487
rect 253 2473 267 2487
rect 373 2473 387 2487
rect 413 2473 427 2487
rect 553 2473 567 2487
rect 593 2473 607 2487
rect 713 2473 727 2487
rect 853 2473 867 2487
rect 933 2473 947 2487
rect 1193 2473 1207 2487
rect 1293 2473 1307 2487
rect 1333 2473 1347 2487
rect 1453 2473 1467 2487
rect 1493 2473 1507 2487
rect 1573 2473 1587 2487
rect 1613 2473 1627 2487
rect 1873 2473 1887 2487
rect 1953 2473 1967 2487
rect 2113 2473 2127 2487
rect 2293 2473 2307 2487
rect 2333 2473 2347 2487
rect 2653 2473 2667 2487
rect 2873 2473 2887 2487
rect 2913 2473 2927 2487
rect 2953 2473 2967 2487
rect 3073 2473 3087 2487
rect 3113 2473 3127 2487
rect 3253 2473 3267 2487
rect 3653 2473 3667 2487
rect 3813 2473 3827 2487
rect 3993 2473 4007 2487
rect 4133 2473 4147 2487
rect 4173 2473 4187 2487
rect 4253 2473 4267 2487
rect 4273 2473 4287 2487
rect 4553 2473 4567 2487
rect 4593 2473 4607 2487
rect 4713 2473 4727 2487
rect 4753 2473 4767 2487
rect 4813 2473 4827 2487
rect 5273 2473 5287 2487
rect 233 2453 247 2467
rect 333 2453 347 2467
rect 693 2453 707 2467
rect 913 2453 927 2467
rect 1013 2453 1027 2467
rect 1173 2453 1187 2467
rect 1673 2453 1687 2467
rect 1833 2453 1847 2467
rect 5333 2472 5347 2486
rect 5413 2473 5427 2487
rect 5453 2473 5467 2487
rect 1913 2453 1927 2467
rect 2073 2453 2087 2467
rect 2393 2453 2407 2467
rect 2553 2453 2567 2467
rect 2693 2453 2707 2467
rect 3013 2453 3027 2467
rect 3293 2453 3307 2467
rect 3493 2453 3507 2467
rect 3533 2453 3547 2467
rect 3713 2453 3727 2467
rect 3953 2453 3967 2467
rect 4353 2453 4367 2467
rect 4433 2453 4447 2467
rect 4473 2453 4487 2467
rect 4893 2453 4907 2467
rect 4993 2453 5007 2467
rect 5033 2453 5047 2467
rect 5213 2453 5227 2467
rect 13 2433 27 2447
rect 113 2433 127 2447
rect 453 2433 467 2447
rect 513 2433 527 2447
rect 573 2433 587 2447
rect 793 2433 807 2447
rect 1073 2433 1087 2447
rect 1313 2433 1327 2447
rect 1353 2433 1367 2447
rect 1433 2433 1447 2447
rect 1473 2433 1487 2447
rect 1513 2433 1527 2447
rect 1553 2433 1567 2447
rect 1633 2433 1647 2447
rect 1993 2433 2007 2447
rect 2213 2433 2227 2447
rect 2313 2433 2327 2447
rect 2773 2433 2787 2447
rect 2813 2433 2827 2447
rect 2893 2433 2907 2447
rect 3093 2433 3107 2447
rect 3153 2433 3167 2447
rect 3373 2433 3387 2447
rect 3613 2433 3627 2447
rect 3833 2433 3847 2447
rect 3873 2433 3887 2447
rect 4153 2433 4167 2447
rect 4193 2433 4207 2447
rect 4233 2433 4247 2447
rect 4533 2433 4547 2447
rect 4573 2433 4587 2447
rect 4613 2433 4627 2447
rect 4693 2433 4707 2447
rect 4733 2433 4747 2447
rect 4833 2433 4847 2447
rect 5113 2433 5127 2447
rect 5353 2433 5367 2447
rect 5393 2433 5407 2447
rect 5433 2433 5447 2447
rect 293 2413 307 2427
rect 1953 2413 1967 2427
rect 2953 2413 2967 2427
rect 3673 2413 3687 2427
rect 4373 2413 4387 2427
rect 5273 2413 5287 2427
rect 4513 2393 4527 2407
rect 1773 2273 1787 2287
rect 2293 2273 2307 2287
rect 3113 2273 3127 2287
rect 3193 2273 3207 2287
rect 4033 2273 4047 2287
rect 5233 2273 5247 2287
rect 5373 2273 5387 2287
rect 193 2253 207 2267
rect 253 2253 267 2267
rect 313 2253 327 2267
rect 553 2254 567 2268
rect 993 2253 1007 2267
rect 1033 2253 1047 2267
rect 1153 2253 1167 2267
rect 1193 2253 1207 2267
rect 1253 2253 1267 2267
rect 1293 2253 1307 2267
rect 1333 2253 1347 2267
rect 1553 2253 1567 2267
rect 1593 2253 1607 2267
rect 1873 2253 1887 2267
rect 1913 2253 1927 2267
rect 2213 2253 2227 2267
rect 2253 2253 2267 2267
rect 2513 2253 2527 2267
rect 2933 2253 2947 2267
rect 2973 2253 2987 2267
rect 3053 2253 3067 2267
rect 3533 2253 3547 2267
rect 3573 2253 3587 2267
rect 3653 2253 3667 2267
rect 3873 2253 3887 2267
rect 4393 2253 4407 2267
rect 4453 2253 4467 2267
rect 4493 2253 4507 2267
rect 4713 2253 4727 2267
rect 4773 2253 4787 2267
rect 4893 2253 4907 2267
rect 4933 2253 4947 2267
rect 4973 2253 4987 2267
rect 5193 2253 5207 2267
rect 33 2233 47 2247
rect 413 2233 427 2247
rect 553 2232 567 2246
rect 733 2233 747 2247
rect 793 2233 807 2247
rect 893 2233 907 2247
rect 1473 2233 1487 2247
rect 1733 2233 1747 2247
rect 1813 2233 1827 2247
rect 1993 2233 2007 2247
rect 2033 2233 2047 2247
rect 2373 2233 2387 2247
rect 2413 2233 2427 2247
rect 2593 2233 2607 2247
rect 2853 2233 2867 2247
rect 3173 2233 3187 2247
rect 3273 2233 3287 2247
rect 3313 2233 3327 2247
rect 3473 2233 3487 2247
rect 3793 2233 3807 2247
rect 3993 2233 4007 2247
rect 4133 2234 4147 2248
rect 4273 2233 4287 2247
rect 4313 2233 4327 2247
rect 4593 2233 4607 2247
rect 4633 2233 4647 2247
rect 5113 2233 5127 2247
rect 5293 2233 5307 2247
rect 5413 2233 5427 2247
rect 253 2213 267 2227
rect 293 2213 307 2227
rect 333 2213 347 2227
rect 393 2213 407 2227
rect 613 2213 627 2227
rect 813 2213 827 2227
rect 1013 2213 1027 2227
rect 1053 2213 1067 2227
rect 1273 2213 1287 2227
rect 1313 2213 1327 2227
rect 1433 2213 1447 2227
rect 1633 2213 1647 2227
rect 1853 2213 1867 2227
rect 2193 2213 2207 2227
rect 2233 2213 2247 2227
rect 2633 2213 2647 2227
rect 2813 2213 2827 2227
rect 3033 2213 3047 2227
rect 3073 2213 3087 2227
rect 3133 2213 3147 2227
rect 3513 2213 3527 2227
rect 3553 2213 3567 2227
rect 3633 2213 3647 2227
rect 3753 2213 3767 2227
rect 3913 2213 3927 2227
rect 4433 2213 4447 2227
rect 4473 2213 4487 2227
rect 4793 2213 4807 2227
rect 4913 2213 4927 2227
rect 4953 2213 4967 2227
rect 5073 2213 5087 2227
rect 5253 2213 5267 2227
rect 5353 2213 5367 2227
rect 53 2193 67 2207
rect 93 2193 107 2207
rect 433 2193 447 2207
rect 533 2193 547 2207
rect 773 2193 787 2207
rect 913 2193 927 2207
rect 953 2193 967 2207
rect 2413 2193 2427 2207
rect 2453 2193 2467 2207
rect 3393 2193 3407 2207
rect 3433 2193 3447 2207
rect 4093 2193 4107 2207
rect 4133 2193 4147 2207
rect 4213 2193 4227 2207
rect 4253 2193 4267 2207
rect 373 2173 387 2187
rect 833 2173 847 2187
rect 493 2153 507 2167
rect 3893 1993 3907 2007
rect 5393 1993 5407 2007
rect 273 1972 287 1986
rect 313 1973 327 1987
rect 2653 1973 2667 1987
rect 2853 1973 2867 1987
rect 2893 1973 2907 1987
rect 3313 1973 3327 1987
rect 3353 1973 3367 1987
rect 3933 1973 3947 1987
rect 5313 1973 5327 1987
rect 93 1953 107 1967
rect 653 1953 667 1967
rect 693 1953 707 1967
rect 773 1953 787 1967
rect 813 1953 827 1967
rect 833 1953 847 1967
rect 873 1953 887 1967
rect 893 1953 907 1967
rect 1073 1953 1087 1967
rect 1273 1953 1287 1967
rect 1493 1952 1507 1966
rect 1693 1953 1707 1967
rect 1853 1953 1867 1967
rect 1933 1953 1947 1967
rect 2093 1953 2107 1967
rect 2133 1953 2147 1967
rect 2473 1953 2487 1967
rect 2513 1953 2527 1967
rect 2613 1953 2627 1967
rect 2753 1953 2767 1967
rect 2793 1953 2807 1967
rect 2973 1953 2987 1967
rect 3013 1954 3027 1968
rect 3193 1953 3207 1967
rect 3493 1953 3507 1967
rect 3533 1953 3547 1967
rect 3573 1953 3587 1967
rect 3773 1953 3787 1967
rect 3813 1953 3827 1967
rect 3993 1953 4007 1967
rect 4113 1953 4127 1967
rect 4213 1953 4227 1967
rect 4253 1953 4267 1967
rect 4373 1953 4387 1967
rect 4413 1953 4427 1967
rect 4513 1953 4527 1967
rect 4673 1953 4687 1967
rect 4713 1953 4727 1967
rect 4833 1953 4847 1967
rect 4873 1953 4887 1967
rect 4973 1953 4987 1967
rect 5013 1953 5027 1967
rect 5053 1953 5067 1967
rect 5173 1954 5187 1968
rect 5433 1953 5447 1967
rect 5473 1953 5487 1967
rect 133 1933 147 1947
rect 273 1933 287 1947
rect 453 1933 467 1947
rect 493 1933 507 1947
rect 1033 1933 1047 1947
rect 1293 1933 1307 1947
rect 1533 1933 1547 1947
rect 1733 1933 1747 1947
rect 1893 1933 1907 1947
rect 1973 1933 1987 1947
rect 2273 1933 2287 1947
rect 2313 1933 2327 1947
rect 2853 1933 2867 1947
rect 3153 1933 3167 1947
rect 3293 1933 3307 1947
rect 3453 1933 3467 1947
rect 3653 1933 3667 1947
rect 3873 1933 3887 1947
rect 4033 1933 4047 1947
rect 4153 1933 4167 1947
rect 4553 1933 4567 1947
rect 4633 1933 4647 1947
rect 4753 1933 4767 1947
rect 5133 1933 5147 1947
rect 5373 1934 5387 1948
rect 213 1913 227 1927
rect 373 1913 387 1927
rect 633 1913 647 1927
rect 673 1913 687 1927
rect 713 1913 727 1927
rect 833 1913 847 1927
rect 913 1913 927 1927
rect 953 1913 967 1927
rect 1373 1913 1387 1927
rect 1613 1913 1627 1927
rect 1673 1913 1687 1927
rect 2153 1913 2167 1927
rect 2193 1913 2207 1927
rect 2453 1913 2467 1927
rect 2493 1913 2507 1927
rect 2593 1913 2607 1927
rect 2672 1913 2686 1927
rect 2693 1913 2707 1927
rect 2813 1913 2827 1927
rect 2953 1913 2967 1927
rect 3013 1914 3027 1928
rect 3073 1913 3087 1927
rect 3553 1913 3567 1927
rect 3593 1913 3607 1927
rect 3693 1913 3707 1927
rect 3753 1913 3767 1927
rect 3833 1913 3847 1927
rect 4233 1913 4247 1927
rect 4352 1913 4366 1927
rect 4373 1913 4387 1927
rect 4433 1913 4447 1927
rect 4473 1913 4487 1927
rect 4813 1913 4827 1927
rect 4853 1913 4867 1927
rect 4893 1913 4907 1927
rect 5033 1913 5047 1927
rect 5173 1913 5187 1927
rect 5413 1913 5427 1927
rect 5453 1913 5467 1927
rect 1713 1893 1727 1907
rect 1953 1893 1967 1907
rect 2053 1893 2067 1907
rect 3513 1893 3527 1907
rect 4093 1893 4107 1907
rect 4173 1893 4187 1907
rect 4773 1892 4787 1906
rect 5133 1893 5147 1907
rect 4573 1873 4587 1887
rect 2913 1773 2927 1787
rect 1553 1753 1567 1767
rect 1733 1753 1747 1767
rect 1773 1753 1787 1767
rect 1913 1753 1927 1767
rect 3773 1773 3787 1787
rect 213 1733 227 1747
rect 93 1713 107 1727
rect 133 1713 147 1727
rect 292 1733 306 1747
rect 313 1733 327 1747
rect 373 1733 387 1747
rect 433 1733 447 1747
rect 533 1733 547 1747
rect 793 1733 807 1747
rect 873 1733 887 1747
rect 1133 1733 1147 1747
rect 1193 1733 1207 1747
rect 1233 1733 1247 1747
rect 1373 1733 1387 1747
rect 1633 1733 1647 1747
rect 1873 1733 1887 1747
rect 2073 1733 2087 1747
rect 2153 1733 2167 1747
rect 2193 1734 2207 1748
rect 3153 1753 3167 1767
rect 4053 1753 4067 1767
rect 4433 1753 4447 1767
rect 5073 1753 5087 1767
rect 2393 1733 2407 1747
rect 2693 1733 2707 1747
rect 2733 1733 2747 1747
rect 2773 1733 2787 1747
rect 2853 1733 2867 1747
rect 3053 1733 3067 1747
rect 3093 1733 3107 1747
rect 3293 1733 3307 1747
rect 3333 1734 3347 1748
rect 3393 1733 3407 1747
rect 3433 1733 3447 1747
rect 3473 1733 3487 1747
rect 3853 1733 3867 1747
rect 3973 1733 3987 1747
rect 4013 1733 4027 1747
rect 4133 1733 4147 1747
rect 4173 1733 4187 1747
rect 4273 1733 4287 1747
rect 4553 1733 4567 1747
rect 4713 1733 4727 1747
rect 4753 1733 4767 1747
rect 5173 1733 5187 1747
rect 5253 1733 5267 1747
rect 5313 1733 5327 1747
rect 713 1713 727 1727
rect 1013 1713 1027 1727
rect 1053 1713 1067 1727
rect 1473 1713 1487 1727
rect 1693 1713 1707 1727
rect 1793 1713 1807 1727
rect 1993 1713 2007 1727
rect 2253 1713 2267 1727
rect 2473 1713 2487 1727
rect 3173 1713 3187 1727
rect 3553 1713 3567 1727
rect 3753 1713 3767 1727
rect 4393 1713 4407 1727
rect 4453 1713 4467 1727
rect 4653 1713 4667 1727
rect 4793 1713 4807 1727
rect 4893 1713 4907 1727
rect 5093 1713 5107 1727
rect 5393 1713 5407 1727
rect 313 1693 327 1707
rect 353 1693 367 1707
rect 453 1693 467 1707
rect 553 1693 567 1707
rect 673 1693 687 1707
rect 893 1693 907 1707
rect 1213 1693 1227 1707
rect 1253 1693 1267 1707
rect 1353 1693 1367 1707
rect 1413 1693 1427 1707
rect 1513 1693 1527 1707
rect 1613 1693 1627 1707
rect 1753 1693 1767 1707
rect 1893 1693 1907 1707
rect 1953 1693 1967 1707
rect 2093 1693 2107 1707
rect 2133 1693 2147 1707
rect 2513 1693 2527 1707
rect 2613 1693 2627 1707
rect 2713 1693 2727 1707
rect 2793 1693 2807 1707
rect 2833 1693 2847 1707
rect 2913 1693 2927 1707
rect 3013 1693 3027 1707
rect 3093 1692 3107 1706
rect 3133 1693 3147 1707
rect 3273 1693 3287 1707
rect 3593 1693 3607 1707
rect 3713 1693 3727 1707
rect 3833 1693 3847 1707
rect 3873 1693 3887 1707
rect 4073 1693 4087 1707
rect 4113 1693 4127 1707
rect 4253 1693 4267 1707
rect 4293 1693 4307 1707
rect 4353 1693 4367 1707
rect 4493 1693 4507 1707
rect 4693 1693 4707 1707
rect 4733 1692 4747 1706
rect 5133 1693 5147 1707
rect 5233 1692 5247 1706
rect 5273 1693 5287 1707
rect 5433 1693 5447 1707
rect 253 1672 267 1686
rect 2173 1673 2187 1687
rect 2293 1673 2307 1687
rect 2333 1673 2347 1687
rect 4033 1673 4047 1687
rect 4573 1673 4587 1687
rect 4613 1673 4627 1687
rect 4833 1673 4847 1687
rect 4873 1673 4887 1687
rect 4953 1673 4967 1687
rect 4993 1673 5007 1687
rect 1373 1653 1387 1667
rect 1413 1653 1427 1667
rect 1713 1473 1727 1487
rect 353 1453 367 1467
rect 393 1453 407 1467
rect 1373 1453 1387 1467
rect 1413 1453 1427 1467
rect 1813 1453 1827 1467
rect 2373 1452 2387 1466
rect 2413 1453 2427 1467
rect 3253 1453 3267 1467
rect 3293 1453 3307 1467
rect 4873 1453 4887 1467
rect 4913 1453 4927 1467
rect 5193 1453 5207 1467
rect 5233 1453 5247 1467
rect 93 1433 107 1447
rect 133 1433 147 1447
rect 273 1433 287 1447
rect 493 1433 507 1447
rect 593 1433 607 1447
rect 693 1433 707 1447
rect 733 1433 747 1447
rect 993 1433 1007 1447
rect 1233 1433 1247 1447
rect 1273 1433 1287 1447
rect 1493 1433 1507 1447
rect 1533 1433 1547 1447
rect 1613 1433 1627 1447
rect 1733 1433 1747 1447
rect 1853 1433 1867 1447
rect 1893 1434 1907 1448
rect 2013 1433 2027 1447
rect 2153 1433 2167 1447
rect 2473 1433 2487 1447
rect 2513 1433 2527 1447
rect 2573 1433 2587 1447
rect 2653 1433 2667 1447
rect 2773 1433 2787 1447
rect 2993 1433 3007 1447
rect 3213 1433 3227 1447
rect 3333 1433 3347 1447
rect 3493 1433 3507 1447
rect 3533 1433 3547 1447
rect 3573 1433 3587 1447
rect 3713 1433 3727 1447
rect 3813 1433 3827 1447
rect 4213 1433 4227 1447
rect 4413 1433 4427 1447
rect 4453 1433 4467 1447
rect 4593 1433 4607 1447
rect 4693 1433 4707 1447
rect 4733 1433 4747 1447
rect 5073 1433 5087 1447
rect 5273 1432 5287 1446
rect 5373 1433 5387 1447
rect 233 1413 247 1427
rect 353 1413 367 1427
rect 453 1413 467 1427
rect 553 1412 567 1426
rect 853 1413 867 1427
rect 893 1413 907 1427
rect 953 1413 967 1427
rect 1033 1413 1047 1427
rect 1113 1413 1127 1427
rect 1153 1413 1167 1427
rect 1313 1413 1327 1427
rect 1573 1413 1587 1427
rect 1753 1413 1767 1427
rect 1973 1413 1987 1427
rect 2193 1413 2207 1427
rect 2353 1413 2367 1427
rect 2813 1413 2827 1427
rect 3013 1413 3027 1427
rect 3253 1413 3267 1427
rect 3413 1413 3427 1427
rect 3753 1413 3767 1427
rect 3953 1413 3967 1427
rect 4113 1413 4127 1427
rect 4253 1413 4267 1427
rect 4553 1413 4567 1427
rect 4653 1413 4667 1427
rect 4813 1413 4827 1427
rect 4893 1413 4907 1427
rect 5033 1413 5047 1427
rect 5193 1412 5207 1426
rect 73 1393 87 1407
rect 113 1393 127 1407
rect 153 1393 167 1407
rect 673 1393 687 1407
rect 713 1393 727 1407
rect 813 1393 827 1407
rect 1213 1393 1227 1407
rect 1353 1393 1367 1407
rect 1473 1393 1487 1407
rect 1513 1393 1527 1407
rect 1713 1393 1727 1407
rect 1873 1393 1887 1407
rect 1933 1392 1947 1406
rect 2053 1393 2067 1407
rect 2273 1393 2287 1407
rect 2453 1393 2467 1407
rect 2493 1393 2507 1407
rect 2533 1393 2547 1407
rect 2673 1393 2687 1407
rect 2753 1393 2767 1407
rect 2853 1393 2867 1407
rect 3093 1393 3107 1407
rect 3213 1393 3227 1407
rect 3513 1393 3527 1407
rect 3553 1393 3567 1407
rect 3653 1393 3667 1407
rect 3833 1393 3847 1407
rect 4373 1393 4387 1407
rect 4433 1393 4447 1407
rect 4753 1393 4767 1407
rect 4953 1393 4967 1407
rect 5313 1393 5327 1407
rect 333 1373 347 1387
rect 533 1373 547 1387
rect 633 1373 647 1387
rect 913 1373 927 1387
rect 1093 1373 1107 1387
rect 1133 1373 1147 1387
rect 3453 1373 3467 1387
rect 3693 1373 3707 1387
rect 4333 1373 4347 1387
rect 4632 1373 4646 1387
rect 4653 1373 4667 1387
rect 5413 1372 5427 1386
rect 2053 1233 2067 1247
rect 2733 1233 2747 1247
rect 4733 1233 4747 1247
rect 4853 1233 4867 1247
rect 73 1213 87 1227
rect 113 1213 127 1227
rect 373 1213 387 1227
rect 413 1213 427 1227
rect 573 1213 587 1227
rect 633 1213 647 1227
rect 673 1213 687 1227
rect 753 1213 767 1227
rect 1013 1213 1027 1227
rect 1133 1213 1147 1227
rect 1173 1213 1187 1227
rect 1413 1213 1427 1227
rect 1453 1213 1467 1227
rect 1793 1213 1807 1227
rect 193 1193 207 1207
rect 233 1193 247 1207
rect 493 1192 507 1206
rect 833 1193 847 1207
rect 1053 1193 1067 1207
rect 1253 1193 1267 1207
rect 1293 1193 1307 1207
rect 1533 1193 1547 1207
rect 1713 1193 1727 1207
rect 53 1173 67 1187
rect 393 1173 407 1187
rect 433 1173 447 1187
rect 613 1173 627 1187
rect 653 1173 667 1187
rect 693 1173 707 1187
rect 873 1173 887 1187
rect 1113 1173 1127 1187
rect 1433 1173 1447 1187
rect 1473 1173 1487 1187
rect 1813 1173 1827 1187
rect 1853 1173 1867 1187
rect 1933 1213 1947 1227
rect 2173 1213 2187 1227
rect 2253 1214 2267 1228
rect 2313 1213 2327 1227
rect 2393 1213 2407 1227
rect 2713 1213 2727 1227
rect 2813 1213 2827 1227
rect 3493 1213 3507 1227
rect 3553 1213 3567 1227
rect 3593 1213 3607 1227
rect 3813 1213 3827 1227
rect 3933 1213 3947 1227
rect 4013 1213 4027 1227
rect 4113 1213 4127 1227
rect 4153 1213 4167 1227
rect 4273 1213 4287 1227
rect 4333 1213 4347 1227
rect 4433 1213 4447 1227
rect 4493 1213 4507 1227
rect 4593 1213 4607 1227
rect 4633 1213 4647 1227
rect 4893 1213 4907 1227
rect 5013 1213 5027 1227
rect 5073 1213 5087 1227
rect 5193 1213 5207 1227
rect 5473 1213 5487 1227
rect 2013 1193 2027 1207
rect 2113 1193 2127 1207
rect 2273 1192 2287 1206
rect 2473 1193 2487 1207
rect 2613 1193 2627 1207
rect 2873 1192 2887 1206
rect 3033 1193 3047 1207
rect 3133 1193 3147 1207
rect 3293 1193 3307 1207
rect 3453 1193 3467 1207
rect 3673 1193 3687 1207
rect 4073 1193 4087 1207
rect 4233 1193 4247 1207
rect 4693 1193 4707 1207
rect 4813 1193 4827 1207
rect 4833 1193 4847 1207
rect 1913 1172 1927 1186
rect 1973 1173 1987 1187
rect 2073 1173 2087 1187
rect 2193 1172 2207 1186
rect 2233 1173 2247 1187
rect 2513 1173 2527 1187
rect 2693 1173 2707 1187
rect 2793 1173 2807 1187
rect 2833 1173 2847 1187
rect 3493 1173 3507 1187
rect 3533 1173 3547 1187
rect 3713 1173 3727 1187
rect 3873 1173 3887 1187
rect 3913 1173 3927 1187
rect 4033 1173 4047 1187
rect 4133 1173 4147 1187
rect 4173 1173 4187 1187
rect 4353 1173 4367 1187
rect 4473 1173 4487 1187
rect 4533 1173 4547 1187
rect 4573 1173 4587 1187
rect 4653 1172 4667 1186
rect 4773 1173 4787 1187
rect 4953 1173 4967 1187
rect 5033 1173 5047 1187
rect 5093 1173 5107 1187
rect 5393 1193 5407 1207
rect 5353 1173 5367 1187
rect 513 1153 527 1167
rect 553 1153 567 1167
rect 3373 1153 3387 1167
rect 3433 1153 3447 1167
rect 5213 1153 5227 1167
rect 2253 1133 2267 1147
rect 2313 1133 2327 1147
rect 5253 1133 5267 1147
rect 2633 953 2647 967
rect 853 933 867 947
rect 893 933 907 947
rect 1053 933 1067 947
rect 1093 933 1107 947
rect 1613 933 1627 947
rect 1653 933 1667 947
rect 1713 933 1727 947
rect 1753 933 1767 947
rect 1833 933 1847 947
rect 1873 933 1887 947
rect 2213 933 2227 947
rect 2253 933 2267 947
rect 2333 933 2347 947
rect 2373 933 2387 947
rect 2593 933 2607 947
rect 4273 933 4287 947
rect 4313 933 4327 947
rect 4593 933 4607 947
rect 4653 933 4667 947
rect 5293 933 5307 947
rect 5433 933 5447 947
rect 5473 933 5487 947
rect 113 913 127 927
rect 373 913 387 927
rect 393 913 407 927
rect 473 912 487 926
rect 513 913 527 927
rect 653 913 667 927
rect 733 913 747 927
rect 773 913 787 927
rect 1013 913 1027 927
rect 1173 913 1187 927
rect 1273 913 1287 927
rect 1313 913 1327 927
rect 1413 913 1427 927
rect 1453 913 1467 927
rect 1493 913 1507 927
rect 1953 913 1967 927
rect 2133 913 2147 927
rect 2173 913 2187 927
rect 2473 913 2487 927
rect 2513 913 2527 927
rect 2733 914 2747 928
rect 2913 913 2927 927
rect 2953 913 2967 927
rect 2993 913 3007 927
rect 3213 913 3227 927
rect 3253 913 3267 927
rect 3413 913 3427 927
rect 3553 913 3567 927
rect 3773 913 3787 927
rect 3933 913 3947 927
rect 3973 913 3987 927
rect 4113 913 4127 927
rect 4153 913 4167 927
rect 4493 913 4507 927
rect 4753 913 4767 927
rect 4793 913 4807 927
rect 4873 913 4887 927
rect 4913 913 4927 927
rect 4993 913 5007 927
rect 5033 913 5047 927
rect 5133 913 5147 927
rect 5173 913 5187 927
rect 5233 913 5247 927
rect 133 893 147 907
rect 253 893 267 907
rect 613 893 627 907
rect 813 893 827 907
rect 953 893 967 907
rect 1073 893 1087 907
rect 1613 893 1627 907
rect 1813 893 1827 907
rect 1853 893 1867 907
rect 2013 893 2027 907
rect 2313 893 2327 907
rect 2413 893 2427 907
rect 2553 893 2567 907
rect 2773 893 2787 907
rect 213 873 227 887
rect 373 873 387 887
rect 453 873 467 887
rect 493 873 507 887
rect 713 873 727 887
rect 753 873 767 887
rect 1193 873 1207 887
rect 1253 873 1267 887
rect 1293 873 1307 887
rect 1433 873 1447 887
rect 1473 873 1487 887
rect 1573 873 1587 887
rect 1973 873 1987 887
rect 2053 873 2067 887
rect 2153 873 2167 887
rect 2453 873 2467 887
rect 2573 873 2587 887
rect 2853 873 2867 887
rect 253 853 267 867
rect 593 853 607 867
rect 893 853 907 867
rect 973 853 987 867
rect 3093 893 3107 907
rect 3393 893 3407 907
rect 3593 893 3607 907
rect 3733 893 3747 907
rect 4013 893 4027 907
rect 4293 893 4307 907
rect 4453 893 4467 907
rect 4713 894 4727 908
rect 5273 893 5287 907
rect 5413 893 5427 907
rect 2933 873 2947 887
rect 2973 873 2987 887
rect 3013 873 3027 887
rect 3153 873 3167 887
rect 3233 873 3247 887
rect 3273 873 3287 887
rect 3313 873 3327 887
rect 3533 873 3547 887
rect 3653 873 3667 887
rect 3893 873 3907 887
rect 3953 873 3967 887
rect 4093 873 4107 887
rect 4373 873 4387 887
rect 2893 852 2907 866
rect 4713 872 4727 886
rect 4813 873 4827 887
rect 4873 873 4887 887
rect 4933 873 4947 887
rect 5013 873 5027 887
rect 5053 873 5067 887
rect 5113 872 5127 886
rect 5193 873 5207 887
rect 5353 873 5367 887
rect 4173 853 4187 867
rect 5233 853 5247 867
rect 5353 833 5367 847
rect 153 713 167 727
rect 253 712 267 726
rect 1193 713 1207 727
rect 2093 713 2107 727
rect 3173 713 3187 727
rect 273 693 287 707
rect 333 693 347 707
rect 433 693 447 707
rect 893 693 907 707
rect 933 693 947 707
rect 993 693 1007 707
rect 1513 693 1527 707
rect 1553 693 1567 707
rect 1633 693 1647 707
rect 1733 693 1747 707
rect 1913 693 1927 707
rect 2133 693 2147 707
rect 2233 693 2247 707
rect 2293 693 2307 707
rect 2393 693 2407 707
rect 2433 693 2447 707
rect 2693 693 2707 707
rect 3253 693 3267 707
rect 3293 693 3307 707
rect 3453 693 3467 707
rect 3773 693 3787 707
rect 3813 693 3827 707
rect 3873 693 3887 707
rect 3913 693 3927 707
rect 3973 693 3987 707
rect 4093 693 4107 707
rect 4233 694 4247 708
rect 4273 693 4287 707
rect 4413 693 4427 707
rect 4453 693 4467 707
rect 4693 693 4707 707
rect 4733 693 4747 707
rect 4773 693 4787 707
rect 4813 693 4827 707
rect 4913 693 4927 707
rect 4993 693 5007 707
rect 5093 693 5107 707
rect 5353 693 5367 707
rect 5393 693 5407 707
rect 73 673 87 687
rect 113 673 127 687
rect 213 673 227 687
rect 513 673 527 687
rect 613 673 627 687
rect 693 673 707 687
rect 833 673 847 687
rect 1153 674 1167 688
rect 1273 673 1287 687
rect 1313 673 1327 687
rect 1433 673 1447 687
rect 1653 673 1667 687
rect 1833 673 1847 687
rect 1973 673 1987 687
rect 2053 673 2067 687
rect 2333 673 2347 687
rect 2613 673 2627 687
rect 2753 674 2767 688
rect 2953 673 2967 687
rect 3033 673 3047 687
rect 3113 673 3127 687
rect 3373 673 3387 687
rect 3533 673 3547 687
rect 3753 673 3767 687
rect 3793 673 3807 687
rect 4073 673 4087 687
rect 4353 673 4367 687
rect 4533 673 4547 687
rect 5033 673 5047 687
rect 5173 673 5187 687
rect 5213 673 5227 687
rect 173 653 187 667
rect 313 653 327 667
rect 353 653 367 667
rect 413 653 427 667
rect 873 653 887 667
rect 913 653 927 667
rect 1053 653 1067 667
rect 1473 653 1487 667
rect 1573 653 1587 667
rect 1613 653 1627 667
rect 1933 653 1947 667
rect 2013 653 2027 667
rect 2153 653 2167 667
rect 2193 653 2207 667
rect 2413 653 2427 667
rect 2453 653 2467 667
rect 2573 653 2587 667
rect 2913 653 2927 667
rect 3173 653 3187 667
rect 3233 653 3247 667
rect 3273 653 3287 667
rect 3313 653 3327 667
rect 3553 653 3567 667
rect 3573 653 3587 667
rect 3853 653 3867 667
rect 3893 653 3907 667
rect 3993 653 4007 667
rect 4033 653 4047 667
rect 4253 653 4267 667
rect 4293 653 4307 667
rect 4573 653 4587 667
rect 4713 653 4727 667
rect 4753 653 4767 667
rect 4893 653 4907 667
rect 4973 653 4987 667
rect 5373 652 5387 666
rect 5413 653 5427 667
rect 533 633 547 647
rect 573 633 587 647
rect 633 633 647 647
rect 673 633 687 647
rect 733 633 747 647
rect 773 633 787 647
rect 1113 633 1127 647
rect 1153 633 1167 647
rect 1713 633 1727 647
rect 2753 633 2767 647
rect 2793 633 2807 647
rect 3413 633 3427 647
rect 3673 633 3687 647
rect 3753 633 3767 647
rect 1613 593 1627 607
rect 4073 632 4087 646
rect 4153 633 4167 647
rect 3353 613 3367 627
rect 873 413 887 427
rect 953 413 967 427
rect 1373 413 1387 427
rect 1433 413 1447 427
rect 1713 413 1727 427
rect 1773 413 1787 427
rect 1933 413 1947 427
rect 2013 413 2027 427
rect 4553 413 4567 427
rect 4593 413 4607 427
rect 4873 413 4887 427
rect 4913 413 4927 427
rect 93 393 107 407
rect 553 393 567 407
rect 593 393 607 407
rect 713 393 727 407
rect 1033 393 1047 407
rect 1073 393 1087 407
rect 1193 393 1207 407
rect 1553 393 1567 407
rect 1853 393 1867 407
rect 1893 393 1907 407
rect 2093 393 2107 407
rect 2133 393 2147 407
rect 2253 393 2267 407
rect 2293 393 2307 407
rect 2333 393 2347 407
rect 2493 393 2507 407
rect 2713 393 2727 407
rect 2753 393 2767 407
rect 2953 393 2967 407
rect 3093 393 3107 407
rect 3193 393 3207 407
rect 3233 393 3247 407
rect 3333 393 3347 407
rect 3373 393 3387 407
rect 3473 393 3487 407
rect 3593 393 3607 407
rect 3813 393 3827 407
rect 3933 393 3947 407
rect 4153 393 4167 407
rect 4193 392 4207 406
rect 4653 393 4667 407
rect 4773 393 4787 407
rect 4813 393 4827 407
rect 5013 393 5027 407
rect 5093 393 5107 407
rect 5153 393 5167 407
rect 5193 393 5207 407
rect 5273 393 5287 407
rect 5373 393 5387 407
rect 133 373 147 387
rect 353 373 367 387
rect 393 373 407 387
rect 753 373 767 387
rect 913 373 927 387
rect 1233 373 1247 387
rect 1353 373 1367 387
rect 1593 373 1607 387
rect 1733 373 1747 387
rect 1953 373 1967 387
rect 2533 373 2547 387
rect 2813 373 2827 387
rect 2893 373 2907 387
rect 2993 373 3007 387
rect 3633 373 3647 387
rect 3973 373 3987 387
rect 4333 373 4347 387
rect 4413 373 4427 387
rect 4573 373 4587 387
rect 4873 373 4887 387
rect 5433 373 5447 387
rect 213 353 227 367
rect 273 353 287 367
rect 533 353 547 367
rect 573 353 587 367
rect 833 353 847 367
rect 1013 353 1027 367
rect 1093 353 1107 367
rect 1313 353 1327 367
rect 1673 353 1687 367
rect 1793 353 1807 367
rect 1913 353 1927 367
rect 2073 353 2087 367
rect 2113 353 2127 367
rect 2153 353 2167 367
rect 2273 353 2287 367
rect 2313 353 2327 367
rect 2393 353 2407 367
rect 2613 353 2627 367
rect 2693 353 2707 367
rect 2733 352 2747 366
rect 2773 353 2787 367
rect 3073 353 3087 367
rect 3173 353 3187 367
rect 3213 353 3227 367
rect 3253 353 3267 367
rect 3393 354 3407 368
rect 3493 353 3507 367
rect 3713 353 3727 367
rect 3793 353 3807 367
rect 4053 353 4067 367
rect 4133 353 4147 367
rect 4213 353 4227 367
rect 4293 353 4307 367
rect 4453 353 4467 367
rect 4613 353 4627 367
rect 4733 353 4747 367
rect 4833 353 4847 367
rect 4993 353 5007 367
rect 5033 353 5047 367
rect 5173 353 5187 367
rect 5213 353 5227 367
rect 5253 353 5267 367
rect 5353 353 5367 367
rect 5473 353 5487 367
rect 2973 333 2987 347
rect 4933 293 4947 307
rect 4973 294 4987 308
rect 253 193 267 207
rect 393 193 407 207
rect 2093 193 2107 207
rect 3593 194 3607 208
rect 4793 193 4807 207
rect 73 173 87 187
rect 293 173 307 187
rect 453 173 467 187
rect 553 173 567 187
rect 593 173 607 187
rect 733 173 747 187
rect 773 173 787 187
rect 853 173 867 187
rect 893 173 907 187
rect 1333 173 1347 187
rect 1413 173 1427 187
rect 1633 173 1647 187
rect 1873 173 1887 187
rect 1953 173 1967 187
rect 1993 173 2007 187
rect 2033 173 2047 187
rect 2193 173 2207 187
rect 2413 173 2427 187
rect 2493 173 2507 187
rect 2733 173 2747 187
rect 2833 173 2847 187
rect 2973 173 2987 187
rect 3013 173 3027 187
rect 3073 173 3087 187
rect 3213 173 3227 187
rect 3253 173 3267 187
rect 3353 173 3367 187
rect 3453 173 3467 187
rect 3553 173 3567 187
rect 3673 173 3687 187
rect 3793 173 3807 187
rect 3933 173 3947 187
rect 4413 173 4427 187
rect 4633 173 4647 187
rect 4733 173 4747 187
rect 5013 173 5027 187
rect 5253 173 5267 187
rect 5333 173 5347 187
rect 113 153 127 167
rect 233 153 247 167
rect 333 153 347 167
rect 1013 153 1027 167
rect 1193 153 1207 167
rect 1253 153 1267 167
rect 1553 153 1567 167
rect 1793 153 1807 167
rect 2113 153 2127 167
rect 2273 153 2287 167
rect 2653 153 2667 167
rect 2913 153 2927 167
rect 3153 153 3167 167
rect 3293 153 3307 167
rect 3393 153 3407 167
rect 3633 153 3647 167
rect 3833 153 3847 167
rect 4013 153 4027 167
rect 4153 153 4167 167
rect 4313 153 4327 167
rect 4493 153 4507 167
rect 4813 153 4827 167
rect 4933 153 4947 167
rect 5093 153 5107 167
rect 5133 153 5147 167
rect 5513 153 5527 167
rect 53 133 67 147
rect 273 133 287 147
rect 413 133 427 147
rect 473 133 487 147
rect 513 133 527 147
rect 673 133 687 147
rect 753 133 767 147
rect 793 133 807 147
rect 833 133 847 147
rect 953 133 967 147
rect 993 133 1007 147
rect 1353 133 1367 147
rect 1393 133 1407 147
rect 1513 133 1527 147
rect 1753 133 1767 147
rect 1973 133 1987 147
rect 2013 133 2027 147
rect 2153 133 2167 147
rect 2313 133 2327 147
rect 2473 133 2487 147
rect 2513 133 2527 147
rect 2613 133 2627 147
rect 2953 133 2967 147
rect 2993 133 3007 147
rect 3193 133 3207 147
rect 3233 133 3247 147
rect 3533 133 3547 147
rect 3593 133 3607 147
rect 3733 133 3747 147
rect 3773 133 3787 147
rect 4053 133 4067 147
rect 4533 133 4547 147
rect 4673 133 4687 147
rect 4713 133 4727 147
rect 4873 133 4887 147
rect 4973 133 4987 147
rect 1073 113 1087 127
rect 1133 113 1147 127
rect 1173 113 1187 127
rect 1213 113 1227 127
rect 1253 113 1267 127
rect 3833 113 3847 127
rect 3873 113 3887 127
rect 4173 113 4187 127
rect 4233 113 4247 127
rect 4333 113 4347 127
rect 4373 113 4387 127
rect 4913 113 4927 127
rect 5373 113 5387 127
rect 5413 113 5427 127
rect 973 93 987 107
rect 4973 93 4987 107
<< metal2 >>
rect 2516 5516 2543 5523
rect 96 5387 103 5413
rect 36 5147 43 5373
rect 116 5347 123 5373
rect 193 5367 207 5373
rect 87 5333 93 5347
rect 227 5333 233 5347
rect 176 5287 183 5313
rect 256 5307 263 5413
rect 396 5387 403 5433
rect 307 5333 313 5347
rect 247 5293 253 5307
rect 336 5227 343 5373
rect 367 5333 373 5347
rect 396 5307 403 5373
rect 413 5327 427 5333
rect 53 5087 67 5093
rect 96 5087 103 5133
rect 296 5087 303 5153
rect 247 5073 253 5087
rect 113 5047 127 5053
rect 76 4863 83 5033
rect 76 4856 93 4863
rect 127 4854 133 4867
rect 120 4853 140 4854
rect 93 4847 107 4853
rect 113 4827 127 4832
rect 76 4587 83 4793
rect 156 4787 163 5013
rect 196 4867 203 5073
rect 227 5033 233 5047
rect 173 4827 187 4833
rect 236 4827 243 4853
rect 296 4847 303 5033
rect 313 5027 327 5033
rect 336 4927 343 5093
rect 396 5047 403 5133
rect 416 5087 423 5213
rect 476 5147 483 5353
rect 516 5347 523 5373
rect 596 5327 603 5353
rect 636 5327 643 5393
rect 753 5367 767 5373
rect 767 5353 773 5367
rect 813 5347 827 5353
rect 587 5316 603 5327
rect 587 5313 600 5316
rect 536 5267 543 5313
rect 496 5127 503 5213
rect 616 5127 623 5153
rect 616 5113 633 5127
rect 567 5103 580 5107
rect 567 5093 583 5103
rect 507 5073 513 5087
rect 427 5033 433 5047
rect 456 5007 463 5073
rect 576 5067 583 5093
rect 533 5047 547 5053
rect 147 4773 153 4787
rect 176 4687 183 4813
rect 316 4747 323 4853
rect 516 4847 523 4913
rect 367 4833 373 4847
rect 407 4813 413 4827
rect 453 4807 467 4813
rect 516 4803 523 4833
rect 556 4827 563 4853
rect 576 4827 583 5053
rect 616 4943 623 5113
rect 656 5088 663 5273
rect 676 5187 683 5333
rect 696 5143 703 5333
rect 736 5267 743 5313
rect 736 5147 743 5253
rect 776 5203 783 5313
rect 876 5247 883 5373
rect 893 5347 907 5353
rect 916 5227 923 5373
rect 1013 5347 1027 5353
rect 776 5196 793 5203
rect 696 5140 723 5143
rect 696 5136 727 5140
rect 713 5127 727 5136
rect 796 5107 803 5193
rect 767 5093 773 5107
rect 640 5084 653 5087
rect 596 4936 623 4943
rect 636 5074 653 5084
rect 636 5073 660 5074
rect 596 4847 603 4936
rect 636 4887 643 5073
rect 660 5066 673 5067
rect 667 5054 673 5066
rect 667 5053 680 5054
rect 676 4903 683 5032
rect 696 5027 703 5093
rect 716 5007 723 5053
rect 836 5023 843 5133
rect 916 5127 923 5213
rect 856 5047 863 5093
rect 876 5067 883 5113
rect 896 5027 903 5093
rect 836 5016 863 5023
rect 676 4896 703 4903
rect 653 4827 667 4833
rect 547 4816 563 4827
rect 547 4813 560 4816
rect 516 4796 543 4803
rect 153 4587 167 4593
rect 216 4587 223 4613
rect 356 4587 363 4793
rect 416 4727 423 4773
rect 127 4583 140 4587
rect 127 4576 153 4583
rect 127 4573 140 4576
rect 76 4547 83 4573
rect 187 4554 193 4567
rect 253 4567 267 4573
rect 476 4567 483 4613
rect 187 4553 200 4554
rect 173 4547 187 4553
rect 96 4383 103 4533
rect 196 4507 203 4532
rect 236 4527 243 4553
rect 76 4376 103 4383
rect 76 4287 83 4376
rect 96 4327 103 4353
rect 136 4287 143 4313
rect 127 4273 143 4287
rect 56 4067 63 4273
rect 107 4053 113 4067
rect 56 3827 63 3993
rect 116 3967 123 4013
rect 136 4007 143 4273
rect 156 3987 163 4273
rect 196 4087 203 4493
rect 213 4307 227 4313
rect 236 4307 243 4513
rect 256 4267 263 4553
rect 316 4507 323 4553
rect 436 4527 443 4553
rect 347 4513 352 4527
rect 376 4387 383 4513
rect 476 4388 483 4553
rect 516 4527 523 4653
rect 536 4527 543 4796
rect 576 4787 583 4813
rect 567 4776 583 4787
rect 567 4773 580 4776
rect 696 4647 703 4896
rect 736 4827 743 4853
rect 756 4827 763 5013
rect 776 4867 783 4933
rect 816 4867 823 4913
rect 856 4867 863 5016
rect 936 4987 943 5333
rect 1047 5313 1053 5327
rect 993 5307 1007 5313
rect 996 5108 1003 5293
rect 1076 5147 1083 5433
rect 2053 5387 2067 5393
rect 1627 5373 1633 5387
rect 1787 5383 1800 5387
rect 1787 5373 1803 5383
rect 2107 5374 2113 5387
rect 2107 5373 2120 5374
rect 1113 5367 1127 5373
rect 1140 5363 1153 5367
rect 1136 5353 1153 5363
rect 807 4813 813 4827
rect 756 4787 763 4813
rect 596 4567 603 4593
rect 673 4567 687 4573
rect 647 4553 653 4567
rect 627 4513 633 4527
rect 316 4267 323 4373
rect 356 4328 363 4353
rect 436 4347 443 4373
rect 473 4347 487 4352
rect 436 4307 443 4333
rect 347 4306 360 4307
rect 347 4293 353 4306
rect 468 4293 473 4307
rect 567 4293 573 4307
rect 233 4067 247 4073
rect 173 4047 187 4053
rect 180 4023 193 4027
rect 176 4013 193 4023
rect 176 3967 183 4013
rect 216 3987 223 4033
rect 76 3787 83 3833
rect 233 3828 247 3833
rect 107 3813 113 3827
rect 127 3773 133 3787
rect 76 3667 83 3773
rect 16 3527 23 3613
rect 36 3307 43 3473
rect 56 3407 63 3553
rect 96 3527 103 3553
rect 136 3527 143 3773
rect 153 3767 167 3773
rect 176 3567 183 3813
rect 196 3727 203 3793
rect 213 3767 227 3773
rect 236 3747 243 3792
rect 276 3703 283 4073
rect 316 4047 323 4073
rect 336 4007 343 4253
rect 336 3867 343 3993
rect 356 3827 363 4053
rect 347 3816 363 3827
rect 347 3813 360 3816
rect 333 3807 347 3813
rect 316 3727 323 3773
rect 353 3767 367 3773
rect 276 3696 303 3703
rect 207 3554 213 3567
rect 207 3553 220 3554
rect 213 3528 227 3532
rect 133 3507 147 3513
rect 133 3500 134 3507
rect 126 3493 127 3500
rect 220 3506 233 3507
rect 113 3487 127 3493
rect 227 3493 233 3506
rect 67 3254 73 3267
rect 133 3267 147 3273
rect 60 3253 80 3254
rect 16 3187 23 3253
rect 93 3247 107 3253
rect 16 3028 23 3113
rect 16 2907 23 2992
rect 36 2787 43 3013
rect 56 3008 63 3232
rect 156 3127 163 3293
rect 216 3227 223 3293
rect 256 3227 263 3533
rect 296 3487 303 3696
rect 316 3607 323 3713
rect 376 3647 383 4273
rect 316 3527 323 3553
rect 353 3493 354 3500
rect 336 3443 343 3493
rect 353 3487 367 3493
rect 376 3467 383 3593
rect 336 3436 363 3443
rect 296 3287 303 3333
rect 356 3267 363 3436
rect 396 3403 403 4033
rect 436 4027 443 4113
rect 476 4087 483 4173
rect 516 4087 523 4293
rect 636 4267 643 4333
rect 467 4033 473 4047
rect 416 3807 423 3853
rect 416 3796 433 3807
rect 420 3793 433 3796
rect 476 3767 483 3993
rect 536 3848 543 4093
rect 556 4047 563 4073
rect 596 4007 603 4033
rect 616 4007 623 4213
rect 656 4047 663 4553
rect 676 4307 683 4513
rect 696 4427 703 4513
rect 716 4487 723 4593
rect 676 4087 683 4293
rect 696 4227 703 4413
rect 716 4307 723 4333
rect 716 4187 723 4293
rect 756 4127 763 4273
rect 736 4067 743 4093
rect 687 4033 693 4047
rect 756 4027 763 4113
rect 776 4067 783 4753
rect 796 4527 803 4673
rect 813 4567 827 4573
rect 836 4347 843 4833
rect 856 4767 863 4853
rect 896 4827 903 4873
rect 896 4747 903 4773
rect 916 4727 923 4913
rect 956 4887 963 5093
rect 1033 5087 1047 5093
rect 993 5067 1007 5072
rect 976 4848 983 5033
rect 856 4547 863 4573
rect 893 4567 907 4573
rect 916 4547 923 4713
rect 936 4687 943 4833
rect 933 4587 947 4593
rect 856 4368 863 4533
rect 876 4347 883 4413
rect 916 4367 923 4473
rect 956 4467 963 4633
rect 976 4387 983 4812
rect 996 4747 1003 4993
rect 1016 4987 1023 5033
rect 1013 4867 1027 4873
rect 1016 4603 1023 4853
rect 996 4596 1023 4603
rect 996 4427 1003 4596
rect 1016 4507 1023 4573
rect 1016 4407 1023 4453
rect 827 4336 843 4347
rect 860 4346 883 4347
rect 827 4333 840 4336
rect 867 4335 883 4346
rect 867 4333 880 4335
rect 847 4293 853 4307
rect 793 4287 807 4293
rect 896 4167 903 4333
rect 853 4067 867 4073
rect 727 4013 733 4027
rect 767 4013 773 4027
rect 616 3947 623 3993
rect 573 3827 587 3833
rect 416 3527 423 3753
rect 436 3527 443 3693
rect 456 3687 463 3753
rect 433 3508 447 3513
rect 396 3396 423 3403
rect 287 3263 300 3267
rect 287 3253 303 3263
rect 76 2987 83 3073
rect 93 3007 107 3013
rect 36 2687 43 2733
rect 16 1447 23 2433
rect 56 2287 63 2972
rect 116 2947 123 3033
rect 156 3007 163 3073
rect 207 3003 220 3007
rect 207 2993 223 3003
rect 173 2967 187 2973
rect 216 2947 223 2993
rect 233 2967 247 2973
rect 136 2787 143 2893
rect 196 2787 203 2853
rect 87 2773 93 2787
rect 256 2767 263 3033
rect 213 2747 227 2753
rect 127 2733 133 2747
rect 167 2733 173 2747
rect 276 2743 283 3093
rect 296 2967 303 3253
rect 316 3207 323 3233
rect 356 3047 363 3253
rect 296 2767 303 2853
rect 316 2787 323 2993
rect 353 2987 367 2993
rect 376 2967 383 3133
rect 396 2787 403 3193
rect 416 2808 423 3396
rect 436 3347 443 3472
rect 436 3147 443 3293
rect 456 3107 463 3633
rect 476 3527 483 3653
rect 536 3527 543 3812
rect 596 3787 603 3873
rect 656 3788 663 3813
rect 696 3807 703 3873
rect 816 3827 823 4053
rect 916 4047 923 4353
rect 976 4328 983 4373
rect 1036 4347 1043 5013
rect 1056 4987 1063 5033
rect 1076 4887 1083 5053
rect 1096 5047 1103 5313
rect 1116 5307 1123 5353
rect 1116 4927 1123 5073
rect 1136 5027 1143 5353
rect 1236 5207 1243 5373
rect 1253 5347 1267 5353
rect 1293 5348 1307 5353
rect 1176 5087 1183 5113
rect 1227 5073 1233 5087
rect 1207 5033 1213 5047
rect 1067 4833 1073 4847
rect 1096 4727 1103 4853
rect 1116 4847 1123 4873
rect 1156 4827 1163 5033
rect 1256 5007 1263 5113
rect 1296 5087 1303 5312
rect 1396 5187 1403 5353
rect 1516 5347 1523 5373
rect 1427 5333 1433 5347
rect 1496 5307 1503 5333
rect 1533 5327 1547 5333
rect 1447 5293 1453 5307
rect 1536 5247 1543 5313
rect 1633 5307 1647 5313
rect 1656 5247 1663 5333
rect 1676 5307 1683 5353
rect 1736 5347 1743 5373
rect 1753 5327 1767 5333
rect 1287 5076 1303 5087
rect 1287 5073 1300 5076
rect 1276 5047 1283 5073
rect 1307 5053 1313 5067
rect 1333 5047 1347 5053
rect 1156 4816 1173 4827
rect 1160 4813 1173 4816
rect 1136 4787 1143 4813
rect 1076 4568 1083 4653
rect 1067 4546 1080 4547
rect 1067 4533 1073 4546
rect 947 4313 953 4327
rect 1013 4308 1027 4313
rect 1036 4308 1043 4333
rect 980 4306 1000 4307
rect 987 4302 1000 4306
rect 987 4293 1003 4302
rect 1026 4300 1027 4308
rect 976 4047 983 4272
rect 916 4040 933 4047
rect 913 4033 933 4040
rect 913 4028 927 4033
rect 913 3987 927 3992
rect 916 3947 923 3973
rect 956 3887 963 3993
rect 727 3773 733 3787
rect 556 3747 563 3773
rect 593 3527 607 3533
rect 656 3527 663 3752
rect 727 3733 733 3747
rect 536 3523 553 3527
rect 516 3516 553 3523
rect 516 3487 523 3516
rect 540 3513 553 3516
rect 507 3476 523 3487
rect 533 3487 547 3492
rect 676 3487 683 3733
rect 736 3527 743 3633
rect 776 3548 783 3813
rect 856 3807 863 3833
rect 827 3773 833 3787
rect 956 3767 963 3833
rect 976 3787 983 3813
rect 996 3807 1003 4293
rect 1056 4287 1063 4473
rect 1096 4447 1103 4593
rect 1136 4547 1143 4573
rect 1156 4487 1163 4733
rect 1196 4707 1203 4973
rect 1236 4867 1243 4893
rect 1273 4847 1287 4853
rect 1096 4307 1103 4393
rect 1136 4287 1143 4413
rect 1176 4407 1183 4673
rect 1196 4547 1203 4593
rect 1216 4567 1223 4833
rect 1296 4827 1303 4933
rect 1376 4908 1383 5093
rect 1416 5087 1423 5233
rect 1676 5187 1683 5293
rect 1453 5087 1467 5093
rect 1536 5088 1543 5173
rect 1533 5047 1547 5052
rect 1476 4967 1483 5033
rect 1316 4827 1323 4893
rect 1247 4813 1253 4827
rect 1336 4787 1343 4853
rect 1236 4607 1243 4633
rect 1276 4567 1283 4593
rect 1316 4567 1323 4613
rect 1356 4607 1363 4793
rect 1213 4547 1227 4553
rect 1293 4527 1307 4533
rect 1156 4327 1163 4373
rect 1176 4287 1183 4393
rect 1216 4287 1223 4313
rect 1040 4286 1063 4287
rect 1047 4275 1063 4286
rect 1047 4273 1060 4275
rect 1016 3927 1023 4272
rect 1036 4007 1043 4173
rect 1076 4147 1083 4273
rect 1056 4047 1063 4093
rect 1136 4047 1143 4273
rect 1176 4187 1183 4273
rect 1107 4033 1113 4047
rect 1056 3983 1063 4033
rect 1036 3976 1063 3983
rect 1073 3987 1087 3993
rect 1036 3827 1043 3976
rect 1116 3947 1123 3993
rect 1076 3807 1083 3913
rect 1116 3847 1123 3933
rect 1136 3823 1143 3953
rect 1116 3816 1143 3823
rect 913 3747 927 3753
rect 507 3473 520 3476
rect 567 3473 573 3487
rect 476 3307 483 3453
rect 516 3267 523 3433
rect 547 3293 553 3307
rect 553 3247 567 3253
rect 436 3027 443 3093
rect 496 3047 503 3133
rect 516 3127 523 3173
rect 596 3167 603 3393
rect 696 3347 703 3513
rect 867 3523 880 3527
rect 867 3513 883 3523
rect 716 3447 723 3493
rect 776 3487 783 3512
rect 813 3507 827 3513
rect 776 3476 793 3487
rect 780 3473 793 3476
rect 756 3407 763 3473
rect 656 3287 663 3333
rect 807 3293 813 3307
rect 533 3007 547 3013
rect 487 2993 493 3007
rect 436 2947 443 2973
rect 453 2967 467 2973
rect 456 2787 463 2913
rect 316 2747 323 2773
rect 256 2736 283 2743
rect 216 2707 223 2733
rect 93 2487 107 2493
rect 147 2473 153 2487
rect 127 2433 133 2447
rect 176 2267 183 2493
rect 236 2467 243 2533
rect 256 2487 263 2736
rect 276 2548 283 2713
rect 327 2693 333 2707
rect 416 2563 423 2772
rect 436 2607 443 2733
rect 476 2727 483 2933
rect 496 2907 503 2953
rect 556 2947 563 3093
rect 616 3007 623 3073
rect 636 3047 643 3233
rect 676 3227 683 3253
rect 693 3227 707 3233
rect 736 3227 743 3293
rect 633 3027 647 3033
rect 593 2987 607 2993
rect 636 2867 643 2953
rect 513 2787 527 2793
rect 516 2727 523 2773
rect 676 2767 683 3093
rect 753 3007 767 3013
rect 713 2983 727 2993
rect 713 2980 743 2983
rect 716 2976 743 2980
rect 736 2787 743 2976
rect 776 2967 783 3293
rect 836 3283 843 3473
rect 876 3407 883 3513
rect 816 3276 843 3283
rect 793 3247 807 3253
rect 816 3087 823 3276
rect 856 3267 863 3333
rect 873 3288 887 3293
rect 847 3256 863 3267
rect 847 3253 860 3256
rect 876 3227 883 3252
rect 896 3207 903 3573
rect 936 3288 943 3633
rect 996 3587 1003 3793
rect 1116 3647 1123 3816
rect 1176 3808 1183 4013
rect 1196 4007 1203 4133
rect 1213 4047 1227 4053
rect 1236 4028 1243 4333
rect 1296 4327 1303 4373
rect 1356 4368 1363 4513
rect 1376 4387 1383 4872
rect 1456 4867 1463 4893
rect 1393 4848 1407 4853
rect 1427 4813 1433 4827
rect 1396 4767 1403 4812
rect 1456 4787 1463 4853
rect 1496 4827 1503 4893
rect 1516 4847 1523 4933
rect 1456 4776 1473 4787
rect 1460 4773 1473 4776
rect 1256 4047 1263 4093
rect 1276 4027 1283 4293
rect 1356 4187 1363 4332
rect 1376 4267 1383 4293
rect 1273 4007 1287 4013
rect 1236 3967 1243 3992
rect 1276 3983 1283 3993
rect 1256 3976 1283 3983
rect 1256 3947 1263 3976
rect 1296 3907 1303 4073
rect 1336 4047 1343 4113
rect 1356 4087 1363 4133
rect 1136 3747 1143 3793
rect 953 3547 967 3553
rect 956 3347 963 3493
rect 976 3307 983 3373
rect 996 3367 1003 3533
rect 1016 3327 1023 3513
rect 1036 3287 1043 3573
rect 933 3247 947 3252
rect 853 3007 867 3013
rect 893 2987 907 2993
rect 827 2953 833 2967
rect 876 2907 883 2953
rect 516 2716 533 2727
rect 520 2713 533 2716
rect 473 2707 487 2713
rect 556 2627 563 2753
rect 716 2747 723 2773
rect 796 2747 803 2813
rect 936 2808 943 2993
rect 1016 2967 1023 3073
rect 1056 3027 1063 3473
rect 1096 3467 1103 3513
rect 1116 3487 1123 3593
rect 1136 3587 1143 3733
rect 1176 3667 1183 3772
rect 1196 3607 1203 3893
rect 1216 3567 1223 3793
rect 1236 3747 1243 3873
rect 1256 3767 1263 3813
rect 1316 3807 1323 3953
rect 1336 3887 1343 4033
rect 1256 3756 1273 3767
rect 1260 3753 1273 3756
rect 1336 3763 1343 3833
rect 1356 3827 1363 3993
rect 1376 3987 1383 4013
rect 1396 3923 1403 4473
rect 1416 4388 1423 4633
rect 1447 4553 1453 4567
rect 1476 4527 1483 4593
rect 1496 4567 1503 4713
rect 1536 4608 1543 4793
rect 1556 4647 1563 5133
rect 1756 5127 1763 5313
rect 1747 5116 1763 5127
rect 1747 5113 1760 5116
rect 1587 5073 1593 5087
rect 1596 4967 1603 5033
rect 1616 4907 1623 5093
rect 1713 5087 1727 5093
rect 1636 4987 1643 5073
rect 1687 5053 1693 5067
rect 1696 5008 1703 5053
rect 1796 5047 1803 5373
rect 1827 5333 1833 5347
rect 1816 5047 1823 5333
rect 1876 5327 1883 5373
rect 1916 5347 1923 5373
rect 1833 5087 1847 5093
rect 1956 5087 1963 5333
rect 2033 5327 2047 5333
rect 1847 5073 1853 5087
rect 1927 5073 1933 5087
rect 1956 5076 1973 5087
rect 1960 5073 1973 5076
rect 1847 5033 1853 5047
rect 1576 4827 1583 4893
rect 1607 4853 1613 4867
rect 1636 4827 1643 4933
rect 1676 4827 1683 4853
rect 1576 4816 1593 4827
rect 1580 4813 1593 4816
rect 1696 4727 1703 4972
rect 1720 4863 1733 4867
rect 1716 4853 1733 4863
rect 1716 4627 1723 4853
rect 1776 4847 1783 5033
rect 1876 5007 1883 5073
rect 2016 5047 2023 5273
rect 2076 5267 2083 5333
rect 2116 5167 2123 5352
rect 2136 5143 2143 5393
rect 2216 5387 2223 5453
rect 2347 5374 2353 5387
rect 2347 5373 2360 5374
rect 2153 5368 2167 5373
rect 2156 5287 2163 5332
rect 2196 5267 2203 5333
rect 2176 5147 2183 5233
rect 2276 5227 2283 5373
rect 2433 5368 2447 5373
rect 2353 5347 2367 5352
rect 2427 5346 2440 5347
rect 2427 5333 2433 5346
rect 2313 5327 2327 5333
rect 2116 5136 2143 5143
rect 2116 5107 2123 5136
rect 2147 5123 2160 5127
rect 2147 5113 2163 5123
rect 2267 5123 2280 5127
rect 2267 5113 2283 5123
rect 1956 5007 1963 5033
rect 2036 4947 2043 5093
rect 2113 5088 2127 5093
rect 2076 5003 2083 5073
rect 2107 5066 2120 5067
rect 2107 5053 2113 5066
rect 2076 4996 2103 5003
rect 1947 4853 1953 4867
rect 1747 4813 1753 4827
rect 1493 4547 1507 4553
rect 1416 4307 1423 4352
rect 1436 4347 1443 4513
rect 1536 4467 1543 4572
rect 1596 4567 1603 4593
rect 1613 4587 1627 4593
rect 1567 4533 1573 4547
rect 1656 4527 1663 4573
rect 1716 4567 1723 4613
rect 1796 4603 1803 4813
rect 1816 4767 1823 4833
rect 1856 4827 1863 4853
rect 1813 4707 1827 4713
rect 1787 4596 1803 4603
rect 1776 4567 1783 4593
rect 1816 4567 1823 4633
rect 1836 4567 1843 4653
rect 1856 4607 1863 4713
rect 1876 4567 1883 4853
rect 1976 4827 1983 4893
rect 1907 4813 1913 4827
rect 1967 4816 1983 4827
rect 1967 4813 1980 4816
rect 1916 4787 1923 4813
rect 1996 4803 2003 4933
rect 2036 4827 2043 4853
rect 2056 4847 2063 4893
rect 2096 4867 2103 4996
rect 1976 4796 2003 4803
rect 1927 4776 1943 4783
rect 1907 4553 1913 4567
rect 1656 4513 1673 4527
rect 1847 4513 1853 4527
rect 1456 4108 1463 4413
rect 1536 4347 1543 4373
rect 1587 4343 1600 4347
rect 1587 4333 1603 4343
rect 1513 4287 1527 4293
rect 1556 4227 1563 4293
rect 1596 4187 1603 4333
rect 1616 4307 1623 4513
rect 1656 4347 1663 4513
rect 1716 4407 1723 4513
rect 1687 4293 1693 4307
rect 1376 3916 1403 3923
rect 1376 3867 1383 3916
rect 1336 3756 1363 3763
rect 1276 3727 1283 3753
rect 1316 3707 1323 3753
rect 1147 3523 1160 3527
rect 1147 3513 1163 3523
rect 1207 3513 1213 3527
rect 1156 3487 1163 3513
rect 1096 3387 1103 3453
rect 1236 3347 1243 3693
rect 1256 3527 1263 3593
rect 1173 3287 1187 3293
rect 1087 3273 1093 3287
rect 1133 3267 1147 3273
rect 1076 3007 1083 3093
rect 1116 3007 1123 3073
rect 1136 3027 1143 3253
rect 1233 3247 1247 3253
rect 1196 3207 1203 3233
rect 1053 2967 1067 2973
rect 813 2787 827 2793
rect 933 2767 947 2772
rect 833 2747 847 2753
rect 707 2736 723 2747
rect 707 2733 720 2736
rect 873 2747 887 2753
rect 573 2707 587 2713
rect 396 2556 423 2563
rect 273 2507 287 2512
rect 276 2467 283 2493
rect 347 2453 353 2467
rect 233 2447 247 2453
rect 376 2447 383 2473
rect 256 2267 263 2373
rect 296 2283 303 2413
rect 396 2367 403 2556
rect 413 2467 427 2473
rect 476 2447 483 2513
rect 467 2436 483 2447
rect 467 2433 480 2436
rect 496 2407 503 2613
rect 513 2447 527 2453
rect 276 2276 303 2283
rect 176 2253 193 2267
rect 36 2067 43 2233
rect 53 2207 67 2213
rect 176 2207 183 2253
rect 276 2247 283 2276
rect 313 2267 327 2273
rect 296 2227 303 2253
rect 336 2227 343 2353
rect 396 2227 403 2273
rect 413 2247 427 2253
rect 536 2227 543 2593
rect 556 2487 563 2533
rect 596 2487 603 2573
rect 636 2487 643 2713
rect 713 2707 727 2713
rect 836 2707 843 2733
rect 653 2507 667 2513
rect 636 2447 643 2473
rect 696 2467 703 2573
rect 733 2527 747 2533
rect 747 2514 753 2527
rect 747 2513 760 2514
rect 713 2487 727 2493
rect 587 2433 593 2447
rect 556 2268 563 2393
rect 560 2246 573 2247
rect 567 2233 573 2246
rect 613 2227 627 2233
rect 267 2216 293 2223
rect 96 2167 103 2193
rect 96 2007 103 2053
rect 36 1907 43 1993
rect 107 1953 113 1967
rect 96 1827 103 1893
rect 136 1887 143 1933
rect 236 1927 243 2053
rect 227 1916 243 1927
rect 256 1987 263 2153
rect 276 2008 283 2193
rect 336 2187 343 2213
rect 433 2207 447 2213
rect 533 2207 547 2213
rect 387 2173 393 2187
rect 493 2167 507 2173
rect 316 1987 323 2033
rect 256 1986 280 1987
rect 256 1973 273 1986
rect 227 1913 240 1916
rect 36 1667 43 1753
rect 96 1727 103 1773
rect 136 1727 143 1873
rect 256 1827 263 1973
rect 356 1967 363 1993
rect 96 1447 103 1653
rect 156 1447 163 1813
rect 276 1763 283 1933
rect 256 1756 283 1763
rect 227 1733 233 1747
rect 256 1708 263 1756
rect 296 1747 303 1953
rect 493 1947 507 1953
rect 367 1913 373 1927
rect 316 1747 323 1773
rect 147 1436 163 1447
rect 147 1433 160 1436
rect 76 1407 83 1433
rect 236 1427 243 1653
rect 256 1467 263 1672
rect 276 1447 283 1733
rect 307 1693 313 1707
rect 336 1667 343 1913
rect 456 1887 463 1933
rect 376 1747 383 1813
rect 456 1767 463 1873
rect 427 1733 433 1747
rect 367 1693 373 1707
rect 456 1487 463 1693
rect 536 1667 543 1733
rect 556 1707 563 1833
rect 347 1453 353 1467
rect 107 1393 113 1407
rect 167 1393 173 1407
rect 16 407 23 1393
rect 87 1213 113 1227
rect 56 1027 63 1173
rect 96 803 103 1213
rect 236 1207 243 1273
rect 196 1047 203 1193
rect 296 1187 303 1213
rect 113 907 127 913
rect 136 907 143 1033
rect 256 907 263 1013
rect 76 796 103 803
rect 76 687 83 796
rect 96 447 103 753
rect 116 687 123 813
rect 36 367 43 433
rect 107 393 113 407
rect 136 387 143 893
rect 227 883 240 887
rect 227 873 243 883
rect 236 827 243 873
rect 256 748 263 853
rect 316 787 323 1393
rect 336 1007 343 1373
rect 356 1167 363 1413
rect 373 1227 387 1233
rect 396 1207 403 1453
rect 496 1447 503 1473
rect 556 1448 563 1693
rect 596 1487 603 2133
rect 656 2047 663 2353
rect 676 2067 683 2333
rect 756 2287 763 2492
rect 796 2447 803 2513
rect 696 1967 703 2273
rect 747 2233 753 2247
rect 787 2233 793 2247
rect 816 2227 823 2593
rect 887 2493 893 2507
rect 936 2487 943 2613
rect 976 2587 983 2773
rect 996 2767 1003 2933
rect 1016 2787 1023 2953
rect 1133 2947 1147 2953
rect 1176 2907 1183 2993
rect 1196 2968 1203 3193
rect 1256 3187 1263 3513
rect 1276 3508 1283 3653
rect 1296 3487 1303 3653
rect 1316 3588 1323 3633
rect 1280 3486 1303 3487
rect 1287 3475 1303 3486
rect 1287 3473 1300 3475
rect 1316 3307 1323 3552
rect 1336 3547 1343 3733
rect 1356 3547 1363 3756
rect 1376 3667 1383 3813
rect 1396 3787 1403 3873
rect 1416 3807 1423 4093
rect 1447 4086 1460 4087
rect 1447 4073 1453 4086
rect 1496 4067 1503 4093
rect 1556 4083 1563 4173
rect 1636 4107 1643 4273
rect 1556 4076 1583 4083
rect 1467 4034 1473 4047
rect 1467 4033 1480 4034
rect 1460 4026 1480 4027
rect 1460 4022 1473 4026
rect 1456 4013 1473 4022
rect 1456 3967 1463 4013
rect 1476 3947 1483 3973
rect 1516 3847 1523 4073
rect 1553 4047 1567 4053
rect 1556 3807 1563 3853
rect 1447 3773 1453 3787
rect 1356 3536 1373 3547
rect 1360 3533 1373 3536
rect 1336 3407 1343 3533
rect 1356 3467 1363 3493
rect 1376 3447 1383 3473
rect 1316 3267 1323 3293
rect 1336 3287 1343 3353
rect 1347 3273 1353 3287
rect 1376 3267 1383 3313
rect 1356 3256 1373 3263
rect 1276 3107 1283 3233
rect 1296 3027 1303 3053
rect 1336 3027 1343 3233
rect 1356 3107 1363 3256
rect 1396 3227 1403 3393
rect 1416 3247 1423 3533
rect 1456 3527 1463 3773
rect 1476 3587 1483 3793
rect 1493 3787 1507 3793
rect 1556 3767 1563 3793
rect 1576 3787 1583 4076
rect 1513 3747 1527 3753
rect 1576 3707 1583 3733
rect 1456 3516 1473 3527
rect 1460 3513 1473 3516
rect 1527 3513 1533 3527
rect 1456 3287 1463 3473
rect 1496 3347 1503 3473
rect 1516 3447 1523 3473
rect 1516 3323 1523 3433
rect 1536 3327 1543 3473
rect 1556 3447 1563 3513
rect 1576 3387 1583 3573
rect 1596 3527 1603 4053
rect 1656 4007 1663 4073
rect 1696 4067 1703 4153
rect 1716 4083 1723 4333
rect 1736 4103 1743 4493
rect 1756 4467 1763 4513
rect 1793 4507 1807 4513
rect 1876 4427 1883 4493
rect 1896 4347 1903 4393
rect 1936 4367 1943 4776
rect 1976 4627 1983 4796
rect 2007 4773 2013 4787
rect 1956 4507 1963 4533
rect 1976 4527 1983 4613
rect 2013 4607 2027 4613
rect 2036 4567 2043 4633
rect 2040 4543 2053 4547
rect 2036 4533 2053 4543
rect 1853 4308 1867 4313
rect 1887 4293 1893 4307
rect 1776 4167 1783 4253
rect 1736 4096 1763 4103
rect 1716 4076 1743 4083
rect 1736 4067 1743 4076
rect 1696 4056 1713 4067
rect 1700 4053 1713 4056
rect 1616 3967 1623 3993
rect 1636 3507 1643 3913
rect 1676 3827 1683 4033
rect 1707 4013 1713 4027
rect 1736 4007 1743 4053
rect 1756 3847 1763 4096
rect 1776 3867 1783 4153
rect 1796 4068 1803 4193
rect 1856 4127 1863 4272
rect 1916 4267 1923 4333
rect 1727 3823 1740 3827
rect 1727 3813 1743 3823
rect 1656 3727 1663 3773
rect 1696 3687 1703 3773
rect 1696 3527 1703 3673
rect 1736 3607 1743 3813
rect 1753 3788 1767 3793
rect 1733 3527 1747 3533
rect 1496 3316 1523 3323
rect 1496 3247 1503 3316
rect 1556 3307 1563 3353
rect 1553 3287 1567 3293
rect 1453 3228 1467 3233
rect 1436 3216 1453 3223
rect 1396 3187 1403 3213
rect 1408 3176 1423 3183
rect 1216 2987 1223 3013
rect 993 2747 1007 2753
rect 1036 2747 1043 2813
rect 1053 2787 1067 2793
rect 1116 2767 1123 2893
rect 1196 2827 1203 2932
rect 853 2467 867 2473
rect 956 2467 963 2513
rect 907 2453 913 2467
rect 1016 2347 1023 2453
rect 1076 2447 1083 2533
rect 1136 2527 1143 2793
rect 1207 2753 1213 2767
rect 1153 2747 1167 2753
rect 1236 2743 1243 3013
rect 1196 2740 1243 2743
rect 1193 2736 1243 2740
rect 1193 2727 1207 2736
rect 1256 2727 1263 2993
rect 1276 2947 1283 2973
rect 1353 2963 1367 2973
rect 1336 2960 1367 2963
rect 1336 2956 1363 2960
rect 1336 2907 1343 2956
rect 1376 2943 1383 3173
rect 1416 3027 1423 3176
rect 1436 3067 1443 3216
rect 1516 3207 1523 3273
rect 1596 3267 1603 3293
rect 1456 3147 1463 3192
rect 1456 3047 1463 3093
rect 1453 3027 1467 3033
rect 1356 2936 1383 2943
rect 1247 2716 1263 2727
rect 1247 2713 1260 2716
rect 1196 2527 1203 2713
rect 1276 2627 1283 2773
rect 1336 2747 1343 2893
rect 1356 2747 1363 2936
rect 1376 2768 1383 2913
rect 1416 2907 1423 2953
rect 1456 2883 1463 3013
rect 1476 2987 1483 3073
rect 1536 2967 1543 3173
rect 1596 3087 1603 3253
rect 1636 3243 1643 3273
rect 1676 3267 1683 3473
rect 1716 3447 1723 3473
rect 1736 3307 1743 3453
rect 1693 3287 1707 3293
rect 1696 3247 1703 3273
rect 1636 3236 1663 3243
rect 1556 3007 1563 3073
rect 1596 3007 1603 3033
rect 1573 2967 1587 2973
rect 1616 2907 1623 2953
rect 1436 2876 1463 2883
rect 1393 2787 1407 2793
rect 1356 2746 1380 2747
rect 1356 2735 1373 2746
rect 1360 2733 1373 2735
rect 1196 2516 1213 2527
rect 1200 2513 1213 2516
rect 987 2253 993 2267
rect 1047 2253 1053 2267
rect 776 1967 783 2193
rect 836 1967 843 2173
rect 876 1967 883 2253
rect 896 2187 903 2233
rect 1013 2227 1027 2233
rect 913 2207 927 2213
rect 1013 2207 1027 2213
rect 967 2193 973 2207
rect 1053 2207 1067 2213
rect 1076 2147 1083 2433
rect 1096 2123 1103 2253
rect 1116 2227 1123 2493
rect 1193 2487 1207 2493
rect 1336 2487 1343 2613
rect 1356 2567 1363 2593
rect 1160 2463 1173 2467
rect 1156 2453 1173 2463
rect 1293 2467 1307 2473
rect 1156 2267 1163 2453
rect 1356 2447 1363 2553
rect 1416 2503 1423 2733
rect 1436 2507 1443 2876
rect 1456 2767 1463 2853
rect 1476 2767 1483 2793
rect 1496 2767 1503 2813
rect 1556 2787 1563 2813
rect 1636 2808 1643 3193
rect 1656 2967 1663 3236
rect 1716 3207 1723 3253
rect 1640 2786 1653 2787
rect 1647 2774 1653 2786
rect 1676 2787 1683 2993
rect 1736 2967 1743 3293
rect 1756 2987 1763 3752
rect 1776 3687 1783 3813
rect 1776 3487 1783 3633
rect 1796 3567 1803 4032
rect 1813 4007 1827 4013
rect 1816 3867 1823 3933
rect 1836 3807 1843 4053
rect 1853 4007 1867 4013
rect 1856 3887 1863 3913
rect 1896 3907 1903 4113
rect 1936 4068 1943 4293
rect 1956 4247 1963 4333
rect 1976 4083 1983 4373
rect 2013 4347 2027 4353
rect 2036 4307 2043 4533
rect 2056 4263 2063 4413
rect 2076 4287 2083 4573
rect 2096 4327 2103 4653
rect 2116 4387 2123 4793
rect 2156 4767 2163 5113
rect 2176 4907 2183 5093
rect 2233 5088 2247 5093
rect 2227 5066 2240 5067
rect 2227 5053 2233 5066
rect 2256 4967 2263 5033
rect 2276 4987 2283 5113
rect 2296 5067 2303 5093
rect 2336 5067 2343 5273
rect 2356 5127 2363 5333
rect 2493 5327 2507 5333
rect 2393 5307 2407 5313
rect 2407 5113 2413 5127
rect 2456 5087 2463 5273
rect 2476 5107 2483 5313
rect 2516 5263 2523 5516
rect 2567 5456 2593 5463
rect 2536 5287 2543 5373
rect 2576 5367 2583 5433
rect 2593 5347 2607 5353
rect 2516 5256 2543 5263
rect 2387 5073 2393 5087
rect 2336 5056 2353 5067
rect 2340 5053 2353 5056
rect 2327 5043 2340 5047
rect 2327 5040 2343 5043
rect 2327 5033 2347 5040
rect 2333 5027 2347 5033
rect 2296 4847 2303 5013
rect 2436 4987 2443 5073
rect 2496 5067 2503 5153
rect 2487 5044 2500 5047
rect 2487 5034 2503 5044
rect 2480 5033 2503 5034
rect 2473 5007 2487 5012
rect 2233 4827 2247 4833
rect 2207 4823 2220 4827
rect 2207 4813 2223 4823
rect 2216 4807 2223 4813
rect 2336 4807 2343 4833
rect 2287 4793 2293 4807
rect 2153 4567 2167 4573
rect 2196 4427 2203 4573
rect 2216 4567 2223 4793
rect 2136 4328 2143 4413
rect 2193 4307 2207 4313
rect 2127 4306 2140 4307
rect 2127 4293 2133 4306
rect 2216 4287 2223 4553
rect 2236 4548 2243 4773
rect 2316 4607 2323 4653
rect 2236 4343 2243 4512
rect 2256 4487 2263 4573
rect 2296 4487 2303 4593
rect 2313 4547 2327 4553
rect 2336 4527 2343 4793
rect 2356 4527 2363 4713
rect 2376 4687 2383 4953
rect 2396 4807 2403 4853
rect 2456 4847 2463 4893
rect 2473 4827 2487 4833
rect 2496 4787 2503 5033
rect 2487 4773 2493 4787
rect 2396 4567 2403 4713
rect 2436 4567 2443 4593
rect 2516 4587 2523 5173
rect 2536 4967 2543 5256
rect 2596 5187 2603 5333
rect 2613 5307 2627 5313
rect 2656 5267 2663 5373
rect 2733 5367 2747 5373
rect 2776 5347 2783 5433
rect 2767 5336 2783 5347
rect 2767 5333 2780 5336
rect 2716 5307 2723 5333
rect 2796 5327 2803 5373
rect 2856 5367 2863 5393
rect 2896 5387 2903 5453
rect 3093 5387 3107 5393
rect 2993 5367 3007 5373
rect 2860 5343 2873 5347
rect 2856 5333 2873 5343
rect 2836 5267 2843 5293
rect 2856 5287 2863 5333
rect 2893 5307 2907 5313
rect 2976 5287 2983 5333
rect 2996 5307 3003 5353
rect 3036 5347 3043 5373
rect 3116 5363 3123 5523
rect 3156 5387 3163 5453
rect 3096 5356 3123 5363
rect 3193 5367 3207 5373
rect 3027 5336 3043 5347
rect 3027 5333 3040 5336
rect 3076 5287 3083 5333
rect 2556 4827 2563 5093
rect 2587 5074 2593 5087
rect 2616 5087 2623 5153
rect 2580 5073 2600 5074
rect 2613 5067 2627 5073
rect 2576 4907 2583 5052
rect 2593 5027 2607 5033
rect 2576 4847 2583 4893
rect 2636 4883 2643 5213
rect 2656 5107 2663 5133
rect 2747 5113 2753 5127
rect 2727 5073 2733 5087
rect 2747 5073 2753 5087
rect 2687 5053 2693 5067
rect 2616 4880 2643 4883
rect 2613 4876 2643 4880
rect 2613 4867 2627 4876
rect 2696 4867 2703 4973
rect 2776 4947 2783 5033
rect 2576 4837 2593 4847
rect 2580 4834 2593 4837
rect 2580 4833 2600 4834
rect 2600 4826 2613 4827
rect 2607 4813 2613 4826
rect 2536 4647 2543 4793
rect 2636 4787 2643 4853
rect 2713 4827 2727 4833
rect 2747 4813 2753 4827
rect 2556 4623 2563 4673
rect 2536 4616 2563 4623
rect 2387 4553 2393 4567
rect 2536 4563 2543 4616
rect 2576 4607 2583 4713
rect 2516 4556 2543 4563
rect 2433 4547 2447 4553
rect 2476 4523 2483 4553
rect 2427 4516 2483 4523
rect 2256 4367 2263 4473
rect 2416 4407 2423 4453
rect 2236 4336 2263 4343
rect 2056 4256 2083 4263
rect 1956 4076 1983 4083
rect 1956 4047 1963 4076
rect 1973 4047 1987 4053
rect 1933 4027 1947 4032
rect 1976 3927 1983 4033
rect 1993 3987 2007 3993
rect 1896 3896 1913 3907
rect 1900 3893 1913 3896
rect 1856 3827 1863 3873
rect 1936 3827 1943 3873
rect 1833 3787 1847 3793
rect 1856 3527 1863 3773
rect 1813 3503 1827 3513
rect 1796 3500 1827 3503
rect 1796 3496 1823 3500
rect 1776 3028 1783 3373
rect 1796 3367 1803 3496
rect 1896 3487 1903 3813
rect 1956 3803 1963 3833
rect 1936 3796 1963 3803
rect 1916 3487 1923 3793
rect 1936 3547 1943 3796
rect 1976 3787 1983 3853
rect 1996 3843 2003 3893
rect 2016 3887 2023 4233
rect 2033 4007 2047 4013
rect 1996 3836 2023 3843
rect 1956 3647 1963 3773
rect 1996 3747 2003 3813
rect 2016 3807 2023 3836
rect 2036 3827 2043 3993
rect 1973 3548 1987 3553
rect 1887 3473 1903 3487
rect 1816 3307 1823 3413
rect 1896 3347 1903 3473
rect 1936 3403 1943 3533
rect 1973 3507 1987 3512
rect 1936 3396 1963 3403
rect 1796 3267 1803 3293
rect 1816 3187 1823 3293
rect 1896 3247 1903 3273
rect 1916 3267 1923 3373
rect 1807 2993 1813 3007
rect 1713 2947 1727 2953
rect 1716 2868 1723 2933
rect 1756 2907 1763 2973
rect 1776 2847 1783 2992
rect 1836 2967 1843 3233
rect 1876 3187 1883 3233
rect 1933 3203 1947 3213
rect 1916 3200 1947 3203
rect 1916 3196 1943 3200
rect 1647 2773 1660 2774
rect 1466 2753 1467 2760
rect 1453 2747 1467 2753
rect 1613 2727 1627 2733
rect 1616 2627 1623 2713
rect 1636 2567 1643 2772
rect 1653 2747 1667 2752
rect 1716 2747 1723 2832
rect 1796 2827 1803 2953
rect 1707 2736 1723 2747
rect 1707 2733 1720 2736
rect 1736 2727 1743 2793
rect 1767 2773 1773 2787
rect 1793 2763 1807 2773
rect 1776 2760 1807 2763
rect 1776 2756 1803 2760
rect 1776 2507 1783 2756
rect 1836 2747 1843 2793
rect 1856 2787 1863 2953
rect 1916 2947 1923 3196
rect 1933 3007 1947 3013
rect 1956 3007 1963 3396
rect 1996 3307 2003 3593
rect 2016 3588 2023 3793
rect 2056 3787 2063 4153
rect 2076 4088 2083 4256
rect 2093 4247 2107 4253
rect 2136 4207 2143 4233
rect 2096 4127 2103 4153
rect 2076 3907 2083 4052
rect 2096 4047 2103 4113
rect 2136 4027 2143 4193
rect 2156 4067 2163 4193
rect 2176 4107 2183 4273
rect 2256 4067 2263 4336
rect 2287 4334 2293 4347
rect 2436 4347 2443 4413
rect 2456 4387 2463 4493
rect 2280 4333 2300 4334
rect 2353 4327 2367 4333
rect 2276 4167 2283 4312
rect 2296 4207 2303 4312
rect 2313 4247 2327 4253
rect 2136 4003 2143 4013
rect 2116 3996 2143 4003
rect 2056 3727 2063 3773
rect 2076 3687 2083 3793
rect 2096 3668 2103 3973
rect 2116 3807 2123 3996
rect 2013 3547 2027 3552
rect 2056 3547 2063 3593
rect 2033 3267 2047 3273
rect 1996 3207 2003 3233
rect 2033 3207 2047 3213
rect 2036 3147 2043 3193
rect 2056 3067 2063 3493
rect 2096 3367 2103 3632
rect 2116 3567 2123 3793
rect 2156 3787 2163 3813
rect 2176 3787 2183 4053
rect 2196 3827 2203 4013
rect 2216 3947 2223 4053
rect 2233 4027 2247 4033
rect 2236 3827 2243 3873
rect 2256 3787 2263 3913
rect 2156 3776 2173 3787
rect 2160 3773 2173 3776
rect 2276 3607 2283 4093
rect 2356 4087 2363 4313
rect 2413 4287 2427 4293
rect 2307 4013 2313 4027
rect 2336 4007 2343 4033
rect 2376 3843 2383 4213
rect 2416 4107 2423 4273
rect 2436 4187 2443 4333
rect 2456 4307 2463 4373
rect 2476 4227 2483 4433
rect 2516 4307 2523 4556
rect 2567 4554 2573 4567
rect 2596 4567 2603 4613
rect 2676 4567 2683 4733
rect 2776 4727 2783 4933
rect 2796 4867 2803 5033
rect 2816 5027 2823 5113
rect 2707 4613 2713 4627
rect 2767 4613 2773 4627
rect 2560 4553 2580 4554
rect 2647 4553 2653 4567
rect 2676 4556 2693 4567
rect 2680 4553 2693 4556
rect 2547 4546 2560 4547
rect 2547 4533 2553 4546
rect 2736 4527 2743 4593
rect 2796 4567 2803 4653
rect 2816 4587 2823 5013
rect 2836 4847 2843 5253
rect 2856 4867 2863 5273
rect 2996 5107 3003 5193
rect 2953 5087 2967 5093
rect 2907 5073 2913 5087
rect 2933 5047 2947 5053
rect 2996 5047 3003 5093
rect 3053 5088 3067 5093
rect 2987 5036 3003 5047
rect 2987 5033 3000 5036
rect 2893 5027 2907 5033
rect 3056 5027 3063 5052
rect 2906 5020 2907 5027
rect 2916 4947 2923 5013
rect 2893 4867 2907 4873
rect 2956 4867 2963 4953
rect 3016 4943 3023 5013
rect 3053 4967 3067 4973
rect 3047 4960 3067 4967
rect 3047 4956 3063 4960
rect 3047 4953 3060 4956
rect 3016 4936 3053 4943
rect 2873 4807 2887 4813
rect 2836 4607 2843 4793
rect 2876 4743 2883 4793
rect 2876 4736 2903 4743
rect 2787 4553 2793 4567
rect 2627 4513 2633 4527
rect 2767 4513 2773 4527
rect 2616 4427 2623 4513
rect 2647 4333 2653 4347
rect 2593 4327 2607 4333
rect 2513 4287 2527 4293
rect 2556 4287 2563 4313
rect 2693 4307 2707 4313
rect 2456 4067 2463 4093
rect 2396 3967 2403 4013
rect 2416 3847 2423 4053
rect 2496 4027 2503 4173
rect 2527 4033 2533 4047
rect 2573 4027 2587 4033
rect 2456 3847 2463 4013
rect 2547 3993 2553 4007
rect 2476 3887 2483 3953
rect 2356 3836 2383 3843
rect 2296 3767 2303 3793
rect 2316 3767 2323 3793
rect 2356 3788 2363 3836
rect 2376 3816 2433 3823
rect 2353 3747 2367 3752
rect 2316 3607 2323 3713
rect 2136 3547 2143 3593
rect 2156 3427 2163 3553
rect 2187 3533 2193 3547
rect 2260 3523 2273 3527
rect 2256 3513 2273 3523
rect 2136 3416 2153 3423
rect 2076 3267 2083 3293
rect 2096 3207 2103 3293
rect 2136 3283 2143 3416
rect 2116 3276 2143 3283
rect 1973 3007 1987 3013
rect 1956 2967 1963 2993
rect 2016 2987 2023 3053
rect 1996 2976 2013 2983
rect 1996 2827 2003 2976
rect 2036 2967 2043 3033
rect 2056 2947 2063 2993
rect 2076 2907 2083 2973
rect 2116 2947 2123 3276
rect 2147 3253 2153 3267
rect 2176 3087 2183 3493
rect 2196 3307 2203 3373
rect 2256 3287 2263 3513
rect 2287 3473 2293 3487
rect 2316 3463 2323 3513
rect 2336 3487 2343 3713
rect 2296 3456 2323 3463
rect 2267 3233 2273 3247
rect 2296 3243 2303 3456
rect 2356 3407 2363 3573
rect 2313 3307 2327 3313
rect 2287 3236 2303 3243
rect 2213 3227 2227 3233
rect 2176 3028 2183 3073
rect 2133 3007 2147 3013
rect 2167 3006 2180 3007
rect 2167 2994 2173 3006
rect 2160 2993 2173 2994
rect 2153 2967 2167 2972
rect 2196 2967 2203 3113
rect 2213 3007 2227 3013
rect 2356 2987 2363 3133
rect 2376 3107 2383 3816
rect 2396 3447 2403 3793
rect 2453 3787 2467 3793
rect 2413 3767 2427 3773
rect 2456 3727 2463 3773
rect 2476 3747 2483 3813
rect 2416 3567 2423 3613
rect 2447 3533 2453 3547
rect 2476 3543 2483 3733
rect 2496 3687 2503 3853
rect 2516 3667 2523 3993
rect 2576 3947 2583 4013
rect 2556 3827 2563 3893
rect 2556 3787 2563 3813
rect 2576 3687 2583 3773
rect 2596 3707 2603 4033
rect 2613 4007 2627 4013
rect 2636 3807 2643 3973
rect 2676 3947 2683 4293
rect 2716 4267 2723 4333
rect 2733 4287 2747 4293
rect 2696 4067 2703 4233
rect 2656 3808 2663 3933
rect 2676 3827 2683 3893
rect 2696 3867 2703 4053
rect 2733 3987 2747 3993
rect 2756 3907 2763 4313
rect 2776 4167 2783 4193
rect 2796 4147 2803 4553
rect 2833 4547 2847 4553
rect 2876 4527 2883 4573
rect 2896 4503 2903 4736
rect 2916 4687 2923 4833
rect 2947 4813 2953 4827
rect 2996 4807 3003 4833
rect 3016 4827 3023 4913
rect 3076 4907 3083 5233
rect 3096 5227 3103 5356
rect 3127 5333 3133 5347
rect 3167 5333 3173 5347
rect 3216 5248 3223 5523
rect 4256 5487 4263 5523
rect 3447 5456 3473 5463
rect 3233 5387 3247 5393
rect 3353 5387 3367 5393
rect 3413 5387 3427 5393
rect 3456 5387 3463 5433
rect 3576 5347 3583 5413
rect 3676 5387 3683 5413
rect 3676 5376 3693 5387
rect 3680 5373 3693 5376
rect 3800 5383 3813 5387
rect 3796 5373 3813 5383
rect 3427 5333 3433 5347
rect 3096 5067 3103 5133
rect 3116 5063 3123 5093
rect 3176 5087 3183 5153
rect 3147 5083 3160 5087
rect 3147 5073 3163 5083
rect 3116 5056 3143 5063
rect 3116 4947 3123 5033
rect 3036 4767 3043 4893
rect 3116 4867 3123 4893
rect 3136 4887 3143 5056
rect 3156 4907 3163 5073
rect 3176 5027 3183 5073
rect 3176 4867 3183 4953
rect 3216 4883 3223 5212
rect 3236 5107 3243 5173
rect 3256 5083 3263 5273
rect 3236 5076 3263 5083
rect 3236 5047 3243 5076
rect 3276 5067 3283 5213
rect 3296 5147 3303 5333
rect 3296 5087 3303 5133
rect 3316 5127 3323 5233
rect 3336 5047 3343 5333
rect 3476 5287 3483 5333
rect 3553 5287 3567 5293
rect 3556 5187 3563 5273
rect 3576 5247 3583 5333
rect 3596 5307 3603 5353
rect 3616 5327 3623 5353
rect 3776 5347 3783 5373
rect 3627 5313 3633 5327
rect 3676 5307 3683 5333
rect 3596 5227 3603 5293
rect 3507 5113 3513 5127
rect 3396 5087 3403 5113
rect 3596 5107 3603 5213
rect 3716 5187 3723 5333
rect 3796 5267 3803 5373
rect 3827 5333 3833 5347
rect 3740 5203 3753 5207
rect 3736 5193 3753 5203
rect 3447 5073 3453 5087
rect 3413 5027 3427 5033
rect 3196 4876 3223 4883
rect 3073 4848 3087 4853
rect 3080 4826 3093 4827
rect 3056 4816 3073 4823
rect 2916 4587 2923 4613
rect 2876 4496 2903 4503
rect 2793 4047 2807 4053
rect 2787 4033 2793 4047
rect 2816 4028 2823 4373
rect 2836 4287 2843 4473
rect 2856 4287 2863 4413
rect 2876 4307 2883 4496
rect 2916 4487 2923 4533
rect 2936 4427 2943 4753
rect 3016 4607 3023 4633
rect 2973 4568 2987 4573
rect 2967 4546 2980 4547
rect 2967 4533 2973 4546
rect 3016 4387 3023 4593
rect 3056 4587 3063 4816
rect 3087 4813 3093 4826
rect 3133 4807 3147 4813
rect 3096 4587 3103 4693
rect 3136 4547 3143 4673
rect 3156 4647 3163 4853
rect 3196 4547 3203 4876
rect 3267 4853 3273 4867
rect 3227 4843 3240 4847
rect 3227 4833 3243 4843
rect 3236 4707 3243 4833
rect 3253 4807 3267 4813
rect 3256 4683 3263 4793
rect 3296 4687 3303 5013
rect 3516 4943 3523 5073
rect 3547 5063 3560 5067
rect 3547 5053 3563 5063
rect 3533 5047 3547 5053
rect 3516 4936 3543 4943
rect 3496 4867 3503 4933
rect 3516 4867 3523 4913
rect 3356 4827 3363 4853
rect 3467 4833 3473 4847
rect 3236 4676 3263 4683
rect 3213 4567 3227 4573
rect 3236 4568 3243 4676
rect 3213 4560 3233 4567
rect 3216 4554 3233 4560
rect 3256 4567 3263 4653
rect 3216 4553 3240 4554
rect 3033 4527 3047 4533
rect 3216 4527 3223 4553
rect 3016 4347 3023 4373
rect 3056 4367 3063 4473
rect 3076 4327 3083 4393
rect 3153 4347 3167 4353
rect 3107 4334 3113 4347
rect 3100 4333 3113 4334
rect 3193 4328 3207 4333
rect 2873 4287 2887 4293
rect 2856 4247 2863 4273
rect 2896 4267 2903 4313
rect 2913 4307 2927 4313
rect 3013 4287 3027 4293
rect 2973 4267 2987 4273
rect 2986 4260 2987 4267
rect 2876 4107 2883 4153
rect 2847 4034 2853 4047
rect 2847 4033 2860 4034
rect 2776 3967 2783 3993
rect 2816 3947 2823 3992
rect 2627 3796 2643 3807
rect 2627 3793 2640 3796
rect 2476 3536 2493 3543
rect 2473 3507 2487 3512
rect 2496 3487 2503 3533
rect 2516 3527 2523 3653
rect 2576 3607 2583 3673
rect 2516 3516 2533 3527
rect 2520 3513 2533 3516
rect 2567 3513 2573 3527
rect 2516 3447 2523 3473
rect 2396 3308 2403 3353
rect 2396 3147 2403 3272
rect 2416 3103 2423 3373
rect 2556 3323 2563 3473
rect 2536 3316 2563 3323
rect 2433 3267 2447 3273
rect 2396 3096 2423 3103
rect 2396 3007 2403 3096
rect 2273 2947 2287 2953
rect 1893 2807 1907 2813
rect 1916 2747 1923 2813
rect 2133 2787 2147 2793
rect 1953 2767 1967 2773
rect 1396 2496 1423 2503
rect 1313 2427 1327 2433
rect 1376 2427 1383 2473
rect 1396 2447 1403 2496
rect 1573 2487 1587 2493
rect 1427 2476 1453 2483
rect 1493 2467 1507 2473
rect 1613 2467 1627 2473
rect 1796 2467 1803 2733
rect 1993 2727 2007 2733
rect 2016 2707 2023 2773
rect 2113 2747 2127 2753
rect 2316 2747 2323 2773
rect 2356 2767 2363 2973
rect 2376 2807 2383 2953
rect 2433 2787 2447 2793
rect 2353 2747 2367 2753
rect 2067 2733 2073 2747
rect 2207 2713 2213 2727
rect 2153 2707 2167 2713
rect 1956 2547 1963 2693
rect 2196 2687 2203 2713
rect 1956 2487 1963 2533
rect 1873 2467 1887 2473
rect 2076 2467 2083 2493
rect 2347 2473 2353 2487
rect 1427 2433 1433 2447
rect 1500 2443 1513 2447
rect 1496 2433 1513 2443
rect 1196 2267 1203 2293
rect 1256 2267 1263 2373
rect 1347 2263 1360 2267
rect 1347 2253 1363 2263
rect 1153 2247 1167 2253
rect 1076 2116 1103 2123
rect 647 1953 653 1967
rect 827 1953 833 1967
rect 907 1954 913 1967
rect 1076 1967 1083 2116
rect 1196 2063 1203 2253
rect 1276 2187 1283 2213
rect 1296 2163 1303 2253
rect 1313 2207 1327 2213
rect 1176 2056 1203 2063
rect 1276 2156 1303 2163
rect 907 1953 920 1954
rect 636 1847 643 1913
rect 656 1827 663 1953
rect 673 1927 687 1933
rect 716 1807 723 1913
rect 676 1707 683 1793
rect 816 1787 823 1953
rect 913 1927 927 1932
rect 736 1727 743 1753
rect 793 1747 807 1753
rect 727 1713 733 1727
rect 596 1447 603 1473
rect 736 1447 743 1473
rect 453 1427 467 1433
rect 456 1307 463 1413
rect 416 1227 423 1273
rect 393 1187 407 1193
rect 433 1167 447 1173
rect 367 913 373 927
rect 387 913 393 927
rect 436 887 443 973
rect 476 948 483 1253
rect 496 1228 503 1433
rect 693 1428 707 1433
rect 536 1207 543 1373
rect 556 1247 563 1412
rect 636 1387 643 1413
rect 776 1407 783 1553
rect 816 1407 823 1773
rect 836 1707 843 1913
rect 867 1733 873 1747
rect 856 1667 863 1733
rect 887 1693 893 1707
rect 876 1527 883 1693
rect 856 1427 863 1473
rect 896 1427 903 1653
rect 936 1607 943 1953
rect 1027 1933 1033 1947
rect 953 1927 967 1933
rect 1016 1727 1023 1753
rect 1036 1727 1043 1933
rect 1133 1727 1147 1733
rect 1047 1713 1053 1727
rect 700 1406 713 1407
rect 676 1307 683 1393
rect 707 1393 713 1406
rect 913 1387 927 1393
rect 496 927 503 1192
rect 513 1167 527 1173
rect 556 1167 563 1233
rect 573 1207 587 1213
rect 596 1187 603 1293
rect 676 1227 683 1253
rect 753 1227 767 1233
rect 627 1213 633 1227
rect 847 1193 853 1207
rect 876 1187 883 1293
rect 956 1267 963 1413
rect 647 1173 653 1187
rect 513 1147 527 1153
rect 516 987 523 1133
rect 460 926 480 927
rect 467 913 473 926
rect 496 916 513 927
rect 500 913 513 916
rect 436 876 453 887
rect 440 873 453 876
rect 376 827 383 873
rect 156 667 163 713
rect 216 687 223 733
rect 253 707 267 712
rect 327 693 333 707
rect 427 693 433 707
rect 213 667 227 673
rect 156 656 173 667
rect 160 653 173 656
rect 276 507 283 693
rect 307 653 313 667
rect 367 653 373 667
rect 427 653 433 667
rect 456 567 463 873
rect 493 867 507 873
rect 516 627 523 673
rect 536 647 543 693
rect 576 667 583 933
rect 596 867 603 953
rect 616 907 623 1173
rect 696 1067 703 1173
rect 656 927 663 993
rect 736 927 743 993
rect 613 887 627 893
rect 776 887 783 913
rect 816 907 823 1053
rect 976 983 983 1593
rect 996 1407 1003 1433
rect 1036 1387 1043 1413
rect 1013 1227 1027 1233
rect 1016 1147 1023 1213
rect 1056 1207 1063 1473
rect 1156 1447 1163 1513
rect 1176 1487 1183 2056
rect 1276 1967 1283 2156
rect 1356 2147 1363 2253
rect 1436 2227 1443 2333
rect 1476 2263 1483 2433
rect 1456 2256 1483 2263
rect 1296 1947 1303 2093
rect 1456 2067 1463 2256
rect 1476 2187 1483 2233
rect 1476 2107 1483 2173
rect 1496 1988 1503 2433
rect 1556 2347 1563 2433
rect 1567 2253 1573 2267
rect 1607 2253 1613 2267
rect 1516 1967 1523 2053
rect 1500 1966 1523 1967
rect 1507 1955 1523 1966
rect 1507 1953 1520 1955
rect 1536 1947 1543 2093
rect 1616 2067 1623 2253
rect 1636 2247 1643 2433
rect 1633 2227 1647 2233
rect 1676 2187 1683 2453
rect 1727 2233 1733 2247
rect 1696 1967 1703 2133
rect 1756 1987 1763 2253
rect 1707 1953 1713 1967
rect 1733 1947 1747 1953
rect 1387 1923 1400 1927
rect 1387 1913 1403 1923
rect 1396 1887 1403 1913
rect 1196 1747 1203 1773
rect 1233 1747 1247 1753
rect 1387 1743 1400 1747
rect 1387 1733 1403 1743
rect 1373 1727 1387 1733
rect 1227 1693 1233 1707
rect 1367 1703 1380 1707
rect 1367 1693 1383 1703
rect 1256 1647 1263 1693
rect 1376 1667 1383 1693
rect 1396 1687 1403 1733
rect 1496 1727 1503 1932
rect 1627 1923 1640 1927
rect 1627 1913 1643 1923
rect 1687 1913 1693 1927
rect 1487 1713 1493 1727
rect 1513 1707 1527 1713
rect 1416 1667 1423 1693
rect 1536 1487 1543 1793
rect 1553 1767 1567 1773
rect 1413 1467 1427 1473
rect 1227 1433 1233 1447
rect 1287 1433 1293 1447
rect 1153 1427 1167 1433
rect 1313 1427 1327 1433
rect 1093 1387 1107 1393
rect 1116 1327 1123 1413
rect 1356 1407 1363 1433
rect 1376 1407 1383 1453
rect 1487 1433 1493 1447
rect 1547 1433 1553 1447
rect 1493 1427 1507 1433
rect 1576 1427 1583 1753
rect 1636 1747 1643 1913
rect 1676 1887 1683 1913
rect 1716 1807 1723 1893
rect 1776 1847 1783 2273
rect 1836 2267 1843 2453
rect 1916 2407 1923 2453
rect 1980 2443 1993 2447
rect 1953 2427 1967 2433
rect 1976 2433 1993 2443
rect 1976 2407 1983 2433
rect 1916 2367 1923 2393
rect 2076 2347 2083 2453
rect 2116 2427 2123 2473
rect 2296 2447 2303 2473
rect 2213 2427 2227 2433
rect 2313 2427 2327 2433
rect 1907 2253 1913 2267
rect 1813 2227 1827 2233
rect 1847 2213 1853 2227
rect 1876 2007 1883 2253
rect 1996 2247 2003 2333
rect 2033 2247 2047 2253
rect 1816 1803 1823 1973
rect 1847 1953 1853 1967
rect 1896 1947 1903 2053
rect 1936 1967 1943 1993
rect 1996 1987 2003 2233
rect 2176 2227 2183 2333
rect 2293 2267 2307 2273
rect 2336 2267 2343 2313
rect 2207 2253 2213 2267
rect 2267 2253 2273 2267
rect 2233 2227 2247 2233
rect 2176 2216 2193 2227
rect 2180 2213 2193 2216
rect 2296 2207 2303 2253
rect 1973 1927 1987 1933
rect 1816 1796 1843 1803
rect 1787 1753 1793 1767
rect 1633 1727 1647 1733
rect 1687 1713 1693 1727
rect 1736 1707 1743 1753
rect 1807 1713 1813 1727
rect 1736 1696 1753 1707
rect 1740 1693 1753 1696
rect 1613 1687 1627 1693
rect 1616 1447 1623 1573
rect 1147 1373 1153 1387
rect 1216 1327 1223 1393
rect 1116 1187 1123 1313
rect 1136 1227 1143 1253
rect 1147 1213 1173 1227
rect 1296 1207 1303 1273
rect 1436 1267 1443 1393
rect 1476 1367 1483 1393
rect 1516 1347 1523 1393
rect 1456 1243 1463 1313
rect 1413 1227 1427 1233
rect 1436 1236 1463 1243
rect 1267 1193 1273 1207
rect 967 976 983 983
rect 853 947 867 953
rect 707 873 713 887
rect 707 673 713 687
rect 573 647 587 653
rect 616 647 623 673
rect 756 647 763 873
rect 816 667 823 893
rect 896 867 903 933
rect 956 907 963 973
rect 1056 947 1063 973
rect 1087 933 1093 947
rect 1013 927 1027 933
rect 1173 927 1187 933
rect 976 723 983 853
rect 976 720 1003 723
rect 976 716 1007 720
rect 993 707 1007 716
rect 887 693 893 707
rect 616 636 633 647
rect 620 633 633 636
rect 747 636 763 647
rect 773 647 787 653
rect 747 633 760 636
rect 673 627 687 633
rect 536 527 543 553
rect 347 373 353 387
rect 133 367 147 373
rect 260 363 273 367
rect 96 307 103 353
rect 213 347 227 353
rect 256 353 273 363
rect 116 187 123 333
rect 136 207 143 293
rect 256 287 263 353
rect 396 347 403 373
rect 87 173 93 187
rect 113 167 127 173
rect 136 147 143 193
rect 253 187 267 193
rect 296 187 303 273
rect 233 147 247 153
rect 296 147 303 173
rect 336 167 343 193
rect 67 133 73 147
rect 273 127 287 133
rect 396 87 403 193
rect 416 147 423 273
rect 516 207 523 493
rect 536 367 543 513
rect 716 407 723 633
rect 836 547 843 673
rect 913 667 927 673
rect 876 627 883 653
rect 936 623 943 693
rect 956 647 963 673
rect 1016 663 1023 813
rect 1056 687 1063 873
rect 996 656 1023 663
rect 1053 667 1067 673
rect 936 616 963 623
rect 556 287 563 393
rect 573 347 587 353
rect 596 267 603 393
rect 756 387 763 453
rect 876 367 883 413
rect 916 387 923 613
rect 956 427 963 616
rect 847 353 853 367
rect 956 347 963 413
rect 996 403 1003 656
rect 1076 647 1083 893
rect 1236 887 1243 1133
rect 1256 903 1263 1193
rect 1436 1187 1443 1236
rect 1476 1227 1483 1273
rect 1467 1216 1483 1227
rect 1467 1213 1480 1216
rect 1556 1207 1563 1353
rect 1527 1193 1533 1207
rect 1476 1127 1483 1173
rect 1273 927 1287 933
rect 1413 927 1427 933
rect 1556 927 1563 1193
rect 1467 913 1473 927
rect 1313 907 1327 913
rect 1256 896 1283 903
rect 1236 876 1253 887
rect 1240 873 1253 876
rect 1196 823 1203 873
rect 1176 816 1203 823
rect 1156 688 1163 733
rect 1176 727 1183 816
rect 1176 716 1193 727
rect 1180 713 1193 716
rect 1276 687 1283 896
rect 1307 883 1320 887
rect 1307 873 1323 883
rect 1316 687 1323 873
rect 1436 727 1443 873
rect 1456 687 1463 913
rect 1496 887 1503 913
rect 1576 887 1583 1413
rect 1616 1343 1623 1433
rect 1616 1336 1643 1343
rect 1616 947 1623 1073
rect 1636 967 1643 1336
rect 1676 947 1683 1673
rect 1700 1483 1713 1487
rect 1696 1473 1713 1483
rect 1696 1347 1703 1473
rect 1756 1468 1763 1693
rect 1836 1547 1843 1796
rect 1876 1747 1883 1773
rect 1873 1727 1887 1733
rect 1896 1627 1903 1693
rect 1916 1587 1923 1753
rect 1956 1747 1963 1893
rect 1956 1707 1963 1733
rect 1996 1727 2003 1833
rect 2036 1687 2043 2193
rect 2356 2087 2363 2473
rect 2396 2467 2403 2573
rect 2387 2453 2393 2467
rect 2376 2247 2383 2293
rect 2416 2247 2423 2333
rect 2456 2307 2463 2633
rect 2476 2243 2483 3093
rect 2536 3007 2543 3316
rect 2576 3307 2583 3433
rect 2616 3367 2623 3793
rect 2713 3787 2727 3793
rect 2660 3786 2673 3787
rect 2667 3773 2673 3786
rect 2776 3767 2783 3813
rect 2833 3807 2847 3813
rect 2856 3783 2863 4012
rect 2876 3927 2883 4053
rect 2896 4027 2903 4253
rect 2936 4103 2943 4253
rect 2936 4096 2963 4103
rect 2936 4027 2943 4053
rect 2956 4007 2963 4096
rect 2996 4007 3003 4253
rect 3096 4207 3103 4312
rect 3236 4307 3243 4532
rect 3256 4527 3263 4553
rect 3316 4527 3323 4753
rect 3356 4727 3363 4813
rect 3373 4807 3387 4813
rect 3376 4767 3383 4793
rect 3416 4707 3423 4833
rect 3493 4807 3507 4813
rect 3416 4667 3423 4693
rect 3376 4547 3383 4633
rect 3516 4583 3523 4853
rect 3496 4580 3523 4583
rect 3453 4567 3467 4573
rect 3447 4553 3453 4567
rect 3493 4576 3523 4580
rect 3493 4567 3507 4576
rect 3276 4307 3283 4433
rect 3316 4347 3323 4513
rect 3356 4427 3363 4473
rect 3376 4467 3383 4533
rect 3416 4407 3423 4513
rect 3347 4403 3360 4407
rect 3347 4400 3363 4403
rect 3347 4393 3367 4400
rect 3353 4387 3367 4393
rect 3307 4336 3323 4347
rect 3333 4347 3347 4353
rect 3307 4333 3320 4336
rect 3393 4307 3407 4313
rect 3187 4304 3200 4307
rect 3187 4294 3203 4304
rect 3180 4293 3203 4294
rect 3133 4287 3147 4293
rect 3013 4047 3027 4053
rect 3036 4023 3043 4193
rect 3176 4061 3183 4272
rect 3196 4127 3203 4293
rect 3276 4147 3283 4293
rect 3053 4047 3067 4053
rect 3016 4016 3043 4023
rect 2996 3967 3003 3993
rect 2836 3780 2863 3783
rect 2833 3776 2863 3780
rect 2833 3767 2847 3776
rect 2796 3687 2803 3753
rect 2833 3747 2847 3753
rect 2736 3507 2743 3553
rect 2693 3487 2707 3493
rect 2560 3303 2573 3307
rect 2556 3293 2573 3303
rect 2556 3207 2563 3293
rect 2596 3267 2603 3333
rect 2613 3287 2627 3293
rect 2673 3267 2687 3273
rect 2647 3253 2653 3267
rect 2716 3247 2723 3333
rect 2496 2767 2503 2953
rect 2516 2947 2523 2973
rect 2556 2967 2563 3193
rect 2696 3107 2703 3173
rect 2716 3167 2723 3233
rect 2673 3007 2687 3013
rect 2736 2987 2743 3493
rect 2836 3487 2843 3733
rect 2876 3667 2883 3813
rect 2916 3807 2923 3833
rect 2956 3807 2963 3873
rect 2976 3827 2983 3913
rect 2913 3787 2927 3793
rect 2953 3787 2967 3793
rect 2876 3656 2893 3667
rect 2880 3653 2893 3656
rect 2896 3547 2903 3613
rect 2933 3527 2947 3533
rect 2827 3476 2843 3487
rect 2827 3473 2840 3476
rect 2816 3247 2823 3393
rect 2887 3273 2893 3287
rect 2916 3248 2923 3333
rect 2936 3243 2943 3513
rect 2993 3267 3007 3273
rect 2936 3236 2953 3243
rect 2753 3227 2767 3233
rect 2713 2967 2727 2973
rect 2816 2967 2823 3233
rect 2853 3227 2867 3233
rect 2807 2956 2823 2967
rect 2807 2953 2820 2956
rect 2556 2807 2563 2893
rect 2653 2767 2667 2773
rect 2493 2747 2507 2753
rect 2656 2587 2663 2753
rect 2707 2713 2713 2727
rect 2756 2687 2763 2713
rect 2836 2687 2843 3053
rect 2860 2983 2873 2987
rect 2856 2973 2873 2983
rect 2856 2947 2863 2973
rect 2916 2967 2923 3212
rect 2956 3067 2963 3233
rect 3016 3167 3023 4016
rect 3073 4008 3087 4013
rect 3033 3987 3047 3993
rect 3056 3827 3063 3913
rect 3056 3543 3063 3813
rect 3076 3787 3083 3972
rect 3116 3967 3123 4053
rect 3196 3987 3203 4073
rect 3336 4067 3343 4193
rect 3356 4167 3363 4193
rect 3293 4047 3307 4053
rect 3213 4007 3227 4013
rect 3256 3967 3263 4013
rect 3296 3967 3303 4033
rect 3336 4007 3343 4053
rect 3393 4023 3407 4033
rect 3367 4020 3407 4023
rect 3367 4016 3403 4020
rect 3156 3887 3163 3933
rect 3056 3536 3083 3543
rect 3047 3514 3053 3527
rect 3040 3513 3053 3514
rect 3033 3487 3047 3492
rect 3076 3487 3083 3536
rect 3096 3487 3103 3773
rect 3156 3767 3163 3833
rect 3176 3827 3183 3893
rect 3216 3807 3223 3873
rect 3247 3813 3253 3827
rect 3193 3747 3207 3753
rect 3196 3687 3203 3733
rect 3236 3663 3243 3813
rect 3276 3787 3283 3933
rect 3296 3847 3303 3953
rect 3356 3907 3363 3973
rect 3327 3773 3333 3787
rect 3196 3656 3243 3663
rect 3173 3507 3187 3513
rect 3096 3476 3113 3487
rect 3100 3473 3113 3476
rect 3076 3427 3083 3473
rect 3036 3247 3043 3353
rect 3096 3287 3103 3433
rect 3156 3307 3163 3393
rect 3196 3347 3203 3656
rect 3356 3647 3363 3833
rect 3376 3827 3383 3993
rect 3396 3907 3403 3973
rect 3416 3848 3423 4353
rect 3433 4347 3447 4353
rect 3456 4323 3463 4473
rect 3476 4347 3483 4533
rect 3536 4527 3543 4936
rect 3556 4547 3563 5053
rect 3636 5027 3643 5153
rect 3680 5103 3693 5107
rect 3676 5093 3693 5103
rect 3656 4928 3663 5093
rect 3676 4947 3683 5093
rect 3713 5047 3727 5053
rect 3713 4983 3727 4993
rect 3696 4980 3727 4983
rect 3696 4976 3723 4980
rect 3696 4907 3703 4976
rect 3736 4967 3743 5193
rect 3776 5167 3783 5213
rect 3753 5087 3767 5093
rect 3796 5087 3803 5133
rect 3753 5067 3767 5073
rect 3766 5060 3767 5067
rect 3773 5053 3774 5060
rect 3773 5047 3787 5053
rect 3816 5047 3823 5113
rect 3856 5063 3863 5353
rect 3873 5327 3887 5333
rect 3916 5327 3923 5413
rect 4153 5387 4167 5393
rect 4107 5373 4113 5387
rect 3956 5287 3963 5373
rect 3836 5056 3863 5063
rect 3656 4867 3663 4892
rect 3796 4867 3803 5013
rect 3836 4883 3843 5056
rect 3856 5007 3863 5033
rect 3876 5003 3883 5133
rect 3896 5107 3903 5173
rect 3956 5087 3963 5213
rect 3996 5187 4003 5353
rect 4016 5347 4023 5373
rect 4293 5367 4307 5373
rect 4016 5227 4023 5333
rect 4033 5307 4047 5313
rect 3976 5087 3983 5133
rect 4036 5087 4043 5293
rect 4007 5073 4013 5087
rect 3913 5067 3927 5073
rect 4013 5047 4027 5052
rect 4076 5047 4083 5213
rect 4096 5187 4103 5333
rect 4133 5327 4147 5333
rect 4176 5207 4183 5313
rect 4196 5128 4203 5353
rect 4316 5327 4323 5473
rect 4376 5427 4383 5523
rect 4416 5467 4423 5523
rect 4436 5516 4463 5523
rect 4416 5387 4423 5413
rect 4227 5313 4233 5327
rect 4116 5047 4123 5113
rect 3867 4996 3883 5003
rect 3936 4967 3943 5033
rect 3976 4967 3983 5033
rect 3816 4876 3843 4883
rect 3613 4847 3627 4853
rect 3596 4836 3613 4843
rect 3576 4787 3583 4813
rect 3576 4547 3583 4693
rect 3596 4527 3603 4836
rect 3633 4807 3647 4813
rect 3673 4807 3687 4813
rect 3676 4687 3683 4713
rect 3696 4667 3703 4853
rect 3747 4833 3753 4847
rect 3816 4827 3823 4876
rect 3807 4816 3823 4827
rect 3807 4813 3820 4816
rect 3793 4807 3807 4813
rect 3776 4796 3793 4803
rect 3736 4703 3743 4733
rect 3716 4696 3743 4703
rect 3616 4568 3623 4593
rect 3653 4547 3667 4553
rect 3556 4447 3563 4493
rect 3596 4487 3603 4513
rect 3616 4507 3623 4532
rect 3696 4527 3703 4653
rect 3716 4547 3723 4696
rect 3736 4587 3743 4653
rect 3776 4607 3783 4796
rect 3836 4667 3843 4853
rect 3856 4787 3863 4953
rect 3896 4867 3903 4933
rect 3773 4587 3787 4593
rect 3687 4516 3703 4527
rect 3687 4513 3700 4516
rect 3633 4503 3647 4513
rect 3633 4500 3663 4503
rect 3636 4496 3663 4500
rect 3436 4316 3463 4323
rect 3436 4048 3443 4316
rect 3516 4307 3523 4333
rect 3456 4247 3463 4293
rect 3493 4287 3507 4293
rect 3516 4267 3523 4293
rect 3436 3987 3443 4012
rect 3456 3927 3463 4093
rect 3496 4047 3503 4133
rect 3536 4107 3543 4393
rect 3567 4293 3573 4307
rect 3556 4147 3563 4233
rect 3576 4047 3583 4153
rect 3596 4048 3603 4433
rect 3616 4287 3623 4313
rect 3636 4307 3643 4473
rect 3656 4447 3663 4496
rect 3696 4407 3703 4453
rect 3716 4427 3723 4533
rect 3656 4307 3663 4353
rect 3687 4333 3693 4347
rect 3736 4323 3743 4573
rect 3813 4527 3827 4533
rect 3876 4527 3883 4753
rect 3896 4587 3903 4793
rect 3936 4707 3943 4793
rect 3956 4747 3963 4893
rect 4016 4867 4023 4993
rect 4036 4907 4043 5013
rect 4196 4967 4203 5092
rect 4216 5027 4223 5193
rect 4236 5007 4243 5093
rect 4053 4867 4067 4873
rect 4236 4868 4243 4913
rect 3973 4847 3987 4853
rect 4036 4767 4043 4813
rect 3916 4567 3923 4593
rect 3996 4567 4003 4593
rect 4076 4567 4083 4813
rect 4136 4707 4143 4833
rect 4173 4807 4187 4813
rect 4236 4767 4243 4832
rect 3787 4494 3793 4507
rect 3780 4493 3800 4494
rect 3796 4387 3803 4472
rect 3816 4347 3823 4393
rect 3836 4387 3843 4493
rect 3876 4447 3883 4513
rect 3736 4316 3763 4323
rect 3656 4296 3673 4307
rect 3660 4293 3673 4296
rect 3673 4287 3687 4293
rect 3616 4247 3623 4273
rect 3636 4240 3683 4243
rect 3633 4236 3683 4240
rect 3633 4227 3647 4236
rect 3567 4036 3583 4047
rect 3567 4033 3580 4036
rect 3420 3826 3440 3827
rect 3427 3813 3433 3826
rect 3476 3783 3483 4033
rect 3536 4007 3543 4033
rect 3616 4027 3623 4113
rect 3676 4107 3683 4236
rect 3696 4087 3703 4253
rect 3716 4147 3723 4293
rect 3756 4283 3763 4316
rect 3736 4280 3763 4283
rect 3733 4276 3763 4280
rect 3796 4283 3803 4333
rect 3867 4313 3873 4327
rect 3833 4287 3847 4293
rect 3896 4287 3903 4533
rect 3956 4527 3963 4553
rect 3927 4513 3933 4527
rect 3796 4280 3823 4283
rect 3796 4276 3827 4280
rect 3733 4267 3747 4276
rect 3813 4267 3827 4276
rect 3916 4267 3923 4373
rect 3956 4327 3963 4513
rect 3933 4287 3947 4293
rect 3976 4287 3983 4413
rect 3996 4307 4003 4453
rect 4036 4387 4043 4553
rect 4156 4527 4163 4653
rect 4200 4564 4213 4567
rect 4196 4554 4213 4564
rect 4196 4553 4220 4554
rect 4176 4528 4183 4553
rect 4107 4513 4113 4527
rect 4076 4487 4083 4513
rect 4056 4447 4063 4473
rect 3693 4067 3707 4073
rect 3633 4027 3647 4033
rect 3496 3827 3503 3993
rect 3556 3887 3563 3973
rect 3596 3907 3603 4012
rect 3556 3827 3563 3873
rect 3516 3787 3523 3813
rect 3616 3803 3623 4013
rect 3656 3947 3663 4053
rect 3716 4047 3723 4133
rect 3753 4087 3767 4093
rect 3773 4027 3787 4033
rect 3636 3827 3643 3893
rect 3616 3796 3643 3803
rect 3447 3776 3483 3783
rect 3396 3727 3403 3753
rect 3216 3507 3223 3553
rect 3196 3307 3203 3333
rect 3127 3253 3133 3267
rect 3173 3247 3187 3253
rect 3076 3207 3083 3233
rect 3236 3167 3243 3633
rect 3293 3487 3307 3493
rect 3336 3487 3343 3593
rect 3356 3507 3363 3553
rect 3447 3493 3453 3507
rect 3336 3343 3343 3413
rect 3416 3387 3423 3493
rect 3476 3487 3483 3776
rect 3607 3774 3613 3787
rect 3600 3773 3613 3774
rect 3496 3667 3503 3773
rect 3533 3767 3547 3773
rect 3533 3487 3547 3493
rect 3316 3336 3343 3343
rect 3273 3267 3287 3273
rect 3296 3243 3303 3293
rect 3316 3267 3323 3336
rect 3436 3307 3443 3353
rect 3347 3293 3353 3307
rect 3296 3236 3323 3243
rect 2536 2467 2543 2493
rect 2547 2453 2553 2467
rect 2556 2347 2563 2453
rect 2513 2247 2527 2253
rect 2476 2236 2503 2243
rect 2456 2207 2463 2233
rect 2407 2193 2413 2207
rect 2456 2067 2463 2193
rect 2496 2167 2503 2236
rect 2127 1953 2133 1967
rect 2096 1927 2103 1953
rect 2276 1947 2283 1973
rect 2516 1967 2523 2013
rect 2467 1953 2473 1967
rect 2147 1913 2153 1927
rect 2187 1913 2193 1927
rect 1720 1443 1733 1447
rect 1716 1433 1733 1443
rect 1716 1407 1723 1433
rect 1753 1427 1767 1432
rect 1716 1207 1723 1313
rect 1716 1167 1723 1193
rect 1756 1147 1763 1413
rect 1776 1327 1783 1533
rect 1796 1227 1803 1453
rect 1816 1307 1823 1453
rect 1896 1448 1903 1513
rect 1847 1433 1853 1447
rect 1867 1393 1873 1407
rect 1813 1187 1827 1193
rect 1896 1187 1903 1412
rect 1916 1208 1923 1473
rect 1936 1428 1943 1613
rect 2007 1433 2013 1447
rect 1956 1407 1963 1433
rect 2056 1423 2063 1893
rect 2073 1747 2087 1753
rect 2196 1748 2203 1833
rect 2276 1767 2283 1933
rect 2313 1927 2327 1933
rect 2467 1923 2480 1927
rect 2467 1913 2483 1923
rect 2507 1913 2513 1927
rect 2476 1847 2483 1913
rect 2153 1728 2167 1733
rect 2147 1706 2160 1707
rect 2147 1693 2153 1706
rect 2096 1627 2103 1693
rect 2173 1687 2187 1693
rect 2196 1527 2203 1712
rect 2256 1647 2263 1713
rect 2287 1673 2293 1687
rect 2167 1433 2173 1447
rect 2036 1416 2063 1423
rect 1940 1406 1963 1407
rect 1947 1396 1963 1406
rect 1947 1393 1960 1396
rect 1936 1227 1943 1333
rect 1976 1307 1983 1413
rect 2036 1367 2043 1416
rect 1976 1187 1983 1233
rect 2013 1207 2027 1213
rect 1867 1173 1873 1187
rect 1681 936 1683 947
rect 1713 947 1727 953
rect 1876 947 1883 1013
rect 1820 943 1833 947
rect 1753 927 1767 933
rect 1816 933 1833 943
rect 1816 907 1823 933
rect 1916 927 1923 1172
rect 1976 1007 1983 1173
rect 2016 1067 2023 1193
rect 2036 1187 2043 1353
rect 2056 1327 2063 1393
rect 2053 1227 2067 1233
rect 2176 1227 2183 1353
rect 2196 1208 2203 1413
rect 2273 1387 2287 1393
rect 2336 1387 2343 1673
rect 2376 1488 2383 1833
rect 2576 1827 2583 2433
rect 2656 2407 2663 2473
rect 2687 2453 2693 2467
rect 2596 2247 2603 2333
rect 2596 2207 2603 2233
rect 2636 2127 2643 2213
rect 2596 1927 2603 2073
rect 2656 1987 2663 2053
rect 2627 1963 2640 1967
rect 2627 1953 2643 1963
rect 2396 1707 2403 1733
rect 2456 1587 2463 1793
rect 2476 1727 2483 1753
rect 2513 1707 2527 1713
rect 2613 1687 2627 1693
rect 2396 1467 2403 1513
rect 2380 1466 2403 1467
rect 2387 1455 2403 1466
rect 2413 1467 2427 1473
rect 2387 1453 2400 1455
rect 2267 1214 2273 1227
rect 2260 1213 2280 1214
rect 2107 1193 2113 1207
rect 2113 1187 2127 1193
rect 2273 1187 2287 1192
rect 2067 1173 2073 1187
rect 2180 1186 2200 1187
rect 2127 1176 2143 1183
rect 1607 893 1613 907
rect 1487 876 1503 887
rect 1487 873 1500 876
rect 1447 676 1463 687
rect 1447 673 1460 676
rect 1116 647 1123 673
rect 1153 647 1167 652
rect 1036 407 1043 533
rect 976 396 1003 403
rect 976 307 983 396
rect 1087 394 1093 407
rect 1087 393 1100 394
rect 1093 367 1107 372
rect 1013 347 1027 353
rect 447 173 453 187
rect 473 147 487 153
rect 516 147 523 193
rect 727 173 733 187
rect 767 173 773 187
rect 413 127 427 133
rect 476 87 483 133
rect 556 87 563 173
rect 593 167 607 173
rect 796 147 803 193
rect 856 187 863 293
rect 893 187 907 193
rect 1027 153 1033 167
rect 953 147 967 153
rect 1116 148 1123 513
rect 1276 507 1283 673
rect 1476 667 1483 873
rect 1553 707 1567 713
rect 1627 693 1633 707
rect 1516 667 1523 693
rect 1653 667 1667 673
rect 1567 653 1573 667
rect 1627 653 1633 667
rect 1736 647 1743 693
rect 1727 636 1743 647
rect 1727 633 1740 636
rect 1236 467 1243 493
rect 1193 387 1207 393
rect 1236 387 1243 453
rect 1313 367 1327 373
rect 1336 347 1343 453
rect 1376 427 1383 553
rect 1436 427 1443 453
rect 1353 387 1367 393
rect 1376 367 1383 413
rect 1556 407 1563 493
rect 1616 407 1623 593
rect 1716 467 1723 633
rect 1756 507 1763 693
rect 1836 567 1843 673
rect 1796 527 1803 553
rect 1856 447 1863 893
rect 1916 707 1923 753
rect 1936 667 1943 993
rect 1953 907 1967 913
rect 1976 887 1983 953
rect 1973 687 1987 693
rect 1996 667 2003 933
rect 2016 907 2023 1013
rect 2136 927 2143 1176
rect 2187 1173 2193 1186
rect 2247 1173 2253 1187
rect 2216 947 2223 1053
rect 2256 947 2263 1133
rect 2296 1087 2303 1173
rect 2316 1147 2323 1213
rect 2356 1127 2363 1413
rect 2456 1407 2463 1573
rect 2476 1527 2483 1673
rect 2636 1647 2643 1953
rect 2676 1927 2683 1953
rect 2696 1927 2703 2113
rect 2716 1767 2723 2673
rect 2776 2447 2783 2473
rect 2816 2407 2823 2433
rect 2836 2407 2843 2493
rect 2856 2463 2863 2933
rect 2936 2803 2943 2993
rect 3036 2808 3043 2973
rect 3073 2967 3087 2973
rect 3176 2967 3183 3153
rect 3236 2987 3243 3053
rect 3296 3027 3303 3193
rect 3316 3147 3323 3236
rect 3336 3047 3343 3093
rect 3356 3087 3363 3193
rect 3396 3187 3403 3293
rect 3456 3267 3463 3433
rect 3556 3367 3563 3513
rect 3596 3507 3603 3752
rect 3636 3561 3643 3796
rect 3656 3627 3663 3933
rect 3736 3887 3743 4013
rect 3753 3827 3767 3833
rect 3696 3727 3703 3813
rect 3776 3787 3783 3853
rect 3796 3827 3803 4013
rect 3836 4007 3843 4233
rect 3856 4067 3863 4133
rect 3836 3867 3843 3993
rect 3876 3848 3883 4173
rect 3916 4067 3923 4213
rect 4016 4147 4023 4313
rect 4056 4307 4063 4333
rect 4093 4327 4107 4333
rect 4116 4307 4123 4373
rect 4156 4363 4163 4513
rect 4176 4407 4183 4492
rect 4196 4407 4203 4553
rect 4213 4527 4227 4532
rect 4236 4447 4243 4673
rect 4136 4356 4163 4363
rect 4096 4296 4113 4303
rect 4076 4267 4083 4293
rect 4013 4067 4027 4073
rect 3967 4053 3973 4067
rect 3913 4047 3927 4053
rect 4056 4027 4063 4093
rect 4096 4067 4103 4296
rect 4136 4263 4143 4356
rect 4167 4333 4173 4347
rect 4236 4327 4243 4393
rect 4256 4367 4263 5253
rect 4276 5207 4283 5313
rect 4356 5307 4363 5373
rect 4276 5067 4283 5153
rect 4293 5107 4307 5113
rect 4296 4847 4303 4953
rect 4276 4487 4283 4813
rect 4296 4807 4303 4833
rect 4336 4827 4343 5093
rect 4356 5067 4363 5293
rect 4393 5087 4407 5093
rect 4396 5007 4403 5073
rect 4416 4987 4423 5373
rect 4436 5267 4443 5516
rect 4436 5067 4443 5113
rect 4393 4867 4407 4873
rect 4327 4813 4333 4827
rect 4393 4807 4407 4813
rect 4433 4807 4447 4813
rect 4356 4607 4363 4733
rect 4296 4407 4303 4573
rect 4347 4553 4353 4567
rect 4313 4527 4327 4533
rect 4396 4527 4403 4593
rect 4456 4547 4463 4833
rect 4476 4647 4483 5453
rect 4796 5440 4843 5443
rect 4793 5436 4843 5440
rect 4793 5427 4807 5436
rect 4806 5420 4807 5427
rect 4813 5413 4814 5420
rect 4696 5387 4703 5413
rect 4813 5407 4827 5413
rect 4836 5403 4843 5436
rect 4836 5396 4903 5403
rect 4896 5387 4903 5396
rect 4936 5387 4943 5413
rect 4587 5373 4593 5387
rect 4896 5376 4913 5387
rect 4900 5373 4913 5376
rect 4733 5367 4747 5373
rect 4533 5348 4547 5353
rect 4733 5347 4747 5353
rect 4496 5267 4503 5313
rect 4533 5307 4547 5312
rect 4576 5267 4583 5333
rect 4496 5167 4503 5253
rect 4533 5107 4547 5113
rect 4493 5087 4507 5093
rect 4553 5067 4567 5073
rect 4493 5027 4507 5033
rect 4576 4927 4583 5173
rect 4516 4827 4523 4913
rect 4596 4867 4603 5093
rect 4616 5027 4623 5333
rect 4773 5327 4787 5333
rect 4807 5313 4813 5327
rect 4776 5187 4783 5313
rect 4836 5148 4843 5353
rect 4876 5327 4883 5373
rect 4916 5347 4923 5373
rect 4936 5347 4943 5373
rect 4976 5367 4983 5433
rect 5336 5416 5433 5423
rect 5196 5400 5253 5403
rect 5193 5396 5253 5400
rect 5193 5387 5207 5396
rect 4973 5347 4987 5353
rect 4867 5316 4883 5327
rect 4867 5313 4880 5316
rect 4753 5087 4767 5093
rect 4633 5067 4647 5073
rect 4676 5047 4683 5073
rect 4727 5033 4733 5047
rect 4556 4827 4563 4853
rect 4573 4847 4587 4853
rect 4476 4547 4483 4573
rect 4416 4523 4423 4539
rect 4447 4533 4463 4547
rect 4416 4516 4443 4523
rect 4436 4347 4443 4516
rect 4456 4427 4463 4533
rect 4496 4387 4503 4733
rect 4520 4603 4533 4607
rect 4516 4593 4533 4603
rect 4516 4507 4523 4593
rect 4616 4587 4623 4893
rect 4636 4707 4643 4853
rect 4656 4747 4663 5033
rect 4693 5027 4707 5033
rect 4696 4887 4703 5013
rect 4696 4767 4703 4873
rect 4756 4827 4763 4973
rect 4796 4887 4803 5073
rect 4716 4627 4723 4813
rect 4776 4687 4783 4853
rect 4816 4787 4823 4853
rect 4836 4827 4843 5112
rect 4996 5107 5003 5373
rect 5056 5347 5063 5373
rect 5076 5347 5083 5373
rect 5233 5367 5247 5373
rect 5336 5367 5343 5416
rect 5356 5368 5363 5393
rect 5373 5347 5387 5353
rect 5227 5343 5240 5347
rect 5227 5333 5243 5343
rect 4873 5087 4887 5093
rect 4976 5096 4993 5103
rect 4853 5047 4867 5053
rect 4896 4947 4903 5033
rect 4816 4727 4823 4773
rect 4673 4588 4687 4593
rect 4540 4564 4553 4567
rect 4536 4554 4553 4564
rect 4680 4566 4693 4567
rect 4536 4553 4560 4554
rect 4536 4347 4543 4553
rect 4687 4554 4693 4566
rect 4687 4553 4700 4554
rect 4560 4546 4573 4547
rect 4567 4533 4573 4546
rect 4700 4546 4713 4547
rect 4707 4533 4713 4546
rect 4487 4333 4493 4347
rect 4136 4256 4163 4263
rect 4156 4167 4163 4256
rect 4156 4067 4163 4153
rect 4196 4087 4203 4273
rect 4147 4056 4163 4067
rect 4147 4053 4160 4056
rect 3813 3787 3827 3793
rect 3776 3727 3783 3773
rect 3836 3747 3843 3813
rect 3876 3747 3883 3812
rect 3896 3787 3903 3993
rect 3916 3827 3923 3973
rect 3976 3827 3983 3873
rect 4016 3827 4023 4013
rect 4176 3987 4183 4053
rect 4196 4007 4203 4073
rect 4216 4067 4223 4293
rect 4267 4273 4273 4287
rect 4276 4067 4283 4193
rect 4213 4047 4227 4053
rect 4316 4047 4323 4273
rect 4353 4047 4367 4053
rect 4307 4033 4313 4047
rect 4233 4027 4247 4033
rect 4016 3816 4033 3827
rect 4020 3813 4033 3816
rect 3936 3787 3943 3813
rect 3896 3776 3913 3787
rect 3900 3773 3913 3776
rect 4007 3773 4013 3787
rect 3953 3767 3967 3773
rect 3656 3547 3663 3573
rect 3656 3536 3673 3547
rect 3660 3533 3673 3536
rect 3716 3508 3723 3673
rect 3596 3367 3603 3493
rect 3716 3447 3723 3472
rect 3516 3267 3523 3333
rect 3567 3273 3573 3287
rect 3427 3253 3433 3267
rect 3596 3247 3603 3313
rect 3167 2953 3173 2967
rect 3076 2827 3083 2953
rect 3256 2907 3263 3013
rect 3296 2987 3303 3013
rect 3376 3007 3383 3093
rect 3416 3007 3423 3053
rect 3353 2967 3367 2973
rect 3396 2887 3403 2953
rect 3436 2947 3443 3153
rect 3476 2967 3483 2993
rect 3496 2967 3503 3093
rect 3616 3047 3623 3253
rect 3636 3207 3643 3293
rect 3656 3267 3663 3413
rect 3696 3227 3703 3293
rect 3736 3267 3743 3713
rect 3756 3527 3763 3613
rect 3776 3588 3783 3713
rect 3776 3527 3783 3552
rect 3796 3487 3803 3733
rect 4076 3687 4083 3973
rect 4196 3963 4203 3993
rect 4176 3956 4203 3963
rect 4136 3827 4143 3873
rect 4107 3793 4113 3807
rect 4176 3787 4183 3956
rect 4236 3927 4243 4013
rect 4396 4007 4403 4333
rect 4436 4207 4443 4333
rect 4556 4307 4563 4373
rect 4607 4333 4613 4347
rect 4656 4307 4663 4413
rect 4736 4307 4743 4573
rect 4756 4527 4763 4573
rect 4796 4487 4803 4593
rect 4796 4347 4803 4473
rect 4816 4407 4823 4553
rect 4753 4327 4767 4333
rect 4836 4328 4843 4533
rect 4876 4307 4883 4393
rect 4896 4363 4903 4693
rect 4916 4667 4923 5073
rect 4947 5033 4953 5047
rect 4976 4963 4983 5096
rect 5036 5087 5043 5313
rect 5116 5287 5123 5333
rect 5076 5087 5083 5113
rect 5007 5033 5013 5047
rect 4956 4956 4983 4963
rect 4956 4847 4963 4956
rect 4976 4867 4983 4933
rect 4976 4827 4983 4853
rect 5056 4843 5063 5033
rect 5096 4847 5103 5153
rect 5116 5127 5123 5273
rect 5176 5007 5183 5093
rect 5196 5088 5203 5293
rect 5236 5148 5243 5333
rect 5360 5346 5373 5347
rect 5293 5327 5307 5333
rect 5367 5333 5373 5346
rect 5416 5347 5423 5393
rect 5496 5387 5503 5413
rect 5453 5367 5467 5373
rect 5416 5336 5433 5347
rect 5420 5333 5433 5336
rect 5473 5327 5487 5333
rect 5336 5167 5343 5313
rect 5393 5307 5407 5313
rect 5220 5126 5240 5127
rect 5227 5113 5233 5126
rect 5296 5087 5303 5133
rect 5336 5087 5343 5113
rect 5207 5074 5213 5087
rect 5200 5073 5213 5074
rect 5293 5067 5307 5073
rect 5193 5047 5207 5052
rect 5316 5047 5323 5073
rect 5376 5047 5383 5073
rect 5396 5047 5403 5293
rect 5447 5073 5453 5087
rect 5507 5083 5520 5087
rect 5507 5073 5523 5083
rect 5176 4867 5183 4993
rect 5436 4967 5443 5033
rect 5036 4836 5063 4843
rect 4933 4807 4947 4813
rect 4936 4587 4943 4793
rect 4913 4563 4927 4573
rect 4976 4567 4983 4813
rect 4996 4667 5003 4773
rect 4913 4560 4953 4563
rect 4916 4556 4953 4560
rect 4976 4556 4993 4567
rect 4980 4553 4993 4556
rect 5016 4527 5023 4573
rect 4927 4513 4933 4527
rect 4987 4513 4993 4527
rect 5036 4503 5043 4836
rect 5067 4813 5073 4827
rect 5067 4773 5073 4787
rect 5080 4543 5093 4547
rect 5076 4540 5093 4543
rect 5073 4533 5093 4540
rect 5073 4527 5087 4533
rect 5116 4527 5123 4793
rect 5176 4787 5183 4853
rect 5247 4833 5253 4847
rect 5287 4833 5293 4847
rect 5207 4813 5213 4827
rect 5336 4807 5343 4893
rect 5476 4848 5483 5033
rect 5516 5007 5523 5073
rect 5467 4834 5473 4847
rect 5467 4833 5480 4834
rect 5496 4827 5503 4893
rect 5480 4826 5503 4827
rect 5487 4815 5503 4826
rect 5487 4813 5500 4815
rect 5476 4803 5483 4812
rect 5456 4796 5483 4803
rect 5176 4776 5193 4787
rect 5180 4773 5193 4776
rect 5276 4587 5283 4793
rect 5373 4787 5387 4793
rect 5416 4587 5423 4793
rect 5266 4573 5267 4580
rect 5347 4573 5353 4587
rect 5407 4576 5423 4587
rect 5407 4573 5420 4576
rect 5253 4567 5267 4573
rect 5147 4553 5153 4567
rect 5393 4567 5407 4573
rect 5436 4567 5443 4773
rect 5213 4547 5227 4553
rect 5187 4513 5193 4527
rect 5036 4496 5063 4503
rect 4896 4356 4923 4363
rect 4893 4327 4907 4333
rect 4473 4287 4487 4293
rect 4656 4296 4673 4307
rect 4660 4293 4673 4296
rect 4513 4287 4527 4293
rect 4633 4287 4647 4293
rect 4836 4267 4843 4292
rect 4836 4256 4853 4267
rect 4840 4253 4853 4256
rect 4456 4047 4463 4093
rect 4476 4047 4483 4193
rect 4507 4043 4520 4047
rect 4507 4033 4523 4043
rect 4476 4007 4483 4033
rect 4327 3993 4333 4007
rect 4193 3787 4207 3793
rect 4236 3783 4243 3813
rect 4336 3807 4343 3913
rect 4436 3827 4443 3973
rect 4516 3927 4523 4033
rect 4367 3813 4373 3827
rect 4236 3776 4263 3783
rect 4153 3767 4167 3773
rect 3816 3287 3823 3573
rect 3836 3567 3843 3653
rect 3836 3487 3843 3513
rect 3856 3347 3863 3513
rect 3873 3487 3887 3493
rect 3896 3363 3903 3613
rect 3916 3547 3923 3593
rect 3936 3567 3943 3633
rect 3953 3527 3967 3533
rect 3927 3493 3933 3507
rect 3996 3467 4003 3533
rect 4036 3483 4043 3653
rect 4087 3533 4093 3547
rect 4016 3476 4043 3483
rect 3887 3356 3903 3363
rect 3876 3307 3883 3353
rect 3867 3296 3883 3307
rect 3867 3293 3880 3296
rect 3787 3273 3793 3287
rect 3916 3267 3923 3453
rect 4016 3427 4023 3476
rect 4036 3327 4043 3453
rect 4056 3447 4063 3533
rect 4156 3523 4163 3753
rect 4176 3607 4183 3773
rect 4233 3747 4247 3753
rect 4196 3527 4203 3713
rect 4256 3587 4263 3776
rect 4296 3767 4303 3793
rect 4233 3527 4247 3533
rect 4147 3516 4163 3523
rect 4133 3507 4147 3513
rect 4253 3487 4267 3493
rect 4176 3407 4183 3473
rect 3736 3107 3743 3253
rect 4036 3247 4043 3313
rect 4176 3307 4183 3353
rect 4053 3287 4067 3293
rect 4116 3247 4123 3293
rect 4133 3267 4147 3273
rect 4176 3267 4183 3293
rect 4276 3283 4283 3673
rect 4396 3627 4403 3773
rect 4433 3767 4447 3773
rect 4396 3547 4403 3613
rect 4353 3507 4367 3513
rect 4436 3507 4443 3713
rect 4476 3647 4483 3793
rect 4536 3687 4543 4153
rect 4593 4087 4607 4093
rect 4607 4034 4613 4047
rect 4600 4033 4613 4034
rect 4593 4007 4607 4012
rect 4636 3927 4643 4013
rect 4576 3707 4583 3813
rect 4616 3727 4623 3753
rect 4476 3547 4483 3573
rect 4316 3367 4323 3493
rect 4393 3487 4407 3493
rect 4373 3307 4387 3313
rect 4333 3287 4347 3293
rect 4436 3287 4443 3493
rect 4496 3307 4503 3533
rect 4516 3507 4523 3533
rect 4556 3527 4563 3573
rect 4573 3487 4587 3493
rect 4276 3276 4303 3283
rect 4193 3267 4207 3273
rect 4267 3254 4273 3267
rect 4267 3253 4280 3254
rect 3967 3233 3973 3247
rect 4027 3236 4043 3247
rect 4027 3233 4040 3236
rect 4153 3227 4167 3233
rect 3876 3007 3883 3093
rect 4276 3047 4283 3232
rect 4253 3007 4267 3013
rect 4207 2993 4213 3007
rect 2916 2800 2943 2803
rect 2873 2787 2887 2793
rect 2913 2796 2943 2800
rect 2913 2787 2927 2796
rect 3036 2743 3043 2772
rect 3233 2767 3247 2773
rect 3016 2740 3043 2743
rect 3013 2736 3043 2740
rect 3053 2747 3067 2753
rect 2896 2687 2903 2733
rect 3013 2727 3027 2736
rect 2976 2663 2983 2713
rect 3016 2667 3023 2713
rect 2956 2656 2983 2663
rect 2873 2487 2887 2493
rect 2956 2487 2963 2656
rect 3136 2647 3143 2753
rect 3207 2733 3213 2747
rect 3253 2727 3267 2733
rect 3276 2667 3283 2773
rect 3416 2767 3423 2813
rect 3436 2787 3443 2933
rect 3616 2927 3623 2993
rect 3656 2807 3663 2973
rect 3747 2953 3753 2967
rect 3493 2767 3507 2773
rect 3613 2767 3627 2773
rect 3707 2753 3713 2767
rect 3373 2747 3387 2753
rect 3593 2727 3607 2733
rect 3633 2727 3647 2733
rect 3136 2567 3143 2633
rect 3267 2473 3273 2487
rect 2856 2456 2883 2463
rect 2816 2227 2823 2273
rect 2876 2267 2883 2456
rect 2893 2447 2907 2453
rect 2916 2447 2923 2473
rect 3027 2453 3033 2467
rect 3076 2427 3083 2473
rect 3093 2447 3107 2453
rect 2953 2407 2967 2413
rect 3076 2367 3083 2413
rect 2973 2267 2987 2273
rect 2947 2263 2960 2267
rect 2947 2253 2963 2263
rect 2856 2207 2863 2233
rect 2856 2107 2863 2193
rect 2876 2127 2883 2253
rect 2956 2207 2963 2253
rect 3036 2227 3043 2293
rect 3053 2247 3067 2253
rect 3096 2247 3103 2433
rect 3116 2347 3123 2473
rect 3156 2447 3163 2473
rect 3296 2467 3303 2513
rect 3113 2287 3127 2293
rect 3196 2287 3203 2333
rect 3187 2233 3193 2247
rect 2747 1953 2753 1967
rect 2776 1847 2783 1973
rect 2836 1963 2843 2013
rect 2853 1987 2867 1993
rect 2836 1960 2863 1963
rect 2836 1956 2867 1960
rect 2796 1887 2803 1953
rect 2853 1947 2867 1956
rect 2827 1913 2833 1927
rect 2696 1687 2703 1733
rect 2716 1647 2723 1693
rect 2636 1640 2723 1647
rect 2716 1567 2723 1640
rect 2736 1587 2743 1733
rect 2773 1727 2787 1733
rect 2836 1707 2843 1873
rect 2856 1747 2863 1793
rect 2847 1694 2853 1707
rect 2847 1693 2860 1694
rect 2793 1687 2807 1693
rect 2476 1447 2483 1473
rect 2527 1443 2540 1447
rect 2527 1433 2543 1443
rect 2496 1407 2503 1433
rect 2536 1407 2543 1433
rect 2456 1267 2463 1393
rect 2576 1387 2583 1433
rect 2656 1407 2663 1433
rect 2716 1407 2723 1553
rect 2787 1433 2793 1447
rect 2816 1427 2823 1593
rect 2836 1487 2843 1693
rect 2856 1587 2863 1672
rect 2876 1647 2883 1913
rect 2896 1907 2903 1973
rect 2916 1863 2923 2113
rect 2936 1927 2943 2073
rect 2967 1953 2973 1967
rect 2936 1916 2953 1927
rect 2940 1913 2953 1916
rect 2896 1856 2923 1863
rect 2896 1607 2903 1856
rect 2956 1783 2963 1913
rect 2956 1776 2983 1783
rect 2913 1767 2927 1773
rect 2927 1693 2933 1707
rect 2747 1393 2753 1407
rect 2376 947 2383 1213
rect 2396 1187 2403 1213
rect 2487 1193 2493 1207
rect 2516 1187 2523 1213
rect 2596 987 2603 1273
rect 2613 1187 2627 1193
rect 2676 1187 2683 1393
rect 2816 1287 2823 1413
rect 2856 1407 2863 1573
rect 2707 1213 2713 1227
rect 2707 1173 2713 1187
rect 2736 1147 2743 1233
rect 2827 1213 2833 1227
rect 2636 967 2643 993
rect 2320 943 2333 947
rect 2316 933 2333 943
rect 2756 943 2763 1193
rect 2856 1187 2863 1393
rect 2876 1228 2883 1573
rect 2956 1543 2963 1753
rect 2976 1587 2983 1776
rect 2996 1667 3003 2153
rect 3016 1968 3023 2013
rect 3013 1928 3027 1932
rect 3056 1923 3063 2133
rect 3076 2087 3083 2213
rect 3133 2207 3147 2213
rect 3236 2147 3243 2353
rect 3316 2307 3323 2433
rect 3373 2427 3387 2433
rect 3316 2247 3323 2293
rect 3416 2267 3423 2653
rect 3536 2467 3543 2513
rect 3496 2287 3503 2453
rect 3656 2447 3663 2473
rect 3713 2447 3727 2453
rect 3627 2433 3633 2447
rect 3533 2267 3547 2273
rect 3656 2267 3663 2433
rect 3567 2253 3573 2267
rect 3036 1916 3063 1923
rect 3016 1707 3023 1892
rect 3036 1807 3043 1916
rect 3073 1907 3087 1913
rect 3136 1867 3143 2013
rect 3156 1947 3163 2093
rect 3193 1947 3207 1953
rect 3156 1867 3163 1933
rect 3276 1887 3283 2233
rect 3416 2207 3423 2253
rect 3473 2227 3487 2233
rect 3507 2213 3513 2227
rect 3553 2207 3567 2213
rect 3387 2193 3393 2207
rect 3416 2196 3433 2207
rect 3420 2193 3433 2196
rect 3633 2207 3647 2213
rect 3367 1973 3373 1987
rect 3056 1747 3063 1853
rect 3147 1753 3153 1767
rect 3093 1728 3107 1733
rect 3133 1707 3147 1713
rect 3087 1706 3100 1707
rect 3087 1693 3093 1706
rect 3076 1567 3083 1693
rect 3173 1707 3187 1713
rect 3133 1687 3147 1693
rect 2956 1536 2983 1543
rect 2896 1323 2903 1433
rect 2896 1316 2923 1323
rect 2880 1206 2893 1207
rect 2887 1194 2893 1206
rect 2887 1193 2900 1194
rect 2861 1176 2863 1187
rect 2796 1147 2803 1173
rect 2876 1007 2883 1053
rect 2756 936 2783 943
rect 2153 887 2167 893
rect 2056 687 2063 873
rect 2176 827 2183 913
rect 2216 907 2223 933
rect 2256 827 2263 933
rect 2316 907 2323 933
rect 2467 914 2473 927
rect 2460 913 2473 914
rect 2527 913 2533 927
rect 2413 907 2427 913
rect 2553 907 2567 913
rect 2596 907 2603 933
rect 2453 887 2467 892
rect 2093 707 2107 713
rect 2127 693 2133 707
rect 2156 667 2163 753
rect 2193 667 2207 673
rect 1933 647 1947 653
rect 2013 647 2027 653
rect 1596 347 1603 373
rect 1676 367 1683 393
rect 1696 387 1703 413
rect 1256 167 1263 253
rect 1336 187 1343 333
rect 1207 156 1233 163
rect 1353 147 1367 153
rect 1396 147 1403 293
rect 1413 167 1427 173
rect 1556 167 1563 333
rect 1716 267 1723 413
rect 1773 407 1787 413
rect 1896 407 1903 433
rect 1916 427 1923 473
rect 2016 427 2023 473
rect 1847 393 1853 407
rect 1736 307 1743 373
rect 1916 367 1923 413
rect 1656 187 1663 253
rect 1796 247 1803 353
rect 1647 173 1663 187
rect 1513 147 1527 153
rect 673 127 687 133
rect 756 107 763 133
rect 833 127 847 133
rect 993 127 1007 133
rect 1213 127 1227 133
rect 1656 127 1663 173
rect 1756 147 1763 233
rect 1936 187 1943 413
rect 2136 407 2143 593
rect 2196 407 2203 653
rect 2236 407 2243 693
rect 2256 667 2263 733
rect 2456 707 2463 873
rect 2573 867 2587 873
rect 2287 693 2293 707
rect 2387 693 2393 707
rect 2276 487 2283 693
rect 2336 587 2343 673
rect 2436 667 2443 693
rect 2476 667 2483 713
rect 2616 687 2623 813
rect 2656 787 2663 933
rect 2747 924 2760 927
rect 2747 914 2763 924
rect 2740 913 2763 914
rect 2407 653 2413 667
rect 2467 656 2483 667
rect 2573 667 2587 673
rect 2467 653 2480 656
rect 2616 507 2623 673
rect 2696 667 2703 693
rect 2293 407 2307 413
rect 2493 407 2507 413
rect 1953 387 1967 393
rect 2236 396 2253 407
rect 2240 393 2253 396
rect 2093 387 2107 393
rect 2153 367 2167 373
rect 2336 367 2343 393
rect 2376 367 2383 393
rect 2536 387 2543 493
rect 2636 367 2643 413
rect 2267 353 2273 367
rect 2327 356 2343 367
rect 2327 353 2340 356
rect 2627 353 2633 367
rect 1956 187 1963 293
rect 2076 227 2083 353
rect 2116 247 2123 353
rect 2156 307 2163 353
rect 2393 347 2407 353
rect 2036 187 2043 213
rect 1887 173 1893 187
rect 1807 153 1813 167
rect 1936 147 1943 173
rect 1967 133 1973 147
rect 1087 113 1093 127
rect 1120 126 1133 127
rect 1127 113 1133 126
rect 967 93 973 107
rect 1176 87 1183 113
rect 1253 107 1267 113
rect 1996 67 2003 173
rect 2096 147 2103 193
rect 2113 167 2127 173
rect 2013 127 2027 133
rect 2116 107 2123 153
rect 2156 147 2163 213
rect 2187 173 2193 187
rect 2296 167 2303 333
rect 2287 153 2293 167
rect 2416 147 2423 173
rect 2256 87 2263 133
rect 2313 127 2327 133
rect 2436 67 2443 93
rect 2456 47 2463 233
rect 2496 187 2503 273
rect 2536 147 2543 213
rect 2616 147 2623 193
rect 2656 167 2663 493
rect 2716 467 2723 773
rect 2713 407 2727 413
rect 2736 388 2743 892
rect 2756 867 2763 913
rect 2776 907 2783 936
rect 2776 827 2783 893
rect 2876 887 2883 993
rect 2896 888 2903 1172
rect 2916 927 2923 1316
rect 2976 987 2983 1536
rect 2996 1447 3003 1493
rect 3016 1367 3023 1413
rect 3116 1407 3123 1453
rect 3107 1396 3123 1407
rect 3107 1393 3120 1396
rect 2953 927 2967 933
rect 2996 927 3003 1053
rect 3016 1047 3023 1253
rect 3036 1167 3043 1193
rect 3136 1167 3143 1193
rect 3156 1107 3163 1653
rect 3196 1443 3203 1873
rect 3296 1763 3303 1933
rect 3316 1847 3323 1973
rect 3316 1783 3323 1833
rect 3316 1776 3333 1783
rect 3276 1756 3303 1763
rect 3276 1707 3283 1756
rect 3336 1748 3343 1773
rect 3376 1747 3383 1973
rect 3493 1967 3507 1973
rect 3547 1963 3560 1967
rect 3547 1953 3563 1963
rect 3587 1953 3593 1967
rect 3556 1943 3563 1953
rect 3616 1947 3623 2073
rect 3656 1947 3663 2173
rect 3676 2067 3683 2413
rect 3756 2287 3763 2793
rect 3816 2767 3823 2953
rect 3813 2747 3827 2753
rect 3836 2667 3843 2993
rect 3856 2927 3863 2953
rect 3853 2787 3867 2793
rect 3916 2787 3923 2953
rect 3976 2947 3983 2973
rect 4096 2827 4103 2973
rect 3913 2767 3927 2773
rect 3867 2733 3873 2747
rect 3796 2247 3803 2513
rect 3816 2327 3823 2473
rect 3867 2433 3873 2447
rect 3833 2427 3847 2433
rect 3936 2427 3943 2793
rect 4096 2767 4103 2813
rect 4087 2756 4103 2767
rect 4153 2767 4167 2773
rect 4087 2753 4100 2756
rect 4056 2647 4063 2733
rect 4076 2527 4083 2753
rect 3956 2467 3963 2513
rect 3996 2387 4003 2473
rect 3873 2247 3887 2253
rect 3556 1936 3583 1943
rect 3453 1927 3467 1933
rect 3456 1887 3463 1913
rect 3516 1907 3523 1933
rect 3547 1913 3553 1927
rect 3473 1747 3487 1753
rect 3216 1447 3223 1673
rect 3247 1453 3253 1467
rect 3176 1436 3203 1443
rect 3016 907 3023 973
rect 2867 876 2883 887
rect 2867 873 2880 876
rect 3013 887 3027 893
rect 2927 873 2933 887
rect 2987 873 2993 887
rect 2900 866 2920 867
rect 2907 862 2920 866
rect 2907 853 2923 862
rect 2756 688 2763 713
rect 2753 647 2767 652
rect 2796 647 2803 733
rect 2836 667 2843 793
rect 2916 667 2923 853
rect 3036 807 3043 913
rect 2953 687 2967 693
rect 3076 687 3083 793
rect 2927 663 2940 667
rect 3033 663 3047 673
rect 2927 653 2943 663
rect 3033 660 3063 663
rect 3036 656 3063 660
rect 2756 407 2763 513
rect 2693 367 2707 373
rect 2813 367 2827 373
rect 2787 353 2793 367
rect 2736 327 2743 352
rect 2776 207 2783 353
rect 2836 343 2843 393
rect 2896 387 2903 453
rect 2936 407 2943 653
rect 3056 507 3063 656
rect 3096 587 3103 893
rect 3156 887 3163 1013
rect 3156 747 3163 873
rect 3176 727 3183 1436
rect 3253 1407 3267 1413
rect 3227 1393 3233 1407
rect 3276 947 3283 1553
rect 3296 1507 3303 1733
rect 3336 1467 3343 1712
rect 3307 1463 3320 1467
rect 3307 1453 3323 1463
rect 3316 1427 3323 1453
rect 3333 1447 3347 1453
rect 3396 1448 3403 1733
rect 3433 1727 3447 1733
rect 3556 1727 3563 1853
rect 3400 1426 3413 1427
rect 3296 1207 3303 1353
rect 3216 887 3223 913
rect 3236 843 3243 873
rect 3216 836 3243 843
rect 2936 393 2953 407
rect 2796 340 2843 343
rect 2793 336 2843 340
rect 2793 327 2807 336
rect 2936 307 2943 393
rect 2993 368 3007 373
rect 3076 367 3083 453
rect 3116 407 3123 673
rect 3187 653 3193 667
rect 3216 647 3223 836
rect 3256 707 3263 913
rect 3296 907 3303 1193
rect 3316 1067 3323 1413
rect 3407 1413 3413 1426
rect 3456 1387 3463 1693
rect 3576 1647 3583 1936
rect 3667 1936 3683 1943
rect 3596 1707 3603 1913
rect 3576 1527 3583 1633
rect 3676 1587 3683 1936
rect 3696 1927 3703 1993
rect 3756 1927 3763 2213
rect 3913 2207 3927 2213
rect 3896 2007 3903 2153
rect 3956 2027 3963 2273
rect 3996 2247 4003 2313
rect 3927 1973 3933 1987
rect 3813 1967 3827 1973
rect 3996 1967 4003 2053
rect 4036 1987 4043 2273
rect 3800 1963 3813 1967
rect 3796 1953 3813 1963
rect 3696 1787 3703 1913
rect 3776 1907 3783 1953
rect 3773 1767 3787 1773
rect 3707 1693 3713 1707
rect 3756 1687 3763 1713
rect 3716 1447 3723 1633
rect 3487 1433 3493 1447
rect 3356 1167 3363 1373
rect 3496 1227 3503 1253
rect 3516 1247 3523 1393
rect 3536 1327 3543 1433
rect 3576 1407 3583 1433
rect 3716 1407 3723 1433
rect 3767 1413 3773 1427
rect 3567 1396 3583 1407
rect 3567 1393 3580 1396
rect 3667 1393 3673 1407
rect 3696 1287 3703 1373
rect 3436 1167 3443 1213
rect 3453 1187 3467 1193
rect 3536 1187 3543 1273
rect 3553 1227 3567 1233
rect 3587 1213 3593 1227
rect 3487 1173 3493 1187
rect 3376 1027 3383 1153
rect 3413 927 3427 933
rect 3316 887 3323 913
rect 3387 893 3393 907
rect 3287 883 3300 887
rect 3287 880 3303 883
rect 3287 873 3307 880
rect 3293 867 3307 873
rect 3396 807 3403 893
rect 3436 747 3443 1153
rect 3516 967 3523 1093
rect 3676 1027 3683 1193
rect 3716 1187 3723 1253
rect 3796 1247 3803 1953
rect 4036 1947 4043 1973
rect 4076 1967 4083 2413
rect 4136 2248 4143 2473
rect 4156 2447 4163 2633
rect 4173 2487 4187 2493
rect 4196 2447 4203 2993
rect 4296 2983 4303 3276
rect 4433 3267 4447 3273
rect 4387 3253 4393 3267
rect 4456 3067 4463 3293
rect 4536 3287 4543 3413
rect 4636 3387 4643 3713
rect 4656 3508 4663 3753
rect 4696 3487 4703 4173
rect 4716 4067 4723 4113
rect 4716 3967 4723 4053
rect 4827 4033 4833 4047
rect 4773 4027 4787 4033
rect 4896 4007 4903 4033
rect 4736 3827 4743 3993
rect 4796 3967 4803 3993
rect 4893 3987 4907 3993
rect 4753 3847 4767 3853
rect 4916 3843 4923 4356
rect 4936 3887 4943 4353
rect 4956 4087 4963 4333
rect 5036 4327 5043 4473
rect 4976 4247 4983 4273
rect 4996 4047 5003 4273
rect 5036 4167 5043 4313
rect 5056 4307 5063 4496
rect 5116 4287 5123 4513
rect 5236 4367 5243 4513
rect 5173 4347 5187 4353
rect 5193 4327 5207 4333
rect 5227 4313 5233 4327
rect 5133 4287 5147 4293
rect 5167 4273 5173 4287
rect 5073 4267 5087 4273
rect 5016 4047 5023 4133
rect 4776 3836 4823 3843
rect 4916 3836 4943 3843
rect 4776 3823 4783 3836
rect 4756 3816 4783 3823
rect 4756 3807 4763 3816
rect 4713 3787 4727 3793
rect 4753 3787 4767 3793
rect 4796 3787 4803 3813
rect 4816 3807 4823 3836
rect 4816 3796 4833 3807
rect 4820 3793 4833 3796
rect 4916 3787 4923 3813
rect 4867 3773 4873 3787
rect 4836 3607 4843 3653
rect 4787 3524 4800 3527
rect 4787 3514 4803 3524
rect 4780 3513 4803 3514
rect 4656 3427 4663 3472
rect 4736 3467 4743 3513
rect 4773 3487 4787 3492
rect 4767 3480 4787 3487
rect 4767 3473 4783 3480
rect 4487 3256 4513 3263
rect 4553 3247 4567 3253
rect 4476 3027 4483 3232
rect 4576 3147 4583 3293
rect 4596 3107 4603 3233
rect 4616 3207 4623 3333
rect 4653 3287 4667 3293
rect 4696 3267 4703 3333
rect 4687 3257 4703 3267
rect 4687 3254 4700 3257
rect 4680 3253 4700 3254
rect 4716 3247 4723 3293
rect 4673 3227 4687 3232
rect 4536 3027 4543 3053
rect 4636 3047 4643 3133
rect 4573 3027 4587 3033
rect 4467 3020 4483 3027
rect 4467 3013 4487 3020
rect 4413 3008 4427 3013
rect 4473 3007 4487 3013
rect 4627 2993 4633 3007
rect 4296 2976 4323 2983
rect 4287 2953 4293 2967
rect 4236 2788 4243 2953
rect 4316 2847 4323 2976
rect 4336 2807 4343 2993
rect 4373 2947 4387 2953
rect 4416 2947 4423 2972
rect 4593 2967 4607 2973
rect 4647 2953 4653 2967
rect 4236 2467 4243 2752
rect 4256 2747 4263 2793
rect 4327 2783 4340 2787
rect 4327 2773 4343 2783
rect 4276 2747 4283 2773
rect 4336 2747 4343 2773
rect 4347 2736 4363 2743
rect 4296 2667 4303 2733
rect 4253 2487 4267 2493
rect 4267 2473 4273 2487
rect 4287 2473 4293 2487
rect 4233 2447 4247 2453
rect 4096 2207 4103 2233
rect 4196 2227 4203 2433
rect 4133 2207 4147 2212
rect 4216 2207 4223 2293
rect 4316 2247 4323 2553
rect 4356 2467 4363 2736
rect 4396 2607 4403 2833
rect 4413 2787 4427 2793
rect 4447 2773 4453 2787
rect 4436 2527 4443 2773
rect 4536 2767 4543 2813
rect 4476 2467 4483 2513
rect 4536 2508 4543 2753
rect 4567 2733 4573 2747
rect 4556 2487 4563 2653
rect 4596 2487 4603 2573
rect 4540 2486 4553 2487
rect 4433 2447 4447 2453
rect 4273 2227 4287 2233
rect 4247 2193 4253 2207
rect 4096 2167 4103 2193
rect 4316 2187 4323 2233
rect 4107 1953 4113 1967
rect 3833 1927 3847 1933
rect 3820 1923 3833 1927
rect 3816 1913 3833 1923
rect 3816 1687 3823 1913
rect 3876 1907 3883 1933
rect 4093 1907 4107 1913
rect 3836 1767 3843 1793
rect 3836 1707 3843 1753
rect 3856 1747 3863 1773
rect 3976 1747 3983 1813
rect 4016 1747 4023 1773
rect 4053 1747 4067 1753
rect 4136 1747 4143 1953
rect 4156 1947 4163 2013
rect 4256 1987 4263 2013
rect 4253 1967 4267 1973
rect 4200 1963 4213 1967
rect 4196 1953 4213 1963
rect 4156 1787 4163 1933
rect 4196 1903 4203 1953
rect 4227 1913 4233 1927
rect 4196 1896 4223 1903
rect 4176 1747 4183 1893
rect 3867 1693 3873 1707
rect 3816 1447 3823 1613
rect 3813 1427 3827 1433
rect 3836 1407 3843 1453
rect 3836 1327 3843 1393
rect 3936 1323 3943 1733
rect 4067 1693 4073 1707
rect 4033 1687 4047 1693
rect 3956 1387 3963 1413
rect 3936 1316 3963 1323
rect 3936 1227 3943 1293
rect 3636 947 3643 1013
rect 3276 667 3283 733
rect 3307 703 3320 707
rect 3307 693 3323 703
rect 3316 681 3323 693
rect 3236 607 3243 653
rect 3196 407 3203 553
rect 3107 393 3123 407
rect 3247 393 3253 407
rect 3116 367 3123 393
rect 3167 353 3173 367
rect 3073 347 3087 353
rect 2987 346 3000 347
rect 2987 333 2993 346
rect 2816 187 2823 293
rect 3013 187 3027 193
rect 3116 187 3123 353
rect 3216 267 3223 353
rect 3256 243 3263 353
rect 3296 347 3303 633
rect 3316 427 3323 653
rect 3356 627 3363 653
rect 3376 607 3383 673
rect 3416 647 3423 713
rect 3516 707 3523 913
rect 3533 867 3547 873
rect 3453 687 3467 693
rect 3536 687 3543 793
rect 3336 467 3343 593
rect 3336 407 3343 453
rect 3396 407 3403 593
rect 3536 507 3543 673
rect 3556 667 3563 913
rect 3716 907 3723 1013
rect 3727 893 3733 907
rect 3596 847 3603 893
rect 3640 883 3653 887
rect 3636 873 3653 883
rect 3636 807 3643 873
rect 3576 527 3583 653
rect 3676 647 3683 793
rect 3676 607 3683 633
rect 3716 627 3723 733
rect 3736 687 3743 713
rect 3756 687 3763 1073
rect 3816 1023 3823 1213
rect 3860 1183 3873 1187
rect 3856 1173 3873 1183
rect 3927 1173 3933 1187
rect 3856 1087 3863 1173
rect 3776 1016 3823 1023
rect 3776 927 3783 1016
rect 3773 707 3787 713
rect 3767 633 3773 647
rect 3387 396 3403 407
rect 3473 407 3487 413
rect 3387 393 3400 396
rect 3393 368 3407 373
rect 3476 367 3483 393
rect 3496 367 3503 493
rect 3593 407 3607 413
rect 3636 387 3643 493
rect 3796 427 3803 673
rect 3816 407 3823 693
rect 3856 667 3863 933
rect 3876 807 3883 1113
rect 3956 943 3963 1316
rect 3976 1247 3983 1313
rect 3976 1103 3983 1233
rect 3996 1127 4003 1513
rect 4016 1347 4023 1573
rect 4036 1267 4043 1553
rect 4016 1187 4023 1213
rect 4036 1187 4043 1213
rect 3976 1096 4003 1103
rect 3956 941 3983 943
rect 3956 936 3973 941
rect 3933 927 3947 933
rect 3967 873 3973 887
rect 3896 747 3903 873
rect 3913 707 3927 713
rect 3976 707 3983 793
rect 3887 693 3893 707
rect 3853 647 3867 653
rect 3896 627 3903 653
rect 3976 547 3983 693
rect 3996 687 4003 1096
rect 4016 727 4023 893
rect 4056 747 4063 1573
rect 4116 1507 4123 1693
rect 4076 1207 4083 1493
rect 4107 1413 4113 1427
rect 4116 1227 4123 1373
rect 4136 1203 4143 1673
rect 4216 1627 4223 1896
rect 4236 1867 4243 1913
rect 4236 1647 4243 1853
rect 4276 1747 4283 1793
rect 4256 1707 4263 1733
rect 4216 1527 4223 1613
rect 4256 1487 4263 1693
rect 4293 1687 4307 1693
rect 4296 1567 4303 1673
rect 4316 1587 4323 1973
rect 4336 1963 4343 1993
rect 4356 1987 4363 2293
rect 4376 2047 4383 2413
rect 4496 2267 4503 2473
rect 4547 2473 4553 2486
rect 4616 2447 4623 2613
rect 4676 2587 4683 2773
rect 4696 2767 4703 3213
rect 4736 3027 4743 3373
rect 4756 3307 4763 3393
rect 4776 3283 4783 3473
rect 4796 3467 4803 3513
rect 4836 3507 4843 3593
rect 4916 3527 4923 3633
rect 4936 3567 4943 3836
rect 4956 3607 4963 4033
rect 5033 4007 5047 4013
rect 4996 3947 5003 3993
rect 5016 3827 5023 3873
rect 4976 3527 4983 3673
rect 4996 3647 5003 3773
rect 5016 3627 5023 3813
rect 5056 3587 5063 4073
rect 5076 4047 5083 4133
rect 5096 3827 5103 4253
rect 5116 4007 5123 4113
rect 5153 4007 5167 4013
rect 5087 3816 5103 3827
rect 5087 3813 5100 3816
rect 5116 3687 5123 3833
rect 5176 3787 5183 3853
rect 5216 3843 5223 4313
rect 5256 4167 5263 4313
rect 5296 4307 5303 4533
rect 5313 4327 5327 4333
rect 5287 4296 5303 4307
rect 5287 4293 5300 4296
rect 5376 4287 5383 4393
rect 5436 4307 5443 4553
rect 5456 4527 5463 4796
rect 5487 4773 5493 4787
rect 5516 4647 5523 4833
rect 5476 4567 5483 4633
rect 5493 4527 5507 4533
rect 5487 4313 5493 4327
rect 5453 4287 5467 4293
rect 5336 4247 5343 4273
rect 5373 4267 5387 4273
rect 5427 4253 5433 4267
rect 5233 4027 5247 4033
rect 5256 3987 5263 4073
rect 5276 4048 5283 4113
rect 5316 4067 5323 4173
rect 5313 4047 5327 4053
rect 5280 4026 5293 4027
rect 5287 4013 5293 4026
rect 5216 3836 5243 3843
rect 5213 3807 5227 3813
rect 4916 3516 4933 3527
rect 4920 3513 4933 3516
rect 4876 3487 4883 3513
rect 4927 3473 4933 3487
rect 4796 3307 4803 3413
rect 4856 3307 4863 3473
rect 4953 3467 4967 3473
rect 4996 3327 5003 3553
rect 5016 3487 5023 3573
rect 5096 3527 5103 3613
rect 5053 3507 5067 3513
rect 5047 3476 5083 3483
rect 5056 3427 5063 3453
rect 5076 3447 5083 3476
rect 5096 3407 5103 3513
rect 5136 3507 5143 3773
rect 5236 3727 5243 3836
rect 5173 3547 5187 3553
rect 5227 3533 5233 3547
rect 5116 3347 5123 3473
rect 5136 3427 5143 3453
rect 4756 3276 4783 3283
rect 4756 3127 4763 3276
rect 4776 3227 4783 3253
rect 4796 3247 4803 3293
rect 4827 3253 4833 3267
rect 4867 3253 4873 3267
rect 4736 2787 4743 2973
rect 4776 2967 4783 3053
rect 4796 3027 4803 3073
rect 4796 2787 4803 3013
rect 4876 3007 4883 3033
rect 4833 2987 4847 2993
rect 4787 2733 4793 2747
rect 4407 2253 4413 2267
rect 4487 2253 4493 2267
rect 4453 2247 4467 2253
rect 4427 2213 4433 2227
rect 4476 2087 4483 2213
rect 4516 2007 4523 2393
rect 4536 2347 4543 2433
rect 4576 2387 4583 2433
rect 4636 2247 4643 2493
rect 4716 2487 4723 2713
rect 4736 2667 4743 2733
rect 4813 2727 4827 2733
rect 4753 2487 4767 2493
rect 4813 2487 4827 2493
rect 4836 2487 4843 2853
rect 4876 2747 4883 2933
rect 4896 2863 4903 3313
rect 4916 3023 4923 3293
rect 4933 3287 4947 3293
rect 4976 3207 4983 3273
rect 4993 3263 5007 3273
rect 5016 3263 5023 3293
rect 5036 3267 5043 3333
rect 5156 3307 5163 3493
rect 5127 3293 5133 3307
rect 5176 3267 5183 3533
rect 4993 3256 5023 3263
rect 4993 3247 5007 3256
rect 5127 3253 5133 3267
rect 5033 3247 5047 3253
rect 5176 3227 5183 3253
rect 5196 3127 5203 3493
rect 5256 3387 5263 3933
rect 5276 3808 5283 3833
rect 5313 3807 5327 3813
rect 5280 3786 5300 3787
rect 5287 3773 5293 3786
rect 5336 3547 5343 3913
rect 5356 3827 5363 4053
rect 5416 4027 5423 4153
rect 5433 4047 5447 4053
rect 5456 3967 5463 4073
rect 5496 3927 5503 4273
rect 5356 3567 5363 3813
rect 5396 3787 5403 3853
rect 5433 3787 5447 3793
rect 5367 3553 5373 3567
rect 5276 3447 5283 3533
rect 5336 3527 5343 3533
rect 5336 3516 5353 3527
rect 5340 3513 5353 3516
rect 5456 3507 5463 3833
rect 5496 3567 5503 3813
rect 5327 3493 5333 3507
rect 5216 3248 5223 3293
rect 4916 3016 4943 3023
rect 4913 2987 4927 2993
rect 4896 2856 4923 2863
rect 4896 2787 4903 2833
rect 4827 2476 4843 2487
rect 4827 2473 4840 2476
rect 4696 2347 4703 2433
rect 4716 2427 4723 2473
rect 4747 2434 4753 2447
rect 4833 2447 4847 2453
rect 4747 2433 4760 2434
rect 4713 2247 4727 2253
rect 4593 2227 4607 2233
rect 4336 1956 4373 1963
rect 4336 1607 4343 1956
rect 4353 1927 4367 1933
rect 4416 1927 4423 1953
rect 4366 1920 4367 1927
rect 4487 1913 4493 1927
rect 4353 1707 4367 1713
rect 4156 1387 4163 1473
rect 4376 1447 4383 1913
rect 4433 1907 4447 1913
rect 4393 1727 4407 1733
rect 4436 1687 4443 1753
rect 4456 1727 4463 1853
rect 4516 1827 4523 1953
rect 4547 1933 4553 1947
rect 4573 1887 4587 1893
rect 4496 1816 4513 1823
rect 4496 1707 4503 1816
rect 4553 1727 4567 1733
rect 4416 1447 4423 1593
rect 4516 1527 4523 1593
rect 4467 1433 4473 1447
rect 4216 1407 4223 1433
rect 4156 1227 4163 1293
rect 4136 1196 4163 1203
rect 4073 1187 4087 1193
rect 4127 1173 4133 1187
rect 4076 887 4083 973
rect 4107 913 4113 927
rect 4087 873 4093 887
rect 4136 807 4143 953
rect 4156 927 4163 1196
rect 4187 1173 4193 1187
rect 4107 703 4120 707
rect 4107 693 4123 703
rect 3993 667 4007 673
rect 4073 668 4087 673
rect 4047 653 4053 667
rect 3993 647 4007 653
rect 3787 353 3793 367
rect 3236 236 3263 243
rect 2967 173 2973 187
rect 3207 173 3213 187
rect 2733 167 2747 173
rect 2527 133 2533 147
rect 2476 87 2483 133
rect 2836 -24 2843 173
rect 2913 167 2927 173
rect 2956 107 2963 133
rect 2993 127 3007 133
rect 3076 -24 3083 173
rect 3153 167 3167 173
rect 3236 147 3243 236
rect 3256 187 3263 213
rect 3296 167 3303 253
rect 3196 47 3203 133
rect 3356 -17 3363 173
rect 3396 167 3403 332
rect 3496 303 3503 353
rect 3713 347 3727 353
rect 3496 296 3523 303
rect 3456 -17 3463 173
rect 3516 167 3523 296
rect 3536 147 3543 273
rect 3593 208 3607 213
rect 3556 -17 3563 173
rect 3647 153 3653 167
rect 3593 147 3607 153
rect 3676 127 3683 173
rect 3736 147 3743 213
rect 3816 187 3823 393
rect 3856 287 3863 533
rect 4076 487 4083 632
rect 3933 407 3947 413
rect 3967 373 3973 387
rect 4076 367 4083 473
rect 4116 427 4123 693
rect 4147 633 4153 647
rect 4176 467 4183 853
rect 4196 428 4203 1173
rect 4216 1067 4223 1273
rect 4236 1207 4243 1333
rect 4256 1027 4263 1413
rect 4447 1393 4453 1407
rect 4347 1383 4360 1387
rect 4347 1373 4363 1383
rect 4276 1187 4283 1213
rect 4296 987 4303 1253
rect 4356 1227 4363 1373
rect 4347 1216 4363 1227
rect 4347 1213 4360 1216
rect 4376 1187 4383 1393
rect 4536 1247 4543 1693
rect 4556 1687 4563 1713
rect 4596 1707 4603 1993
rect 4627 1933 4633 1947
rect 4656 1887 4663 2133
rect 4716 1967 4723 2073
rect 4676 1867 4683 1953
rect 4676 1827 4683 1853
rect 4713 1727 4727 1733
rect 4736 1728 4743 2353
rect 4756 2187 4763 2412
rect 4776 2127 4783 2253
rect 4796 2087 4803 2213
rect 4756 1947 4763 1973
rect 4776 1928 4783 2033
rect 4796 1927 4803 2073
rect 4856 2007 4863 2573
rect 4876 2447 4883 2593
rect 4876 2227 4883 2333
rect 4896 2267 4903 2453
rect 4916 2307 4923 2856
rect 4936 2587 4943 3016
rect 4996 3007 5003 3113
rect 5116 3007 5123 3113
rect 4993 2987 5007 2993
rect 5067 2993 5073 3007
rect 5033 2983 5047 2993
rect 5033 2980 5063 2983
rect 5036 2976 5067 2980
rect 4956 2627 4963 2933
rect 4996 2847 5003 2973
rect 5053 2967 5067 2976
rect 5156 2967 5163 2993
rect 5196 2967 5203 3073
rect 5216 3007 5223 3212
rect 5236 3167 5243 3313
rect 5316 3307 5323 3493
rect 5496 3487 5503 3513
rect 5316 3263 5323 3293
rect 5376 3287 5383 3413
rect 5436 3327 5443 3473
rect 5467 3293 5473 3307
rect 5296 3260 5323 3263
rect 5253 3247 5267 3253
rect 5293 3256 5323 3260
rect 5293 3247 5307 3256
rect 5407 3256 5433 3263
rect 5300 3043 5313 3047
rect 5296 3033 5313 3043
rect 5107 2953 5113 2967
rect 5196 2956 5213 2967
rect 5200 2953 5213 2956
rect 5136 2867 5143 2953
rect 4973 2787 4987 2793
rect 5273 2787 5287 2793
rect 5067 2783 5080 2787
rect 5067 2773 5083 2783
rect 5013 2767 5027 2773
rect 4987 2733 4993 2747
rect 5033 2727 5047 2733
rect 5076 2707 5083 2773
rect 5153 2747 5167 2753
rect 5036 2467 5043 2513
rect 4993 2447 5007 2453
rect 5036 2347 5043 2453
rect 5127 2443 5140 2447
rect 5127 2433 5143 2443
rect 5136 2407 5143 2433
rect 5156 2367 5163 2573
rect 5196 2527 5203 2753
rect 5216 2467 5223 2693
rect 5296 2667 5303 3033
rect 5327 2993 5333 3007
rect 5356 2987 5363 3233
rect 5407 3213 5413 3227
rect 4987 2263 5000 2267
rect 4987 2253 5003 2263
rect 4933 2247 4947 2253
rect 4907 2213 4913 2227
rect 4956 2187 4963 2213
rect 4833 1967 4847 1973
rect 4887 1963 4900 1967
rect 4887 1953 4903 1963
rect 4896 1927 4903 1953
rect 4796 1916 4813 1927
rect 4800 1913 4813 1916
rect 4776 1767 4783 1892
rect 4726 1720 4727 1727
rect 4556 1676 4573 1687
rect 4560 1673 4573 1676
rect 4627 1673 4633 1687
rect 4636 1647 4643 1673
rect 4656 1527 4663 1713
rect 4556 1427 4563 1453
rect 4596 1447 4603 1513
rect 4676 1507 4683 1653
rect 4696 1607 4703 1693
rect 4733 1687 4747 1692
rect 4756 1667 4763 1733
rect 4433 1227 4447 1233
rect 4593 1227 4607 1233
rect 4367 1176 4383 1187
rect 4367 1173 4380 1176
rect 4467 1173 4473 1187
rect 4356 947 4363 1173
rect 4496 1107 4503 1213
rect 4573 1187 4587 1193
rect 4527 1173 4533 1187
rect 4576 1087 4583 1173
rect 4616 1167 4623 1473
rect 4727 1433 4733 1447
rect 4653 1427 4667 1433
rect 4640 1423 4653 1427
rect 4636 1413 4653 1423
rect 4636 1387 4643 1413
rect 4696 1387 4703 1433
rect 4753 1387 4767 1393
rect 4636 1187 4643 1213
rect 4656 1208 4663 1373
rect 4696 1227 4703 1333
rect 4693 1207 4707 1213
rect 4736 1187 4743 1233
rect 4776 1223 4783 1713
rect 4796 1407 4803 1713
rect 4836 1687 4843 1793
rect 4856 1707 4863 1913
rect 4936 1767 4943 1993
rect 4956 1907 4963 2173
rect 4976 1967 4983 2013
rect 4996 1987 5003 2253
rect 5116 2247 5123 2333
rect 5236 2327 5243 2593
rect 5276 2487 5283 2533
rect 5316 2503 5323 2813
rect 5347 2773 5353 2787
rect 5336 2508 5343 2773
rect 5356 2707 5363 2733
rect 5376 2683 5383 3013
rect 5356 2676 5383 2683
rect 5356 2607 5363 2676
rect 5296 2496 5323 2503
rect 5193 2247 5207 2253
rect 5073 2227 5087 2233
rect 5056 1967 5063 2113
rect 5013 1947 5027 1953
rect 5056 1927 5063 1953
rect 5047 1916 5063 1927
rect 5047 1913 5060 1916
rect 4896 1687 4903 1713
rect 4887 1676 4903 1687
rect 4953 1687 4967 1693
rect 4887 1673 4900 1676
rect 4996 1647 5003 1673
rect 5016 1607 5023 1893
rect 4876 1487 4883 1593
rect 4873 1467 4887 1473
rect 5036 1467 5043 1753
rect 5056 1467 5063 1773
rect 5076 1767 5083 1853
rect 5096 1787 5103 2013
rect 5136 1947 5143 2233
rect 5173 1968 5187 1973
rect 5147 1933 5153 1947
rect 5236 1943 5243 2273
rect 5276 2247 5283 2413
rect 5296 2263 5303 2496
rect 5356 2487 5363 2533
rect 5340 2486 5363 2487
rect 5316 2307 5323 2473
rect 5347 2475 5363 2486
rect 5347 2473 5360 2475
rect 5376 2447 5383 2653
rect 5396 2627 5403 3173
rect 5416 2587 5423 3073
rect 5456 2907 5463 2953
rect 5496 2827 5503 3373
rect 5516 3187 5523 4313
rect 5536 3827 5543 4613
rect 5536 3707 5543 3773
rect 5536 3087 5543 3553
rect 5516 2967 5523 2993
rect 5416 2487 5423 2533
rect 5436 2507 5443 2693
rect 5456 2667 5463 2713
rect 5493 2707 5507 2713
rect 5516 2643 5523 2753
rect 5496 2636 5523 2643
rect 5496 2527 5503 2636
rect 5456 2487 5463 2513
rect 5433 2447 5447 2453
rect 5376 2436 5393 2447
rect 5380 2433 5393 2436
rect 5356 2407 5363 2433
rect 5296 2256 5323 2263
rect 5253 2227 5267 2233
rect 5276 2233 5293 2247
rect 5236 1936 5263 1943
rect 5173 1927 5187 1932
rect 5093 1727 5107 1733
rect 5136 1707 5143 1893
rect 4893 1427 4907 1433
rect 4756 1216 4783 1223
rect 4636 1186 4660 1187
rect 4636 1175 4653 1186
rect 4640 1173 4653 1175
rect 4267 933 4273 947
rect 4327 933 4333 947
rect 4236 708 4243 933
rect 4493 927 4507 933
rect 4220 704 4233 707
rect 4216 694 4233 704
rect 4216 693 4240 694
rect 4216 527 4223 693
rect 4233 667 4247 672
rect 4233 660 4253 667
rect 4236 656 4253 660
rect 4240 653 4253 656
rect 4276 567 4283 693
rect 4296 667 4303 893
rect 4367 873 4373 887
rect 4356 847 4363 873
rect 4433 803 4447 813
rect 4416 800 4447 803
rect 4416 796 4443 800
rect 4416 707 4423 796
rect 4456 787 4463 893
rect 4596 887 4603 933
rect 4636 923 4643 1033
rect 4656 947 4663 1152
rect 4756 967 4763 1216
rect 4816 1207 4823 1413
rect 4916 1407 4923 1453
rect 4916 1287 4923 1393
rect 4773 1187 4787 1193
rect 4667 943 4680 947
rect 4667 933 4683 943
rect 4636 916 4663 923
rect 4616 867 4623 913
rect 4433 723 4447 733
rect 4433 721 4463 723
rect 4433 720 4453 721
rect 4436 716 4453 720
rect 4536 707 4543 773
rect 4533 687 4547 693
rect 4356 587 4363 673
rect 4067 356 4083 367
rect 4067 353 4080 356
rect 4136 247 4143 353
rect 3787 173 3793 187
rect 3776 107 3783 133
rect 3796 127 3803 173
rect 3836 167 3843 213
rect 3933 167 3947 173
rect 3867 160 3923 163
rect 3867 156 3927 160
rect 3913 147 3927 156
rect 4013 167 4027 173
rect 4056 147 4063 233
rect 4156 167 4163 393
rect 4193 387 4207 392
rect 4213 347 4227 353
rect 3873 127 3887 133
rect 4176 127 4183 153
rect 3827 113 3833 127
rect 4227 113 4233 127
rect 4173 107 4187 113
rect 4256 27 4263 453
rect 4296 367 4303 393
rect 4336 387 4343 413
rect 4356 407 4363 573
rect 4536 467 4543 673
rect 4573 667 4587 673
rect 4413 387 4427 393
rect 4453 347 4467 353
rect 4316 87 4323 153
rect 4336 127 4343 333
rect 4496 187 4503 453
rect 4556 427 4563 473
rect 4593 427 4607 433
rect 4656 407 4663 916
rect 4676 827 4683 933
rect 4696 707 4703 953
rect 4747 913 4753 927
rect 4713 908 4727 913
rect 4713 867 4727 872
rect 4776 747 4783 1093
rect 4796 927 4803 953
rect 4836 927 4843 1193
rect 4856 967 4863 1233
rect 4893 1207 4907 1213
rect 4936 1203 4943 1453
rect 5073 1427 5087 1433
rect 5027 1413 5033 1427
rect 4953 1387 4967 1393
rect 5016 1227 5023 1253
rect 5036 1227 5043 1413
rect 5156 1347 5163 1713
rect 5060 1223 5073 1227
rect 5056 1213 5073 1223
rect 4916 1196 4943 1203
rect 4916 1127 4923 1196
rect 4916 927 4923 1073
rect 4956 967 4963 1173
rect 4860 923 4873 927
rect 4856 913 4873 923
rect 4827 873 4833 887
rect 4733 687 4747 693
rect 4773 688 4787 693
rect 4816 667 4823 693
rect 4767 666 4780 667
rect 4767 653 4773 666
rect 4713 647 4727 653
rect 4576 307 4583 373
rect 4413 167 4427 173
rect 4493 167 4507 173
rect 4376 127 4383 153
rect 4533 147 4547 153
rect 4616 47 4623 353
rect 4716 347 4723 633
rect 4836 527 4843 773
rect 4773 407 4787 413
rect 4813 407 4827 413
rect 4836 367 4843 473
rect 4856 447 4863 913
rect 4956 887 4963 953
rect 5036 927 5043 1173
rect 5056 1047 5063 1213
rect 5096 1187 5103 1313
rect 5176 1267 5183 1733
rect 5216 1707 5223 1793
rect 5236 1747 5243 1913
rect 5256 1763 5263 1936
rect 5276 1807 5283 2233
rect 5316 2087 5323 2256
rect 5336 2027 5343 2313
rect 5356 2227 5363 2393
rect 5376 2247 5383 2273
rect 5416 2247 5423 2293
rect 5476 2227 5483 2493
rect 5313 1967 5327 1973
rect 5296 1956 5313 1963
rect 5256 1756 5283 1763
rect 5236 1740 5253 1747
rect 5233 1733 5253 1740
rect 5233 1728 5247 1733
rect 5276 1707 5283 1756
rect 5216 1706 5240 1707
rect 5216 1695 5233 1706
rect 5220 1693 5233 1695
rect 5276 1468 5283 1693
rect 5227 1453 5233 1467
rect 5193 1448 5207 1453
rect 5200 1426 5213 1427
rect 5207 1413 5213 1426
rect 5093 1167 5107 1173
rect 4987 913 4993 927
rect 5116 908 5123 993
rect 5136 927 5143 1253
rect 5156 947 5163 1233
rect 5193 1207 5207 1213
rect 5207 1153 5213 1167
rect 5256 1163 5263 1393
rect 5276 1247 5283 1432
rect 5296 1327 5303 1956
rect 5336 1827 5343 1973
rect 5356 1847 5363 2073
rect 5396 2007 5403 2213
rect 5376 1948 5383 1993
rect 5393 1987 5407 1993
rect 5456 1967 5463 1993
rect 5427 1953 5433 1967
rect 5456 1956 5473 1967
rect 5460 1953 5473 1956
rect 5407 1913 5413 1927
rect 5376 1887 5383 1912
rect 5313 1747 5327 1753
rect 5316 1407 5323 1453
rect 5376 1447 5383 1873
rect 5396 1227 5403 1713
rect 5416 1408 5423 1833
rect 5456 1823 5463 1913
rect 5436 1816 5463 1823
rect 5436 1707 5443 1816
rect 5416 1247 5423 1372
rect 5393 1207 5407 1213
rect 5473 1207 5487 1213
rect 5353 1187 5367 1193
rect 5256 1156 5283 1163
rect 5176 927 5183 1073
rect 5256 1027 5263 1133
rect 5247 1003 5260 1007
rect 5247 993 5263 1003
rect 5256 963 5263 993
rect 5276 987 5283 1156
rect 5256 960 5303 963
rect 5256 956 5307 960
rect 5236 927 5243 953
rect 5293 947 5307 956
rect 5276 907 5283 933
rect 5193 887 5207 893
rect 4887 873 4893 887
rect 4947 876 4963 887
rect 4947 873 4960 876
rect 4913 707 4927 713
rect 4893 647 4907 653
rect 4936 567 4943 793
rect 4976 667 4983 733
rect 4996 727 5003 873
rect 5013 867 5027 873
rect 4993 707 5007 713
rect 5027 673 5033 687
rect 4876 427 4883 453
rect 4916 387 4923 413
rect 4867 373 4873 387
rect 4736 223 4743 353
rect 4716 216 4743 223
rect 4636 147 4643 173
rect 4716 147 4723 216
rect 4787 193 4793 207
rect 4733 187 4747 193
rect 4936 167 4943 293
rect 4956 247 4963 453
rect 4976 308 4983 513
rect 4996 367 5003 473
rect 5056 427 5063 873
rect 5273 887 5287 893
rect 5316 887 5323 973
rect 5116 787 5123 872
rect 5247 853 5253 867
rect 5176 707 5183 793
rect 5080 703 5093 707
rect 5076 693 5093 703
rect 5013 407 5027 413
rect 5033 367 5047 373
rect 5076 367 5083 693
rect 5173 687 5187 693
rect 5216 687 5223 713
rect 5336 707 5343 933
rect 5356 847 5363 873
rect 5336 693 5353 707
rect 5107 393 5113 407
rect 5187 393 5193 407
rect 4976 167 4983 272
rect 5013 167 5027 173
rect 4827 153 4833 167
rect 5093 167 5107 173
rect 5136 167 5143 333
rect 5156 307 5163 393
rect 5216 367 5223 433
rect 5267 393 5273 407
rect 5173 347 5187 353
rect 5256 287 5263 353
rect 4973 147 4987 153
rect 4676 87 4683 133
rect 4876 107 4883 133
rect 4916 87 4923 113
rect 5196 107 5203 193
rect 4967 93 4973 107
rect 5216 87 5223 233
rect 5256 187 5263 233
rect 5296 167 5303 673
rect 5316 127 5323 493
rect 5336 447 5343 693
rect 5376 688 5383 1113
rect 5396 807 5403 1193
rect 5416 1027 5423 1193
rect 5476 947 5483 1013
rect 5427 933 5433 947
rect 5393 707 5407 713
rect 5416 667 5423 893
rect 5376 487 5383 652
rect 5376 407 5383 473
rect 5336 187 5343 313
rect 5356 207 5363 353
rect 5396 247 5403 553
rect 5456 527 5463 873
rect 5436 387 5443 433
rect 5476 367 5483 393
rect 5416 127 5423 153
rect 5367 113 5373 127
rect 5496 47 5503 1233
rect 5516 167 5523 2613
rect 5536 327 5543 3033
rect 3336 -24 3363 -17
rect 3436 -24 3463 -17
rect 3536 -24 3563 -17
rect 4676 -24 4683 33
rect 5396 -24 5403 33
rect 5436 -24 5443 13
<< m3contact >>
rect 2213 5453 2227 5467
rect 393 5433 407 5447
rect 1073 5433 1087 5447
rect 93 5413 107 5427
rect 253 5413 267 5427
rect 113 5373 127 5387
rect 193 5373 207 5387
rect 93 5333 107 5347
rect 233 5333 247 5347
rect 293 5333 307 5347
rect 253 5293 267 5307
rect 173 5273 187 5287
rect 373 5333 387 5347
rect 413 5313 427 5327
rect 393 5293 407 5307
rect 333 5213 347 5227
rect 413 5213 427 5227
rect 293 5153 307 5167
rect 33 5133 47 5147
rect 93 5133 107 5147
rect 53 5093 67 5107
rect 393 5133 407 5147
rect 333 5093 347 5107
rect 107 5073 121 5087
rect 233 5073 247 5087
rect 113 5053 127 5067
rect 93 4853 107 4867
rect 113 4854 127 4868
rect 113 4832 127 4846
rect 213 5033 227 5047
rect 313 5033 327 5047
rect 193 4853 207 4867
rect 233 4853 247 4867
rect 173 4833 187 4847
rect 593 5353 607 5367
rect 513 5333 527 5347
rect 753 5373 767 5387
rect 773 5353 787 5367
rect 813 5353 827 5367
rect 673 5333 687 5347
rect 633 5313 647 5327
rect 653 5273 667 5287
rect 533 5253 547 5267
rect 493 5213 507 5227
rect 473 5133 487 5147
rect 613 5153 627 5167
rect 467 5073 481 5087
rect 493 5073 507 5087
rect 393 5033 407 5047
rect 413 5033 427 5047
rect 573 5053 587 5067
rect 533 5033 547 5047
rect 453 4993 467 5007
rect 333 4913 347 4927
rect 513 4913 527 4927
rect 293 4833 307 4847
rect 153 4773 167 4787
rect 353 4833 367 4847
rect 413 4813 427 4827
rect 453 4813 467 4827
rect 673 5173 687 5187
rect 733 5253 747 5267
rect 893 5353 907 5367
rect 873 5233 887 5247
rect 933 5333 947 5347
rect 1013 5333 1027 5347
rect 913 5213 927 5227
rect 793 5193 807 5207
rect 733 5133 747 5147
rect 713 5113 727 5127
rect 833 5133 847 5147
rect 773 5093 787 5107
rect 653 5052 667 5066
rect 673 5032 687 5046
rect 693 5013 707 5027
rect 753 5013 767 5027
rect 873 5113 887 5127
rect 913 5113 927 5127
rect 853 5033 867 5047
rect 713 4993 727 5007
rect 593 4833 607 4847
rect 653 4833 667 4847
rect 313 4733 327 4747
rect 173 4673 187 4687
rect 213 4613 227 4627
rect 413 4713 427 4727
rect 513 4653 527 4667
rect 473 4613 487 4627
rect 153 4573 167 4587
rect 253 4573 267 4587
rect 353 4573 367 4587
rect 193 4554 207 4568
rect 233 4553 247 4567
rect 73 4533 87 4547
rect 173 4533 187 4547
rect 193 4493 207 4507
rect 93 4353 107 4367
rect 133 4313 147 4327
rect 113 4053 127 4067
rect 53 3993 67 4007
rect 133 3993 147 4007
rect 213 4293 227 4307
rect 333 4513 347 4527
rect 433 4513 447 4527
rect 313 4493 327 4507
rect 773 4933 787 4947
rect 813 4913 827 4927
rect 893 5013 907 5027
rect 1053 5313 1067 5327
rect 993 5293 1007 5307
rect 2053 5393 2067 5407
rect 2133 5393 2147 5407
rect 1633 5373 1647 5387
rect 1733 5373 1747 5387
rect 2113 5374 2127 5388
rect 1113 5353 1127 5367
rect 1093 5313 1107 5327
rect 1073 5133 1087 5147
rect 953 5093 967 5107
rect 993 5094 1007 5108
rect 1033 5093 1047 5107
rect 933 4973 947 4987
rect 913 4913 927 4927
rect 893 4873 907 4887
rect 833 4833 847 4847
rect 733 4813 747 4827
rect 813 4813 827 4827
rect 753 4773 767 4787
rect 773 4753 787 4767
rect 693 4633 707 4647
rect 593 4593 607 4607
rect 713 4593 727 4607
rect 653 4553 667 4567
rect 673 4553 687 4567
rect 633 4513 647 4527
rect 313 4373 327 4387
rect 373 4373 387 4387
rect 433 4373 447 4387
rect 473 4374 487 4388
rect 353 4353 367 4367
rect 473 4352 487 4366
rect 353 4292 367 4306
rect 432 4293 446 4307
rect 454 4293 468 4307
rect 553 4293 567 4307
rect 193 4073 207 4087
rect 273 4073 287 4087
rect 313 4073 327 4087
rect 233 4053 247 4067
rect 173 4033 187 4047
rect 153 3973 167 3987
rect 213 3973 227 3987
rect 73 3833 87 3847
rect 233 3833 247 3847
rect 113 3813 127 3827
rect 173 3813 187 3827
rect 133 3773 147 3787
rect 153 3773 167 3787
rect 73 3653 87 3667
rect 13 3613 27 3627
rect 53 3553 67 3567
rect 93 3553 107 3567
rect 13 3513 27 3527
rect 233 3792 247 3806
rect 213 3753 227 3767
rect 193 3713 207 3727
rect 333 3853 347 3867
rect 333 3793 347 3807
rect 353 3753 367 3767
rect 313 3713 327 3727
rect 213 3554 227 3568
rect 213 3532 227 3546
rect 112 3493 126 3507
rect 134 3493 148 3507
rect 213 3492 227 3506
rect 53 3393 67 3407
rect 13 3253 27 3267
rect 73 3254 87 3268
rect 133 3253 147 3267
rect 53 3232 67 3246
rect 93 3233 107 3247
rect 13 3173 27 3187
rect 13 3113 27 3127
rect 13 3014 27 3028
rect 13 2992 27 3006
rect 13 2893 27 2907
rect 473 4173 487 4187
rect 433 4113 447 4127
rect 393 4033 407 4047
rect 373 3633 387 3647
rect 313 3593 327 3607
rect 373 3593 387 3607
rect 313 3553 327 3567
rect 332 3493 346 3507
rect 354 3493 368 3507
rect 293 3473 307 3487
rect 373 3453 387 3467
rect 293 3333 307 3347
rect 633 4253 647 4267
rect 613 4213 627 4227
rect 533 4093 547 4107
rect 513 4073 527 4087
rect 473 4033 487 4047
rect 413 3853 427 3867
rect 553 4073 567 4087
rect 673 4513 687 4527
rect 713 4473 727 4487
rect 693 4413 707 4427
rect 713 4293 727 4307
rect 693 4213 707 4227
rect 753 4273 767 4287
rect 713 4173 727 4187
rect 753 4113 767 4127
rect 733 4093 747 4107
rect 687 4073 701 4087
rect 653 4033 667 4047
rect 673 4033 687 4047
rect 793 4673 807 4687
rect 813 4573 827 4587
rect 893 4773 907 4787
rect 853 4753 867 4767
rect 893 4733 907 4747
rect 993 5053 1007 5067
rect 1073 5053 1087 5067
rect 993 4993 1007 5007
rect 947 4833 961 4847
rect 973 4834 987 4848
rect 913 4713 927 4727
rect 853 4573 867 4587
rect 893 4553 907 4567
rect 933 4673 947 4687
rect 953 4633 967 4647
rect 933 4593 947 4607
rect 913 4473 927 4487
rect 873 4413 887 4427
rect 853 4354 867 4368
rect 1033 5013 1047 5027
rect 1013 4973 1027 4987
rect 1013 4873 1027 4887
rect 993 4733 1007 4747
rect 1013 4493 1027 4507
rect 993 4413 1007 4427
rect 1013 4393 1027 4407
rect 973 4373 987 4387
rect 893 4333 907 4347
rect 853 4293 867 4307
rect 793 4273 807 4287
rect 893 4153 907 4167
rect 853 4073 867 4087
rect 773 4053 787 4067
rect 733 4013 747 4027
rect 753 4013 767 4027
rect 593 3993 607 4007
rect 613 3933 627 3947
rect 593 3873 607 3887
rect 693 3873 707 3887
rect 533 3834 547 3848
rect 573 3833 587 3847
rect 473 3753 487 3767
rect 433 3693 447 3707
rect 453 3673 467 3687
rect 473 3653 487 3667
rect 453 3633 467 3647
rect 413 3513 427 3527
rect 433 3494 447 3508
rect 153 3113 167 3127
rect 273 3093 287 3107
rect 73 3073 87 3087
rect 153 3073 167 3087
rect 53 2994 67 3008
rect 93 3013 107 3027
rect 53 2972 67 2986
rect 33 2773 47 2787
rect 33 2733 47 2747
rect 33 2673 47 2687
rect 253 3033 267 3047
rect 173 2973 187 2987
rect 233 2973 247 2987
rect 113 2933 127 2947
rect 213 2933 227 2947
rect 133 2893 147 2907
rect 193 2853 207 2867
rect 73 2773 87 2787
rect 213 2753 227 2767
rect 253 2753 267 2767
rect 133 2733 147 2747
rect 153 2733 167 2747
rect 313 3193 327 3207
rect 393 3193 407 3207
rect 373 3133 387 3147
rect 353 3033 367 3047
rect 293 2853 307 2867
rect 353 2973 367 2987
rect 433 3333 447 3347
rect 433 3133 447 3147
rect 1053 4973 1067 4987
rect 1113 5293 1127 5307
rect 1253 5353 1267 5367
rect 1293 5334 1307 5348
rect 1233 5193 1247 5207
rect 1173 5113 1187 5127
rect 1239 5113 1253 5127
rect 1233 5073 1247 5087
rect 1213 5033 1227 5047
rect 1133 5013 1147 5027
rect 1113 4913 1127 4927
rect 1073 4873 1087 4887
rect 1113 4873 1127 4887
rect 1073 4833 1087 4847
rect 1113 4833 1127 4847
rect 1433 5333 1447 5347
rect 1513 5333 1527 5347
rect 1639 5333 1653 5347
rect 1533 5313 1547 5327
rect 1633 5313 1647 5327
rect 1453 5293 1467 5307
rect 1493 5293 1507 5307
rect 1753 5333 1767 5347
rect 1673 5293 1687 5307
rect 1413 5233 1427 5247
rect 1533 5233 1547 5247
rect 1653 5233 1667 5247
rect 1393 5173 1407 5187
rect 1313 5053 1327 5067
rect 1333 5053 1347 5067
rect 1273 5033 1287 5047
rect 1253 4993 1267 5007
rect 1193 4973 1207 4987
rect 1173 4799 1187 4813
rect 1133 4773 1147 4787
rect 1153 4733 1167 4747
rect 1093 4713 1107 4727
rect 1073 4653 1087 4667
rect 1073 4532 1087 4546
rect 1053 4473 1067 4487
rect 1033 4333 1047 4347
rect 953 4313 967 4327
rect 973 4314 987 4328
rect 1012 4294 1026 4308
rect 1034 4294 1048 4308
rect 973 4272 987 4286
rect 913 4014 927 4028
rect 913 3973 927 3987
rect 913 3933 927 3947
rect 953 3873 967 3887
rect 853 3833 867 3847
rect 953 3833 967 3847
rect 653 3774 667 3788
rect 733 3773 747 3787
rect 553 3733 567 3747
rect 593 3533 607 3547
rect 673 3733 687 3747
rect 713 3733 727 3747
rect 653 3513 667 3527
rect 533 3492 547 3506
rect 733 3633 747 3647
rect 833 3773 847 3787
rect 1133 4533 1147 4547
rect 1293 4933 1307 4947
rect 1233 4893 1247 4907
rect 1213 4833 1227 4847
rect 1273 4833 1287 4847
rect 1193 4693 1207 4707
rect 1173 4673 1187 4687
rect 1153 4473 1167 4487
rect 1093 4433 1107 4447
rect 1133 4413 1147 4427
rect 1093 4393 1107 4407
rect 1093 4293 1107 4307
rect 1193 4593 1207 4607
rect 1533 5173 1547 5187
rect 1673 5173 1687 5187
rect 1453 5093 1467 5107
rect 1553 5133 1567 5147
rect 1533 5052 1547 5066
rect 1473 4953 1487 4967
rect 1513 4933 1527 4947
rect 1313 4893 1327 4907
rect 1373 4894 1387 4908
rect 1453 4893 1467 4907
rect 1493 4893 1507 4907
rect 1373 4872 1387 4886
rect 1333 4853 1347 4867
rect 1233 4813 1247 4827
rect 1313 4813 1327 4827
rect 1333 4773 1347 4787
rect 1233 4633 1247 4647
rect 1313 4613 1327 4627
rect 1273 4593 1287 4607
rect 1353 4593 1367 4607
rect 1213 4533 1227 4547
rect 1293 4533 1307 4547
rect 1173 4393 1187 4407
rect 1153 4373 1167 4387
rect 1293 4373 1307 4387
rect 1013 4272 1027 4286
rect 1213 4273 1227 4287
rect 1033 4173 1047 4187
rect 1073 4133 1087 4147
rect 1053 4093 1067 4107
rect 1173 4173 1187 4187
rect 1193 4133 1207 4147
rect 1113 4033 1127 4047
rect 1133 4033 1147 4047
rect 1173 4013 1187 4027
rect 1013 3913 1027 3927
rect 1073 3973 1087 3987
rect 1133 3953 1147 3967
rect 1113 3933 1127 3947
rect 1073 3913 1087 3927
rect 1113 3833 1127 3847
rect 973 3773 987 3787
rect 913 3733 927 3747
rect 933 3633 947 3647
rect 893 3573 907 3587
rect 773 3534 787 3548
rect 553 3473 567 3487
rect 473 3453 487 3467
rect 513 3433 527 3447
rect 593 3393 607 3407
rect 553 3293 567 3307
rect 553 3233 567 3247
rect 513 3173 527 3187
rect 493 3133 507 3147
rect 432 3093 446 3107
rect 454 3093 468 3107
rect 713 3493 727 3507
rect 813 3493 827 3507
rect 713 3433 727 3447
rect 753 3393 767 3407
rect 653 3333 667 3347
rect 693 3333 707 3347
rect 733 3293 747 3307
rect 793 3293 807 3307
rect 593 3153 607 3167
rect 513 3113 527 3127
rect 553 3093 567 3107
rect 493 2993 507 3007
rect 533 2993 547 3007
rect 433 2973 447 2987
rect 453 2953 467 2967
rect 493 2953 507 2967
rect 433 2933 447 2947
rect 473 2933 487 2947
rect 453 2913 467 2927
rect 413 2794 427 2808
rect 313 2773 327 2787
rect 213 2693 227 2707
rect 233 2533 247 2547
rect 93 2493 107 2507
rect 153 2473 167 2487
rect 133 2433 147 2447
rect 53 2273 67 2287
rect 313 2693 327 2707
rect 613 3073 627 3087
rect 693 3233 707 3247
rect 673 3213 687 3227
rect 733 3213 747 3227
rect 673 3093 687 3107
rect 633 3013 647 3027
rect 593 2993 607 3007
rect 553 2933 567 2947
rect 493 2893 507 2907
rect 633 2853 647 2867
rect 513 2793 527 2807
rect 753 3013 767 3027
rect 699 2993 713 3007
rect 873 3393 887 3407
rect 853 3333 867 3347
rect 793 3233 807 3247
rect 873 3274 887 3288
rect 873 3213 887 3227
rect 1213 4053 1227 4067
rect 1393 4853 1407 4867
rect 1453 4853 1467 4867
rect 1393 4812 1407 4826
rect 1433 4813 1447 4827
rect 1479 4813 1493 4827
rect 1393 4753 1407 4767
rect 1493 4713 1507 4727
rect 1413 4633 1427 4647
rect 1393 4473 1407 4487
rect 1373 4373 1387 4387
rect 1353 4354 1367 4368
rect 1273 4293 1287 4307
rect 1253 4093 1267 4107
rect 1233 4014 1247 4028
rect 1373 4253 1387 4267
rect 1353 4173 1367 4187
rect 1353 4133 1367 4147
rect 1333 4113 1347 4127
rect 1293 4073 1307 4087
rect 1273 4013 1287 4027
rect 1233 3953 1247 3967
rect 1253 3933 1267 3947
rect 1353 4073 1367 4087
rect 1313 3953 1327 3967
rect 1193 3893 1207 3907
rect 1293 3893 1307 3907
rect 1173 3794 1187 3808
rect 1133 3733 1147 3747
rect 1113 3633 1127 3647
rect 1113 3593 1127 3607
rect 953 3553 967 3567
rect 973 3373 987 3387
rect 953 3333 967 3347
rect 1013 3513 1027 3527
rect 993 3353 1007 3367
rect 933 3274 947 3288
rect 1033 3273 1047 3287
rect 933 3233 947 3247
rect 893 3193 907 3207
rect 813 3073 827 3087
rect 1013 3073 1027 3087
rect 853 3013 867 3027
rect 893 2973 907 2987
rect 813 2953 827 2967
rect 773 2939 787 2953
rect 873 2893 887 2907
rect 793 2813 807 2827
rect 713 2773 727 2787
rect 473 2693 487 2707
rect 1173 3653 1187 3667
rect 1233 3873 1247 3887
rect 1213 3793 1227 3807
rect 1193 3593 1207 3607
rect 1133 3573 1147 3587
rect 1373 4013 1387 4027
rect 1333 3873 1347 3887
rect 1333 3833 1347 3847
rect 1373 3973 1387 3987
rect 1473 4593 1487 4607
rect 1433 4553 1447 4567
rect 1713 5093 1727 5107
rect 1593 5073 1607 5087
rect 1593 4953 1607 4967
rect 1633 5073 1647 5087
rect 1673 5053 1687 5067
rect 1813 5333 1827 5347
rect 2113 5352 2127 5366
rect 1913 5333 1927 5347
rect 1873 5313 1887 5327
rect 1833 5093 1847 5107
rect 2033 5313 2047 5327
rect 2013 5273 2027 5287
rect 1853 5073 1867 5087
rect 1913 5073 1927 5087
rect 1793 5033 1807 5047
rect 1813 5033 1827 5047
rect 1833 5033 1847 5047
rect 1693 4994 1707 5008
rect 1633 4973 1647 4987
rect 1693 4972 1707 4986
rect 1633 4933 1647 4947
rect 1573 4893 1587 4907
rect 1613 4893 1627 4907
rect 1593 4853 1607 4867
rect 1673 4813 1687 4827
rect 1693 4713 1707 4727
rect 1553 4633 1567 4647
rect 2073 5253 2087 5267
rect 2113 5153 2127 5167
rect 2213 5373 2227 5387
rect 2353 5374 2367 5388
rect 2433 5373 2447 5387
rect 2153 5354 2167 5368
rect 2153 5273 2167 5287
rect 2193 5253 2207 5267
rect 2173 5233 2187 5247
rect 2353 5352 2367 5366
rect 2313 5313 2327 5327
rect 2333 5273 2347 5287
rect 2273 5213 2287 5227
rect 2173 5133 2187 5147
rect 2113 5093 2127 5107
rect 1873 4993 1887 5007
rect 1953 4993 1967 5007
rect 2073 5073 2087 5087
rect 2113 5052 2127 5066
rect 1993 4933 2007 4947
rect 2033 4933 2047 4947
rect 1973 4893 1987 4907
rect 1953 4853 1967 4867
rect 1773 4833 1787 4847
rect 1813 4833 1827 4847
rect 1733 4813 1747 4827
rect 1713 4613 1727 4627
rect 1533 4594 1547 4608
rect 1593 4593 1607 4607
rect 1493 4533 1507 4547
rect 1413 4374 1427 4388
rect 1413 4352 1427 4366
rect 1613 4573 1627 4587
rect 1653 4573 1667 4587
rect 1553 4533 1567 4547
rect 1773 4593 1787 4607
rect 1853 4813 1867 4827
rect 1813 4753 1827 4767
rect 1813 4693 1827 4707
rect 1833 4653 1847 4667
rect 1813 4633 1827 4647
rect 1853 4593 1867 4607
rect 1893 4813 1907 4827
rect 2053 4893 2067 4907
rect 2033 4853 2047 4867
rect 1913 4773 1927 4787
rect 1833 4553 1847 4567
rect 1873 4553 1887 4567
rect 1893 4553 1907 4567
rect 1613 4513 1627 4527
rect 1713 4513 1727 4527
rect 1853 4513 1867 4527
rect 1533 4453 1547 4467
rect 1453 4413 1467 4427
rect 1533 4373 1547 4387
rect 1513 4273 1527 4287
rect 1553 4213 1567 4227
rect 1733 4493 1747 4507
rect 1713 4393 1727 4407
rect 1693 4293 1707 4307
rect 1553 4173 1567 4187
rect 1593 4173 1607 4187
rect 1413 4093 1427 4107
rect 1453 4094 1467 4108
rect 1493 4093 1507 4107
rect 1393 3873 1407 3887
rect 1373 3853 1387 3867
rect 1233 3733 1247 3747
rect 1273 3713 1287 3727
rect 1333 3733 1347 3747
rect 1233 3693 1247 3707
rect 1313 3693 1327 3707
rect 1213 3553 1227 3567
rect 1193 3513 1207 3527
rect 1093 3453 1107 3467
rect 1093 3373 1107 3387
rect 1272 3653 1286 3667
rect 1294 3653 1308 3667
rect 1253 3593 1267 3607
rect 1233 3333 1247 3347
rect 1073 3273 1087 3287
rect 1133 3273 1147 3287
rect 1173 3273 1187 3287
rect 1233 3253 1247 3267
rect 1073 3093 1087 3107
rect 1053 3013 1067 3027
rect 1113 3073 1127 3087
rect 1193 3193 1207 3207
rect 1133 3013 1147 3027
rect 1053 2973 1067 2987
rect 993 2933 1007 2947
rect 813 2793 827 2807
rect 933 2794 947 2808
rect 833 2753 847 2767
rect 933 2753 947 2767
rect 873 2733 887 2747
rect 713 2713 727 2727
rect 573 2693 587 2707
rect 493 2613 507 2627
rect 553 2613 567 2627
rect 433 2593 447 2607
rect 273 2534 287 2548
rect 273 2493 287 2507
rect 253 2459 267 2473
rect 276 2453 290 2467
rect 353 2453 367 2467
rect 233 2433 247 2447
rect 373 2433 387 2447
rect 253 2373 267 2387
rect 473 2513 487 2527
rect 413 2453 427 2467
rect 533 2593 547 2607
rect 513 2453 527 2467
rect 493 2393 507 2407
rect 333 2353 347 2367
rect 393 2353 407 2367
rect 53 2213 67 2227
rect 313 2273 327 2287
rect 293 2253 307 2267
rect 273 2233 287 2247
rect 393 2273 407 2287
rect 413 2253 427 2267
rect 593 2573 607 2587
rect 553 2533 567 2547
rect 833 2693 847 2707
rect 933 2613 947 2627
rect 813 2593 827 2607
rect 693 2573 707 2587
rect 653 2513 667 2527
rect 633 2473 647 2487
rect 733 2533 747 2547
rect 753 2514 767 2528
rect 793 2513 807 2527
rect 713 2493 727 2507
rect 753 2492 767 2506
rect 593 2433 607 2447
rect 633 2433 647 2447
rect 553 2393 567 2407
rect 653 2353 667 2367
rect 573 2233 587 2247
rect 613 2233 627 2247
rect 433 2213 447 2227
rect 173 2193 187 2207
rect 273 2193 287 2207
rect 93 2153 107 2167
rect 253 2153 267 2167
rect 33 2053 47 2067
rect 93 2053 107 2067
rect 233 2053 247 2067
rect 33 1993 47 2007
rect 93 1993 107 2007
rect 113 1953 127 1967
rect 33 1893 47 1907
rect 93 1893 107 1907
rect 533 2213 547 2227
rect 333 2173 347 2187
rect 393 2173 407 2187
rect 493 2173 507 2187
rect 593 2133 607 2147
rect 313 2033 327 2047
rect 273 1994 287 2008
rect 353 1993 367 2007
rect 133 1873 147 1887
rect 93 1813 107 1827
rect 93 1773 107 1787
rect 33 1753 47 1767
rect 293 1953 307 1967
rect 353 1953 367 1967
rect 493 1953 507 1967
rect 153 1813 167 1827
rect 253 1813 267 1827
rect 33 1653 47 1667
rect 93 1653 107 1667
rect 233 1733 247 1747
rect 333 1913 347 1927
rect 353 1913 367 1927
rect 313 1773 327 1787
rect 272 1733 286 1747
rect 253 1694 267 1708
rect 233 1653 247 1667
rect 13 1433 27 1447
rect 73 1433 87 1447
rect 253 1453 267 1467
rect 293 1693 307 1707
rect 453 1873 467 1887
rect 373 1813 387 1827
rect 553 1833 567 1847
rect 453 1753 467 1767
rect 413 1733 427 1747
rect 373 1693 387 1707
rect 440 1693 453 1707
rect 453 1693 454 1707
rect 333 1653 347 1667
rect 533 1653 547 1667
rect 453 1473 467 1487
rect 493 1473 507 1487
rect 333 1453 347 1467
rect 13 1393 27 1407
rect 93 1393 107 1407
rect 173 1393 187 1407
rect 313 1393 327 1407
rect 233 1273 247 1287
rect 67 1173 81 1187
rect 53 1013 67 1027
rect 293 1213 307 1227
rect 293 1173 307 1187
rect 133 1033 147 1047
rect 193 1033 207 1047
rect 253 1013 267 1027
rect 113 893 127 907
rect 113 813 127 827
rect 93 753 107 767
rect 33 433 47 447
rect 93 433 107 447
rect 13 393 27 407
rect 113 393 127 407
rect 233 813 247 827
rect 373 1233 387 1247
rect 673 2333 687 2347
rect 693 2273 707 2287
rect 753 2273 767 2287
rect 673 2053 687 2067
rect 653 2033 667 2047
rect 753 2233 767 2247
rect 773 2233 787 2247
rect 893 2493 907 2507
rect 1133 2933 1147 2947
rect 1273 3494 1287 3508
rect 1313 3633 1327 3647
rect 1313 3574 1327 3588
rect 1313 3552 1327 3566
rect 1453 4072 1467 4086
rect 1513 4073 1527 4087
rect 1693 4153 1707 4167
rect 1633 4093 1647 4107
rect 1473 4034 1487 4048
rect 1473 3973 1487 3987
rect 1453 3953 1467 3967
rect 1473 3933 1487 3947
rect 1553 4033 1567 4047
rect 1553 3853 1567 3867
rect 1413 3793 1427 3807
rect 1473 3793 1487 3807
rect 1553 3793 1567 3807
rect 1453 3773 1467 3787
rect 1373 3653 1387 3667
rect 1373 3473 1387 3487
rect 1353 3453 1367 3467
rect 1373 3433 1387 3447
rect 1333 3393 1347 3407
rect 1393 3393 1407 3407
rect 1333 3353 1347 3367
rect 1313 3293 1327 3307
rect 1373 3313 1387 3327
rect 1333 3273 1347 3287
rect 1313 3253 1327 3267
rect 1333 3233 1347 3247
rect 1253 3173 1267 3187
rect 1273 3093 1287 3107
rect 1293 3053 1307 3067
rect 1493 3773 1507 3787
rect 1593 4053 1607 4067
rect 1573 3773 1587 3787
rect 1513 3733 1527 3747
rect 1573 3733 1587 3747
rect 1573 3693 1587 3707
rect 1473 3573 1487 3587
rect 1573 3573 1587 3587
rect 1533 3513 1547 3527
rect 1553 3513 1567 3527
rect 1513 3473 1527 3487
rect 1513 3433 1527 3447
rect 1493 3333 1507 3347
rect 1553 3433 1567 3447
rect 1793 4493 1807 4507
rect 1753 4453 1767 4467
rect 1873 4413 1887 4427
rect 1893 4393 1907 4407
rect 1993 4773 2007 4787
rect 2093 4653 2107 4667
rect 2033 4633 2047 4647
rect 1973 4613 1987 4627
rect 2013 4613 2027 4627
rect 1973 4513 1987 4527
rect 1953 4493 1967 4507
rect 1973 4373 1987 4387
rect 1933 4353 1947 4367
rect 1893 4333 1907 4347
rect 1853 4294 1867 4308
rect 1873 4293 1887 4307
rect 1793 4193 1807 4207
rect 1773 4153 1787 4167
rect 1733 4053 1747 4067
rect 1613 3953 1627 3967
rect 1633 3913 1647 3927
rect 1593 3513 1607 3527
rect 1713 4013 1727 4027
rect 1733 3993 1747 4007
rect 1913 4253 1927 4267
rect 1853 4113 1867 4127
rect 1893 4113 1907 4127
rect 1793 4032 1807 4046
rect 1773 3853 1787 3867
rect 1753 3833 1767 3847
rect 1653 3713 1667 3727
rect 1693 3673 1707 3687
rect 1753 3793 1767 3807
rect 1753 3752 1767 3766
rect 1733 3593 1747 3607
rect 1733 3533 1747 3547
rect 1573 3373 1587 3387
rect 1553 3353 1567 3367
rect 1533 3313 1547 3327
rect 1593 3293 1607 3307
rect 1553 3273 1567 3287
rect 1413 3233 1427 3247
rect 1372 3173 1386 3187
rect 1394 3173 1408 3187
rect 1353 3093 1367 3107
rect 1213 3013 1227 3027
rect 1193 2954 1207 2968
rect 1113 2893 1127 2907
rect 1173 2893 1187 2907
rect 1033 2813 1047 2827
rect 1013 2773 1027 2787
rect 993 2753 1007 2767
rect 1053 2793 1067 2807
rect 1193 2813 1207 2827
rect 973 2573 987 2587
rect 1073 2533 1087 2547
rect 853 2453 867 2467
rect 893 2453 907 2467
rect 953 2453 967 2467
rect 1153 2753 1167 2767
rect 1213 2753 1227 2767
rect 1253 2993 1267 3007
rect 1273 2933 1287 2947
rect 1453 3214 1467 3228
rect 1453 3192 1467 3206
rect 1513 3193 1527 3207
rect 1533 3173 1547 3187
rect 1453 3133 1467 3147
rect 1453 3093 1467 3107
rect 1433 3053 1447 3067
rect 1473 3073 1487 3087
rect 1453 3033 1467 3047
rect 1413 2953 1427 2967
rect 1333 2893 1347 2907
rect 1373 2913 1387 2927
rect 1413 2893 1427 2907
rect 1473 2973 1487 2987
rect 1733 3453 1747 3467
rect 1713 3433 1727 3447
rect 1733 3293 1747 3307
rect 1693 3273 1707 3287
rect 1633 3193 1647 3207
rect 1553 3073 1567 3087
rect 1593 3073 1607 3087
rect 1593 3033 1607 3047
rect 1566 2993 1567 3007
rect 1567 2993 1580 3007
rect 1573 2973 1587 2987
rect 1613 2893 1627 2907
rect 1393 2793 1407 2807
rect 1373 2754 1387 2768
rect 1413 2733 1427 2747
rect 1273 2613 1287 2627
rect 1333 2613 1347 2627
rect 1133 2513 1147 2527
rect 1193 2493 1207 2507
rect 1013 2333 1027 2347
rect 873 2253 887 2267
rect 973 2253 987 2267
rect 1053 2253 1067 2267
rect 813 1967 827 1981
rect 1013 2233 1027 2247
rect 913 2213 927 2227
rect 973 2193 987 2207
rect 1013 2193 1027 2207
rect 1053 2193 1067 2207
rect 893 2173 907 2187
rect 1093 2253 1107 2267
rect 1073 2133 1087 2147
rect 1353 2593 1367 2607
rect 1353 2553 1367 2567
rect 1173 2467 1187 2481
rect 1293 2453 1307 2467
rect 1453 2853 1467 2867
rect 1493 2813 1507 2827
rect 1553 2813 1567 2827
rect 1693 3233 1707 3247
rect 1713 3193 1727 3207
rect 1633 2794 1647 2808
rect 1653 2774 1667 2788
rect 1773 3673 1787 3687
rect 1773 3633 1787 3647
rect 1813 3993 1827 4007
rect 1813 3933 1827 3947
rect 1813 3853 1827 3867
rect 1853 4013 1867 4027
rect 1853 3913 1867 3927
rect 1953 4233 1967 4247
rect 2013 4353 2027 4367
rect 2053 4413 2067 4427
rect 2233 5093 2247 5107
rect 2233 5052 2247 5066
rect 2433 5332 2447 5346
rect 2493 5333 2507 5347
rect 2393 5313 2407 5327
rect 2453 5273 2467 5287
rect 2353 5113 2367 5127
rect 2413 5113 2427 5127
rect 2553 5453 2567 5467
rect 2593 5453 2607 5467
rect 2893 5453 2907 5467
rect 2573 5433 2587 5447
rect 2773 5433 2787 5447
rect 2533 5373 2547 5387
rect 2593 5353 2607 5367
rect 2533 5273 2547 5287
rect 2513 5173 2527 5187
rect 2493 5153 2507 5167
rect 2473 5093 2487 5107
rect 2393 5073 2407 5087
rect 2453 5073 2467 5087
rect 2293 5053 2307 5067
rect 2293 5013 2307 5027
rect 2333 5013 2347 5027
rect 2273 4973 2287 4987
rect 2253 4953 2267 4967
rect 2173 4893 2187 4907
rect 2493 5053 2507 5067
rect 2473 5012 2487 5026
rect 2433 4973 2447 4987
rect 2373 4953 2387 4967
rect 2333 4833 2347 4847
rect 2233 4813 2247 4827
rect 2213 4793 2227 4807
rect 2273 4793 2287 4807
rect 2153 4753 2167 4767
rect 2153 4553 2167 4567
rect 2233 4773 2247 4787
rect 2213 4553 2227 4567
rect 2133 4413 2147 4427
rect 2193 4413 2207 4427
rect 2113 4373 2127 4387
rect 2093 4313 2107 4327
rect 2133 4292 2147 4306
rect 2193 4293 2207 4307
rect 2313 4653 2327 4667
rect 2293 4593 2307 4607
rect 2233 4512 2247 4526
rect 2313 4553 2327 4567
rect 2353 4713 2367 4727
rect 2453 4893 2467 4907
rect 2393 4853 2407 4867
rect 2473 4833 2487 4847
rect 2473 4773 2487 4787
rect 2393 4713 2407 4727
rect 2373 4673 2387 4687
rect 2433 4593 2447 4607
rect 2613 5313 2627 5327
rect 2733 5353 2747 5367
rect 2853 5393 2867 5407
rect 2793 5373 2807 5387
rect 3093 5393 3107 5407
rect 2993 5353 3007 5367
rect 2713 5293 2727 5307
rect 2833 5293 2847 5307
rect 2893 5313 2907 5327
rect 3153 5453 3167 5467
rect 2993 5293 3007 5307
rect 2853 5273 2867 5287
rect 2973 5273 2987 5287
rect 3073 5273 3087 5287
rect 2653 5253 2667 5267
rect 2833 5253 2847 5267
rect 2633 5213 2647 5227
rect 2593 5173 2607 5187
rect 2613 5153 2627 5167
rect 2553 5093 2567 5107
rect 2533 4953 2547 4967
rect 2593 5074 2607 5088
rect 2573 5052 2587 5066
rect 2613 5053 2627 5067
rect 2593 5013 2607 5027
rect 2573 4893 2587 4907
rect 2653 5133 2667 5147
rect 2753 5113 2767 5127
rect 2813 5113 2827 5127
rect 2733 5073 2747 5087
rect 2753 5073 2767 5087
rect 2673 5053 2687 5067
rect 2793 5033 2807 5047
rect 2693 4973 2707 4987
rect 2773 4933 2787 4947
rect 2613 4853 2627 4867
rect 2553 4813 2567 4827
rect 2593 4812 2607 4826
rect 2713 4833 2727 4847
rect 2733 4813 2747 4827
rect 2673 4733 2687 4747
rect 2573 4713 2587 4727
rect 2553 4673 2567 4687
rect 2533 4633 2547 4647
rect 2373 4553 2387 4567
rect 2473 4553 2487 4567
rect 2593 4613 2607 4627
rect 2433 4533 2447 4547
rect 2333 4513 2347 4527
rect 2453 4493 2467 4507
rect 2253 4473 2267 4487
rect 2293 4473 2307 4487
rect 2413 4453 2427 4467
rect 2433 4413 2447 4427
rect 2413 4393 2427 4407
rect 2253 4353 2267 4367
rect 2073 4273 2087 4287
rect 2173 4273 2187 4287
rect 2013 4233 2027 4247
rect 1933 4054 1947 4068
rect 1973 4053 1987 4067
rect 1953 4033 1967 4047
rect 1933 4013 1947 4027
rect 1993 3973 2007 3987
rect 1973 3913 1987 3927
rect 1913 3893 1927 3907
rect 1993 3893 2007 3907
rect 1853 3873 1867 3887
rect 1933 3873 1947 3887
rect 1973 3853 1987 3867
rect 1953 3833 1967 3847
rect 1833 3793 1847 3807
rect 1853 3773 1867 3787
rect 1793 3553 1807 3567
rect 1773 3373 1787 3387
rect 1913 3793 1927 3807
rect 2053 4153 2067 4167
rect 2033 4013 2047 4027
rect 2013 3873 2027 3887
rect 1993 3813 2007 3827
rect 2033 3813 2047 3827
rect 1993 3733 2007 3747
rect 1953 3633 1967 3647
rect 1993 3593 2007 3607
rect 1973 3553 1987 3567
rect 1913 3473 1927 3487
rect 1813 3413 1827 3427
rect 1793 3353 1807 3367
rect 1973 3512 1987 3526
rect 1913 3373 1927 3387
rect 1893 3333 1907 3347
rect 1793 3293 1807 3307
rect 1833 3233 1847 3247
rect 1893 3233 1907 3247
rect 1813 3173 1827 3187
rect 1773 3014 1787 3028
rect 1773 2992 1787 3006
rect 1813 2993 1827 3007
rect 1733 2953 1747 2967
rect 1713 2933 1727 2947
rect 1753 2893 1767 2907
rect 1713 2854 1727 2868
rect 1873 3173 1887 3187
rect 1713 2832 1727 2846
rect 1773 2833 1787 2847
rect 1673 2773 1687 2787
rect 1452 2753 1466 2767
rect 1474 2753 1488 2767
rect 1613 2733 1627 2747
rect 1613 2613 1627 2627
rect 1653 2752 1667 2766
rect 1793 2813 1807 2827
rect 1733 2793 1747 2807
rect 1833 2793 1847 2807
rect 1773 2773 1787 2787
rect 1733 2713 1747 2727
rect 1633 2553 1647 2567
rect 1933 3013 1947 3027
rect 2093 4233 2107 4247
rect 2133 4233 2147 4247
rect 2132 4193 2146 4207
rect 2154 4193 2168 4207
rect 2093 4153 2107 4167
rect 2093 4113 2107 4127
rect 2073 4074 2087 4088
rect 2073 4052 2087 4066
rect 2173 4093 2187 4107
rect 2293 4334 2307 4348
rect 2473 4433 2487 4447
rect 2453 4373 2467 4387
rect 2353 4333 2367 4347
rect 2272 4312 2286 4326
rect 2294 4312 2308 4326
rect 2313 4233 2327 4247
rect 2293 4193 2307 4207
rect 2273 4153 2287 4167
rect 2273 4093 2287 4107
rect 2153 4053 2167 4067
rect 2093 3973 2107 3987
rect 2073 3893 2087 3907
rect 2073 3793 2087 3807
rect 2053 3713 2067 3727
rect 2073 3673 2087 3687
rect 2113 3793 2127 3807
rect 2093 3654 2107 3668
rect 2093 3632 2107 3646
rect 2053 3593 2067 3607
rect 2013 3574 2027 3588
rect 2013 3552 2027 3566
rect 1993 3293 2007 3307
rect 2033 3253 2047 3267
rect 2033 3213 2047 3227
rect 1993 3193 2007 3207
rect 2033 3133 2047 3147
rect 2193 4013 2207 4027
rect 2233 4033 2247 4047
rect 2213 3933 2227 3947
rect 2253 3913 2267 3927
rect 2233 3873 2247 3887
rect 2413 4293 2427 4307
rect 2373 4213 2387 4227
rect 2293 4013 2307 4027
rect 2333 3993 2347 4007
rect 2573 4554 2587 4568
rect 2813 5013 2827 5027
rect 2773 4713 2787 4727
rect 2793 4653 2807 4667
rect 2693 4613 2707 4627
rect 2773 4613 2787 4627
rect 2733 4593 2747 4607
rect 2593 4553 2607 4567
rect 2633 4553 2647 4567
rect 2553 4532 2567 4546
rect 3073 5233 3087 5247
rect 2993 5193 3007 5207
rect 2953 5093 2967 5107
rect 2893 5073 2907 5087
rect 2933 5053 2947 5067
rect 3053 5074 3067 5088
rect 2892 5013 2906 5027
rect 2914 5013 2928 5027
rect 3013 5013 3027 5027
rect 3053 5013 3067 5027
rect 2953 4953 2967 4967
rect 2913 4933 2927 4947
rect 3053 4973 3067 4987
rect 3033 4953 3047 4967
rect 3053 4933 3067 4947
rect 3013 4913 3027 4927
rect 2853 4853 2867 4867
rect 2893 4853 2907 4867
rect 2953 4853 2967 4867
rect 2913 4833 2927 4847
rect 2873 4813 2887 4827
rect 2847 4793 2861 4807
rect 2813 4573 2827 4587
rect 2873 4573 2887 4587
rect 2773 4553 2787 4567
rect 2613 4513 2627 4527
rect 2753 4513 2767 4527
rect 2613 4413 2627 4427
rect 2593 4333 2607 4347
rect 2633 4333 2647 4347
rect 2553 4313 2567 4327
rect 2693 4313 2707 4327
rect 2513 4293 2527 4307
rect 2673 4293 2687 4307
rect 2473 4213 2487 4227
rect 2433 4173 2447 4187
rect 2493 4173 2507 4187
rect 2413 4093 2427 4107
rect 2453 4093 2467 4107
rect 2393 3953 2407 3967
rect 2513 4033 2527 4047
rect 2593 4033 2607 4047
rect 2453 4013 2467 4027
rect 2493 4013 2507 4027
rect 2573 4013 2587 4027
rect 2533 3993 2547 4007
rect 2473 3953 2487 3967
rect 2473 3873 2487 3887
rect 2493 3853 2507 3867
rect 2313 3793 2327 3807
rect 2413 3833 2427 3847
rect 2453 3833 2467 3847
rect 2353 3774 2367 3788
rect 2293 3753 2307 3767
rect 2353 3733 2367 3747
rect 2312 3713 2326 3727
rect 2334 3713 2348 3727
rect 2133 3593 2147 3607
rect 2273 3593 2287 3607
rect 2313 3593 2327 3607
rect 2113 3553 2127 3567
rect 2153 3553 2167 3567
rect 2193 3533 2207 3547
rect 2093 3353 2107 3367
rect 2073 3293 2087 3307
rect 2153 3413 2167 3427
rect 2093 3193 2107 3207
rect 2013 3053 2027 3067
rect 2053 3053 2067 3067
rect 1973 3013 1987 3027
rect 1953 2993 1967 3007
rect 1913 2933 1927 2947
rect 2013 2973 2027 2987
rect 2053 2933 2067 2947
rect 2133 3253 2147 3267
rect 2193 3373 2207 3387
rect 2273 3473 2287 3487
rect 2353 3573 2367 3587
rect 2273 3233 2287 3247
rect 2353 3393 2367 3407
rect 2313 3313 2327 3327
rect 2213 3213 2227 3227
rect 2353 3133 2367 3147
rect 2193 3113 2207 3127
rect 2173 3073 2187 3087
rect 2173 3014 2187 3028
rect 2133 2993 2147 3007
rect 2153 2994 2167 3008
rect 2153 2972 2167 2986
rect 2213 3013 2227 3027
rect 2393 3793 2407 3807
rect 2453 3793 2467 3807
rect 2413 3753 2427 3767
rect 2473 3733 2487 3747
rect 2453 3713 2467 3727
rect 2413 3613 2427 3627
rect 2433 3533 2447 3547
rect 2493 3673 2507 3687
rect 2573 3933 2587 3947
rect 2553 3893 2567 3907
rect 2553 3773 2567 3787
rect 2613 4013 2627 4027
rect 2633 3973 2647 3987
rect 2733 4273 2747 4287
rect 2693 4233 2707 4247
rect 2652 3933 2666 3947
rect 2674 3933 2688 3947
rect 2673 3893 2687 3907
rect 2733 3973 2747 3987
rect 2773 4193 2787 4207
rect 2773 4153 2787 4167
rect 2833 4533 2847 4547
rect 2933 4813 2947 4827
rect 3193 5353 3207 5367
rect 3133 5333 3147 5347
rect 3153 5333 3167 5347
rect 4253 5473 4267 5487
rect 4313 5473 4327 5487
rect 3433 5453 3447 5467
rect 3473 5453 3487 5467
rect 3453 5433 3467 5447
rect 3233 5393 3247 5407
rect 3353 5393 3367 5407
rect 3413 5393 3427 5407
rect 3573 5413 3587 5427
rect 3673 5413 3687 5427
rect 3913 5413 3927 5427
rect 3613 5353 3627 5367
rect 3347 5333 3361 5347
rect 3413 5333 3427 5347
rect 3253 5273 3267 5287
rect 3213 5234 3227 5248
rect 3093 5213 3107 5227
rect 3213 5212 3227 5226
rect 3173 5153 3187 5167
rect 3093 5133 3107 5147
rect 3113 5093 3127 5107
rect 3093 5053 3107 5067
rect 3113 4933 3127 4947
rect 3033 4893 3047 4907
rect 3073 4893 3087 4907
rect 3113 4893 3127 4907
rect 3013 4813 3027 4827
rect 2993 4793 3007 4807
rect 3173 5013 3187 5027
rect 3173 4953 3187 4967
rect 3153 4893 3167 4907
rect 3133 4873 3147 4887
rect 3233 5173 3247 5187
rect 3273 5213 3287 5227
rect 3313 5233 3327 5247
rect 3293 5133 3307 5147
rect 3473 5273 3487 5287
rect 3553 5273 3567 5287
rect 3773 5333 3787 5347
rect 3613 5313 3627 5327
rect 3593 5293 3607 5307
rect 3673 5293 3687 5307
rect 3573 5233 3587 5247
rect 3593 5213 3607 5227
rect 3553 5173 3567 5187
rect 3393 5113 3407 5127
rect 3513 5113 3527 5127
rect 3853 5353 3867 5367
rect 3813 5333 3827 5347
rect 3793 5253 3807 5267
rect 3773 5213 3787 5227
rect 3753 5193 3767 5207
rect 3713 5173 3727 5187
rect 3633 5153 3647 5167
rect 3453 5073 3467 5087
rect 3499 5073 3513 5087
rect 3293 5013 3307 5027
rect 3413 5013 3427 5027
rect 3073 4834 3087 4848
rect 2933 4753 2947 4767
rect 3033 4753 3047 4767
rect 2913 4673 2927 4687
rect 2913 4613 2927 4627
rect 2833 4473 2847 4487
rect 2813 4373 2827 4387
rect 2793 4133 2807 4147
rect 2793 4053 2807 4067
rect 2773 4033 2787 4047
rect 2853 4413 2867 4427
rect 2913 4473 2927 4487
rect 3013 4633 3027 4647
rect 2973 4573 2987 4587
rect 2973 4532 2987 4546
rect 2933 4413 2947 4427
rect 3073 4812 3087 4826
rect 3133 4793 3147 4807
rect 3093 4693 3107 4707
rect 3133 4673 3147 4687
rect 3153 4633 3167 4647
rect 3273 4853 3287 4867
rect 3213 4819 3227 4833
rect 3253 4793 3267 4807
rect 3233 4693 3247 4707
rect 3493 4933 3507 4947
rect 3533 5033 3547 5047
rect 3513 4913 3527 4927
rect 3493 4853 3507 4867
rect 3473 4833 3487 4847
rect 3353 4813 3367 4827
rect 3313 4753 3327 4767
rect 3213 4573 3227 4587
rect 3293 4673 3307 4687
rect 3253 4653 3267 4667
rect 3253 4553 3267 4567
rect 3033 4533 3047 4547
rect 3193 4533 3207 4547
rect 3233 4532 3247 4546
rect 3053 4473 3067 4487
rect 3013 4373 3027 4387
rect 3073 4393 3087 4407
rect 3053 4353 3067 4367
rect 3013 4333 3027 4347
rect 3153 4353 3167 4367
rect 3093 4334 3107 4348
rect 2913 4313 2927 4327
rect 2873 4293 2887 4307
rect 2853 4273 2867 4287
rect 3093 4312 3107 4326
rect 3193 4314 3207 4328
rect 3013 4293 3027 4307
rect 2893 4253 2907 4267
rect 2972 4253 2986 4267
rect 2994 4253 3008 4267
rect 2853 4233 2867 4247
rect 2873 4153 2887 4167
rect 2873 4093 2887 4107
rect 2853 4034 2867 4048
rect 2813 4014 2827 4028
rect 2853 4012 2867 4026
rect 2773 3953 2787 3967
rect 2813 3933 2827 3947
rect 2753 3893 2767 3907
rect 2693 3853 2707 3867
rect 2833 3813 2847 3827
rect 2653 3794 2667 3808
rect 2713 3793 2727 3807
rect 2593 3693 2607 3707
rect 2573 3673 2587 3687
rect 2513 3653 2527 3667
rect 2493 3533 2507 3547
rect 2473 3512 2487 3526
rect 2573 3593 2587 3607
rect 2553 3513 2567 3527
rect 2393 3433 2407 3447
rect 2513 3433 2527 3447
rect 2413 3373 2427 3387
rect 2393 3353 2407 3367
rect 2393 3294 2407 3308
rect 2393 3133 2407 3147
rect 2373 3093 2387 3107
rect 2573 3433 2587 3447
rect 2433 3273 2447 3287
rect 2473 3093 2487 3107
rect 2113 2933 2127 2947
rect 2273 2933 2287 2947
rect 2073 2893 2087 2907
rect 1913 2813 1927 2827
rect 1993 2813 2007 2827
rect 1893 2793 1907 2807
rect 1953 2773 1967 2787
rect 2133 2773 2147 2787
rect 2313 2773 2327 2787
rect 1373 2473 1387 2487
rect 1433 2493 1447 2507
rect 1573 2493 1587 2507
rect 1773 2493 1787 2507
rect 1413 2473 1427 2487
rect 1493 2453 1507 2467
rect 1993 2713 2007 2727
rect 2373 2953 2387 2967
rect 2373 2793 2387 2807
rect 2433 2773 2447 2787
rect 2053 2733 2067 2747
rect 2113 2733 2127 2747
rect 2353 2733 2367 2747
rect 2193 2713 2207 2727
rect 1953 2693 1967 2707
rect 2013 2693 2027 2707
rect 2153 2693 2167 2707
rect 2193 2673 2207 2687
rect 2453 2633 2467 2647
rect 2393 2573 2407 2587
rect 1953 2533 1967 2547
rect 2073 2493 2087 2507
rect 1967 2473 1981 2487
rect 2353 2473 2367 2487
rect 1613 2453 1627 2467
rect 1793 2453 1807 2467
rect 1873 2453 1887 2467
rect 1393 2433 1407 2447
rect 1413 2433 1427 2447
rect 1313 2413 1327 2427
rect 1373 2413 1387 2427
rect 1253 2373 1267 2387
rect 1193 2293 1207 2307
rect 1433 2333 1447 2347
rect 1153 2233 1167 2247
rect 1113 2213 1127 2227
rect 633 1953 647 1967
rect 913 1954 927 1968
rect 1273 2173 1287 2187
rect 1313 2193 1327 2207
rect 933 1953 947 1967
rect 633 1833 647 1847
rect 673 1933 687 1947
rect 653 1813 667 1827
rect 673 1793 687 1807
rect 713 1793 727 1807
rect 913 1932 927 1946
rect 813 1773 827 1787
rect 733 1753 747 1767
rect 793 1753 807 1767
rect 733 1713 747 1727
rect 773 1553 787 1567
rect 593 1473 607 1487
rect 733 1473 747 1487
rect 453 1433 467 1447
rect 553 1434 567 1448
rect 453 1293 467 1307
rect 413 1273 427 1287
rect 473 1253 487 1267
rect 393 1193 407 1207
rect 353 1153 367 1167
rect 433 1153 447 1167
rect 333 993 347 1007
rect 433 973 447 987
rect 353 913 367 927
rect 633 1413 647 1427
rect 693 1414 707 1428
rect 493 1214 507 1228
rect 853 1733 867 1747
rect 833 1693 847 1707
rect 873 1693 887 1707
rect 853 1653 867 1667
rect 893 1653 907 1667
rect 873 1513 887 1527
rect 853 1473 867 1487
rect 953 1933 967 1947
rect 1013 1933 1027 1947
rect 1013 1753 1027 1767
rect 1033 1713 1047 1727
rect 1133 1713 1147 1727
rect 933 1593 947 1607
rect 973 1593 987 1607
rect 693 1392 707 1406
rect 773 1393 787 1407
rect 913 1393 927 1407
rect 593 1293 607 1307
rect 673 1293 687 1307
rect 873 1293 887 1307
rect 553 1233 567 1247
rect 533 1193 547 1207
rect 473 934 487 948
rect 513 1173 527 1187
rect 573 1193 587 1207
rect 673 1253 687 1267
rect 753 1233 767 1247
rect 613 1213 627 1227
rect 853 1193 867 1207
rect 953 1253 967 1267
rect 593 1173 607 1187
rect 633 1173 647 1187
rect 513 1133 527 1147
rect 513 973 527 987
rect 593 953 607 967
rect 573 933 587 947
rect 453 912 467 926
rect 373 813 387 827
rect 313 773 327 787
rect 213 733 227 747
rect 253 734 267 748
rect 253 693 267 707
rect 313 693 327 707
rect 413 693 427 707
rect 213 653 227 667
rect 293 653 307 667
rect 373 653 387 667
rect 433 653 447 667
rect 493 853 507 867
rect 533 693 547 707
rect 693 1053 707 1067
rect 813 1053 827 1067
rect 653 993 667 1007
rect 733 993 747 1007
rect 953 973 967 987
rect 1153 1513 1167 1527
rect 1053 1473 1067 1487
rect 993 1393 1007 1407
rect 1033 1373 1047 1387
rect 1013 1233 1027 1247
rect 1353 2133 1367 2147
rect 1293 2093 1307 2107
rect 1473 2173 1487 2187
rect 1473 2093 1487 2107
rect 1453 2053 1467 2067
rect 1553 2333 1567 2347
rect 1573 2253 1587 2267
rect 1613 2253 1627 2267
rect 1533 2093 1547 2107
rect 1513 2053 1527 2067
rect 1493 1974 1507 1988
rect 1633 2233 1647 2247
rect 1753 2253 1767 2267
rect 1713 2233 1727 2247
rect 1673 2173 1687 2187
rect 1693 2133 1707 2147
rect 1613 2053 1627 2067
rect 1753 1973 1767 1987
rect 1713 1953 1727 1967
rect 1733 1953 1747 1967
rect 1279 1933 1293 1947
rect 1493 1932 1507 1946
rect 1393 1873 1407 1887
rect 1193 1773 1207 1787
rect 1233 1753 1247 1767
rect 1373 1713 1387 1727
rect 1233 1693 1247 1707
rect 1340 1693 1353 1707
rect 1353 1693 1354 1707
rect 1693 1913 1707 1927
rect 1533 1793 1547 1807
rect 1493 1713 1507 1727
rect 1513 1713 1527 1727
rect 1393 1673 1407 1687
rect 1253 1633 1267 1647
rect 1553 1773 1567 1787
rect 1573 1753 1587 1767
rect 1173 1473 1187 1487
rect 1413 1473 1427 1487
rect 1533 1473 1547 1487
rect 1153 1433 1167 1447
rect 1213 1433 1227 1447
rect 1293 1433 1307 1447
rect 1313 1433 1327 1447
rect 1353 1433 1367 1447
rect 1093 1393 1107 1407
rect 1473 1433 1487 1447
rect 1553 1433 1567 1447
rect 1673 1873 1687 1887
rect 1953 2433 1967 2447
rect 1913 2393 1927 2407
rect 1973 2393 1987 2407
rect 1913 2353 1927 2367
rect 2293 2433 2307 2447
rect 2113 2413 2127 2427
rect 2213 2413 2227 2427
rect 2313 2413 2327 2427
rect 1993 2333 2007 2347
rect 2073 2333 2087 2347
rect 2173 2333 2187 2347
rect 1873 2267 1887 2281
rect 1833 2253 1847 2267
rect 1893 2253 1907 2267
rect 1813 2213 1827 2227
rect 1833 2213 1847 2227
rect 2033 2253 2047 2267
rect 1893 2053 1907 2067
rect 1873 1993 1887 2007
rect 1813 1973 1827 1987
rect 1773 1833 1787 1847
rect 1713 1793 1727 1807
rect 1833 1953 1847 1967
rect 1933 1993 1947 2007
rect 2333 2313 2347 2327
rect 2193 2253 2207 2267
rect 2273 2253 2287 2267
rect 2293 2253 2307 2267
rect 2333 2253 2347 2267
rect 2233 2233 2247 2247
rect 2033 2193 2047 2207
rect 2293 2193 2307 2207
rect 1993 1973 2007 1987
rect 1973 1913 1987 1927
rect 1793 1753 1807 1767
rect 1633 1713 1647 1727
rect 1673 1713 1687 1727
rect 1813 1713 1827 1727
rect 1613 1673 1627 1687
rect 1673 1673 1687 1687
rect 1613 1573 1627 1587
rect 1493 1413 1507 1427
rect 1373 1393 1387 1407
rect 1433 1393 1447 1407
rect 1153 1373 1167 1387
rect 1113 1313 1127 1327
rect 1213 1313 1227 1327
rect 1293 1273 1307 1287
rect 1133 1253 1147 1267
rect 1473 1353 1487 1367
rect 1553 1353 1567 1367
rect 1513 1333 1527 1347
rect 1453 1313 1467 1327
rect 1433 1253 1447 1267
rect 1413 1233 1427 1247
rect 1473 1273 1487 1287
rect 1273 1193 1287 1207
rect 1013 1133 1027 1147
rect 1233 1133 1247 1147
rect 1053 973 1067 987
rect 853 953 867 967
rect 613 873 627 887
rect 693 873 707 887
rect 773 873 787 887
rect 713 673 727 687
rect 573 653 587 667
rect 1013 933 1027 947
rect 1073 933 1087 947
rect 1173 933 1187 947
rect 1053 873 1067 887
rect 1013 813 1027 827
rect 873 693 887 707
rect 913 673 927 687
rect 713 633 727 647
rect 773 653 787 667
rect 813 653 827 667
rect 513 613 527 627
rect 673 613 687 627
rect 453 553 467 567
rect 533 553 547 567
rect 533 513 547 527
rect 273 493 287 507
rect 513 493 527 507
rect 333 373 347 387
rect 33 353 47 367
rect 93 353 107 367
rect 133 353 147 367
rect 113 333 127 347
rect 213 333 227 347
rect 93 293 107 307
rect 133 293 147 307
rect 393 333 407 347
rect 253 273 267 287
rect 293 273 307 287
rect 413 273 427 287
rect 133 193 147 207
rect 93 173 107 187
rect 113 173 127 187
rect 333 193 347 207
rect 253 173 267 187
rect 73 133 87 147
rect 133 133 147 147
rect 233 133 247 147
rect 293 133 307 147
rect 273 113 287 127
rect 873 613 887 627
rect 913 613 927 627
rect 953 673 967 687
rect 1053 673 1067 687
rect 953 633 967 647
rect 833 533 847 547
rect 753 453 767 467
rect 573 333 587 347
rect 553 273 567 287
rect 886 413 887 427
rect 887 413 900 427
rect 739 373 753 387
rect 853 353 867 367
rect 873 353 887 367
rect 1513 1193 1527 1207
rect 1553 1193 1567 1207
rect 1473 1113 1487 1127
rect 1273 933 1287 947
rect 1413 933 1427 947
rect 1473 913 1487 927
rect 1553 913 1567 927
rect 1153 733 1167 747
rect 1113 673 1127 687
rect 1313 893 1327 907
rect 1433 713 1447 727
rect 1613 1073 1627 1087
rect 1633 953 1647 967
rect 1873 1773 1887 1787
rect 1873 1713 1887 1727
rect 1893 1613 1907 1627
rect 1993 1833 2007 1847
rect 1953 1733 1967 1747
rect 2373 2453 2387 2467
rect 2413 2333 2427 2347
rect 2373 2293 2387 2307
rect 2453 2293 2467 2307
rect 2453 2233 2467 2247
rect 2653 3772 2667 3786
rect 2933 4013 2947 4027
rect 3373 4793 3387 4807
rect 3373 4753 3387 4767
rect 3353 4713 3367 4727
rect 3493 4793 3507 4807
rect 3413 4693 3427 4707
rect 3413 4653 3427 4667
rect 3373 4633 3387 4647
rect 3453 4573 3467 4587
rect 3433 4553 3447 4567
rect 3473 4533 3487 4547
rect 3273 4433 3287 4447
rect 3353 4473 3367 4487
rect 3373 4453 3387 4467
rect 3353 4413 3367 4427
rect 3453 4473 3467 4487
rect 3333 4393 3347 4407
rect 3413 4393 3427 4407
rect 3353 4373 3367 4387
rect 3333 4353 3347 4367
rect 3413 4353 3427 4367
rect 3393 4293 3407 4307
rect 3133 4273 3147 4287
rect 3173 4272 3187 4286
rect 3033 4193 3047 4207
rect 3093 4193 3107 4207
rect 3013 4053 3027 4067
rect 3053 4053 3067 4067
rect 3113 4053 3127 4067
rect 3332 4193 3346 4207
rect 3354 4193 3368 4207
rect 3273 4133 3287 4147
rect 3193 4113 3207 4127
rect 3193 4073 3207 4087
rect 2953 3993 2967 4007
rect 2993 3953 3007 3967
rect 2873 3913 2887 3927
rect 2973 3913 2987 3927
rect 2953 3873 2967 3887
rect 2913 3833 2927 3847
rect 2773 3753 2787 3767
rect 2833 3733 2847 3747
rect 2793 3673 2807 3687
rect 2733 3553 2747 3567
rect 2693 3473 2707 3487
rect 2613 3353 2627 3367
rect 2593 3333 2607 3347
rect 2713 3333 2727 3347
rect 2613 3273 2627 3287
rect 2653 3253 2667 3267
rect 2673 3253 2687 3267
rect 2553 3193 2567 3207
rect 2533 2993 2547 3007
rect 2493 2953 2507 2967
rect 2693 3173 2707 3187
rect 2713 3153 2727 3167
rect 2693 3093 2707 3107
rect 2673 3013 2687 3027
rect 2913 3793 2927 3807
rect 2953 3793 2967 3807
rect 2893 3653 2907 3667
rect 2893 3613 2907 3627
rect 2933 3513 2947 3527
rect 2813 3393 2827 3407
rect 2913 3333 2927 3347
rect 2893 3273 2907 3287
rect 2993 3253 3007 3267
rect 2967 3233 2981 3247
rect 2753 3213 2767 3227
rect 2853 3213 2867 3227
rect 2913 3212 2927 3226
rect 2833 3053 2847 3067
rect 2713 2953 2727 2967
rect 2513 2933 2527 2947
rect 2553 2893 2567 2907
rect 2553 2793 2567 2807
rect 2653 2773 2667 2787
rect 2493 2733 2507 2747
rect 2693 2713 2707 2727
rect 3073 4013 3087 4027
rect 3033 3973 3047 3987
rect 3073 3972 3087 3986
rect 3053 3913 3067 3927
rect 3173 4047 3187 4061
rect 3353 4153 3367 4167
rect 3293 4033 3307 4047
rect 3213 3993 3227 4007
rect 3193 3973 3207 3987
rect 3333 3993 3347 4007
rect 3373 3993 3387 4007
rect 3353 3973 3367 3987
rect 3113 3953 3127 3967
rect 3253 3953 3267 3967
rect 3293 3953 3307 3967
rect 3153 3933 3167 3947
rect 3273 3933 3287 3947
rect 3173 3893 3187 3907
rect 3153 3873 3167 3887
rect 3153 3833 3167 3847
rect 3033 3514 3047 3528
rect 3033 3492 3047 3506
rect 3213 3873 3227 3887
rect 3173 3813 3187 3827
rect 3233 3813 3247 3827
rect 3193 3733 3207 3747
rect 3193 3673 3207 3687
rect 3353 3893 3367 3907
rect 3293 3833 3307 3847
rect 3353 3833 3367 3847
rect 3333 3773 3347 3787
rect 3173 3513 3187 3527
rect 3113 3473 3127 3487
rect 3093 3433 3107 3447
rect 3073 3413 3087 3427
rect 3033 3353 3047 3367
rect 3153 3393 3167 3407
rect 3393 3893 3407 3907
rect 3433 4333 3447 4347
rect 3633 5013 3647 5027
rect 3713 5053 3727 5067
rect 3713 4993 3727 5007
rect 3673 4933 3687 4947
rect 3653 4914 3667 4928
rect 3773 5153 3787 5167
rect 3793 5133 3807 5147
rect 3753 5093 3767 5107
rect 3813 5113 3827 5127
rect 3752 5053 3766 5067
rect 3774 5053 3788 5067
rect 4153 5393 4167 5407
rect 4013 5373 4027 5387
rect 4093 5373 4107 5387
rect 3873 5313 3887 5327
rect 3953 5273 3967 5287
rect 3953 5213 3967 5227
rect 3893 5173 3907 5187
rect 3873 5133 3887 5147
rect 3793 5013 3807 5027
rect 3733 4953 3747 4967
rect 3653 4892 3667 4906
rect 3693 4893 3707 4907
rect 3853 4993 3867 5007
rect 3893 5093 3907 5107
rect 4293 5353 4307 5367
rect 4033 5313 4047 5327
rect 4013 5213 4027 5227
rect 3993 5173 4007 5187
rect 3973 5133 3987 5147
rect 4073 5213 4087 5227
rect 3973 5073 3987 5087
rect 4013 5073 4027 5087
rect 4033 5073 4047 5087
rect 3913 5053 3927 5067
rect 4013 5052 4027 5066
rect 4133 5313 4147 5327
rect 4173 5313 4187 5327
rect 4173 5193 4187 5207
rect 4093 5173 4107 5187
rect 4413 5453 4427 5467
rect 4373 5413 4387 5427
rect 4413 5413 4427 5427
rect 4353 5373 4367 5387
rect 4213 5313 4227 5327
rect 4253 5253 4267 5267
rect 4213 5193 4227 5207
rect 4113 5113 4127 5127
rect 4193 5114 4207 5128
rect 4033 5013 4047 5027
rect 4013 4993 4027 5007
rect 3853 4953 3867 4967
rect 3933 4953 3947 4967
rect 3973 4953 3987 4967
rect 3573 4813 3587 4827
rect 3573 4773 3587 4787
rect 3573 4693 3587 4707
rect 3573 4533 3587 4547
rect 3613 4833 3627 4847
rect 3633 4793 3647 4807
rect 3673 4793 3687 4807
rect 3673 4713 3687 4727
rect 3673 4673 3687 4687
rect 3733 4833 3747 4847
rect 3833 4853 3847 4867
rect 3733 4733 3747 4747
rect 3693 4653 3707 4667
rect 3613 4593 3627 4607
rect 3613 4532 3627 4546
rect 3653 4533 3667 4547
rect 3733 4653 3747 4667
rect 3793 4793 3807 4807
rect 3893 4933 3907 4947
rect 3953 4893 3967 4907
rect 3893 4853 3907 4867
rect 3907 4793 3921 4807
rect 3853 4773 3867 4787
rect 3873 4753 3887 4767
rect 3833 4653 3847 4667
rect 3773 4593 3787 4607
rect 3713 4533 3727 4547
rect 3613 4493 3627 4507
rect 3593 4473 3607 4487
rect 3633 4473 3647 4487
rect 3553 4433 3567 4447
rect 3593 4433 3607 4447
rect 3533 4393 3547 4407
rect 3513 4293 3527 4307
rect 3493 4273 3507 4287
rect 3513 4253 3527 4267
rect 3453 4233 3467 4247
rect 3493 4133 3507 4147
rect 3453 4093 3467 4107
rect 3433 4034 3447 4048
rect 3433 3973 3447 3987
rect 3553 4293 3567 4307
rect 3553 4233 3567 4247
rect 3573 4153 3587 4167
rect 3553 4133 3567 4147
rect 3533 4093 3547 4107
rect 3693 4453 3707 4467
rect 3653 4433 3667 4447
rect 3713 4413 3727 4427
rect 3693 4393 3707 4407
rect 3673 4333 3687 4347
rect 4213 5013 4227 5027
rect 4233 4993 4247 5007
rect 4193 4953 4207 4967
rect 4233 4913 4247 4927
rect 4033 4893 4047 4907
rect 4053 4873 4067 4887
rect 3973 4833 3987 4847
rect 4033 4753 4047 4767
rect 3953 4733 3967 4747
rect 3933 4693 3947 4707
rect 3913 4593 3927 4607
rect 3993 4593 4007 4607
rect 3893 4573 3907 4587
rect 4233 4832 4247 4846
rect 4173 4793 4187 4807
rect 4233 4753 4247 4767
rect 4133 4693 4147 4707
rect 4233 4673 4247 4687
rect 4153 4653 4167 4667
rect 3893 4533 3907 4547
rect 3813 4513 3827 4527
rect 3773 4494 3787 4508
rect 3793 4472 3807 4486
rect 3813 4393 3827 4407
rect 3793 4373 3807 4387
rect 3873 4433 3887 4447
rect 3833 4373 3847 4387
rect 3793 4333 3807 4347
rect 3633 4293 3647 4307
rect 3613 4273 3627 4287
rect 3673 4273 3687 4287
rect 3693 4253 3707 4267
rect 3613 4233 3627 4247
rect 3633 4213 3647 4227
rect 3613 4113 3627 4127
rect 3473 4033 3487 4047
rect 3533 4033 3547 4047
rect 3593 4034 3607 4048
rect 3453 3913 3467 3927
rect 3413 3834 3427 3848
rect 3433 3812 3447 3826
rect 3673 4093 3687 4107
rect 3873 4313 3887 4327
rect 3913 4513 3927 4527
rect 3953 4513 3967 4527
rect 3913 4373 3927 4387
rect 3733 4253 3747 4267
rect 3833 4273 3847 4287
rect 3993 4453 4007 4467
rect 3973 4413 3987 4427
rect 3933 4293 3947 4307
rect 4093 4513 4107 4527
rect 4173 4514 4187 4528
rect 4052 4473 4066 4487
rect 4074 4473 4088 4487
rect 4053 4433 4067 4447
rect 4033 4373 4047 4387
rect 4113 4373 4127 4387
rect 4013 4313 4027 4327
rect 3993 4293 4007 4307
rect 3913 4253 3927 4267
rect 3833 4233 3847 4247
rect 3713 4133 3727 4147
rect 3693 4073 3707 4087
rect 3633 4033 3647 4047
rect 3613 4013 3627 4027
rect 3553 3973 3567 3987
rect 3593 3893 3607 3907
rect 3553 3873 3567 3887
rect 3493 3813 3507 3827
rect 3753 4093 3767 4107
rect 3713 4033 3727 4047
rect 3773 4013 3787 4027
rect 3653 3933 3667 3947
rect 3633 3893 3647 3907
rect 3393 3753 3407 3767
rect 3393 3713 3407 3727
rect 3233 3633 3247 3647
rect 3353 3633 3367 3647
rect 3213 3553 3227 3567
rect 3193 3333 3207 3347
rect 3113 3253 3127 3267
rect 3173 3233 3187 3247
rect 3073 3193 3087 3207
rect 3333 3593 3347 3607
rect 3293 3493 3307 3507
rect 3353 3553 3367 3567
rect 3353 3493 3367 3507
rect 3433 3493 3447 3507
rect 3333 3473 3347 3487
rect 3333 3413 3347 3427
rect 3513 3773 3527 3787
rect 3593 3774 3607 3788
rect 3533 3753 3547 3767
rect 3593 3752 3607 3766
rect 3493 3653 3507 3667
rect 3553 3513 3567 3527
rect 3533 3493 3547 3507
rect 3473 3473 3487 3487
rect 3453 3433 3467 3447
rect 3413 3373 3427 3387
rect 3433 3353 3447 3367
rect 3273 3273 3287 3287
rect 3353 3293 3367 3307
rect 3379 3293 3393 3307
rect 3293 3193 3307 3207
rect 3013 3153 3027 3167
rect 3173 3153 3187 3167
rect 3233 3153 3247 3167
rect 2953 3053 2967 3067
rect 2933 2993 2947 3007
rect 2853 2933 2867 2947
rect 2713 2673 2727 2687
rect 2753 2673 2767 2687
rect 2833 2673 2847 2687
rect 2653 2573 2667 2587
rect 2533 2493 2547 2507
rect 2533 2453 2547 2467
rect 2573 2433 2587 2447
rect 2553 2333 2567 2347
rect 2393 2193 2407 2207
rect 2353 2073 2367 2087
rect 2513 2233 2527 2247
rect 2493 2153 2507 2167
rect 2453 2053 2467 2067
rect 2513 2013 2527 2027
rect 2273 1973 2287 1987
rect 2113 1953 2127 1967
rect 2453 1953 2467 1967
rect 2093 1913 2107 1927
rect 2133 1913 2147 1927
rect 2173 1913 2187 1927
rect 2033 1673 2047 1687
rect 1933 1613 1947 1627
rect 1913 1573 1927 1587
rect 1773 1533 1787 1547
rect 1833 1533 1847 1547
rect 1753 1454 1767 1468
rect 1753 1432 1767 1446
rect 1713 1379 1727 1393
rect 1693 1333 1707 1347
rect 1713 1313 1727 1327
rect 1713 1153 1727 1167
rect 1893 1513 1907 1527
rect 1793 1453 1807 1467
rect 1773 1313 1787 1327
rect 1913 1473 1927 1487
rect 1833 1433 1847 1447
rect 1893 1412 1907 1426
rect 1853 1393 1867 1407
rect 1813 1293 1827 1307
rect 1813 1193 1827 1207
rect 1953 1433 1967 1447
rect 1993 1433 2007 1447
rect 1933 1414 1947 1428
rect 2193 1833 2207 1847
rect 2073 1753 2087 1767
rect 2313 1913 2327 1927
rect 2513 1913 2527 1927
rect 2373 1833 2387 1847
rect 2473 1833 2487 1847
rect 2273 1753 2287 1767
rect 2153 1714 2167 1728
rect 2193 1712 2207 1726
rect 2153 1692 2167 1706
rect 2173 1693 2187 1707
rect 2093 1613 2107 1627
rect 2273 1673 2287 1687
rect 2253 1633 2267 1647
rect 2193 1513 2207 1527
rect 2173 1433 2187 1447
rect 1933 1333 1947 1347
rect 2033 1353 2047 1367
rect 1973 1293 1987 1307
rect 1973 1233 1987 1247
rect 1913 1194 1927 1208
rect 2013 1213 2027 1227
rect 1873 1173 1887 1187
rect 1893 1173 1907 1187
rect 1753 1133 1767 1147
rect 1873 1013 1887 1027
rect 1667 933 1681 947
rect 1713 953 1727 967
rect 1753 913 1767 927
rect 2173 1353 2187 1367
rect 2053 1313 2067 1327
rect 2053 1213 2067 1227
rect 2673 2453 2687 2467
rect 2653 2393 2667 2407
rect 2593 2333 2607 2347
rect 2593 2193 2607 2207
rect 2633 2113 2647 2127
rect 2693 2113 2707 2127
rect 2593 2073 2607 2087
rect 2653 2053 2667 2067
rect 2673 1953 2687 1967
rect 2573 1813 2587 1827
rect 2453 1793 2467 1807
rect 2393 1693 2407 1707
rect 2473 1753 2487 1767
rect 2513 1713 2527 1727
rect 2473 1673 2487 1687
rect 2613 1673 2627 1687
rect 2453 1573 2467 1587
rect 2393 1513 2407 1527
rect 2373 1474 2387 1488
rect 2413 1473 2427 1487
rect 2273 1373 2287 1387
rect 2333 1373 2347 1387
rect 2273 1214 2287 1228
rect 2093 1193 2107 1207
rect 2193 1194 2207 1208
rect 2033 1173 2047 1187
rect 2053 1173 2067 1187
rect 2113 1173 2127 1187
rect 2013 1053 2027 1067
rect 2013 1013 2027 1027
rect 1933 993 1947 1007
rect 1973 993 1987 1007
rect 1913 913 1927 927
rect 1593 893 1607 907
rect 1153 652 1167 666
rect 1073 633 1087 647
rect 1033 533 1047 547
rect 1113 513 1127 527
rect 953 333 967 347
rect 1093 394 1107 408
rect 1093 372 1107 386
rect 1013 333 1027 347
rect 853 293 867 307
rect 973 293 987 307
rect 593 253 607 267
rect 513 193 527 207
rect 793 193 807 207
rect 433 173 447 187
rect 473 153 487 167
rect 713 173 727 187
rect 753 173 767 187
rect 413 113 427 127
rect 593 153 607 167
rect 893 193 907 207
rect 953 153 967 167
rect 1033 153 1047 167
rect 1553 713 1567 727
rect 1613 693 1627 707
rect 1753 693 1767 707
rect 1513 653 1527 667
rect 1553 653 1567 667
rect 1633 653 1647 667
rect 1653 653 1667 667
rect 1626 593 1627 607
rect 1627 593 1640 607
rect 1373 553 1387 567
rect 1233 493 1247 507
rect 1273 493 1287 507
rect 1233 453 1247 467
rect 1333 453 1347 467
rect 1193 373 1207 387
rect 1313 373 1327 387
rect 1553 493 1567 507
rect 1433 453 1447 467
rect 1353 393 1367 407
rect 1793 553 1807 567
rect 1833 553 1847 567
rect 1793 513 1807 527
rect 1753 493 1767 507
rect 1713 453 1727 467
rect 1913 753 1927 767
rect 1973 953 1987 967
rect 1953 893 1967 907
rect 1993 933 2007 947
rect 1973 693 1987 707
rect 2173 1172 2187 1186
rect 2253 1173 2267 1187
rect 2273 1173 2287 1187
rect 2294 1173 2308 1187
rect 2239 1133 2253 1147
rect 2213 1053 2227 1067
rect 2833 2493 2847 2507
rect 2773 2473 2787 2487
rect 2873 2793 2887 2807
rect 3233 3053 3247 3067
rect 3353 3193 3367 3207
rect 3313 3133 3327 3147
rect 3333 3093 3347 3107
rect 3733 3873 3747 3887
rect 3773 3853 3787 3867
rect 3753 3833 3767 3847
rect 3913 4213 3927 4227
rect 3873 4173 3887 4187
rect 3853 4133 3867 4147
rect 3833 3853 3847 3867
rect 4093 4313 4107 4327
rect 4173 4492 4187 4506
rect 4213 4532 4227 4546
rect 4233 4433 4247 4447
rect 4172 4393 4186 4407
rect 4194 4393 4208 4407
rect 4233 4393 4247 4407
rect 4053 4293 4067 4307
rect 4073 4253 4087 4267
rect 4013 4133 4027 4147
rect 4053 4093 4067 4107
rect 4013 4073 4027 4087
rect 3913 4053 3927 4067
rect 3953 4053 3967 4067
rect 4153 4333 4167 4347
rect 4353 5293 4367 5307
rect 4273 5193 4287 5207
rect 4273 5153 4287 5167
rect 4293 5113 4307 5127
rect 4293 4953 4307 4967
rect 4273 4813 4287 4827
rect 4393 5093 4407 5107
rect 4393 4993 4407 5007
rect 4473 5453 4487 5467
rect 4433 5253 4447 5267
rect 4433 5113 4447 5127
rect 4413 4973 4427 4987
rect 4393 4853 4407 4867
rect 4453 4833 4467 4847
rect 4313 4813 4327 4827
rect 4393 4813 4407 4827
rect 4293 4793 4307 4807
rect 4433 4813 4447 4827
rect 4353 4733 4367 4747
rect 4273 4473 4287 4487
rect 4353 4553 4367 4567
rect 4413 4539 4427 4553
rect 4693 5413 4707 5427
rect 4792 5413 4806 5427
rect 4814 5413 4828 5427
rect 4973 5433 4987 5447
rect 4933 5413 4947 5427
rect 4573 5373 4587 5387
rect 4733 5373 4747 5387
rect 4873 5373 4887 5387
rect 4933 5373 4947 5387
rect 4533 5334 4547 5348
rect 4733 5333 4747 5347
rect 4533 5293 4547 5307
rect 4493 5253 4507 5267
rect 4573 5253 4587 5267
rect 4573 5173 4587 5187
rect 4493 5153 4507 5167
rect 4533 5113 4547 5127
rect 4493 5073 4507 5087
rect 4553 5073 4567 5087
rect 4493 5033 4507 5047
rect 4593 5093 4607 5107
rect 4513 4913 4527 4927
rect 4573 4913 4587 4927
rect 4773 5313 4787 5327
rect 4793 5313 4807 5327
rect 4773 5173 4787 5187
rect 5253 5393 5267 5407
rect 5073 5373 5087 5387
rect 5233 5373 5247 5387
rect 4973 5353 4987 5367
rect 4913 5333 4927 5347
rect 4833 5134 4847 5148
rect 4833 5112 4847 5126
rect 4753 5093 4767 5107
rect 4633 5053 4647 5067
rect 4673 5033 4687 5047
rect 4713 5033 4727 5047
rect 4613 5013 4627 5027
rect 4613 4893 4627 4907
rect 4553 4853 4567 4867
rect 4593 4853 4607 4867
rect 4573 4833 4587 4847
rect 4493 4733 4507 4747
rect 4473 4633 4487 4647
rect 4313 4513 4327 4527
rect 4393 4513 4407 4527
rect 4473 4533 4487 4547
rect 4293 4393 4307 4407
rect 4253 4353 4267 4367
rect 4453 4413 4467 4427
rect 4693 5013 4707 5027
rect 4753 4973 4767 4987
rect 4693 4873 4707 4887
rect 4793 4873 4807 4887
rect 4693 4753 4707 4767
rect 4653 4733 4667 4747
rect 4633 4693 4647 4707
rect 5433 5413 5447 5427
rect 5493 5413 5507 5427
rect 5353 5393 5367 5407
rect 5413 5393 5427 5407
rect 5333 5353 5347 5367
rect 5373 5353 5387 5367
rect 5053 5333 5067 5347
rect 5033 5313 5047 5327
rect 4873 5093 4887 5107
rect 4853 5053 4867 5067
rect 4893 4933 4907 4947
rect 4813 4773 4827 4787
rect 4813 4713 4827 4727
rect 4893 4693 4907 4707
rect 4773 4673 4787 4687
rect 4713 4613 4727 4627
rect 4673 4574 4687 4588
rect 4733 4573 4747 4587
rect 4567 4554 4581 4568
rect 4513 4493 4527 4507
rect 4493 4373 4507 4387
rect 4673 4552 4687 4566
rect 4553 4532 4567 4546
rect 4693 4532 4707 4546
rect 4653 4413 4667 4427
rect 4553 4373 4567 4387
rect 4393 4333 4407 4347
rect 4473 4333 4487 4347
rect 4193 4273 4207 4287
rect 4153 4153 4167 4167
rect 4173 4053 4187 4067
rect 3893 3993 3907 4007
rect 3873 3834 3887 3848
rect 3793 3813 3807 3827
rect 3833 3813 3847 3827
rect 3813 3793 3827 3807
rect 3913 3973 3927 3987
rect 3973 3873 3987 3887
rect 4253 4273 4267 4287
rect 4273 4193 4287 4207
rect 4213 4053 4227 4067
rect 4353 4053 4367 4067
rect 4233 4033 4247 4047
rect 4293 4033 4307 4047
rect 4193 3993 4207 4007
rect 4073 3973 4087 3987
rect 4173 3973 4187 3987
rect 3913 3813 3927 3827
rect 3933 3773 3947 3787
rect 3993 3773 4007 3787
rect 3953 3753 3967 3767
rect 3793 3733 3807 3747
rect 3833 3733 3847 3747
rect 3873 3733 3887 3747
rect 3693 3713 3707 3727
rect 3733 3713 3747 3727
rect 3773 3713 3787 3727
rect 3713 3673 3727 3687
rect 3653 3613 3667 3627
rect 3653 3573 3667 3587
rect 3633 3547 3647 3561
rect 3713 3472 3727 3486
rect 3713 3433 3727 3447
rect 3653 3413 3667 3427
rect 3553 3353 3567 3367
rect 3593 3353 3607 3367
rect 3513 3333 3527 3347
rect 3573 3273 3587 3287
rect 3433 3253 3447 3267
rect 3499 3253 3513 3267
rect 3593 3233 3607 3247
rect 3393 3173 3407 3187
rect 3433 3153 3447 3167
rect 3373 3093 3387 3107
rect 3353 3073 3367 3087
rect 3333 3033 3347 3047
rect 3073 2953 3087 2967
rect 3173 2953 3187 2967
rect 3413 3053 3427 3067
rect 3386 2993 3387 3007
rect 3387 2993 3400 3007
rect 3293 2973 3307 2987
rect 3353 2973 3367 2987
rect 3253 2893 3267 2907
rect 3493 3093 3507 3107
rect 3753 3613 3767 3627
rect 3773 3574 3787 3588
rect 3773 3552 3787 3566
rect 3773 3513 3787 3527
rect 4133 3873 4147 3887
rect 4113 3793 4127 3807
rect 4593 4333 4607 4347
rect 4753 4513 4767 4527
rect 4793 4473 4807 4487
rect 4813 4393 4827 4407
rect 4873 4393 4887 4407
rect 4753 4313 4767 4327
rect 4833 4314 4847 4328
rect 4933 5033 4947 5047
rect 4993 5093 5007 5107
rect 5113 5273 5127 5287
rect 5093 5153 5107 5167
rect 5073 5113 5087 5127
rect 4993 5033 5007 5047
rect 4973 4933 4987 4947
rect 4973 4853 4987 4867
rect 5113 5113 5127 5127
rect 5293 5333 5307 5347
rect 5353 5332 5367 5346
rect 5453 5353 5467 5367
rect 5393 5313 5407 5327
rect 5473 5313 5487 5327
rect 5333 5153 5347 5167
rect 5233 5134 5247 5148
rect 5293 5133 5307 5147
rect 5213 5112 5227 5126
rect 5193 5074 5207 5088
rect 5333 5113 5347 5127
rect 5313 5073 5327 5087
rect 5373 5073 5387 5087
rect 5293 5053 5307 5067
rect 5433 5073 5447 5087
rect 5193 5033 5207 5047
rect 5173 4993 5187 5007
rect 5433 4953 5447 4967
rect 5333 4893 5347 4907
rect 5173 4853 5187 4867
rect 4933 4813 4947 4827
rect 4913 4653 4927 4667
rect 4933 4573 4947 4587
rect 4993 4653 5007 4667
rect 5013 4573 5027 4587
rect 4913 4513 4927 4527
rect 4993 4513 5007 4527
rect 5053 4813 5067 4827
rect 5073 4773 5087 4787
rect 5253 4833 5267 4847
rect 5273 4833 5287 4847
rect 5193 4813 5207 4827
rect 5513 4993 5527 5007
rect 5493 4893 5507 4907
rect 5473 4834 5487 4848
rect 5513 4833 5527 4847
rect 5373 4773 5387 4787
rect 5433 4773 5447 4787
rect 5252 4573 5266 4587
rect 5274 4573 5288 4587
rect 5333 4573 5347 4587
rect 5153 4553 5167 4567
rect 5393 4553 5407 4567
rect 5213 4533 5227 4547
rect 5073 4513 5087 4527
rect 5113 4513 5127 4527
rect 5173 4513 5187 4527
rect 4893 4333 4907 4347
rect 4473 4273 4487 4287
rect 4513 4273 4527 4287
rect 4633 4273 4647 4287
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4453 4093 4467 4107
rect 4693 4173 4707 4187
rect 4533 4153 4547 4167
rect 4473 4033 4487 4047
rect 4313 3993 4327 4007
rect 4433 3973 4447 3987
rect 4233 3913 4247 3927
rect 4333 3913 4347 3927
rect 4193 3793 4207 3807
rect 4173 3773 4187 3787
rect 4513 3913 4527 3927
rect 4353 3813 4367 3827
rect 4293 3793 4307 3807
rect 4153 3753 4167 3767
rect 4073 3673 4087 3687
rect 3833 3653 3847 3667
rect 4033 3653 4047 3667
rect 3813 3573 3827 3587
rect 3933 3633 3947 3647
rect 3893 3613 3907 3627
rect 3833 3513 3847 3527
rect 3873 3473 3887 3487
rect 3873 3353 3887 3367
rect 3913 3593 3927 3607
rect 3933 3553 3947 3567
rect 3953 3513 3967 3527
rect 3913 3493 3927 3507
rect 4073 3533 4087 3547
rect 3913 3453 3927 3467
rect 3993 3453 4007 3467
rect 3793 3273 3807 3287
rect 3813 3273 3827 3287
rect 4033 3453 4047 3467
rect 4013 3413 4027 3427
rect 4133 3513 4147 3527
rect 4233 3733 4247 3747
rect 4193 3713 4207 3727
rect 4173 3593 4187 3607
rect 4273 3673 4287 3687
rect 4253 3573 4267 3587
rect 4233 3533 4247 3547
rect 4253 3493 4267 3507
rect 4053 3433 4067 3447
rect 4173 3393 4187 3407
rect 4173 3353 4187 3367
rect 4033 3313 4047 3327
rect 3693 3213 3707 3227
rect 3633 3193 3647 3207
rect 4053 3293 4067 3307
rect 4173 3293 4187 3307
rect 4133 3273 4147 3287
rect 4433 3753 4447 3767
rect 4433 3713 4447 3727
rect 4393 3613 4407 3627
rect 4393 3533 4407 3547
rect 4593 4093 4607 4107
rect 4593 4034 4607 4048
rect 4593 4012 4607 4026
rect 4633 3913 4647 3927
rect 4612 3713 4626 3727
rect 4634 3713 4648 3727
rect 4573 3693 4587 3707
rect 4533 3673 4547 3687
rect 4473 3633 4487 3647
rect 4473 3573 4487 3587
rect 4553 3573 4567 3587
rect 4493 3533 4507 3547
rect 4353 3493 4367 3507
rect 4393 3493 4407 3507
rect 4313 3353 4327 3367
rect 4373 3313 4387 3327
rect 4513 3493 4527 3507
rect 4573 3493 4587 3507
rect 4533 3413 4547 3427
rect 4193 3253 4207 3267
rect 4253 3253 4267 3267
rect 3953 3233 3967 3247
rect 4113 3233 4127 3247
rect 4153 3233 4167 3247
rect 3733 3093 3747 3107
rect 3873 3093 3887 3107
rect 3613 3033 3627 3047
rect 3833 3007 3847 3021
rect 4273 3033 4287 3047
rect 4253 3013 4267 3027
rect 4193 2993 4207 3007
rect 3473 2953 3487 2967
rect 3433 2933 3447 2947
rect 3393 2873 3407 2887
rect 3073 2813 3087 2827
rect 3413 2813 3427 2827
rect 3033 2794 3047 2808
rect 3233 2753 3247 2767
rect 3053 2733 3067 2747
rect 2893 2673 2907 2687
rect 2873 2493 2887 2507
rect 3013 2653 3027 2667
rect 3193 2733 3207 2747
rect 3253 2713 3267 2727
rect 3613 2913 3627 2927
rect 3753 2953 3767 2967
rect 3653 2793 3667 2807
rect 3433 2773 3447 2787
rect 3493 2753 3507 2767
rect 3613 2753 3627 2767
rect 3713 2753 3727 2767
rect 3373 2733 3387 2747
rect 3593 2713 3607 2727
rect 3633 2713 3647 2727
rect 3273 2653 3287 2667
rect 3413 2653 3427 2667
rect 3133 2633 3147 2647
rect 3133 2553 3147 2567
rect 3293 2513 3307 2527
rect 2939 2473 2953 2487
rect 3153 2473 3167 2487
rect 3273 2473 3287 2487
rect 2812 2393 2826 2407
rect 2834 2393 2848 2407
rect 2813 2273 2827 2287
rect 2893 2453 2907 2467
rect 3033 2453 3047 2467
rect 2913 2433 2927 2447
rect 3093 2453 3107 2467
rect 3073 2413 3087 2427
rect 2953 2393 2967 2407
rect 3073 2353 3087 2367
rect 3033 2293 3047 2307
rect 2973 2273 2987 2287
rect 2873 2253 2887 2267
rect 2853 2193 2867 2207
rect 3313 2433 3327 2447
rect 3233 2353 3247 2367
rect 3113 2333 3127 2347
rect 3193 2333 3207 2347
rect 3113 2293 3127 2307
rect 3053 2233 3067 2247
rect 3093 2233 3107 2247
rect 3193 2233 3207 2247
rect 2953 2193 2967 2207
rect 2993 2153 3007 2167
rect 2873 2113 2887 2127
rect 2913 2113 2927 2127
rect 2853 2093 2867 2107
rect 2833 2013 2847 2027
rect 2773 1973 2787 1987
rect 2733 1953 2747 1967
rect 2807 1953 2821 1967
rect 2853 1993 2867 2007
rect 2833 1913 2847 1927
rect 2873 1913 2887 1927
rect 2793 1873 2807 1887
rect 2833 1873 2847 1887
rect 2773 1833 2787 1847
rect 2713 1753 2727 1767
rect 2693 1673 2707 1687
rect 2773 1713 2787 1727
rect 2853 1793 2867 1807
rect 2853 1694 2867 1708
rect 2793 1673 2807 1687
rect 2813 1593 2827 1607
rect 2733 1573 2747 1587
rect 2713 1553 2727 1567
rect 2473 1513 2487 1527
rect 2473 1473 2487 1487
rect 2493 1433 2507 1447
rect 2793 1433 2807 1447
rect 2853 1672 2867 1686
rect 2893 1893 2907 1907
rect 2933 2073 2947 2087
rect 2953 1953 2967 1967
rect 2873 1633 2887 1647
rect 2913 1753 2927 1767
rect 2953 1753 2967 1767
rect 2933 1693 2947 1707
rect 2893 1593 2907 1607
rect 2852 1573 2866 1587
rect 2874 1573 2888 1587
rect 2833 1473 2847 1487
rect 2653 1393 2667 1407
rect 2713 1393 2727 1407
rect 2733 1393 2747 1407
rect 2573 1373 2587 1387
rect 2593 1273 2607 1287
rect 2453 1253 2467 1267
rect 2373 1213 2387 1227
rect 2513 1213 2527 1227
rect 2353 1113 2367 1127
rect 2293 1073 2307 1087
rect 2493 1193 2507 1207
rect 2393 1173 2407 1187
rect 2813 1273 2827 1287
rect 2693 1213 2707 1227
rect 2613 1173 2627 1187
rect 2673 1173 2687 1187
rect 2713 1173 2727 1187
rect 2833 1213 2847 1227
rect 2753 1193 2767 1207
rect 2733 1133 2747 1147
rect 2633 993 2647 1007
rect 2593 973 2607 987
rect 2653 933 2667 947
rect 3053 2133 3067 2147
rect 3013 2013 3027 2027
rect 3013 1932 3027 1946
rect 3133 2193 3147 2207
rect 3373 2413 3387 2427
rect 3313 2293 3327 2307
rect 3273 2247 3287 2261
rect 3533 2513 3547 2527
rect 3633 2433 3647 2447
rect 3653 2433 3667 2447
rect 3713 2433 3727 2447
rect 3493 2273 3507 2287
rect 3533 2273 3547 2287
rect 3413 2253 3427 2267
rect 3553 2253 3567 2267
rect 3233 2133 3247 2147
rect 3153 2093 3167 2107
rect 3073 2073 3087 2087
rect 3133 2013 3147 2027
rect 3013 1892 3027 1906
rect 3073 1893 3087 1907
rect 3193 1933 3207 1947
rect 3473 2213 3487 2227
rect 3493 2213 3507 2227
rect 3373 2193 3387 2207
rect 3553 2193 3567 2207
rect 3633 2193 3647 2207
rect 3653 2173 3667 2187
rect 3613 2073 3627 2087
rect 3373 1973 3387 1987
rect 3493 1973 3507 1987
rect 3193 1873 3207 1887
rect 3273 1873 3287 1887
rect 3053 1853 3067 1867
rect 3132 1853 3146 1867
rect 3154 1853 3168 1867
rect 3033 1793 3047 1807
rect 3133 1753 3147 1767
rect 3093 1714 3107 1728
rect 3133 1713 3147 1727
rect 3073 1693 3087 1707
rect 2993 1653 3007 1667
rect 2973 1573 2987 1587
rect 3173 1693 3187 1707
rect 3133 1673 3147 1687
rect 3153 1653 3167 1667
rect 3073 1553 3087 1567
rect 2893 1433 2907 1447
rect 2873 1214 2887 1228
rect 2893 1194 2907 1208
rect 2847 1173 2861 1187
rect 2893 1172 2907 1186
rect 2793 1133 2807 1147
rect 2873 1053 2887 1067
rect 2873 993 2887 1007
rect 2153 893 2167 907
rect 2213 893 2227 907
rect 2413 913 2427 927
rect 2453 914 2467 928
rect 2533 913 2547 927
rect 2553 913 2567 927
rect 2453 892 2467 906
rect 2593 893 2607 907
rect 2173 813 2187 827
rect 2253 813 2267 827
rect 2153 753 2167 767
rect 2093 693 2107 707
rect 2113 693 2127 707
rect 2039 673 2053 687
rect 2253 733 2267 747
rect 2193 673 2207 687
rect 1993 653 2007 667
rect 1933 633 1947 647
rect 2013 633 2027 647
rect 2133 593 2147 607
rect 1913 473 1927 487
rect 2013 473 2027 487
rect 1853 433 1867 447
rect 1893 433 1907 447
rect 1693 413 1707 427
rect 1613 393 1627 407
rect 1673 393 1687 407
rect 1373 353 1387 367
rect 1693 373 1707 387
rect 1333 333 1347 347
rect 1553 333 1567 347
rect 1593 333 1607 347
rect 1253 253 1267 267
rect 1393 293 1407 307
rect 1233 153 1247 167
rect 1353 153 1367 167
rect 1113 134 1127 148
rect 1913 413 1927 427
rect 1773 393 1787 407
rect 1833 393 1847 407
rect 1733 293 1747 307
rect 1653 253 1667 267
rect 1713 253 1727 267
rect 1753 233 1767 247
rect 1793 233 1807 247
rect 1413 153 1427 167
rect 1513 153 1527 167
rect 1566 153 1567 167
rect 1567 153 1580 167
rect 673 113 687 127
rect 833 113 847 127
rect 1213 133 1227 147
rect 2573 853 2587 867
rect 2613 813 2627 827
rect 2473 713 2487 727
rect 2273 693 2287 707
rect 2373 693 2387 707
rect 2453 693 2467 707
rect 2253 653 2267 667
rect 2733 892 2747 906
rect 2653 773 2667 787
rect 2713 773 2727 787
rect 2393 653 2407 667
rect 2433 653 2447 667
rect 2573 673 2587 687
rect 2333 573 2347 587
rect 2693 653 2707 667
rect 2533 493 2547 507
rect 2613 493 2627 507
rect 2653 493 2667 507
rect 2273 473 2287 487
rect 2293 413 2307 427
rect 2493 413 2507 427
rect 1953 393 1967 407
rect 2193 393 2207 407
rect 2373 393 2387 407
rect 2093 373 2107 387
rect 2153 373 2167 387
rect 2633 413 2647 427
rect 2253 353 2267 367
rect 2372 353 2386 367
rect 2633 353 2647 367
rect 1953 293 1967 307
rect 2293 333 2307 347
rect 2393 333 2407 347
rect 2153 293 2167 307
rect 2113 233 2127 247
rect 2033 213 2047 227
rect 2073 213 2087 227
rect 2153 213 2167 227
rect 1893 173 1907 187
rect 1933 173 1947 187
rect 1813 153 1827 167
rect 1933 133 1947 147
rect 1953 133 1967 147
rect 993 113 1007 127
rect 1093 113 1107 127
rect 1113 112 1127 126
rect 1653 113 1667 127
rect 753 93 767 107
rect 953 93 967 107
rect 1253 93 1267 107
rect 393 73 407 87
rect 473 73 487 87
rect 553 73 567 87
rect 1173 73 1187 87
rect 2113 173 2127 187
rect 2093 133 2107 147
rect 2013 113 2027 127
rect 2173 173 2187 187
rect 2493 273 2507 287
rect 2453 233 2467 247
rect 2293 153 2307 167
rect 2253 133 2267 147
rect 2413 133 2427 147
rect 2113 93 2127 107
rect 2313 113 2327 127
rect 2433 93 2447 107
rect 2253 73 2267 87
rect 1993 53 2007 67
rect 2433 53 2447 67
rect 2533 213 2547 227
rect 2613 193 2627 207
rect 2713 453 2727 467
rect 2713 413 2727 427
rect 2753 853 2767 867
rect 2993 1493 3007 1507
rect 3113 1453 3127 1467
rect 3013 1353 3027 1367
rect 3013 1253 3027 1267
rect 2993 1053 3007 1067
rect 2973 973 2987 987
rect 2953 933 2967 947
rect 3033 1153 3047 1167
rect 3133 1153 3147 1167
rect 3313 1833 3327 1847
rect 3333 1773 3347 1787
rect 3593 1953 3607 1967
rect 3513 1933 3527 1947
rect 3813 2753 3827 2767
rect 3913 2953 3927 2967
rect 3853 2913 3867 2927
rect 3973 2933 3987 2947
rect 4093 2813 4107 2827
rect 3853 2773 3867 2787
rect 3913 2773 3927 2787
rect 3873 2733 3887 2747
rect 3833 2653 3847 2667
rect 3793 2513 3807 2527
rect 3753 2273 3767 2287
rect 3853 2433 3867 2447
rect 4153 2753 4167 2767
rect 4053 2633 4067 2647
rect 4153 2633 4167 2647
rect 3953 2513 3967 2527
rect 4073 2513 4087 2527
rect 3833 2413 3847 2427
rect 3933 2413 3947 2427
rect 4073 2413 4087 2427
rect 3993 2373 4007 2387
rect 3813 2313 3827 2327
rect 3993 2313 4007 2327
rect 3953 2273 3967 2287
rect 3873 2233 3887 2247
rect 3673 2053 3687 2067
rect 3693 1993 3707 2007
rect 3453 1913 3467 1927
rect 3533 1913 3547 1927
rect 3453 1873 3467 1887
rect 3553 1853 3567 1867
rect 3473 1753 3487 1767
rect 3373 1733 3387 1747
rect 3213 1673 3227 1687
rect 3273 1553 3287 1567
rect 3233 1453 3247 1467
rect 3153 1093 3167 1107
rect 3013 1033 3027 1047
rect 3153 1013 3167 1027
rect 3013 973 3027 987
rect 3033 913 3047 927
rect 3013 893 3027 907
rect 2893 874 2907 888
rect 2913 873 2927 887
rect 2993 873 3007 887
rect 2773 813 2787 827
rect 2833 793 2847 807
rect 2793 733 2807 747
rect 2753 713 2767 727
rect 2753 652 2767 666
rect 3033 793 3047 807
rect 3073 793 3087 807
rect 2953 693 2967 707
rect 3073 673 3087 687
rect 2833 653 2847 667
rect 2753 513 2767 527
rect 2893 453 2907 467
rect 2833 393 2847 407
rect 2693 373 2707 387
rect 2733 374 2747 388
rect 2793 353 2807 367
rect 2813 353 2827 367
rect 2733 313 2747 327
rect 3153 733 3167 747
rect 3233 1393 3247 1407
rect 3253 1393 3267 1407
rect 3333 1712 3347 1726
rect 3293 1493 3307 1507
rect 3333 1453 3347 1467
rect 3433 1713 3447 1727
rect 3453 1693 3467 1707
rect 3393 1434 3407 1448
rect 3313 1413 3327 1427
rect 3293 1353 3307 1367
rect 3273 933 3287 947
rect 3213 873 3227 887
rect 3093 573 3107 587
rect 3053 493 3067 507
rect 3073 453 3087 467
rect 2793 313 2807 327
rect 2993 354 3007 368
rect 3193 653 3207 667
rect 3393 1412 3407 1426
rect 3613 1933 3627 1947
rect 3573 1633 3587 1647
rect 3913 2193 3927 2207
rect 3893 2153 3907 2167
rect 3993 2053 4007 2067
rect 3953 2013 3967 2027
rect 3813 1973 3827 1987
rect 3913 1973 3927 1987
rect 4033 1973 4047 1987
rect 3773 1893 3787 1907
rect 3693 1773 3707 1787
rect 3773 1753 3787 1767
rect 3693 1693 3707 1707
rect 3753 1673 3767 1687
rect 3713 1633 3727 1647
rect 3673 1573 3687 1587
rect 3573 1513 3587 1527
rect 3473 1433 3487 1447
rect 3353 1373 3367 1387
rect 3493 1253 3507 1267
rect 3773 1413 3787 1427
rect 3673 1393 3687 1407
rect 3713 1393 3727 1407
rect 3533 1313 3547 1327
rect 3533 1273 3547 1287
rect 3693 1273 3707 1287
rect 3513 1233 3527 1247
rect 3433 1213 3447 1227
rect 3713 1253 3727 1267
rect 3553 1233 3567 1247
rect 3573 1213 3587 1227
rect 3453 1173 3467 1187
rect 3473 1173 3487 1187
rect 3353 1153 3367 1167
rect 3313 1053 3327 1067
rect 3373 1013 3387 1027
rect 3413 933 3427 947
rect 3313 913 3327 927
rect 3293 893 3307 907
rect 3373 893 3387 907
rect 3293 853 3307 867
rect 3393 793 3407 807
rect 3513 1093 3527 1107
rect 4173 2493 4187 2507
rect 4333 3273 4347 3287
rect 4433 3273 4447 3287
rect 4373 3253 4387 3267
rect 4713 4113 4727 4127
rect 4833 4033 4847 4047
rect 4893 4033 4907 4047
rect 4773 4013 4787 4027
rect 4713 3953 4727 3967
rect 4893 3973 4907 3987
rect 4793 3953 4807 3967
rect 4753 3853 4767 3867
rect 4933 4353 4947 4367
rect 4953 4333 4967 4347
rect 4973 4233 4987 4247
rect 4953 4073 4967 4087
rect 5067 4293 5081 4307
rect 5233 4353 5247 4367
rect 5173 4333 5187 4347
rect 5193 4313 5207 4327
rect 5213 4313 5227 4327
rect 5253 4313 5267 4327
rect 5133 4293 5147 4307
rect 5073 4273 5087 4287
rect 5113 4273 5127 4287
rect 5153 4273 5167 4287
rect 5033 4153 5047 4167
rect 5013 4133 5027 4147
rect 5073 4133 5087 4147
rect 5053 4073 5067 4087
rect 4953 4033 4967 4047
rect 4993 4033 5007 4047
rect 4933 3873 4947 3887
rect 4733 3813 4747 3827
rect 4793 3813 4807 3827
rect 4713 3773 4727 3787
rect 4753 3773 4767 3787
rect 4807 3773 4821 3787
rect 4853 3773 4867 3787
rect 4913 3773 4927 3787
rect 4833 3653 4847 3667
rect 4913 3633 4927 3647
rect 4833 3593 4847 3607
rect 4693 3473 4707 3487
rect 4773 3492 4787 3506
rect 4733 3453 4747 3467
rect 4653 3413 4667 3427
rect 4753 3393 4767 3407
rect 4633 3373 4647 3387
rect 4733 3373 4747 3387
rect 4613 3333 4627 3347
rect 4693 3333 4707 3347
rect 4533 3273 4547 3287
rect 4473 3254 4487 3268
rect 4473 3232 4487 3246
rect 4553 3233 4567 3247
rect 4453 3053 4467 3067
rect 4573 3133 4587 3147
rect 4653 3293 4667 3307
rect 4713 3293 4727 3307
rect 4673 3232 4687 3246
rect 4713 3233 4727 3247
rect 4613 3193 4627 3207
rect 4633 3133 4647 3147
rect 4593 3093 4607 3107
rect 4533 3053 4547 3067
rect 4573 3033 4587 3047
rect 4633 3033 4647 3047
rect 4439 3013 4453 3027
rect 4413 2994 4427 3008
rect 4473 2993 4487 3007
rect 4613 2993 4627 3007
rect 4293 2953 4307 2967
rect 4313 2833 4327 2847
rect 4593 2953 4607 2967
rect 4633 2953 4647 2967
rect 4373 2933 4387 2947
rect 4413 2933 4427 2947
rect 4393 2833 4407 2847
rect 4253 2793 4267 2807
rect 4333 2793 4347 2807
rect 4233 2752 4247 2766
rect 4273 2733 4287 2747
rect 4293 2653 4307 2667
rect 4313 2553 4327 2567
rect 4253 2493 4267 2507
rect 4293 2473 4307 2487
rect 4233 2453 4247 2467
rect 4273 2459 4287 2473
rect 4093 2233 4107 2247
rect 4213 2293 4227 2307
rect 4133 2212 4147 2226
rect 4193 2213 4207 2227
rect 4533 2813 4547 2827
rect 4413 2793 4427 2807
rect 4433 2773 4447 2787
rect 4393 2593 4407 2607
rect 4433 2513 4447 2527
rect 4473 2513 4487 2527
rect 4553 2733 4567 2747
rect 4553 2653 4567 2667
rect 4533 2494 4547 2508
rect 4613 2613 4627 2627
rect 4593 2573 4607 2587
rect 4493 2473 4507 2487
rect 4433 2433 4447 2447
rect 4353 2293 4367 2307
rect 4273 2213 4287 2227
rect 4233 2193 4247 2207
rect 4313 2173 4327 2187
rect 4093 2153 4107 2167
rect 4153 2013 4167 2027
rect 4253 2013 4267 2027
rect 4073 1953 4087 1967
rect 4093 1953 4107 1967
rect 4133 1953 4147 1967
rect 3833 1933 3847 1947
rect 4093 1913 4107 1927
rect 3873 1893 3887 1907
rect 3973 1813 3987 1827
rect 3833 1793 3847 1807
rect 3853 1773 3867 1787
rect 3833 1753 3847 1767
rect 4013 1773 4027 1787
rect 4333 1993 4347 2007
rect 4253 1973 4267 1987
rect 4313 1973 4327 1987
rect 4213 1913 4227 1927
rect 4153 1773 4167 1787
rect 3933 1733 3947 1747
rect 4053 1733 4067 1747
rect 3853 1693 3867 1707
rect 3813 1673 3827 1687
rect 3813 1613 3827 1627
rect 3833 1453 3847 1467
rect 3813 1413 3827 1427
rect 3833 1313 3847 1327
rect 4033 1693 4047 1707
rect 4053 1693 4067 1707
rect 4013 1573 4027 1587
rect 4053 1573 4067 1587
rect 3993 1513 4007 1527
rect 3953 1373 3967 1387
rect 3933 1293 3947 1307
rect 3793 1233 3807 1247
rect 3753 1073 3767 1087
rect 3633 1013 3647 1027
rect 3673 1013 3687 1027
rect 3713 1013 3727 1027
rect 3513 953 3527 967
rect 3633 933 3647 947
rect 3513 913 3527 927
rect 3273 733 3287 747
rect 3433 733 3447 747
rect 3413 713 3427 727
rect 3313 667 3327 681
rect 3353 653 3367 667
rect 3213 633 3227 647
rect 3293 633 3307 647
rect 3233 593 3247 607
rect 3193 553 3207 567
rect 3253 393 3267 407
rect 3113 353 3127 367
rect 3153 353 3167 367
rect 2993 332 3007 346
rect 3073 333 3087 347
rect 2813 293 2827 307
rect 2933 293 2947 307
rect 2773 193 2787 207
rect 3013 193 3027 207
rect 3213 253 3227 267
rect 3533 853 3547 867
rect 3533 793 3547 807
rect 3513 693 3527 707
rect 3453 673 3467 687
rect 3333 593 3347 607
rect 3372 593 3386 607
rect 3394 593 3408 607
rect 3333 453 3347 467
rect 3313 413 3327 427
rect 3713 893 3727 907
rect 3593 833 3607 847
rect 3633 793 3647 807
rect 3673 793 3687 807
rect 3713 733 3727 747
rect 3733 713 3747 727
rect 3933 1173 3947 1187
rect 3873 1113 3887 1127
rect 3853 1073 3867 1087
rect 3853 933 3867 947
rect 3773 713 3787 727
rect 3733 673 3747 687
rect 3773 633 3787 647
rect 3713 613 3727 627
rect 3673 593 3687 607
rect 3573 513 3587 527
rect 3493 493 3507 507
rect 3533 493 3547 507
rect 3633 493 3647 507
rect 3473 413 3487 427
rect 3393 373 3407 387
rect 3593 413 3607 427
rect 3793 413 3807 427
rect 3933 933 3947 947
rect 3973 1313 3987 1327
rect 3973 1233 3987 1247
rect 4033 1553 4047 1567
rect 4013 1333 4027 1347
rect 4033 1253 4047 1267
rect 4033 1213 4047 1227
rect 4013 1173 4027 1187
rect 3993 1113 4007 1127
rect 3973 927 3987 941
rect 3973 873 3987 887
rect 3873 793 3887 807
rect 3973 793 3987 807
rect 3893 733 3907 747
rect 3913 713 3927 727
rect 3893 693 3907 707
rect 3853 633 3867 647
rect 3893 613 3907 627
rect 4133 1673 4147 1687
rect 4073 1493 4087 1507
rect 4113 1493 4127 1507
rect 4093 1413 4107 1427
rect 4113 1373 4127 1387
rect 4100 1213 4113 1227
rect 4113 1213 4114 1227
rect 4233 1853 4247 1867
rect 4273 1793 4287 1807
rect 4253 1733 4267 1747
rect 4233 1633 4247 1647
rect 4213 1613 4227 1627
rect 4213 1513 4227 1527
rect 4293 1673 4307 1687
rect 4533 2472 4547 2486
rect 5033 4013 5047 4027
rect 4993 3933 5007 3947
rect 5013 3873 5027 3887
rect 4973 3673 4987 3687
rect 4953 3593 4967 3607
rect 4933 3553 4947 3567
rect 4993 3633 5007 3647
rect 5013 3613 5027 3627
rect 5113 4113 5127 4127
rect 5153 4013 5167 4027
rect 5173 3853 5187 3867
rect 5373 4393 5387 4407
rect 5313 4313 5327 4327
rect 5473 4773 5487 4787
rect 5473 4633 5487 4647
rect 5513 4633 5527 4647
rect 5533 4613 5547 4627
rect 5493 4533 5507 4547
rect 5493 4313 5507 4327
rect 5513 4313 5527 4327
rect 5346 4273 5347 4287
rect 5347 4273 5360 4287
rect 5453 4273 5467 4287
rect 5373 4253 5387 4267
rect 5413 4253 5427 4267
rect 5333 4233 5347 4247
rect 5313 4173 5327 4187
rect 5253 4153 5267 4167
rect 5273 4113 5287 4127
rect 5233 4013 5247 4027
rect 5413 4153 5427 4167
rect 5313 4033 5327 4047
rect 5273 4012 5287 4026
rect 5253 3973 5267 3987
rect 5253 3933 5267 3947
rect 5213 3813 5227 3827
rect 5113 3673 5127 3687
rect 5093 3613 5107 3627
rect 5013 3573 5027 3587
rect 5053 3573 5067 3587
rect 4993 3553 5007 3567
rect 4852 3473 4866 3487
rect 4874 3473 4888 3487
rect 4933 3473 4947 3487
rect 4793 3413 4807 3427
rect 4953 3453 4967 3467
rect 5053 3493 5067 3507
rect 5033 3473 5047 3487
rect 5053 3453 5067 3467
rect 5073 3433 5087 3447
rect 5053 3413 5067 3427
rect 5233 3713 5247 3727
rect 5173 3553 5187 3567
rect 5233 3533 5247 3547
rect 5133 3493 5147 3507
rect 5093 3393 5107 3407
rect 5133 3453 5147 3467
rect 5133 3413 5147 3427
rect 5033 3333 5047 3347
rect 5113 3333 5127 3347
rect 4893 3313 4907 3327
rect 4993 3313 5007 3327
rect 4853 3293 4867 3307
rect 4833 3253 4847 3267
rect 4853 3253 4867 3267
rect 4793 3233 4807 3247
rect 4773 3213 4787 3227
rect 4753 3113 4767 3127
rect 4793 3073 4807 3087
rect 4773 3053 4787 3067
rect 4733 3013 4747 3027
rect 4873 3033 4887 3047
rect 4793 3013 4807 3027
rect 4833 2973 4847 2987
rect 4833 2853 4847 2867
rect 4733 2773 4747 2787
rect 4793 2733 4807 2747
rect 4813 2733 4827 2747
rect 4713 2713 4727 2727
rect 4673 2573 4687 2587
rect 4633 2493 4647 2507
rect 4413 2253 4427 2267
rect 4473 2253 4487 2267
rect 4453 2233 4467 2247
rect 4413 2213 4427 2227
rect 4473 2073 4487 2087
rect 4373 2033 4387 2047
rect 4573 2373 4587 2387
rect 4533 2333 4547 2347
rect 4733 2653 4747 2667
rect 4753 2493 4767 2507
rect 4813 2493 4827 2507
rect 4913 3293 4927 3307
rect 5013 3293 5027 3307
rect 4933 3273 4947 3287
rect 4993 3273 5007 3287
rect 5133 3293 5147 3307
rect 5153 3293 5167 3307
rect 5193 3493 5207 3507
rect 5033 3253 5047 3267
rect 5113 3253 5127 3267
rect 5173 3213 5187 3227
rect 4973 3193 4987 3207
rect 5333 3913 5347 3927
rect 5313 3813 5327 3827
rect 5273 3794 5287 3808
rect 5293 3772 5307 3786
rect 5433 4053 5447 4067
rect 5453 3953 5467 3967
rect 5493 3913 5507 3927
rect 5393 3853 5407 3867
rect 5353 3813 5367 3827
rect 5433 3773 5447 3787
rect 5353 3553 5367 3567
rect 5333 3533 5347 3547
rect 5493 3813 5507 3827
rect 5493 3553 5507 3567
rect 5493 3513 5507 3527
rect 5313 3493 5327 3507
rect 5453 3493 5467 3507
rect 5273 3433 5287 3447
rect 5253 3373 5267 3387
rect 5233 3313 5247 3327
rect 5213 3234 5227 3248
rect 4993 3113 5007 3127
rect 5113 3113 5127 3127
rect 5193 3113 5207 3127
rect 4913 2993 4927 3007
rect 4893 2833 4907 2847
rect 4873 2733 4887 2747
rect 4873 2593 4887 2607
rect 4853 2573 4867 2587
rect 4833 2453 4847 2467
rect 4753 2434 4767 2448
rect 4713 2413 4727 2427
rect 4753 2412 4767 2426
rect 4733 2353 4747 2367
rect 4693 2333 4707 2347
rect 4713 2233 4727 2247
rect 4593 2213 4607 2227
rect 4653 2133 4667 2147
rect 4513 1993 4527 2007
rect 4593 1993 4607 2007
rect 4353 1973 4367 1987
rect 4353 1933 4367 1947
rect 4413 1913 4427 1927
rect 4493 1913 4507 1927
rect 4353 1713 4367 1727
rect 4333 1593 4347 1607
rect 4313 1573 4327 1587
rect 4293 1553 4307 1567
rect 4153 1473 4167 1487
rect 4253 1473 4267 1487
rect 4433 1893 4447 1907
rect 4453 1853 4467 1867
rect 4393 1733 4407 1747
rect 4533 1933 4547 1947
rect 4573 1893 4587 1907
rect 4513 1813 4527 1827
rect 4553 1713 4567 1727
rect 4533 1693 4547 1707
rect 4433 1673 4447 1687
rect 4413 1593 4427 1607
rect 4513 1593 4527 1607
rect 4513 1513 4527 1527
rect 4373 1433 4387 1447
rect 4473 1433 4487 1447
rect 4213 1393 4227 1407
rect 4153 1373 4167 1387
rect 4233 1333 4247 1347
rect 4153 1293 4167 1307
rect 4213 1273 4227 1287
rect 4073 1173 4087 1187
rect 4113 1173 4127 1187
rect 4073 973 4087 987
rect 4133 953 4147 967
rect 4093 913 4107 927
rect 4073 873 4087 887
rect 4193 1173 4207 1187
rect 4133 793 4147 807
rect 4053 733 4067 747
rect 4013 713 4027 727
rect 3993 673 4007 687
rect 4053 653 4067 667
rect 4073 654 4087 668
rect 3993 633 4007 647
rect 3853 533 3867 547
rect 3973 533 3987 547
rect 3647 373 3661 387
rect 3473 353 3487 367
rect 3773 353 3787 367
rect 3293 333 3307 347
rect 3393 332 3407 346
rect 3293 253 3307 267
rect 2813 173 2827 187
rect 2913 173 2927 187
rect 2953 173 2967 187
rect 3113 173 3127 187
rect 3153 173 3167 187
rect 3193 173 3207 187
rect 2639 153 2653 167
rect 2733 153 2747 167
rect 2533 133 2547 147
rect 2599 133 2613 147
rect 2473 73 2487 87
rect 2453 33 2467 47
rect 2993 113 3007 127
rect 2953 93 2967 107
rect 3253 213 3267 227
rect 3193 33 3207 47
rect 3713 333 3727 347
rect 3533 273 3547 287
rect 3513 153 3527 167
rect 3593 213 3607 227
rect 3733 213 3747 227
rect 3593 153 3607 167
rect 3653 153 3667 167
rect 4073 473 4087 487
rect 3933 413 3947 427
rect 3953 373 3967 387
rect 4133 633 4147 647
rect 4173 453 4187 467
rect 4213 1053 4227 1067
rect 4453 1393 4467 1407
rect 4293 1253 4307 1267
rect 4273 1173 4287 1187
rect 4253 1013 4267 1027
rect 4613 1933 4627 1947
rect 4713 2073 4727 2087
rect 4653 1873 4667 1887
rect 4673 1853 4687 1867
rect 4673 1813 4687 1827
rect 4773 2267 4787 2281
rect 4753 2173 4767 2187
rect 4773 2113 4787 2127
rect 4793 2073 4807 2087
rect 4773 2033 4787 2047
rect 4753 1973 4767 1987
rect 4773 1914 4787 1928
rect 4873 2433 4887 2447
rect 4873 2333 4887 2347
rect 5193 3073 5207 3087
rect 4993 2993 5007 3007
rect 5053 2993 5067 3007
rect 5373 3413 5387 3427
rect 5313 3293 5327 3307
rect 5253 3253 5267 3267
rect 5493 3373 5507 3387
rect 5433 3313 5447 3327
rect 5453 3293 5467 3307
rect 5233 3153 5247 3167
rect 5213 2993 5227 3007
rect 5113 2953 5127 2967
rect 5153 2953 5167 2967
rect 5133 2853 5147 2867
rect 4993 2833 5007 2847
rect 4973 2793 4987 2807
rect 5273 2793 5287 2807
rect 5013 2753 5027 2767
rect 4973 2733 4987 2747
rect 5033 2713 5047 2727
rect 5153 2753 5167 2767
rect 5073 2693 5087 2707
rect 4953 2613 4967 2627
rect 4933 2573 4947 2587
rect 5153 2573 5167 2587
rect 5033 2513 5047 2527
rect 4993 2433 5007 2447
rect 5133 2393 5147 2407
rect 5213 2693 5227 2707
rect 5193 2513 5207 2527
rect 5313 2993 5327 3007
rect 5393 3213 5407 3227
rect 5393 3173 5407 3187
rect 5313 2813 5327 2827
rect 5293 2653 5307 2667
rect 5233 2593 5247 2607
rect 5153 2353 5167 2367
rect 5033 2333 5047 2347
rect 5113 2333 5127 2347
rect 4913 2293 4927 2307
rect 4933 2233 4947 2247
rect 4873 2213 4887 2227
rect 4893 2213 4907 2227
rect 4953 2173 4967 2187
rect 4853 1993 4867 2007
rect 4933 1993 4947 2007
rect 4833 1973 4847 1987
rect 4833 1793 4847 1807
rect 4773 1753 4787 1767
rect 4712 1713 4726 1727
rect 4734 1714 4748 1728
rect 4593 1693 4607 1707
rect 4633 1673 4647 1687
rect 4633 1633 4647 1647
rect 4673 1653 4687 1667
rect 4593 1513 4607 1527
rect 4653 1513 4667 1527
rect 4553 1453 4567 1467
rect 4733 1673 4747 1687
rect 4773 1713 4787 1727
rect 4753 1653 4767 1667
rect 4693 1593 4707 1607
rect 4673 1493 4687 1507
rect 4613 1473 4627 1487
rect 4433 1233 4447 1247
rect 4533 1233 4547 1247
rect 4593 1233 4607 1247
rect 4453 1173 4467 1187
rect 4293 973 4307 987
rect 4573 1193 4587 1207
rect 4513 1173 4527 1187
rect 4493 1093 4507 1107
rect 4653 1433 4667 1447
rect 4713 1433 4727 1447
rect 4693 1373 4707 1387
rect 4753 1373 4767 1387
rect 4693 1333 4707 1347
rect 4693 1213 4707 1227
rect 4653 1194 4667 1208
rect 4973 2013 4987 2027
rect 5273 2533 5287 2547
rect 5353 2773 5367 2787
rect 5353 2693 5367 2707
rect 5373 2653 5387 2667
rect 5353 2593 5367 2607
rect 5353 2533 5367 2547
rect 5233 2313 5247 2327
rect 5073 2233 5087 2247
rect 5133 2233 5147 2247
rect 5193 2233 5207 2247
rect 5053 2113 5067 2127
rect 4993 1973 5007 1987
rect 5093 2013 5107 2027
rect 5013 1933 5027 1947
rect 4953 1893 4967 1907
rect 5013 1893 5027 1907
rect 4933 1753 4947 1767
rect 4853 1693 4867 1707
rect 4953 1693 4967 1707
rect 4993 1633 5007 1647
rect 5073 1853 5087 1867
rect 5053 1773 5067 1787
rect 5033 1753 5047 1767
rect 4873 1593 4887 1607
rect 5013 1593 5027 1607
rect 4873 1473 4887 1487
rect 5173 1973 5187 1987
rect 5153 1933 5167 1947
rect 5173 1932 5187 1946
rect 5333 2494 5347 2508
rect 5313 2473 5327 2487
rect 5413 3073 5427 3087
rect 5393 2613 5407 2627
rect 5453 2893 5467 2907
rect 5533 3813 5547 3827
rect 5533 3773 5547 3787
rect 5533 3693 5547 3707
rect 5533 3553 5547 3567
rect 5513 3173 5527 3187
rect 5533 3073 5547 3087
rect 5533 3033 5547 3047
rect 5513 2993 5527 3007
rect 5493 2813 5507 2827
rect 5433 2693 5447 2707
rect 5413 2573 5427 2587
rect 5413 2533 5427 2547
rect 5493 2693 5507 2707
rect 5453 2653 5467 2667
rect 5513 2613 5527 2627
rect 5433 2493 5447 2507
rect 5473 2493 5487 2507
rect 5433 2453 5447 2467
rect 5353 2393 5367 2407
rect 5333 2313 5347 2327
rect 5313 2293 5327 2307
rect 5253 2233 5267 2247
rect 5233 1913 5247 1927
rect 5093 1773 5107 1787
rect 5093 1733 5107 1747
rect 5213 1793 5227 1807
rect 5153 1713 5167 1727
rect 4933 1453 4947 1467
rect 5032 1453 5046 1467
rect 5054 1453 5068 1467
rect 4893 1433 4907 1447
rect 4793 1393 4807 1407
rect 4733 1173 4747 1187
rect 4613 1153 4627 1167
rect 4653 1152 4667 1166
rect 4573 1073 4587 1087
rect 4633 1033 4647 1047
rect 4233 933 4247 947
rect 4253 933 4267 947
rect 4333 933 4347 947
rect 4353 933 4367 947
rect 4493 933 4507 947
rect 4233 672 4247 686
rect 4353 873 4367 887
rect 4353 833 4367 847
rect 4433 813 4447 827
rect 4613 913 4627 927
rect 4913 1393 4927 1407
rect 4913 1273 4927 1287
rect 4773 1193 4787 1207
rect 4773 1093 4787 1107
rect 4693 953 4707 967
rect 4753 953 4767 967
rect 4593 873 4607 887
rect 4613 853 4627 867
rect 4453 773 4467 787
rect 4533 773 4547 787
rect 4433 733 4447 747
rect 4453 707 4467 721
rect 4533 693 4547 707
rect 4573 673 4587 687
rect 4353 573 4367 587
rect 4273 553 4287 567
rect 4213 513 4227 527
rect 4253 453 4267 467
rect 4113 413 4127 427
rect 4193 414 4207 428
rect 3853 273 3867 287
rect 4053 233 4067 247
rect 4133 233 4147 247
rect 3833 213 3847 227
rect 3773 173 3787 187
rect 3813 173 3827 187
rect 3673 113 3687 127
rect 3853 153 3867 167
rect 3933 153 3947 167
rect 4013 173 4027 187
rect 4193 373 4207 387
rect 4213 333 4227 347
rect 4173 153 4187 167
rect 3873 133 3887 147
rect 3913 133 3927 147
rect 3793 113 3807 127
rect 3813 113 3827 127
rect 4213 113 4227 127
rect 3773 93 3787 107
rect 4173 93 4187 107
rect 4333 413 4347 427
rect 4293 393 4307 407
rect 4553 473 4567 487
rect 4493 453 4507 467
rect 4533 453 4547 467
rect 4353 393 4367 407
rect 4413 393 4427 407
rect 4333 333 4347 347
rect 4453 333 4467 347
rect 4593 433 4607 447
rect 4673 813 4687 827
rect 4713 913 4727 927
rect 4733 913 4747 927
rect 4713 853 4727 867
rect 4793 953 4807 967
rect 4893 1193 4907 1207
rect 5013 1413 5027 1427
rect 5073 1413 5087 1427
rect 4953 1373 4967 1387
rect 5013 1253 5027 1267
rect 5153 1333 5167 1347
rect 5093 1313 5107 1327
rect 5033 1213 5047 1227
rect 4913 1113 4927 1127
rect 4913 1073 4927 1087
rect 4853 953 4867 967
rect 4953 953 4967 967
rect 4833 913 4847 927
rect 4833 873 4847 887
rect 4833 773 4847 787
rect 4773 733 4787 747
rect 4733 673 4747 687
rect 4773 674 4787 688
rect 4773 652 4787 666
rect 4813 653 4827 667
rect 4713 633 4727 647
rect 4573 293 4587 307
rect 4373 153 4387 167
rect 4413 153 4427 167
rect 4493 173 4507 187
rect 4533 153 4547 167
rect 4333 99 4347 113
rect 4313 73 4327 87
rect 4833 513 4847 527
rect 4833 473 4847 487
rect 4773 413 4787 427
rect 4813 413 4827 427
rect 5313 2073 5327 2087
rect 5413 2293 5427 2307
rect 5373 2233 5387 2247
rect 5393 2213 5407 2227
rect 5473 2213 5487 2227
rect 5353 2073 5367 2087
rect 5333 2013 5347 2027
rect 5333 1973 5347 1987
rect 5273 1793 5287 1807
rect 5233 1714 5247 1728
rect 5213 1453 5227 1467
rect 5273 1454 5287 1468
rect 5193 1434 5207 1448
rect 5213 1413 5227 1427
rect 5253 1393 5267 1407
rect 5133 1253 5147 1267
rect 5173 1253 5187 1267
rect 5093 1153 5107 1167
rect 5053 1033 5067 1047
rect 5113 993 5127 1007
rect 4973 913 4987 927
rect 5153 1233 5167 1247
rect 5193 1193 5207 1207
rect 5193 1153 5207 1167
rect 5313 1953 5327 1967
rect 5373 1993 5387 2007
rect 5453 1993 5467 2007
rect 5393 1973 5407 1987
rect 5413 1953 5427 1967
rect 5373 1912 5387 1926
rect 5393 1913 5407 1927
rect 5373 1873 5387 1887
rect 5353 1833 5367 1847
rect 5333 1813 5347 1827
rect 5313 1753 5327 1767
rect 5313 1453 5327 1467
rect 5413 1833 5427 1847
rect 5293 1313 5307 1327
rect 5273 1233 5287 1247
rect 5413 1394 5427 1408
rect 5413 1233 5427 1247
rect 5493 1233 5507 1247
rect 5393 1213 5407 1227
rect 5353 1193 5367 1207
rect 5413 1193 5427 1207
rect 5473 1193 5487 1207
rect 5173 1073 5187 1087
rect 5153 933 5167 947
rect 5253 1013 5267 1027
rect 5233 993 5247 1007
rect 5233 953 5247 967
rect 5373 1113 5387 1127
rect 5273 973 5287 987
rect 5313 973 5327 987
rect 5273 933 5287 947
rect 5113 894 5127 908
rect 5193 893 5207 907
rect 4893 873 4907 887
rect 4993 873 5007 887
rect 4933 793 4947 807
rect 4913 713 4927 727
rect 4893 633 4907 647
rect 4973 733 4987 747
rect 5013 853 5027 867
rect 4993 713 5007 727
rect 5013 673 5027 687
rect 4933 553 4947 567
rect 4973 513 4987 527
rect 4873 453 4887 467
rect 4953 453 4967 467
rect 4853 433 4867 447
rect 4853 373 4867 387
rect 4913 373 4927 387
rect 4713 333 4727 347
rect 4733 193 4747 207
rect 4773 193 4787 207
rect 4993 473 5007 487
rect 5333 933 5347 947
rect 5273 873 5287 887
rect 5313 873 5327 887
rect 5253 853 5267 867
rect 5173 793 5187 807
rect 5113 773 5127 787
rect 5213 713 5227 727
rect 5173 693 5187 707
rect 5013 413 5027 427
rect 5053 413 5067 427
rect 5033 373 5047 387
rect 5293 673 5307 687
rect 5213 433 5227 447
rect 5113 393 5127 407
rect 5173 393 5187 407
rect 5073 353 5087 367
rect 5133 333 5147 347
rect 4973 272 4987 286
rect 4953 233 4967 247
rect 4833 153 4847 167
rect 4919 153 4933 167
rect 4973 153 4987 167
rect 5013 153 5027 167
rect 5093 173 5107 187
rect 5253 393 5267 407
rect 5173 333 5187 347
rect 5153 293 5167 307
rect 5253 273 5267 287
rect 5213 233 5227 247
rect 5253 233 5267 247
rect 5193 193 5207 207
rect 4633 133 4647 147
rect 4873 93 4887 107
rect 4953 93 4967 107
rect 5193 93 5207 107
rect 5313 493 5327 507
rect 5293 153 5307 167
rect 5413 1013 5427 1027
rect 5473 1013 5487 1027
rect 5413 933 5427 947
rect 5393 793 5407 807
rect 5393 713 5407 727
rect 5373 674 5387 688
rect 5453 873 5467 887
rect 5393 553 5407 567
rect 5373 473 5387 487
rect 5333 433 5347 447
rect 5339 353 5353 367
rect 5333 313 5347 327
rect 5453 513 5467 527
rect 5433 433 5447 447
rect 5473 393 5487 407
rect 5393 233 5407 247
rect 5353 193 5367 207
rect 5413 153 5427 167
rect 5313 113 5327 127
rect 5353 113 5367 127
rect 4673 73 4687 87
rect 4913 73 4927 87
rect 5213 73 5227 87
rect 5533 313 5547 327
rect 4613 33 4627 47
rect 4673 33 4687 47
rect 5393 33 5407 47
rect 5493 33 5507 47
rect 4253 13 4267 27
rect 5433 13 5447 27
<< metal3 >>
rect 4267 5476 4313 5484
rect 2227 5456 2553 5464
rect 2607 5456 2893 5464
rect 3167 5456 3433 5464
rect 3487 5456 4344 5464
rect 407 5436 1073 5444
rect 2587 5436 2773 5444
rect 2787 5436 3453 5444
rect 4336 5444 4344 5456
rect 4427 5456 4473 5464
rect 4336 5436 4973 5444
rect 107 5416 253 5424
rect 3587 5416 3673 5424
rect 3687 5416 3913 5424
rect 4387 5416 4413 5424
rect 4707 5416 4792 5424
rect 4828 5416 4933 5424
rect 5447 5416 5493 5424
rect 2067 5396 2133 5404
rect 2867 5396 3093 5404
rect 3107 5396 3233 5404
rect 3367 5396 3413 5404
rect 3427 5396 4153 5404
rect 5267 5396 5353 5404
rect 5367 5396 5413 5404
rect 127 5376 193 5384
rect 207 5376 753 5384
rect 1647 5376 1733 5384
rect 2127 5376 2213 5384
rect 2367 5376 2433 5384
rect 2447 5376 2533 5384
rect 2547 5376 2793 5384
rect 4027 5376 4093 5384
rect 4367 5376 4573 5384
rect 4747 5376 4873 5384
rect 4947 5376 5073 5384
rect 607 5356 744 5364
rect 107 5336 233 5344
rect 247 5336 293 5344
rect 307 5336 373 5344
rect 527 5336 673 5344
rect 427 5316 633 5324
rect 736 5324 744 5356
rect 787 5356 813 5364
rect 1127 5356 1253 5364
rect 893 5344 907 5353
rect 2127 5356 2153 5364
rect 2607 5356 2733 5364
rect 3007 5356 3193 5364
rect 3207 5356 3613 5364
rect 3867 5356 4293 5364
rect 5233 5364 5247 5373
rect 4987 5360 5247 5364
rect 4987 5356 5244 5360
rect 5256 5356 5333 5364
rect 893 5340 933 5344
rect 896 5336 933 5340
rect 976 5336 1013 5344
rect 976 5324 984 5336
rect 1096 5336 1293 5344
rect 1096 5327 1104 5336
rect 1447 5336 1513 5344
rect 1527 5336 1639 5344
rect 1767 5336 1813 5344
rect 1827 5336 1913 5344
rect 2353 5344 2367 5352
rect 2353 5340 2433 5344
rect 2356 5336 2433 5340
rect 2447 5336 2493 5344
rect 3147 5333 3153 5347
rect 3361 5336 3413 5344
rect 3787 5336 3813 5344
rect 4547 5336 4733 5344
rect 4927 5336 5053 5344
rect 5256 5344 5264 5356
rect 5387 5356 5453 5364
rect 5076 5336 5264 5344
rect 736 5316 984 5324
rect 1067 5316 1093 5324
rect 1547 5316 1633 5324
rect 1887 5316 2033 5324
rect 2047 5316 2313 5324
rect 2327 5316 2393 5324
rect 2627 5316 2724 5324
rect 2716 5307 2724 5316
rect 3627 5316 3873 5324
rect 4047 5316 4133 5324
rect 4187 5316 4213 5324
rect 4787 5313 4793 5327
rect 5076 5324 5084 5336
rect 5307 5336 5353 5344
rect 5047 5316 5084 5324
rect 5407 5316 5473 5324
rect 267 5296 393 5304
rect 1007 5296 1113 5304
rect 1467 5296 1493 5304
rect 1507 5296 1673 5304
rect 2727 5296 2833 5304
rect 2893 5304 2907 5313
rect 2893 5300 2993 5304
rect 2896 5296 2993 5300
rect 3607 5296 3673 5304
rect 4367 5296 4533 5304
rect 187 5276 653 5284
rect 2027 5276 2153 5284
rect 2167 5276 2333 5284
rect 2467 5276 2533 5284
rect 2867 5276 2973 5284
rect 2987 5276 3073 5284
rect 3267 5276 3473 5284
rect 3487 5276 3553 5284
rect 3967 5276 5113 5284
rect 547 5256 733 5264
rect 2087 5256 2193 5264
rect 2207 5256 2653 5264
rect 2847 5256 3793 5264
rect 4267 5256 4433 5264
rect 4507 5256 4573 5264
rect 887 5236 1413 5244
rect 1427 5236 1533 5244
rect 1667 5236 2173 5244
rect 3087 5236 3213 5244
rect 3327 5236 3573 5244
rect 347 5216 413 5224
rect 427 5216 493 5224
rect 507 5216 913 5224
rect 2287 5216 2633 5224
rect 3107 5216 3213 5224
rect 3287 5216 3593 5224
rect 3787 5216 3953 5224
rect 4027 5216 4073 5224
rect 807 5196 1233 5204
rect 1247 5196 2993 5204
rect 3767 5196 4173 5204
rect 4227 5196 4273 5204
rect 687 5176 1393 5184
rect 1407 5176 1533 5184
rect 1687 5176 2513 5184
rect 2607 5176 3233 5184
rect 3567 5176 3713 5184
rect 3907 5176 3993 5184
rect 4007 5176 4093 5184
rect 4587 5176 4773 5184
rect 307 5156 613 5164
rect 2127 5156 2493 5164
rect 2627 5156 3173 5164
rect 3647 5156 3773 5164
rect 4287 5156 4493 5164
rect 5107 5156 5333 5164
rect 47 5136 93 5144
rect 407 5136 473 5144
rect 747 5136 833 5144
rect 1087 5136 1553 5144
rect 2187 5136 2653 5144
rect 3107 5136 3293 5144
rect 3807 5136 3873 5144
rect 3987 5136 4284 5144
rect 727 5116 764 5124
rect 756 5107 764 5116
rect 887 5116 913 5124
rect 1187 5116 1239 5124
rect 2367 5116 2413 5124
rect 2767 5116 2813 5124
rect 3407 5116 3513 5124
rect 3527 5116 3813 5124
rect 3827 5116 4113 5124
rect 4127 5116 4193 5124
rect 4276 5127 4284 5136
rect 4847 5136 5233 5144
rect 5247 5136 5293 5144
rect 4276 5116 4293 5127
rect 4280 5113 4293 5116
rect 4307 5116 4433 5124
rect 4447 5116 4533 5124
rect 4847 5116 5073 5124
rect 5127 5116 5213 5124
rect 5227 5116 5333 5124
rect 67 5096 333 5104
rect 756 5096 773 5107
rect 760 5093 773 5096
rect 787 5096 953 5104
rect 1007 5096 1033 5104
rect 1727 5096 1833 5104
rect 2127 5096 2233 5104
rect 2487 5096 2553 5104
rect 3056 5100 3113 5104
rect 121 5076 233 5084
rect 481 5076 493 5084
rect 1453 5084 1467 5093
rect 1247 5076 1304 5084
rect 1453 5080 1593 5084
rect 1456 5076 1593 5080
rect 587 5056 653 5064
rect 113 5044 127 5053
rect 1007 5056 1073 5064
rect 1296 5064 1304 5076
rect 1607 5076 1633 5084
rect 1867 5076 1913 5084
rect 1927 5076 2073 5084
rect 2407 5076 2453 5084
rect 2607 5076 2733 5084
rect 2747 5073 2753 5087
rect 2767 5076 2893 5084
rect 2953 5084 2967 5093
rect 3053 5096 3113 5100
rect 3053 5088 3067 5096
rect 3767 5096 3893 5104
rect 4407 5100 4504 5104
rect 4407 5096 4507 5100
rect 2953 5080 3053 5084
rect 2956 5076 3053 5080
rect 4493 5087 4507 5096
rect 4607 5096 4753 5104
rect 4887 5096 4993 5104
rect 3467 5076 3499 5084
rect 3896 5076 3973 5084
rect 1296 5056 1313 5064
rect 1327 5053 1333 5067
rect 1547 5056 1673 5064
rect 2127 5056 2233 5064
rect 2247 5056 2293 5064
rect 2507 5056 2573 5064
rect 2627 5056 2673 5064
rect 2947 5056 3093 5064
rect 3727 5056 3752 5064
rect 3896 5064 3904 5076
rect 4027 5073 4033 5087
rect 4567 5080 4644 5084
rect 4567 5076 4647 5080
rect 4633 5067 4647 5076
rect 4896 5076 5193 5084
rect 3788 5056 3904 5064
rect 3927 5056 4013 5064
rect 4896 5064 4904 5076
rect 5207 5076 5313 5084
rect 5387 5076 5433 5084
rect 4867 5056 4904 5064
rect 5196 5060 5293 5064
rect 5193 5056 5293 5060
rect 5193 5047 5207 5056
rect 113 5040 213 5044
rect 116 5036 213 5040
rect 227 5036 313 5044
rect 407 5033 413 5047
rect 427 5036 533 5044
rect 687 5036 853 5044
rect 1227 5036 1273 5044
rect 1827 5033 1833 5047
rect 2807 5036 3224 5044
rect 3416 5040 3533 5044
rect 707 5016 753 5024
rect 907 5016 964 5024
rect 467 4996 713 5004
rect 956 5004 964 5016
rect 1047 5016 1133 5024
rect 1793 5024 1807 5033
rect 1296 5016 2293 5024
rect 956 4996 993 5004
rect 1296 5004 1304 5016
rect 2347 5016 2473 5024
rect 2607 5016 2813 5024
rect 2827 5016 2892 5024
rect 2928 5016 3013 5024
rect 3067 5016 3173 5024
rect 3216 5024 3224 5036
rect 3413 5036 3533 5040
rect 3413 5027 3427 5036
rect 4507 5036 4673 5044
rect 4687 5036 4713 5044
rect 4947 5036 4993 5044
rect 3216 5016 3293 5024
rect 3647 5016 3793 5024
rect 4047 5016 4213 5024
rect 4627 5016 4693 5024
rect 1267 4996 1304 5004
rect 1707 4996 1873 5004
rect 1887 4996 1953 5004
rect 3727 4996 3853 5004
rect 4027 4996 4233 5004
rect 4247 4996 4393 5004
rect 5187 4996 5513 5004
rect 947 4976 1013 4984
rect 1067 4976 1193 4984
rect 1647 4976 1693 4984
rect 2287 4976 2433 4984
rect 2447 4976 2693 4984
rect 3067 4976 4413 4984
rect 4767 4976 5164 4984
rect 1487 4956 1593 4964
rect 1607 4956 2253 4964
rect 2387 4956 2533 4964
rect 2967 4956 3033 4964
rect 3187 4956 3733 4964
rect 3867 4956 3933 4964
rect 3987 4956 4193 4964
rect 4207 4956 4293 4964
rect 5156 4964 5164 4976
rect 5156 4956 5433 4964
rect 787 4936 1293 4944
rect 1307 4936 1513 4944
rect 1527 4936 1633 4944
rect 2007 4936 2033 4944
rect 2787 4936 2913 4944
rect 3067 4936 3113 4944
rect 3507 4936 3673 4944
rect 3687 4936 3893 4944
rect 4907 4936 4973 4944
rect 347 4916 513 4924
rect 827 4916 913 4924
rect 1127 4916 3013 4924
rect 3527 4916 3653 4924
rect 4247 4916 4513 4924
rect 4527 4916 4573 4924
rect 1247 4896 1313 4904
rect 1387 4896 1453 4904
rect 1507 4896 1573 4904
rect 1587 4896 1613 4904
rect 1987 4896 2053 4904
rect 2067 4896 2173 4904
rect 2467 4896 2573 4904
rect 3047 4896 3073 4904
rect 3127 4896 3153 4904
rect 3667 4896 3693 4904
rect 3967 4896 4033 4904
rect 4627 4896 5333 4904
rect 5347 4896 5493 4904
rect 907 4876 1013 4884
rect 1027 4876 1073 4884
rect 1127 4876 1373 4884
rect 1387 4876 2964 4884
rect 107 4856 113 4864
rect 2956 4867 2964 4876
rect 3147 4884 3160 4887
rect 3147 4873 3164 4884
rect 127 4864 140 4867
rect 127 4856 144 4864
rect 127 4854 140 4856
rect 120 4853 140 4854
rect 207 4856 233 4864
rect 1347 4856 1393 4864
rect 1467 4856 1593 4864
rect 1967 4856 2033 4864
rect 2047 4856 2393 4864
rect 2627 4860 2724 4864
rect 2627 4856 2727 4860
rect 127 4836 173 4844
rect 307 4836 353 4844
rect 607 4836 653 4844
rect 667 4836 833 4844
rect 961 4836 973 4844
rect 2713 4847 2727 4856
rect 2867 4856 2893 4864
rect 2916 4860 2953 4864
rect 2913 4856 2953 4860
rect 1087 4836 1113 4844
rect 1227 4836 1273 4844
rect 1787 4836 1813 4844
rect 2236 4840 2333 4844
rect 2233 4836 2333 4840
rect 2233 4827 2247 4836
rect 2913 4847 2927 4856
rect 3156 4864 3164 4873
rect 4707 4876 4793 4884
rect 3156 4856 3273 4864
rect 3287 4856 3493 4864
rect 3847 4856 3893 4864
rect 4053 4864 4067 4873
rect 3907 4860 4067 4864
rect 3907 4856 4064 4860
rect 4407 4856 4553 4864
rect 4567 4856 4593 4864
rect 4987 4856 5173 4864
rect 3460 4844 3473 4847
rect 3087 4836 3213 4844
rect 3456 4836 3473 4844
rect 427 4816 453 4824
rect 747 4816 813 4824
rect 1184 4816 1233 4824
rect 1184 4813 1193 4816
rect 1327 4816 1393 4824
rect 1187 4799 1193 4813
rect 1447 4816 1479 4824
rect 1687 4816 1733 4824
rect 1867 4816 1893 4824
rect 2473 4824 2487 4833
rect 2473 4820 2553 4824
rect 2476 4816 2553 4820
rect 2567 4816 2593 4824
rect 2607 4816 2733 4824
rect 2887 4816 2933 4824
rect 3027 4816 3073 4824
rect 3205 4819 3213 4836
rect 3460 4833 3473 4836
rect 3487 4836 3613 4844
rect 3627 4836 3733 4844
rect 3987 4836 4233 4844
rect 4467 4836 4573 4844
rect 5267 4833 5273 4847
rect 5487 4836 5513 4844
rect 3367 4816 3573 4824
rect 4287 4816 4313 4824
rect 4327 4816 4393 4824
rect 4947 4816 5053 4824
rect 5067 4816 5193 4824
rect 2227 4796 2273 4804
rect 2861 4796 2993 4804
rect 3147 4796 3253 4804
rect 3387 4796 3493 4804
rect 3507 4796 3633 4804
rect 3687 4796 3793 4804
rect 3921 4796 4173 4804
rect 4433 4804 4447 4813
rect 4307 4800 4447 4804
rect 4307 4796 4444 4800
rect 167 4776 753 4784
rect 907 4776 1133 4784
rect 1147 4776 1333 4784
rect 1927 4776 1993 4784
rect 2247 4776 2473 4784
rect 3587 4776 3853 4784
rect 4827 4776 5073 4784
rect 5387 4776 5433 4784
rect 5447 4776 5473 4784
rect 787 4756 853 4764
rect 1407 4756 1813 4764
rect 2236 4764 2244 4773
rect 2167 4756 2244 4764
rect 2947 4756 3033 4764
rect 3327 4756 3373 4764
rect 3887 4756 4033 4764
rect 4247 4756 4693 4764
rect 327 4736 893 4744
rect 1007 4736 1153 4744
rect 2687 4736 2804 4744
rect 427 4716 913 4724
rect 1107 4716 1493 4724
rect 1707 4716 2353 4724
rect 2407 4716 2573 4724
rect 2587 4716 2773 4724
rect 2796 4724 2804 4736
rect 3747 4736 3953 4744
rect 4367 4736 4493 4744
rect 4507 4736 4653 4744
rect 2796 4716 3353 4724
rect 3687 4716 4813 4724
rect 1207 4696 1344 4704
rect 187 4676 793 4684
rect 947 4676 1173 4684
rect 1336 4684 1344 4696
rect 1716 4696 1813 4704
rect 1716 4684 1724 4696
rect 3107 4696 3233 4704
rect 3247 4696 3413 4704
rect 3587 4696 3933 4704
rect 3947 4696 4133 4704
rect 4647 4696 4893 4704
rect 1336 4676 1724 4684
rect 2387 4676 2553 4684
rect 2927 4676 3133 4684
rect 3307 4676 3673 4684
rect 4247 4676 4773 4684
rect 527 4656 1073 4664
rect 1847 4656 2093 4664
rect 2107 4656 2313 4664
rect 2807 4656 3253 4664
rect 3427 4656 3693 4664
rect 3707 4656 3733 4664
rect 3847 4656 4153 4664
rect 4776 4664 4784 4673
rect 4776 4656 4913 4664
rect 4927 4656 4993 4664
rect 707 4636 953 4644
rect 1247 4636 1324 4644
rect 1316 4627 1324 4636
rect 1427 4636 1553 4644
rect 1827 4636 2033 4644
rect 2047 4636 2533 4644
rect 3027 4636 3153 4644
rect 3387 4636 4473 4644
rect 5487 4636 5513 4644
rect 227 4616 473 4624
rect 1327 4616 1713 4624
rect 1987 4616 2013 4624
rect 2607 4616 2693 4624
rect 2787 4616 2913 4624
rect 4727 4616 5533 4624
rect 607 4596 713 4604
rect 1207 4596 1273 4604
rect 1287 4596 1353 4604
rect 1487 4596 1533 4604
rect 1547 4596 1593 4604
rect 1607 4596 1773 4604
rect 1867 4596 2293 4604
rect 2447 4596 2733 4604
rect 3627 4596 3773 4604
rect 3927 4596 3993 4604
rect 167 4576 253 4584
rect 267 4576 353 4584
rect 933 4584 947 4593
rect 867 4580 947 4584
rect 867 4576 944 4580
rect 1627 4576 1653 4584
rect 2827 4576 2873 4584
rect 2987 4576 3213 4584
rect 3467 4576 3624 4584
rect 207 4556 233 4564
rect 667 4553 673 4567
rect 813 4564 827 4573
rect 813 4560 893 4564
rect 816 4556 893 4560
rect 907 4564 920 4567
rect 907 4553 924 4564
rect 1616 4564 1624 4573
rect 1447 4556 1624 4564
rect 1716 4556 1833 4564
rect 87 4536 173 4544
rect 916 4544 924 4553
rect 916 4536 1044 4544
rect 347 4516 433 4524
rect 647 4516 673 4524
rect 1036 4524 1044 4536
rect 1087 4536 1133 4544
rect 1227 4536 1293 4544
rect 1507 4536 1553 4544
rect 1716 4527 1724 4556
rect 1887 4553 1893 4567
rect 2167 4556 2213 4564
rect 2327 4556 2373 4564
rect 2487 4556 2573 4564
rect 2587 4554 2593 4567
rect 2580 4553 2593 4554
rect 2647 4556 2773 4564
rect 3267 4556 3433 4564
rect 2447 4536 2553 4544
rect 2847 4536 2973 4544
rect 2987 4536 3033 4544
rect 3207 4536 3233 4544
rect 3487 4536 3573 4544
rect 3616 4546 3624 4576
rect 4687 4576 4733 4584
rect 4947 4576 5013 4584
rect 5266 4573 5267 4580
rect 5288 4576 5333 4584
rect 3896 4547 3904 4573
rect 4367 4556 4417 4564
rect 4407 4553 4417 4556
rect 4581 4556 4673 4564
rect 3667 4536 3713 4544
rect 4227 4540 4324 4544
rect 4227 4536 4327 4540
rect 4407 4539 4413 4553
rect 5253 4564 5267 4573
rect 5167 4556 5224 4564
rect 5253 4560 5393 4564
rect 5255 4556 5393 4560
rect 5216 4547 5224 4556
rect 1036 4516 1613 4524
rect 1867 4516 1973 4524
rect 2247 4516 2333 4524
rect 2627 4516 2753 4524
rect 3827 4516 3913 4524
rect 3967 4516 4093 4524
rect 4107 4516 4173 4524
rect 4313 4527 4327 4536
rect 4487 4536 4553 4544
rect 4567 4536 4693 4544
rect 5227 4536 5493 4544
rect 4327 4516 4393 4524
rect 4767 4516 4913 4524
rect 4980 4524 4993 4527
rect 4976 4516 4993 4524
rect 4980 4513 4993 4516
rect 5007 4516 5073 4524
rect 5127 4516 5173 4524
rect 207 4496 313 4504
rect 1027 4496 1733 4504
rect 1807 4496 1953 4504
rect 2356 4496 2453 4504
rect 727 4476 913 4484
rect 1067 4476 1153 4484
rect 1167 4476 1393 4484
rect 1407 4476 2253 4484
rect 2356 4484 2364 4496
rect 3627 4496 3773 4504
rect 4187 4496 4513 4504
rect 2307 4476 2364 4484
rect 2847 4476 2913 4484
rect 3067 4476 3353 4484
rect 3467 4476 3593 4484
rect 3607 4476 3633 4484
rect 3807 4476 4052 4484
rect 4088 4476 4273 4484
rect 4516 4484 4524 4493
rect 4516 4476 4793 4484
rect 1547 4456 1753 4464
rect 2427 4456 3373 4464
rect 3707 4456 3993 4464
rect 1536 4444 1544 4453
rect 1107 4436 1544 4444
rect 2487 4436 3273 4444
rect 3567 4436 3593 4444
rect 3667 4436 3873 4444
rect 4067 4436 4233 4444
rect 707 4416 873 4424
rect 1007 4416 1133 4424
rect 1467 4416 1873 4424
rect 2067 4416 2133 4424
rect 2147 4416 2193 4424
rect 2447 4416 2613 4424
rect 2867 4416 2933 4424
rect 3367 4416 3713 4424
rect 3727 4416 3973 4424
rect 4467 4416 4653 4424
rect 1027 4396 1093 4404
rect 1187 4396 1713 4404
rect 1907 4396 2413 4404
rect 3087 4396 3333 4404
rect 3427 4396 3533 4404
rect 3547 4396 3693 4404
rect 3827 4396 4172 4404
rect 4208 4396 4233 4404
rect 4307 4396 4813 4404
rect 4827 4396 4873 4404
rect 4887 4396 5373 4404
rect 327 4376 373 4384
rect 447 4376 473 4384
rect 987 4376 1153 4384
rect 1307 4376 1373 4384
rect 1427 4376 1533 4384
rect 1987 4376 2113 4384
rect 2467 4376 2813 4384
rect 2827 4376 3013 4384
rect 3367 4376 3793 4384
rect 3847 4376 3913 4384
rect 4047 4376 4113 4384
rect 4507 4376 4553 4384
rect 107 4356 353 4364
rect 367 4356 473 4364
rect 1367 4356 1413 4364
rect 853 4344 867 4354
rect 1947 4356 2013 4364
rect 2267 4356 3053 4364
rect 3167 4356 3333 4364
rect 3427 4356 4253 4364
rect 4947 4356 5233 4364
rect 853 4340 893 4344
rect 856 4336 893 4340
rect 1047 4336 1893 4344
rect 2307 4336 2353 4344
rect 2607 4336 2633 4344
rect 3027 4336 3093 4344
rect 3336 4344 3344 4353
rect 3336 4336 3433 4344
rect 3496 4336 3673 4344
rect 147 4320 224 4324
rect 147 4316 227 4320
rect 213 4307 227 4316
rect 967 4314 973 4327
rect 967 4313 980 4314
rect 2107 4316 2272 4324
rect 2308 4316 2553 4324
rect 2707 4316 2913 4324
rect 3107 4316 3193 4324
rect 3496 4324 3504 4336
rect 3687 4336 3793 4344
rect 4096 4340 4153 4344
rect 4093 4336 4153 4340
rect 4093 4327 4107 4336
rect 4407 4336 4473 4344
rect 4487 4336 4593 4344
rect 4967 4336 5173 4344
rect 3476 4316 3504 4324
rect 367 4296 432 4304
rect 468 4296 553 4304
rect 727 4296 853 4304
rect 867 4296 1012 4304
rect 767 4276 793 4284
rect 973 4286 987 4296
rect 1033 4294 1034 4300
rect 1033 4287 1047 4294
rect 1107 4296 1273 4304
rect 1707 4296 1853 4304
rect 1867 4294 1873 4307
rect 1860 4293 1873 4294
rect 2147 4296 2193 4304
rect 2427 4296 2513 4304
rect 2687 4300 2744 4304
rect 2687 4296 2747 4300
rect 2733 4287 2747 4296
rect 2887 4296 3013 4304
rect 3476 4304 3484 4316
rect 3887 4316 4013 4324
rect 4767 4316 4833 4324
rect 4893 4324 4907 4333
rect 4847 4320 4907 4324
rect 4847 4316 4904 4320
rect 5207 4313 5213 4327
rect 5267 4316 5313 4324
rect 5507 4313 5513 4327
rect 3407 4296 3484 4304
rect 3527 4296 3553 4304
rect 3647 4296 3933 4304
rect 4007 4296 4053 4304
rect 5081 4296 5133 4304
rect 1020 4286 1047 4287
rect 1027 4280 1047 4286
rect 1027 4276 1044 4280
rect 1027 4273 1040 4276
rect 1227 4276 1513 4284
rect 2087 4276 2173 4284
rect 2867 4276 3133 4284
rect 3147 4276 3173 4284
rect 3507 4276 3613 4284
rect 3687 4276 3833 4284
rect 4207 4276 4253 4284
rect 4487 4276 4513 4284
rect 4527 4276 4633 4284
rect 5087 4276 5113 4284
rect 5127 4276 5153 4284
rect 5360 4276 5453 4284
rect 647 4256 1373 4264
rect 1927 4260 2104 4264
rect 1927 4256 2107 4260
rect 2093 4247 2107 4256
rect 2907 4256 2972 4264
rect 3008 4256 3513 4264
rect 3707 4256 3733 4264
rect 3927 4256 4073 4264
rect 5387 4256 5413 4264
rect 1967 4236 2013 4244
rect 2147 4236 2313 4244
rect 2707 4236 2853 4244
rect 3467 4236 3553 4244
rect 3627 4236 3833 4244
rect 4987 4236 5333 4244
rect 627 4216 693 4224
rect 1567 4216 2373 4224
rect 2387 4216 2473 4224
rect 3336 4216 3633 4224
rect 3336 4207 3344 4216
rect 3856 4216 3913 4224
rect 1807 4196 2132 4204
rect 2168 4196 2293 4204
rect 2787 4196 3033 4204
rect 3047 4196 3093 4204
rect 3107 4196 3332 4204
rect 3856 4204 3864 4216
rect 3368 4196 3864 4204
rect 4287 4196 4433 4204
rect 4447 4196 4473 4204
rect 487 4176 713 4184
rect 1047 4176 1173 4184
rect 1367 4176 1553 4184
rect 1607 4176 2433 4184
rect 2447 4176 2493 4184
rect 2507 4176 3873 4184
rect 4707 4176 5313 4184
rect 907 4156 1693 4164
rect 1787 4156 2053 4164
rect 2067 4156 2093 4164
rect 2287 4156 2773 4164
rect 2887 4156 3353 4164
rect 3587 4156 4153 4164
rect 4547 4156 5033 4164
rect 5267 4156 5413 4164
rect 1087 4136 1193 4144
rect 1207 4136 1284 4144
rect 447 4116 753 4124
rect 1276 4124 1284 4136
rect 1367 4136 2793 4144
rect 3287 4136 3493 4144
rect 3567 4136 3713 4144
rect 3867 4136 4013 4144
rect 5027 4136 5073 4144
rect 1276 4116 1333 4124
rect 1347 4116 1853 4124
rect 1867 4116 1893 4124
rect 2107 4116 3193 4124
rect 3207 4116 3613 4124
rect 4727 4116 5113 4124
rect 5127 4116 5273 4124
rect 547 4096 733 4104
rect 1067 4096 1253 4104
rect 1427 4096 1453 4104
rect 1507 4096 1633 4104
rect 2187 4096 2273 4104
rect 2427 4096 2453 4104
rect 2467 4096 2873 4104
rect 3467 4096 3533 4104
rect 3687 4096 3753 4104
rect 4067 4096 4453 4104
rect 4467 4096 4593 4104
rect 136 4076 193 4084
rect 136 4067 144 4076
rect 207 4076 273 4084
rect 327 4076 513 4084
rect 567 4076 687 4084
rect 1307 4076 1353 4084
rect 127 4056 144 4067
rect 127 4053 140 4056
rect 316 4064 324 4073
rect 247 4056 324 4064
rect 853 4064 867 4073
rect 1467 4076 1513 4084
rect 2087 4076 2184 4084
rect 787 4060 867 4064
rect 787 4056 864 4060
rect 1607 4056 1733 4064
rect 1947 4056 1973 4064
rect 187 4036 393 4044
rect 487 4036 653 4044
rect 667 4033 673 4047
rect 1127 4033 1133 4047
rect 1213 4044 1227 4053
rect 2087 4056 2153 4064
rect 2176 4064 2184 4076
rect 3207 4076 3693 4084
rect 4967 4076 5053 4084
rect 2176 4056 2224 4064
rect 1147 4040 1227 4044
rect 1147 4036 1224 4040
rect 2216 4047 2224 4056
rect 2807 4056 3013 4064
rect 3067 4056 3113 4064
rect 1487 4036 1553 4044
rect 1807 4036 1953 4044
rect 2216 4036 2233 4047
rect 2220 4033 2233 4036
rect 2527 4036 2593 4044
rect 2607 4036 2773 4044
rect 3927 4056 3953 4064
rect 4013 4064 4027 4073
rect 4013 4060 4173 4064
rect 4016 4056 4173 4060
rect 4227 4056 4353 4064
rect 3178 4044 3187 4047
rect 2867 4036 2944 4044
rect 3178 4036 3293 4044
rect 747 4013 753 4027
rect 776 4016 913 4024
rect 67 3996 133 4004
rect 776 4004 784 4016
rect 1187 4016 1233 4024
rect 1287 4016 1373 4024
rect 1727 4016 1853 4024
rect 1947 4016 2033 4024
rect 2207 4016 2293 4024
rect 2467 4016 2493 4024
rect 2587 4016 2613 4024
rect 2936 4027 2944 4036
rect 3447 4036 3473 4044
rect 3547 4036 3593 4044
rect 3647 4036 3713 4044
rect 4247 4036 4293 4044
rect 4487 4036 4593 4044
rect 4847 4036 4893 4044
rect 4967 4036 4993 4044
rect 5433 4044 5447 4053
rect 5327 4040 5447 4044
rect 5327 4036 5444 4040
rect 2827 4016 2853 4024
rect 2947 4016 3073 4024
rect 3627 4016 3773 4024
rect 4607 4016 4773 4024
rect 4787 4016 5033 4024
rect 5047 4016 5153 4024
rect 5247 4016 5273 4024
rect 607 3996 784 4004
rect 1747 3996 1813 4004
rect 2347 3996 2533 4004
rect 2547 4004 2560 4007
rect 2547 3996 2564 4004
rect 2547 3993 2560 3996
rect 2967 4000 3044 4004
rect 2967 3996 3047 4000
rect 3033 3987 3047 3996
rect 3227 3996 3333 4004
rect 3387 3996 3893 4004
rect 4207 3996 4313 4004
rect 167 3976 213 3984
rect 927 3976 1073 3984
rect 1387 3976 1473 3984
rect 2007 3976 2093 3984
rect 2647 3976 2733 3984
rect 3087 3976 3193 3984
rect 3367 3976 3433 3984
rect 3567 3976 3913 3984
rect 4087 3976 4173 3984
rect 4447 3976 4893 3984
rect 4907 3976 5253 3984
rect 1147 3956 1233 3964
rect 1327 3956 1453 3964
rect 1627 3956 2393 3964
rect 2487 3956 2773 3964
rect 2787 3956 2993 3964
rect 3127 3956 3253 3964
rect 3307 3956 3564 3964
rect 627 3936 913 3944
rect 1127 3936 1253 3944
rect 1487 3936 1813 3944
rect 2227 3936 2573 3944
rect 2596 3936 2652 3944
rect 1027 3916 1073 3924
rect 1087 3916 1633 3924
rect 1867 3916 1973 3924
rect 1987 3916 2253 3924
rect 2596 3924 2604 3936
rect 2688 3936 2813 3944
rect 3167 3936 3273 3944
rect 3556 3944 3564 3956
rect 4727 3956 4793 3964
rect 5316 3956 5453 3964
rect 3556 3936 3653 3944
rect 3956 3936 4064 3944
rect 2267 3916 2604 3924
rect 2656 3916 2873 3924
rect 1207 3896 1293 3904
rect 1927 3896 1993 3904
rect 2007 3896 2073 3904
rect 2656 3904 2664 3916
rect 2987 3916 3053 3924
rect 3067 3916 3453 3924
rect 3956 3924 3964 3936
rect 3696 3916 3964 3924
rect 4056 3924 4064 3936
rect 5007 3936 5253 3944
rect 5316 3944 5324 3956
rect 5267 3936 5324 3944
rect 4056 3916 4233 3924
rect 2567 3896 2664 3904
rect 2687 3896 2753 3904
rect 3187 3896 3353 3904
rect 3407 3896 3593 3904
rect 3696 3904 3704 3916
rect 4347 3916 4513 3924
rect 4527 3916 4633 3924
rect 5347 3916 5493 3924
rect 3647 3896 3704 3904
rect 607 3876 693 3884
rect 707 3876 953 3884
rect 1247 3876 1333 3884
rect 1407 3876 1853 3884
rect 1947 3876 2013 3884
rect 2027 3876 2233 3884
rect 2247 3876 2473 3884
rect 2967 3876 3153 3884
rect 3227 3876 3553 3884
rect 3747 3876 3973 3884
rect 3987 3876 4133 3884
rect 4947 3876 5013 3884
rect 347 3856 413 3864
rect 1360 3864 1373 3867
rect 1356 3853 1373 3864
rect 1567 3856 1773 3864
rect 1827 3856 1973 3864
rect 2507 3856 2693 3864
rect 3787 3856 3833 3864
rect 4767 3856 5173 3864
rect 5187 3856 5393 3864
rect 87 3836 233 3844
rect 1356 3847 1364 3853
rect 547 3836 573 3844
rect 867 3836 953 3844
rect 967 3836 1113 3844
rect 1347 3836 1364 3847
rect 1347 3833 1360 3836
rect 1767 3836 1953 3844
rect 2927 3836 3044 3844
rect 127 3816 173 3824
rect 2007 3816 2033 3824
rect 247 3796 333 3804
rect 2416 3807 2424 3833
rect 2456 3807 2464 3833
rect 3036 3824 3044 3836
rect 3167 3836 3293 3844
rect 3367 3836 3413 3844
rect 3767 3836 3873 3844
rect 3036 3816 3173 3824
rect 3247 3816 3433 3824
rect 1187 3796 1213 3804
rect 1427 3796 1473 3804
rect 1567 3796 1753 3804
rect 1847 3796 1913 3804
rect 1927 3796 2073 3804
rect 2127 3796 2313 3804
rect 2407 3796 2424 3807
rect 2407 3793 2420 3796
rect 2667 3796 2713 3804
rect 2833 3804 2847 3813
rect 3447 3816 3493 3824
rect 3807 3816 3833 3824
rect 3927 3816 4353 3824
rect 4747 3816 4793 3824
rect 5327 3816 5353 3824
rect 5507 3816 5533 3824
rect 2833 3800 2913 3804
rect 2836 3796 2913 3800
rect 4100 3804 4113 3807
rect 3827 3796 3944 3804
rect 4096 3796 4113 3804
rect 147 3773 153 3787
rect 667 3776 733 3784
rect 847 3776 973 3784
rect 227 3756 353 3764
rect 367 3756 473 3764
rect 916 3747 924 3776
rect 1467 3776 1493 3784
rect 1587 3780 1764 3784
rect 1587 3776 1767 3780
rect 1753 3766 1767 3776
rect 1867 3776 2353 3784
rect 2567 3776 2653 3784
rect 2716 3784 2724 3793
rect 2953 3784 2967 3793
rect 2716 3780 2967 3784
rect 2716 3776 2964 3780
rect 3347 3776 3444 3784
rect 2307 3756 2413 3764
rect 2787 3756 3393 3764
rect 3436 3764 3444 3776
rect 3527 3776 3593 3784
rect 3936 3787 3944 3796
rect 4100 3793 4113 3796
rect 4127 3796 4193 3804
rect 4207 3796 4293 3804
rect 5213 3804 5227 3813
rect 5213 3800 5273 3804
rect 5216 3796 5273 3800
rect 3947 3776 3993 3784
rect 4187 3780 4444 3784
rect 4187 3776 4447 3780
rect 4433 3767 4447 3776
rect 4727 3776 4753 3784
rect 4821 3776 4853 3784
rect 4927 3776 5293 3784
rect 5307 3776 5433 3784
rect 5547 3776 5584 3784
rect 3436 3756 3533 3764
rect 3547 3756 3593 3764
rect 3967 3756 4153 3764
rect 567 3736 673 3744
rect 687 3736 713 3744
rect 1147 3736 1233 3744
rect 1347 3736 1513 3744
rect 1587 3736 1993 3744
rect 2367 3736 2473 3744
rect 2847 3736 3193 3744
rect 3807 3736 3833 3744
rect 3887 3736 4233 3744
rect 207 3716 313 3724
rect 1287 3716 1653 3724
rect 2067 3716 2312 3724
rect 2348 3716 2453 3724
rect 3407 3716 3693 3724
rect 3707 3716 3733 3724
rect 3787 3716 4193 3724
rect 4447 3716 4612 3724
rect 4648 3716 5233 3724
rect 447 3696 1233 3704
rect 1327 3696 1573 3704
rect 2036 3696 2593 3704
rect 1316 3684 1324 3693
rect 467 3676 1324 3684
rect 1707 3676 1773 3684
rect 2036 3684 2044 3696
rect 4587 3696 5533 3704
rect 1787 3676 2044 3684
rect 2087 3676 2493 3684
rect 2587 3676 2793 3684
rect 3207 3676 3713 3684
rect 3727 3676 4073 3684
rect 4287 3676 4533 3684
rect 4987 3676 5113 3684
rect 87 3656 473 3664
rect 1187 3656 1272 3664
rect 1308 3656 1373 3664
rect 1387 3656 2093 3664
rect 2107 3656 2513 3664
rect 2907 3656 3493 3664
rect 3507 3656 3833 3664
rect 4047 3656 4833 3664
rect 387 3636 453 3644
rect 747 3636 933 3644
rect 947 3636 1113 3644
rect 1327 3636 1773 3644
rect 1967 3636 2093 3644
rect 3247 3636 3353 3644
rect 3947 3636 4473 3644
rect 4927 3636 4993 3644
rect 27 3616 2413 3624
rect 2427 3616 2893 3624
rect 3667 3616 3753 3624
rect 3907 3616 4393 3624
rect 5027 3616 5093 3624
rect 327 3596 373 3604
rect 1127 3596 1184 3604
rect 907 3576 1133 3584
rect 1176 3584 1184 3596
rect 1207 3596 1253 3604
rect 1747 3596 1993 3604
rect 2067 3596 2133 3604
rect 2147 3596 2273 3604
rect 2327 3596 2573 3604
rect 3347 3596 3404 3604
rect 1176 3576 1313 3584
rect 1487 3576 1573 3584
rect 2027 3576 2353 3584
rect 3396 3584 3404 3596
rect 3927 3596 4173 3604
rect 4847 3596 4953 3604
rect 3396 3576 3653 3584
rect 3787 3576 3813 3584
rect 4267 3576 4473 3584
rect 4487 3576 4553 3584
rect 5027 3576 5053 3584
rect -24 3556 53 3564
rect 107 3556 213 3564
rect 227 3556 313 3564
rect 1227 3556 1313 3564
rect 115 3536 213 3544
rect -24 3516 13 3524
rect 115 3507 123 3536
rect 227 3536 593 3544
rect 953 3544 967 3553
rect 1807 3556 1973 3564
rect 1987 3556 2013 3564
rect 2127 3556 2153 3564
rect 2747 3556 3213 3564
rect 3227 3556 3353 3564
rect 3787 3556 3933 3564
rect 4947 3556 4993 3564
rect 5187 3556 5353 3564
rect 5507 3556 5533 3564
rect 787 3536 1184 3544
rect 336 3520 413 3524
rect 333 3516 413 3520
rect 333 3507 347 3516
rect 593 3524 607 3533
rect 1176 3527 1184 3536
rect 2180 3544 2193 3547
rect 593 3520 653 3524
rect 596 3516 653 3520
rect 816 3520 1013 3524
rect 813 3516 1013 3520
rect 148 3496 213 3504
rect 346 3500 347 3507
rect 368 3496 433 3504
rect 813 3507 827 3516
rect 1176 3516 1193 3527
rect 1180 3513 1193 3516
rect 1547 3513 1553 3527
rect 1733 3524 1747 3533
rect 2176 3533 2193 3544
rect 2447 3536 2493 3544
rect 3638 3544 3647 3547
rect 3638 3536 4073 3544
rect 4407 3536 4493 3544
rect 5247 3536 5333 3544
rect 1607 3520 1747 3524
rect 1607 3516 1744 3520
rect 2176 3524 2184 3533
rect 1987 3516 2184 3524
rect 2487 3516 2553 3524
rect 2947 3516 3033 3524
rect 3567 3516 3773 3524
rect 3847 3516 3953 3524
rect 4233 3524 4247 3533
rect 4147 3520 4247 3524
rect 4147 3516 4244 3520
rect 5507 3516 5584 3524
rect 447 3496 533 3504
rect 727 3496 813 3504
rect 307 3476 553 3484
rect 1273 3484 1287 3494
rect 3173 3504 3187 3513
rect 3047 3500 3187 3504
rect 3047 3496 3184 3500
rect 3367 3496 3433 3504
rect 3876 3500 3913 3504
rect 1273 3480 1373 3484
rect 1276 3476 1373 3480
rect 1527 3476 1913 3484
rect 2287 3476 2693 3484
rect 3293 3484 3307 3493
rect 3127 3476 3333 3484
rect 3533 3484 3547 3493
rect 3873 3496 3913 3500
rect 3873 3487 3887 3496
rect 4267 3496 4353 3504
rect 4407 3496 4513 3504
rect 4527 3496 4573 3504
rect 4787 3496 5053 3504
rect 5147 3496 5193 3504
rect 5327 3496 5453 3504
rect 3487 3476 3713 3484
rect 4707 3476 4852 3484
rect 4888 3476 4933 3484
rect 4947 3476 5033 3484
rect 387 3456 473 3464
rect 1107 3456 1353 3464
rect 1747 3456 2284 3464
rect 527 3436 713 3444
rect 1387 3436 1513 3444
rect 1567 3436 1713 3444
rect 2276 3444 2284 3456
rect 3927 3456 3993 3464
rect 4007 3456 4033 3464
rect 4747 3456 4953 3464
rect 5067 3456 5133 3464
rect 2276 3436 2393 3444
rect 2527 3436 2573 3444
rect 3107 3436 3453 3444
rect 3727 3436 4053 3444
rect 5087 3436 5273 3444
rect 1827 3416 2153 3424
rect 3087 3416 3333 3424
rect 3667 3416 4013 3424
rect 4547 3416 4653 3424
rect 4807 3416 5053 3424
rect 5147 3416 5373 3424
rect 67 3396 593 3404
rect 767 3396 873 3404
rect 887 3396 984 3404
rect 976 3387 984 3396
rect 1347 3396 1393 3404
rect 2367 3396 2813 3404
rect 3336 3404 3344 3413
rect 3167 3396 3224 3404
rect 3336 3396 4173 3404
rect 987 3376 1093 3384
rect 1587 3376 1773 3384
rect 1787 3376 1913 3384
rect 2207 3376 2413 3384
rect 3216 3384 3224 3396
rect 4767 3396 5093 3404
rect 3216 3376 3413 3384
rect 4647 3376 4733 3384
rect 5267 3376 5493 3384
rect 1007 3356 1333 3364
rect 1567 3356 1793 3364
rect 2107 3356 2393 3364
rect 2407 3356 2613 3364
rect 2627 3356 3033 3364
rect 3447 3356 3553 3364
rect 3607 3356 3873 3364
rect 4187 3356 4313 3364
rect 307 3336 433 3344
rect 667 3336 693 3344
rect 707 3336 853 3344
rect 867 3336 953 3344
rect 1247 3336 1493 3344
rect 1907 3336 2593 3344
rect 2727 3336 2913 3344
rect 3207 3336 3513 3344
rect 4627 3336 4693 3344
rect 5047 3336 5113 3344
rect 1387 3316 1533 3324
rect 4047 3316 4373 3324
rect 4907 3316 4993 3324
rect 5247 3316 5433 3324
rect 567 3296 733 3304
rect 747 3296 793 3304
rect 1327 3296 1593 3304
rect 1696 3300 1733 3304
rect 1693 3296 1733 3300
rect 887 3276 933 3284
rect 1693 3287 1707 3296
rect 1807 3296 1993 3304
rect 2007 3296 2073 3304
rect 2313 3304 2327 3313
rect 2313 3300 2393 3304
rect 2316 3296 2393 3300
rect 3367 3296 3379 3304
rect 4067 3296 4173 3304
rect 4667 3296 4713 3304
rect 4867 3296 4913 3304
rect 5027 3296 5133 3304
rect 5147 3293 5153 3307
rect 5327 3296 5453 3304
rect 1047 3276 1073 3284
rect 1147 3276 1173 3284
rect 1347 3276 1553 3284
rect 2447 3276 2613 3284
rect 2907 3276 3273 3284
rect 3587 3276 3793 3284
rect 3807 3273 3813 3287
rect 4147 3276 4304 3284
rect -24 3256 13 3264
rect 87 3256 133 3264
rect 1247 3256 1313 3264
rect 2047 3256 2133 3264
rect 2667 3253 2673 3267
rect 3007 3256 3113 3264
rect 3447 3256 3499 3264
rect 4207 3256 4253 3264
rect 4296 3264 4304 3276
rect 4347 3276 4433 3284
rect 4496 3276 4533 3284
rect 4296 3256 4373 3264
rect 4387 3256 4473 3264
rect 4496 3247 4504 3276
rect 4947 3276 4993 3284
rect 4847 3253 4853 3267
rect 5047 3256 5113 3264
rect 67 3236 93 3244
rect 567 3236 693 3244
rect 707 3236 793 3244
rect 807 3236 933 3244
rect 1347 3236 1413 3244
rect 1456 3240 1693 3244
rect 1453 3236 1693 3240
rect 1453 3228 1467 3236
rect 1847 3236 1893 3244
rect 2287 3236 2967 3244
rect 2981 3236 3173 3244
rect 3607 3236 3953 3244
rect 3967 3236 4113 3244
rect 4127 3236 4153 3244
rect 4480 3246 4504 3247
rect 4487 3236 4504 3246
rect 4487 3233 4500 3236
rect 4567 3236 4673 3244
rect 4727 3236 4793 3244
rect 5253 3244 5267 3253
rect 5227 3240 5267 3244
rect 5227 3236 5264 3240
rect 687 3216 733 3224
rect 747 3216 873 3224
rect 2047 3216 2213 3224
rect 2767 3216 2853 3224
rect 2867 3216 2913 3224
rect 3707 3216 4773 3224
rect 5187 3216 5393 3224
rect 327 3196 393 3204
rect 907 3196 1193 3204
rect 1467 3196 1513 3204
rect 1647 3196 1713 3204
rect 2007 3196 2093 3204
rect 2107 3196 2553 3204
rect 2916 3204 2924 3212
rect 2916 3196 3073 3204
rect 3087 3196 3293 3204
rect 3367 3196 3633 3204
rect 4627 3196 4973 3204
rect 27 3176 513 3184
rect 1267 3176 1372 3184
rect 1408 3176 1533 3184
rect 1547 3176 1813 3184
rect 1887 3176 2693 3184
rect 3296 3184 3304 3193
rect 3296 3176 3393 3184
rect 5407 3176 5513 3184
rect 607 3156 2713 3164
rect 3027 3156 3173 3164
rect 3247 3156 3433 3164
rect 3456 3156 5233 3164
rect 387 3136 433 3144
rect 447 3136 493 3144
rect 507 3136 1453 3144
rect 1476 3136 2033 3144
rect 27 3116 153 3124
rect 1476 3124 1484 3136
rect 2367 3136 2393 3144
rect 3456 3144 3464 3156
rect 3327 3136 3464 3144
rect 4587 3136 4633 3144
rect 527 3116 1484 3124
rect 2207 3116 4753 3124
rect 4767 3116 4993 3124
rect 5127 3116 5193 3124
rect 287 3096 432 3104
rect 468 3096 553 3104
rect 687 3096 1073 3104
rect 1087 3096 1273 3104
rect 1367 3096 1453 3104
rect 2387 3096 2473 3104
rect 2707 3096 3333 3104
rect 3387 3096 3493 3104
rect 3507 3096 3733 3104
rect 3887 3096 4593 3104
rect 87 3076 153 3084
rect 167 3076 613 3084
rect 627 3076 813 3084
rect 1027 3076 1113 3084
rect 1127 3076 1473 3084
rect 1567 3076 1593 3084
rect 2187 3076 3353 3084
rect 4807 3076 5193 3084
rect 5427 3076 5533 3084
rect 1307 3056 1433 3064
rect 2027 3056 2053 3064
rect 2847 3056 2953 3064
rect 3247 3056 3413 3064
rect 4467 3056 4533 3064
rect 4576 3056 4773 3064
rect 4576 3047 4584 3056
rect 267 3036 353 3044
rect 1467 3036 1593 3044
rect 3347 3036 3613 3044
rect 4287 3036 4573 3044
rect 4647 3036 4873 3044
rect 5547 3036 5584 3044
rect 0 3024 13 3027
rect -4 3014 13 3024
rect -4 3013 20 3014
rect 107 3016 633 3024
rect -4 2984 4 3013
rect 27 2996 53 3004
rect 176 2987 184 3016
rect 767 3016 853 3024
rect 867 3016 1053 3024
rect 1147 3016 1213 3024
rect 1787 3016 1933 3024
rect 1987 3016 2144 3024
rect 2136 3007 2144 3016
rect 2187 3016 2213 3024
rect 507 2996 533 3004
rect 607 2996 699 3004
rect 1267 2996 1566 3004
rect 1787 2996 1813 3004
rect 1827 2996 1953 3004
rect 2147 2994 2153 3007
rect 2147 2993 2160 2994
rect 2673 3004 2687 3013
rect 4267 3016 4439 3024
rect 4747 3016 4793 3024
rect 2547 3000 2687 3004
rect 2547 2996 2684 3000
rect 2947 2996 3386 3004
rect 3838 3004 3847 3007
rect 3838 2996 4193 3004
rect -4 2976 53 2984
rect 247 2976 353 2984
rect 447 2976 893 2984
rect 907 2976 1053 2984
rect 1487 2976 1573 2984
rect 2027 2976 2153 2984
rect 3307 2976 3353 2984
rect 467 2956 493 2964
rect 779 2956 813 2964
rect 779 2953 787 2956
rect 1207 2956 1413 2964
rect 1747 2956 2373 2964
rect 2507 2956 2713 2964
rect 2727 2956 3073 2964
rect 3187 2956 3473 2964
rect 3767 2956 3913 2964
rect 4416 2964 4424 2994
rect 4487 2996 4613 3004
rect 5007 2996 5053 3004
rect 5227 2996 5313 3004
rect 5527 2996 5584 3004
rect 4913 2984 4927 2993
rect 4847 2980 4927 2984
rect 4847 2976 4924 2980
rect 4307 2956 4593 2964
rect 4607 2956 4633 2964
rect 5127 2956 5153 2964
rect 127 2936 213 2944
rect 227 2936 433 2944
rect 487 2936 553 2944
rect 1007 2936 1133 2944
rect 1147 2936 1273 2944
rect 1727 2936 1913 2944
rect 1927 2936 2053 2944
rect 2127 2936 2273 2944
rect 2527 2936 2853 2944
rect 3447 2936 3973 2944
rect 4387 2936 4413 2944
rect 467 2916 1373 2924
rect 3627 2916 3853 2924
rect 27 2896 133 2904
rect 507 2896 873 2904
rect 1127 2896 1173 2904
rect 1187 2896 1333 2904
rect 1427 2896 1613 2904
rect 1767 2896 2073 2904
rect 2567 2896 3253 2904
rect 3876 2896 5453 2904
rect 3876 2884 3884 2896
rect 3407 2876 3884 2884
rect 207 2856 293 2864
rect 307 2856 633 2864
rect 1467 2856 1713 2864
rect 4847 2856 5133 2864
rect 1727 2836 1773 2844
rect 4327 2836 4393 2844
rect 4907 2836 4993 2844
rect 807 2816 1033 2824
rect 1047 2816 1193 2824
rect 1507 2816 1553 2824
rect 1567 2816 1793 2824
rect 1927 2816 1993 2824
rect 3087 2816 3413 2824
rect 4107 2816 4533 2824
rect 5327 2816 5493 2824
rect 427 2796 513 2804
rect 827 2796 933 2804
rect 1407 2796 1633 2804
rect 1647 2796 1733 2804
rect 1847 2796 1893 2804
rect 2387 2796 2553 2804
rect 47 2776 73 2784
rect 87 2776 313 2784
rect 816 2784 824 2793
rect 727 2776 824 2784
rect 1053 2784 1067 2793
rect 1027 2780 1067 2784
rect 1027 2776 1064 2780
rect 2433 2787 2447 2796
rect 2887 2796 3033 2804
rect 3416 2804 3424 2813
rect 3416 2796 3653 2804
rect 4267 2796 4333 2804
rect 4413 2787 4427 2793
rect 1667 2774 1673 2787
rect 1660 2773 1673 2774
rect 1787 2776 1953 2784
rect 2147 2776 2313 2784
rect 2667 2776 3433 2784
rect 3867 2776 3913 2784
rect 4413 2780 4433 2787
rect 4416 2776 4433 2780
rect 4420 2773 4433 2776
rect 4973 2784 4987 2793
rect 4747 2780 4987 2784
rect 5273 2784 5287 2793
rect 5273 2780 5353 2784
rect 4747 2776 4984 2780
rect 5276 2776 5353 2780
rect 227 2756 253 2764
rect 947 2756 993 2764
rect 1167 2756 1213 2764
rect 1387 2756 1452 2764
rect 1473 2753 1474 2760
rect -24 2736 33 2744
rect 147 2733 153 2747
rect 833 2744 847 2753
rect 833 2740 873 2744
rect 836 2736 873 2740
rect 1473 2744 1487 2753
rect 3247 2760 3384 2764
rect 3247 2756 3387 2760
rect 1427 2740 1487 2744
rect 1427 2736 1484 2740
rect 1653 2744 1667 2752
rect 3373 2747 3387 2756
rect 3507 2756 3613 2764
rect 3727 2756 3813 2764
rect 4167 2756 4233 2764
rect 1627 2740 1667 2744
rect 1627 2736 1664 2740
rect 2067 2736 2113 2744
rect 2367 2736 2493 2744
rect 3067 2736 3193 2744
rect 3613 2744 3627 2753
rect 5027 2756 5153 2764
rect 3613 2740 3873 2744
rect 3616 2736 3873 2740
rect 4287 2736 4553 2744
rect 4807 2733 4813 2747
rect 4887 2736 4973 2744
rect 1747 2716 1993 2724
rect 2207 2716 2693 2724
rect 3267 2716 3593 2724
rect 3607 2716 3633 2724
rect 4727 2716 5033 2724
rect 227 2696 313 2704
rect 487 2696 573 2704
rect 713 2704 727 2713
rect 713 2700 833 2704
rect 716 2696 833 2700
rect 1967 2696 2013 2704
rect 2027 2696 2153 2704
rect 5087 2696 5213 2704
rect 5227 2696 5353 2704
rect 5447 2696 5493 2704
rect 47 2676 2193 2684
rect 2727 2676 2753 2684
rect 2767 2676 2833 2684
rect 2847 2676 2893 2684
rect 3027 2656 3273 2664
rect 3287 2656 3413 2664
rect 3427 2656 3833 2664
rect 4307 2656 4553 2664
rect 4567 2656 4733 2664
rect 4747 2656 5293 2664
rect 5307 2656 5373 2664
rect 5387 2656 5453 2664
rect 2467 2636 3133 2644
rect 4067 2636 4153 2644
rect 507 2616 553 2624
rect 947 2616 1273 2624
rect 1347 2616 1613 2624
rect 4627 2616 4953 2624
rect 5407 2616 5513 2624
rect 447 2596 533 2604
rect 827 2596 1353 2604
rect 4407 2596 4873 2604
rect 5247 2596 5353 2604
rect 607 2576 693 2584
rect 707 2576 973 2584
rect 2407 2576 2653 2584
rect 4607 2576 4673 2584
rect 4867 2576 4933 2584
rect 5167 2576 5413 2584
rect 1367 2556 1633 2564
rect 3147 2556 4313 2564
rect 247 2536 273 2544
rect 567 2536 733 2544
rect 1087 2536 1953 2544
rect 5287 2536 5353 2544
rect 5367 2536 5413 2544
rect 487 2516 653 2524
rect 767 2516 793 2524
rect 807 2516 1133 2524
rect 3307 2516 3533 2524
rect 3547 2516 3793 2524
rect 3807 2516 3953 2524
rect 3967 2516 4073 2524
rect 4447 2516 4473 2524
rect 4636 2516 5033 2524
rect 107 2496 273 2504
rect 167 2476 261 2484
rect 253 2473 261 2476
rect 713 2484 727 2493
rect 767 2496 893 2504
rect 1207 2496 1433 2504
rect 1587 2496 1773 2504
rect 2087 2496 2533 2504
rect 2847 2496 2873 2504
rect 4187 2496 4253 2504
rect 4636 2507 4644 2516
rect 5047 2516 5193 2524
rect 4547 2496 4633 2504
rect 4767 2496 4813 2504
rect 5320 2504 5333 2507
rect 5316 2500 5333 2504
rect 5313 2494 5333 2500
rect 5313 2493 5340 2494
rect 5447 2496 5473 2504
rect 5313 2487 5327 2493
rect 647 2480 727 2484
rect 647 2476 724 2480
rect 1387 2476 1413 2484
rect 1981 2476 2353 2484
rect 2787 2476 2939 2484
rect 3167 2476 3273 2484
rect 4273 2473 4293 2487
rect 4507 2476 4533 2484
rect 290 2456 353 2464
rect 367 2456 413 2464
rect 867 2456 893 2464
rect 1173 2464 1187 2467
rect 967 2456 1293 2464
rect 1307 2456 1493 2464
rect 1507 2456 1613 2464
rect 1627 2456 1793 2464
rect 1887 2456 2373 2464
rect 2547 2456 2673 2464
rect 2907 2456 3033 2464
rect 3047 2456 3093 2464
rect 147 2436 233 2444
rect 513 2444 527 2453
rect 387 2440 527 2444
rect 387 2436 524 2440
rect 607 2436 633 2444
rect 1407 2433 1413 2447
rect 1967 2436 2293 2444
rect 2587 2436 2913 2444
rect 3327 2440 3384 2444
rect 3327 2436 3387 2440
rect 3373 2427 3387 2436
rect 3647 2433 3653 2447
rect 3840 2444 3853 2447
rect 3727 2436 3853 2444
rect 3833 2433 3853 2436
rect 4233 2444 4247 2453
rect 4233 2440 4433 2444
rect 4236 2436 4433 2440
rect 4833 2444 4847 2453
rect 4767 2436 4873 2444
rect 5433 2444 5447 2453
rect 5007 2440 5447 2444
rect 5007 2436 5444 2440
rect 1327 2416 1373 2424
rect 2127 2416 2213 2424
rect 2327 2416 3073 2424
rect 3833 2427 3847 2433
rect 3947 2416 4073 2424
rect 4727 2416 4753 2424
rect 507 2396 553 2404
rect 1927 2396 1973 2404
rect 2667 2396 2812 2404
rect 2848 2396 2953 2404
rect 5147 2396 5353 2404
rect 267 2376 1253 2384
rect 4007 2376 4573 2384
rect 347 2356 393 2364
rect 667 2356 1913 2364
rect 3087 2356 3233 2364
rect 4747 2356 5153 2364
rect 687 2336 1013 2344
rect 1027 2336 1224 2344
rect 1216 2324 1224 2336
rect 1447 2336 1553 2344
rect 2007 2336 2073 2344
rect 2187 2336 2413 2344
rect 2567 2336 2593 2344
rect 3127 2336 3193 2344
rect 3996 2336 4533 2344
rect 3996 2327 4004 2336
rect 4707 2336 4873 2344
rect 5047 2336 5113 2344
rect 1216 2316 2333 2324
rect 3827 2316 3993 2324
rect 5247 2316 5333 2324
rect 1207 2296 2373 2304
rect 2387 2296 2453 2304
rect 3047 2296 3113 2304
rect 3327 2296 4213 2304
rect 4367 2296 4913 2304
rect 5327 2296 5413 2304
rect 67 2276 313 2284
rect 327 2276 393 2284
rect 707 2276 753 2284
rect 2827 2276 2973 2284
rect 3507 2276 3533 2284
rect 3767 2276 3953 2284
rect 307 2256 413 2264
rect 887 2256 973 2264
rect 1067 2256 1093 2264
rect 1587 2256 1613 2264
rect 1767 2256 1833 2264
rect 1879 2253 1893 2267
rect 2047 2256 2193 2264
rect 2287 2253 2293 2267
rect 2347 2256 2873 2264
rect 3427 2256 3553 2264
rect 4427 2256 4473 2264
rect 4773 2264 4781 2267
rect 4716 2260 4781 2264
rect 4713 2256 4781 2260
rect 4713 2247 4727 2256
rect 587 2236 613 2244
rect 767 2233 773 2247
rect 1027 2236 1153 2244
rect 1647 2236 1713 2244
rect 2467 2236 2513 2244
rect 3067 2236 3093 2244
rect 3107 2236 3193 2244
rect 3273 2244 3281 2247
rect 3207 2236 3281 2244
rect 3887 2236 4093 2244
rect 4467 2240 4604 2244
rect 4467 2236 4607 2240
rect 53 2204 67 2213
rect 276 2207 284 2233
rect 447 2216 533 2224
rect 547 2216 913 2224
rect 1056 2220 1113 2224
rect 1053 2216 1113 2220
rect 1053 2207 1067 2216
rect 1827 2213 1833 2227
rect 2233 2224 2247 2233
rect 4593 2227 4607 2236
rect 4947 2236 5073 2244
rect 5147 2236 5193 2244
rect 5267 2236 5373 2244
rect 1847 2220 2247 2224
rect 1847 2216 2244 2220
rect 3487 2213 3493 2227
rect 4147 2216 4193 2224
rect 4287 2216 4413 2224
rect 4887 2213 4893 2227
rect 5407 2216 5473 2224
rect 53 2200 173 2204
rect 56 2196 173 2200
rect 987 2196 1013 2204
rect 1327 2196 2033 2204
rect 2047 2196 2293 2204
rect 2307 2196 2393 2204
rect 2607 2196 2853 2204
rect 2967 2196 3133 2204
rect 3147 2196 3373 2204
rect 3567 2196 3633 2204
rect 3647 2196 3913 2204
rect 4136 2204 4144 2212
rect 4136 2196 4233 2204
rect 347 2176 393 2184
rect 407 2176 493 2184
rect 907 2176 1273 2184
rect 1487 2176 1673 2184
rect 3667 2176 4313 2184
rect 4767 2176 4953 2184
rect 107 2156 253 2164
rect 2507 2156 2993 2164
rect 3907 2156 4093 2164
rect 607 2136 1073 2144
rect 1367 2136 1693 2144
rect 3067 2136 3233 2144
rect 3247 2136 4653 2144
rect 2647 2116 2693 2124
rect 2887 2116 2913 2124
rect 4787 2116 5053 2124
rect 1307 2096 1473 2104
rect 1487 2096 1533 2104
rect 2867 2096 3153 2104
rect 2367 2076 2593 2084
rect 2947 2076 3073 2084
rect 3087 2076 3613 2084
rect 4487 2076 4713 2084
rect 4727 2076 4793 2084
rect 5327 2076 5353 2084
rect 47 2056 93 2064
rect 247 2056 673 2064
rect 1467 2056 1513 2064
rect 1627 2056 1893 2064
rect 2467 2056 2653 2064
rect 3687 2056 3993 2064
rect 327 2036 653 2044
rect 4387 2036 4773 2044
rect 2527 2016 2833 2024
rect 3027 2016 3133 2024
rect 3967 2016 4153 2024
rect 4267 2016 4973 2024
rect 5107 2016 5333 2024
rect 47 1996 93 2004
rect 287 1996 353 2004
rect 1887 1996 1933 2004
rect 3707 1996 4333 2004
rect 4527 1996 4593 2004
rect 4867 1996 4933 2004
rect 5387 1996 5453 2004
rect -24 1956 113 1964
rect 307 1956 353 1964
rect 813 1964 821 1967
rect 647 1956 821 1964
rect 927 1954 933 1967
rect 920 1953 933 1954
rect 493 1944 507 1953
rect 493 1940 673 1944
rect 496 1936 673 1940
rect 347 1913 353 1927
rect 913 1924 927 1932
rect 1027 1936 1279 1944
rect 1496 1946 1504 1974
rect 1767 1976 1813 1984
rect 2007 1976 2273 1984
rect 2853 1984 2867 1993
rect 2787 1980 2867 1984
rect 2787 1976 2864 1980
rect 3387 1976 3493 1984
rect 3827 1976 3913 1984
rect 4047 1976 4253 1984
rect 4327 1976 4353 1984
rect 4767 1976 4833 1984
rect 4847 1976 4993 1984
rect 5007 1976 5173 1984
rect 5347 1976 5393 1984
rect 1727 1953 1733 1967
rect 1847 1956 2113 1964
rect 2127 1956 2453 1964
rect 2687 1956 2733 1964
rect 2821 1956 2953 1964
rect 3580 1964 3593 1967
rect 3576 1953 3593 1964
rect 4087 1953 4093 1967
rect 4107 1956 4133 1964
rect 5327 1956 5413 1964
rect 953 1924 967 1933
rect 3027 1936 3193 1944
rect 3576 1944 3584 1953
rect 3527 1936 3584 1944
rect 3627 1936 3833 1944
rect 4367 1936 4533 1944
rect 4547 1936 4613 1944
rect 5027 1936 5153 1944
rect 5167 1946 5180 1947
rect 5167 1933 5173 1946
rect 913 1920 967 1924
rect 916 1916 964 1920
rect 1707 1916 1973 1924
rect 2107 1916 2133 1924
rect 2147 1916 2173 1924
rect 2327 1916 2513 1924
rect 2847 1916 2873 1924
rect 3467 1916 3533 1924
rect 4107 1916 4213 1924
rect 4427 1916 4493 1924
rect 4787 1916 5233 1924
rect 5380 1926 5393 1927
rect 5387 1913 5393 1926
rect 47 1896 93 1904
rect 2907 1896 3013 1904
rect 3027 1896 3073 1904
rect 3787 1896 3873 1904
rect 4447 1896 4573 1904
rect 4967 1896 5013 1904
rect 147 1876 453 1884
rect 1407 1876 1673 1884
rect 2807 1876 2833 1884
rect 3207 1876 3273 1884
rect 3287 1876 3453 1884
rect 4667 1876 5373 1884
rect 3067 1856 3132 1864
rect 3168 1856 3553 1864
rect 4247 1856 4453 1864
rect 4687 1856 5073 1864
rect 567 1836 633 1844
rect 1787 1836 1993 1844
rect 2007 1836 2193 1844
rect 2387 1836 2473 1844
rect 2487 1836 2773 1844
rect 2787 1836 3313 1844
rect 5367 1836 5413 1844
rect 56 1816 93 1824
rect 56 1804 64 1816
rect 167 1816 253 1824
rect 267 1816 373 1824
rect 387 1816 653 1824
rect 3987 1816 4464 1824
rect 36 1796 64 1804
rect 36 1767 44 1796
rect 687 1796 713 1804
rect 1547 1796 1713 1804
rect 2573 1804 2587 1813
rect 2467 1800 2587 1804
rect 2467 1796 2584 1800
rect 2867 1796 3033 1804
rect 3847 1796 4273 1804
rect 4456 1804 4464 1816
rect 4527 1816 4673 1824
rect 5320 1824 5333 1827
rect 5316 1813 5333 1824
rect 4456 1796 4833 1804
rect 5227 1796 5273 1804
rect 107 1776 313 1784
rect 827 1776 1193 1784
rect 1567 1776 1873 1784
rect 3347 1776 3693 1784
rect 3867 1776 4013 1784
rect 4027 1776 4153 1784
rect 5067 1776 5093 1784
rect 5316 1767 5324 1813
rect 467 1756 733 1764
rect 1027 1756 1233 1764
rect 1587 1756 1793 1764
rect 2287 1756 2473 1764
rect 2727 1756 2913 1764
rect 2927 1756 2953 1764
rect 2967 1756 3133 1764
rect 3787 1756 3833 1764
rect 4787 1756 4924 1764
rect 247 1736 272 1744
rect 286 1736 413 1744
rect 793 1744 807 1753
rect 793 1740 853 1744
rect 796 1736 853 1740
rect 2073 1744 2087 1753
rect 1967 1740 2087 1744
rect 1967 1736 2084 1740
rect 3473 1744 3487 1753
rect 3387 1740 3487 1744
rect 3387 1736 3484 1740
rect 3947 1736 4053 1744
rect 4267 1736 4393 1744
rect 4916 1744 4924 1756
rect 4947 1756 5033 1764
rect 4916 1736 5093 1744
rect 747 1716 1033 1724
rect 1147 1716 1373 1724
rect 1507 1713 1513 1727
rect 1647 1716 1673 1724
rect 1827 1716 1873 1724
rect 2167 1716 2193 1724
rect 2527 1716 2773 1724
rect 3107 1716 3133 1724
rect 3347 1716 3433 1724
rect 4567 1716 4712 1724
rect 4748 1716 4773 1724
rect 5167 1716 5233 1724
rect 267 1696 293 1704
rect 387 1696 440 1704
rect 847 1696 873 1704
rect 1247 1696 1340 1704
rect 2160 1706 2173 1707
rect 2167 1693 2173 1706
rect 2867 1696 2933 1704
rect 3087 1696 3173 1704
rect 3467 1696 3693 1704
rect 3756 1696 3853 1704
rect 1407 1676 1613 1684
rect 1687 1676 2033 1684
rect 2047 1676 2273 1684
rect 2393 1684 2407 1693
rect 3756 1687 3764 1696
rect 4047 1693 4053 1707
rect 4353 1704 4367 1713
rect 4296 1700 4367 1704
rect 4293 1696 4364 1700
rect 4293 1687 4307 1696
rect 4547 1696 4593 1704
rect 4756 1696 4853 1704
rect 4756 1687 4764 1696
rect 4867 1696 4953 1704
rect 2393 1680 2473 1684
rect 2396 1676 2473 1680
rect 2487 1676 2613 1684
rect 2707 1676 2793 1684
rect 2867 1676 3133 1684
rect 3227 1676 3753 1684
rect 3827 1676 4133 1684
rect 4447 1676 4633 1684
rect 4747 1676 4764 1687
rect 4747 1673 4760 1676
rect 47 1656 93 1664
rect 247 1656 333 1664
rect 347 1656 533 1664
rect 867 1656 893 1664
rect 3007 1656 3153 1664
rect 4687 1656 4753 1664
rect 1267 1636 2253 1644
rect 2887 1636 3573 1644
rect 3727 1636 4233 1644
rect 4647 1636 4993 1644
rect 1907 1616 1933 1624
rect 1947 1616 2093 1624
rect 3827 1616 4213 1624
rect 947 1596 973 1604
rect 2827 1596 2893 1604
rect 4347 1596 4413 1604
rect 4527 1596 4693 1604
rect 4887 1596 5013 1604
rect 1627 1576 1913 1584
rect 2136 1576 2453 1584
rect 2136 1564 2144 1576
rect 2747 1576 2852 1584
rect 2888 1576 2973 1584
rect 3687 1576 4013 1584
rect 4067 1576 4313 1584
rect 787 1556 2144 1564
rect 2727 1556 3073 1564
rect 3676 1564 3684 1573
rect 3287 1556 3684 1564
rect 4047 1556 4293 1564
rect 1787 1536 1833 1544
rect 887 1516 1153 1524
rect 1907 1516 2193 1524
rect 2407 1516 2473 1524
rect 3587 1516 3993 1524
rect 4227 1516 4513 1524
rect 4607 1516 4653 1524
rect 3007 1496 3293 1504
rect 4087 1496 4113 1504
rect 4127 1496 4673 1504
rect 467 1476 493 1484
rect 607 1476 733 1484
rect 867 1476 1053 1484
rect 1067 1476 1173 1484
rect 1427 1476 1533 1484
rect 1547 1476 1913 1484
rect 2387 1476 2413 1484
rect 2487 1476 2833 1484
rect 4167 1476 4253 1484
rect 4627 1476 4873 1484
rect 267 1456 333 1464
rect 1767 1456 1793 1464
rect 3127 1456 3233 1464
rect 3247 1456 3333 1464
rect 3847 1456 4553 1464
rect 4947 1456 5032 1464
rect 5068 1456 5213 1464
rect 5287 1456 5313 1464
rect 27 1436 73 1444
rect 467 1436 553 1444
rect 1167 1436 1213 1444
rect 1307 1433 1313 1447
rect 1367 1436 1473 1444
rect 1567 1436 1753 1444
rect 1820 1444 1833 1447
rect 1816 1433 1833 1444
rect 1967 1436 1993 1444
rect 2187 1436 2493 1444
rect 2807 1436 2893 1444
rect 3407 1436 3473 1444
rect 4387 1436 4473 1444
rect 4667 1436 4713 1444
rect 4907 1436 5193 1444
rect 647 1416 693 1424
rect 1816 1424 1824 1433
rect 1507 1416 1824 1424
rect 1907 1416 1933 1424
rect 3327 1416 3393 1424
rect 3787 1416 3813 1424
rect 4107 1416 5013 1424
rect 5087 1416 5213 1424
rect 27 1396 93 1404
rect 187 1396 313 1404
rect 707 1396 773 1404
rect 927 1396 993 1404
rect 1107 1396 1373 1404
rect 1387 1396 1433 1404
rect 1720 1396 1853 1404
rect 1720 1393 1729 1396
rect 2667 1396 2713 1404
rect 2727 1393 2733 1407
rect 3247 1393 3253 1407
rect 3687 1396 3713 1404
rect 4227 1396 4453 1404
rect 4756 1400 4793 1404
rect 4753 1396 4793 1400
rect 1047 1376 1153 1384
rect 1727 1386 1729 1393
rect 4753 1387 4767 1396
rect 4927 1400 4964 1404
rect 4927 1396 4967 1400
rect 2287 1376 2333 1384
rect 2347 1376 2573 1384
rect 3367 1376 3953 1384
rect 4127 1376 4153 1384
rect 4707 1376 4753 1384
rect 4953 1387 4967 1396
rect 5267 1396 5413 1404
rect 1487 1356 1553 1364
rect 2047 1356 2173 1364
rect 3027 1356 3293 1364
rect 1527 1336 1693 1344
rect 1707 1336 1933 1344
rect 4027 1336 4233 1344
rect 4707 1336 5153 1344
rect 1127 1316 1213 1324
rect 1227 1316 1453 1324
rect 1727 1316 1773 1324
rect 2067 1316 3533 1324
rect 3547 1316 3833 1324
rect 3987 1316 5093 1324
rect 5107 1316 5293 1324
rect 467 1296 593 1304
rect 687 1296 873 1304
rect 1827 1296 1973 1304
rect 3947 1296 4153 1304
rect 247 1276 413 1284
rect 1307 1276 1473 1284
rect 2607 1276 2813 1284
rect 3547 1276 3693 1284
rect 4227 1276 4913 1284
rect 487 1256 673 1264
rect 967 1256 1133 1264
rect 1447 1264 1460 1267
rect 1447 1253 1464 1264
rect 2467 1256 3013 1264
rect 3507 1256 3713 1264
rect 4047 1256 4293 1264
rect 5027 1256 5133 1264
rect 5147 1256 5173 1264
rect 567 1236 753 1244
rect 1027 1236 1413 1244
rect 1456 1244 1464 1253
rect 1456 1236 1973 1244
rect 3527 1236 3553 1244
rect 3807 1236 3973 1244
rect 4547 1236 4593 1244
rect 5167 1236 5273 1244
rect 5427 1236 5493 1244
rect 373 1224 387 1233
rect 307 1220 387 1224
rect 307 1216 384 1220
rect 507 1216 613 1224
rect 2027 1216 2053 1224
rect 2287 1216 2373 1224
rect 2527 1216 2693 1224
rect 2707 1224 2720 1227
rect 2707 1216 2724 1224
rect 2707 1213 2720 1216
rect 2847 1216 2873 1224
rect 3447 1216 3573 1224
rect 4047 1216 4100 1224
rect 4433 1224 4447 1233
rect 4433 1220 4693 1224
rect 4436 1216 4693 1220
rect 5047 1216 5393 1224
rect 547 1196 573 1204
rect 867 1196 1273 1204
rect 1287 1196 1513 1204
rect 1567 1196 1813 1204
rect 1927 1196 2093 1204
rect 2207 1196 2493 1204
rect 2507 1196 2753 1204
rect 2767 1196 2893 1204
rect 4587 1196 4653 1204
rect 4787 1196 4893 1204
rect 5207 1196 5353 1204
rect 5427 1196 5473 1204
rect 81 1176 293 1184
rect 393 1184 407 1193
rect 393 1180 513 1184
rect 396 1176 513 1180
rect 607 1176 633 1184
rect 1887 1173 1893 1187
rect 2047 1173 2053 1187
rect 2127 1176 2173 1184
rect 2267 1173 2273 1187
rect 2308 1176 2393 1184
rect 2407 1176 2613 1184
rect 2687 1176 2713 1184
rect 2727 1176 2847 1184
rect 2861 1176 2893 1184
rect 3467 1173 3473 1187
rect 3947 1176 4013 1184
rect 4087 1176 4113 1184
rect 4207 1176 4273 1184
rect 4467 1176 4513 1184
rect 4773 1184 4787 1193
rect 4747 1180 4787 1184
rect 4747 1176 4784 1180
rect 367 1156 433 1164
rect 1727 1156 3033 1164
rect 3047 1156 3133 1164
rect 3147 1156 3353 1164
rect 4627 1156 4653 1164
rect 5107 1156 5193 1164
rect 527 1136 1013 1144
rect 1027 1136 1233 1144
rect 1767 1136 2239 1144
rect 2747 1136 2793 1144
rect 1487 1116 2353 1124
rect 3887 1116 3993 1124
rect 4927 1116 5373 1124
rect 3167 1096 3513 1104
rect 4507 1096 4773 1104
rect 1627 1076 2293 1084
rect 3767 1076 3853 1084
rect 4587 1076 4913 1084
rect 4927 1076 5173 1084
rect 707 1056 813 1064
rect 2027 1056 2213 1064
rect 2887 1056 2993 1064
rect 3327 1056 4213 1064
rect 147 1036 193 1044
rect 3027 1036 4633 1044
rect 4647 1036 5053 1044
rect 67 1016 253 1024
rect 1887 1016 2013 1024
rect 3167 1016 3373 1024
rect 3387 1016 3633 1024
rect 3687 1016 3713 1024
rect 3727 1016 4253 1024
rect 5267 1016 5413 1024
rect 5427 1016 5473 1024
rect 347 996 653 1004
rect 667 996 733 1004
rect 1947 996 1973 1004
rect 2647 996 2873 1004
rect 5127 996 5233 1004
rect 447 976 513 984
rect 967 976 1053 984
rect 2607 976 2664 984
rect 607 956 853 964
rect 1647 956 1713 964
rect 1727 956 1973 964
rect 2656 947 2664 976
rect 2987 976 3013 984
rect 4087 976 4293 984
rect 5287 976 5313 984
rect 3527 956 4133 964
rect 4707 956 4753 964
rect 4807 956 4853 964
rect 4967 956 5233 964
rect 487 936 573 944
rect 1027 936 1073 944
rect 1087 936 1173 944
rect 1187 936 1273 944
rect 1427 936 1667 944
rect 1681 936 1993 944
rect 3287 940 3324 944
rect 3287 936 3327 940
rect 367 924 387 927
rect 367 916 453 924
rect 367 913 387 916
rect 1487 916 1553 924
rect 1767 916 1913 924
rect 1927 920 1964 924
rect 1927 916 1967 920
rect 1953 907 1967 916
rect 2427 916 2453 924
rect 2547 913 2553 927
rect 2953 924 2967 933
rect 3313 927 3327 936
rect 2953 920 3033 924
rect 2956 916 3033 920
rect 3647 936 3853 944
rect 3867 936 3933 944
rect 3413 924 3427 933
rect 4247 933 4253 947
rect 4347 933 4353 947
rect 5167 936 5273 944
rect 5347 936 5413 944
rect 3413 920 3513 924
rect 3416 916 3513 920
rect 3979 924 3987 927
rect 3979 916 4093 924
rect 4493 924 4507 933
rect 4493 920 4613 924
rect 4496 916 4613 920
rect 4727 913 4733 927
rect 4847 916 4973 924
rect 127 896 344 904
rect 336 884 344 896
rect 1327 896 1593 904
rect 2167 896 2213 904
rect 2467 896 2593 904
rect 2747 896 3013 904
rect 3307 896 3373 904
rect 3387 896 3713 904
rect 5127 896 5193 904
rect 336 876 444 884
rect 436 864 444 876
rect 627 876 693 884
rect 787 876 1053 884
rect 2907 874 2913 887
rect 2900 873 2913 874
rect 2980 884 2993 887
rect 2976 876 2993 884
rect 2980 873 2993 876
rect 3007 876 3213 884
rect 3987 876 4073 884
rect 4367 876 4593 884
rect 4847 876 4893 884
rect 5007 876 5273 884
rect 5327 876 5453 884
rect 436 856 493 864
rect 2587 856 2753 864
rect 3307 856 3533 864
rect 4627 856 4713 864
rect 5027 856 5253 864
rect 3607 836 4353 844
rect 127 816 233 824
rect 247 816 373 824
rect 1027 816 2173 824
rect 2187 816 2253 824
rect 2627 816 2773 824
rect 4447 816 4673 824
rect 2847 796 3033 804
rect 3087 796 3393 804
rect 3407 796 3533 804
rect 3647 796 3673 804
rect 3887 796 3973 804
rect 4147 796 4933 804
rect 5187 796 5393 804
rect 236 776 313 784
rect 236 764 244 776
rect 2667 776 2713 784
rect 4467 776 4533 784
rect 4847 776 5113 784
rect 107 756 244 764
rect 1927 756 2153 764
rect 227 736 253 744
rect 1167 736 2253 744
rect 2807 736 3153 744
rect 3287 736 3433 744
rect 3727 736 3893 744
rect 4067 736 4433 744
rect 4787 736 4973 744
rect 1447 716 1553 724
rect 2487 716 2753 724
rect 3427 716 3733 724
rect 3927 716 4013 724
rect 267 696 313 704
rect 327 696 413 704
rect 427 696 533 704
rect 887 700 964 704
rect 887 696 967 700
rect 953 687 967 696
rect 1627 696 1753 704
rect 2107 693 2113 707
rect 2287 696 2373 704
rect 2387 696 2453 704
rect 727 676 913 684
rect 1067 676 1113 684
rect 1973 684 1987 693
rect 1973 680 2039 684
rect 1976 676 2039 680
rect 227 656 293 664
rect 387 656 433 664
rect 447 656 573 664
rect 787 656 813 664
rect 1527 656 1553 664
rect 1647 653 1653 667
rect 2193 664 2207 673
rect 2953 684 2967 693
rect 3456 696 3513 704
rect 3456 687 3464 696
rect 3773 704 3787 713
rect 4927 716 4993 724
rect 5227 716 5393 724
rect 3773 700 3893 704
rect 3776 696 3893 700
rect 4453 704 4462 707
rect 4236 700 4462 704
rect 4233 696 4462 700
rect 2953 680 3073 684
rect 2956 676 3073 680
rect 2007 660 2207 664
rect 2007 656 2204 660
rect 2267 656 2393 664
rect 2573 664 2587 673
rect 3376 676 3453 684
rect 3376 667 3384 676
rect 3747 676 3993 684
rect 4233 686 4247 696
rect 4547 696 5173 704
rect 4587 676 4733 684
rect 4787 676 5013 684
rect 5027 684 5040 687
rect 5027 676 5044 684
rect 5027 673 5040 676
rect 5307 676 5373 684
rect 2447 660 2587 664
rect 2447 656 2584 660
rect 2707 656 2753 664
rect 2767 656 2833 664
rect 3313 664 3321 667
rect 3207 656 3321 664
rect 3367 656 3384 667
rect 3367 653 3380 656
rect 4067 654 4073 667
rect 4067 653 4080 654
rect 4787 656 4813 664
rect 727 636 953 644
rect 1153 644 1167 652
rect 1087 640 1167 644
rect 1087 636 1164 640
rect 1947 636 2013 644
rect 3227 636 3293 644
rect 3787 636 3853 644
rect 4007 636 4133 644
rect 4727 636 4893 644
rect 527 616 673 624
rect 887 616 913 624
rect 3727 616 3893 624
rect 1640 596 2133 604
rect 3247 596 3333 604
rect 3347 596 3372 604
rect 3408 596 3673 604
rect 2347 576 3093 584
rect 3107 576 4353 584
rect 467 556 533 564
rect 1387 556 1793 564
rect 2336 564 2344 573
rect 1847 556 2344 564
rect 3207 556 4273 564
rect 4947 556 5393 564
rect 847 536 1033 544
rect 3867 536 3973 544
rect 547 516 1113 524
rect 1807 516 2753 524
rect 3496 516 3573 524
rect 3496 507 3504 516
rect 3587 516 4213 524
rect 4847 516 4973 524
rect 5356 516 5453 524
rect 287 496 513 504
rect 1247 496 1273 504
rect 1567 496 1753 504
rect 2547 496 2613 504
rect 2627 496 2653 504
rect 3067 496 3493 504
rect 3547 496 3633 504
rect 5356 504 5364 516
rect 5327 496 5364 504
rect 1927 476 2013 484
rect 2027 476 2273 484
rect 4087 476 4553 484
rect 4847 476 4993 484
rect 5007 476 5373 484
rect 767 456 1233 464
rect 1347 456 1433 464
rect 1447 456 1713 464
rect 2727 456 2893 464
rect 3087 456 3333 464
rect 4187 456 4253 464
rect 4507 456 4533 464
rect 4887 456 4953 464
rect 47 436 93 444
rect 1867 436 1893 444
rect 900 416 1693 424
rect 1776 420 1913 424
rect 1773 416 1913 420
rect 27 396 113 404
rect 1773 407 1787 416
rect 1107 396 1353 404
rect 1627 396 1673 404
rect 1847 396 1953 404
rect 2293 404 2307 413
rect 2647 416 2713 424
rect 3327 416 3473 424
rect 3607 416 3793 424
rect 3947 416 4113 424
rect 4207 416 4333 424
rect 4593 424 4607 433
rect 4776 436 4853 444
rect 4776 427 4784 436
rect 4867 436 5213 444
rect 5227 436 5333 444
rect 5347 436 5433 444
rect 4347 416 4773 424
rect 4827 416 5013 424
rect 5027 416 5053 424
rect 2207 400 2307 404
rect 2207 396 2304 400
rect 2493 404 2507 413
rect 2387 400 2507 404
rect 2387 396 2504 400
rect 2847 396 3253 404
rect 4307 396 4353 404
rect 4367 396 4413 404
rect 5127 396 5173 404
rect 5187 396 5253 404
rect 5487 396 5584 404
rect 136 380 333 384
rect 133 376 333 380
rect 133 367 147 376
rect 347 376 739 384
rect 1107 376 1193 384
rect 1707 376 2093 384
rect 2167 376 2693 384
rect 2707 376 2733 384
rect 3661 376 3953 384
rect 4207 376 4853 384
rect 4867 384 4880 387
rect 4867 376 4884 384
rect 4867 373 4880 376
rect 4927 376 5033 384
rect 47 356 93 364
rect 867 353 873 367
rect 1313 364 1327 373
rect 1313 360 1373 364
rect 1316 356 1373 360
rect 2267 356 2372 364
rect 2396 360 2633 364
rect 2393 356 2633 360
rect 2393 347 2407 356
rect 2807 353 2813 367
rect 2827 356 2993 364
rect 3127 356 3153 364
rect 3393 364 3407 373
rect 3393 360 3473 364
rect 3396 356 3473 360
rect 3716 360 3773 364
rect 3713 356 3773 360
rect 3713 347 3727 356
rect 5087 356 5339 364
rect 127 336 213 344
rect 407 336 573 344
rect 967 336 1013 344
rect 1027 336 1333 344
rect 1567 336 1593 344
rect 1607 336 2293 344
rect 3007 336 3073 344
rect 3307 336 3393 344
rect 4227 336 4333 344
rect 4347 336 4453 344
rect 4467 336 4713 344
rect 5147 336 5173 344
rect 2747 316 2793 324
rect 5347 316 5533 324
rect 107 296 133 304
rect 867 296 973 304
rect 1407 296 1733 304
rect 1967 296 2153 304
rect 2827 296 2933 304
rect 4587 296 5153 304
rect 267 276 293 284
rect 427 276 553 284
rect 2507 276 3533 284
rect 3547 276 3853 284
rect 4987 276 5253 284
rect 607 256 1253 264
rect 1667 256 1713 264
rect 3227 256 3293 264
rect 1767 236 1793 244
rect 2127 236 2453 244
rect 4067 236 4133 244
rect 4967 236 5213 244
rect 5267 236 5393 244
rect 2047 216 2073 224
rect 2087 216 2153 224
rect 2167 216 2533 224
rect 3267 216 3593 224
rect 3747 216 3833 224
rect 147 196 333 204
rect 527 196 793 204
rect 807 196 893 204
rect 2627 196 2773 204
rect 4747 196 4773 204
rect 5207 196 5353 204
rect 107 173 113 187
rect 267 176 433 184
rect 447 176 713 184
rect 727 176 753 184
rect 1907 176 1933 184
rect 2127 176 2173 184
rect 2736 180 2813 184
rect 2733 176 2813 180
rect 2733 167 2747 176
rect 2927 176 2953 184
rect 3013 184 3027 193
rect 3013 180 3113 184
rect 3016 176 3113 180
rect 3167 176 3193 184
rect 3596 176 3773 184
rect 3596 167 3604 176
rect 3827 176 3884 184
rect 487 156 593 164
rect 967 156 1033 164
rect 1247 156 1353 164
rect 1427 156 1513 164
rect 1580 156 1813 164
rect 2307 156 2639 164
rect 3527 156 3593 164
rect 3667 156 3853 164
rect 87 136 133 144
rect 247 136 293 144
rect 3876 147 3884 176
rect 4027 176 4493 184
rect 4507 176 5093 184
rect 3947 156 4173 164
rect 4387 156 4413 164
rect 4847 156 4919 164
rect 4987 156 5013 164
rect 5307 156 5413 164
rect 1127 136 1213 144
rect 1947 133 1953 147
rect 2107 136 2253 144
rect 2316 140 2413 144
rect 2313 136 2413 140
rect 2313 127 2327 136
rect 2547 136 2599 144
rect 4376 144 4384 153
rect 3927 136 4384 144
rect 4533 144 4547 153
rect 4533 140 4633 144
rect 4536 136 4633 140
rect 287 116 413 124
rect 687 116 833 124
rect 847 116 993 124
rect 1107 126 1120 127
rect 1107 113 1113 126
rect 1667 116 2013 124
rect 3007 116 3673 124
rect 3807 113 3813 127
rect 4227 116 4341 124
rect 4333 113 4341 116
rect 5327 116 5353 124
rect 767 96 953 104
rect 1267 96 2113 104
rect 2447 96 2953 104
rect 3787 96 4173 104
rect 4887 96 4953 104
rect 4967 96 5193 104
rect 407 76 473 84
rect 567 76 1173 84
rect 2267 76 2473 84
rect 4327 76 4673 84
rect 4927 76 5213 84
rect 2007 56 2433 64
rect 2467 36 3193 44
rect 4627 36 4673 44
rect 5407 36 5493 44
rect 4267 16 5433 24
use NOR2X1  _760_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727424219
transform 1 0 3550 0 1 790
box -12 -8 92 272
use INVX1  _761_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727401709
transform -1 0 3510 0 1 270
box -12 -8 72 272
use NOR2X1  _762_
timestamp 1727424219
transform 1 0 2950 0 1 270
box -12 -8 92 272
use OAI21X1  _763_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727399082
transform -1 0 3310 0 -1 790
box -12 -8 112 272
use INVX2  _764_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727401709
transform -1 0 2790 0 1 1310
box -12 -8 72 272
use NOR2X1  _765_
timestamp 1727424219
transform 1 0 3130 0 -1 1830
box -12 -8 92 272
use AOI22X1  _766_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727401709
transform 1 0 2930 0 1 790
box -14 -8 132 272
use OAI21X1  _767_
timestamp 1727399082
transform -1 0 3290 0 1 790
box -12 -8 112 272
use INVX1  _768_
timestamp 1727401709
transform 1 0 3070 0 1 270
box -12 -8 72 272
use INVX1  _769_
timestamp 1727401709
transform 1 0 4330 0 -1 1310
box -12 -8 72 272
use NAND2X1  _770_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727424219
transform 1 0 4270 0 1 790
box -12 -8 92 272
use OAI21X1  _771_
timestamp 1727399082
transform 1 0 4230 0 -1 790
box -12 -8 112 272
use AOI22X1  _772_
timestamp 1727401709
transform -1 0 2790 0 1 270
box -14 -8 132 272
use OAI21X1  _773_
timestamp 1727399082
transform 1 0 3170 0 1 270
box -12 -8 112 272
use NOR2X1  _774_
timestamp 1727424219
transform 1 0 3590 0 -1 270
box -12 -8 92 272
use OAI21X1  _775_
timestamp 1727399082
transform -1 0 3410 0 1 270
box -12 -8 112 272
use AOI22X1  _776_
timestamp 1727401709
transform 1 0 2070 0 1 270
box -14 -8 132 272
use OAI21X1  _777_
timestamp 1727399082
transform -1 0 3270 0 -1 270
box -12 -8 112 272
use INVX1  _778_
timestamp 1727401709
transform 1 0 3790 0 1 270
box -12 -8 72 272
use NAND2X1  _779_
timestamp 1727424219
transform 1 0 3830 0 -1 270
box -12 -8 92 272
use OAI21X1  _780_
timestamp 1727399082
transform -1 0 3810 0 -1 270
box -12 -8 112 272
use AOI22X1  _781_
timestamp 1727401709
transform -1 0 2050 0 -1 270
box -14 -8 132 272
use OAI21X1  _782_
timestamp 1727399082
transform -1 0 3030 0 -1 270
box -12 -8 112 272
use INVX2  _783_
timestamp 1727401709
transform 1 0 3470 0 1 2870
box -12 -8 72 272
use NAND2X1  _784_
timestamp 1727424219
transform -1 0 3310 0 1 2870
box -12 -8 92 272
use OAI21X1  _785_
timestamp 1727399082
transform 1 0 3350 0 1 2870
box -12 -8 112 272
use INVX2  _786_
timestamp 1727401709
transform -1 0 2470 0 -1 4430
box -12 -8 72 272
use NAND2X1  _787_
timestamp 1727424219
transform -1 0 2370 0 -1 3910
box -12 -8 92 272
use OAI21X1  _788_
timestamp 1727399082
transform -1 0 2490 0 -1 3910
box -12 -8 112 272
use INVX2  _789_
timestamp 1727401709
transform -1 0 3090 0 -1 3910
box -12 -8 72 272
use NAND2X1  _790_
timestamp 1727424219
transform -1 0 2870 0 -1 3390
box -12 -8 92 272
use OAI21X1  _791_
timestamp 1727399082
transform -1 0 3350 0 -1 3390
box -12 -8 112 272
use INVX2  _792_
timestamp 1727401709
transform -1 0 3450 0 -1 3910
box -12 -8 72 272
use NAND2X1  _793_
timestamp 1727424219
transform -1 0 3090 0 -1 3390
box -12 -8 92 272
use OAI21X1  _794_
timestamp 1727399082
transform 1 0 3390 0 -1 3390
box -12 -8 112 272
use NAND2X1  _795_
timestamp 1727424219
transform 1 0 2710 0 -1 2870
box -12 -8 92 272
use OAI21X1  _796_
timestamp 1727399082
transform -1 0 2930 0 -1 2870
box -12 -8 112 272
use NAND2X1  _797_
timestamp 1727424219
transform 1 0 2210 0 -1 3390
box -12 -8 92 272
use OAI21X1  _798_
timestamp 1727399082
transform -1 0 2350 0 1 3390
box -12 -8 112 272
use NAND2X1  _799_
timestamp 1727424219
transform 1 0 2890 0 1 3390
box -12 -8 92 272
use OAI21X1  _800_
timestamp 1727399082
transform -1 0 3090 0 1 3390
box -12 -8 112 272
use NAND2X1  _801_
timestamp 1727424219
transform 1 0 2910 0 -1 3390
box -12 -8 92 272
use OAI21X1  _802_
timestamp 1727399082
transform -1 0 3210 0 -1 3390
box -12 -8 112 272
use INVX1  _803_
timestamp 1727401709
transform -1 0 1210 0 1 790
box -12 -8 72 272
use NAND2X1  _804_
timestamp 1727424219
transform 1 0 1610 0 1 790
box -12 -8 92 272
use OAI21X1  _805_
timestamp 1727399082
transform 1 0 1250 0 1 790
box -12 -8 112 272
use INVX1  _806_
timestamp 1727401709
transform 1 0 430 0 -1 1830
box -12 -8 72 272
use NAND2X1  _807_
timestamp 1727424219
transform 1 0 270 0 1 1830
box -12 -8 92 272
use OAI21X1  _808_
timestamp 1727399082
transform -1 0 390 0 -1 1830
box -12 -8 112 272
use INVX1  _809_
timestamp 1727401709
transform 1 0 370 0 1 790
box -12 -8 72 272
use NAND2X1  _810_
timestamp 1727424219
transform 1 0 510 0 -1 1310
box -12 -8 92 272
use OAI21X1  _811_
timestamp 1727399082
transform 1 0 450 0 1 790
box -12 -8 112 272
use INVX1  _812_
timestamp 1727401709
transform -1 0 310 0 -1 270
box -12 -8 72 272
use NAND2X1  _813_
timestamp 1727424219
transform 1 0 1210 0 -1 270
box -12 -8 92 272
use OAI21X1  _814_
timestamp 1727399082
transform 1 0 530 0 1 270
box -12 -8 112 272
use INVX1  _815_
timestamp 1727401709
transform -1 0 2170 0 1 1830
box -12 -8 72 272
use NAND2X1  _816_
timestamp 1727424219
transform 1 0 2850 0 1 1830
box -12 -8 92 272
use OAI21X1  _817_
timestamp 1727399082
transform 1 0 2450 0 1 1830
box -12 -8 112 272
use INVX1  _818_
timestamp 1727401709
transform -1 0 1150 0 -1 1310
box -12 -8 72 272
use NAND2X1  _819_
timestamp 1727424219
transform -1 0 2430 0 1 1310
box -12 -8 92 272
use OAI21X1  _820_
timestamp 1727399082
transform 1 0 1410 0 -1 1310
box -12 -8 112 272
use INVX1  _821_
timestamp 1727401709
transform -1 0 1390 0 -1 1830
box -12 -8 72 272
use NAND2X1  _822_
timestamp 1727424219
transform 1 0 2290 0 -1 1830
box -12 -8 92 272
use OAI21X1  _823_
timestamp 1727399082
transform 1 0 1190 0 -1 1830
box -12 -8 112 272
use INVX1  _824_
timestamp 1727401709
transform -1 0 1890 0 -1 2350
box -12 -8 72 272
use NAND2X1  _825_
timestamp 1727424219
transform 1 0 2410 0 -1 2350
box -12 -8 92 272
use OAI21X1  _826_
timestamp 1727399082
transform -1 0 2270 0 -1 2350
box -12 -8 112 272
use INVX1  _827_
timestamp 1727401709
transform -1 0 3670 0 -1 2350
box -12 -8 72 272
use NAND2X1  _828_
timestamp 1727424219
transform -1 0 3450 0 -1 2350
box -12 -8 92 272
use OAI21X1  _829_
timestamp 1727399082
transform -1 0 3590 0 -1 2350
box -12 -8 112 272
use INVX1  _830_
timestamp 1727401709
transform 1 0 4770 0 -1 2350
box -12 -8 72 272
use NAND2X1  _831_
timestamp 1727424219
transform -1 0 4270 0 -1 2350
box -12 -8 92 272
use OAI21X1  _832_
timestamp 1727399082
transform -1 0 4510 0 -1 2350
box -12 -8 112 272
use INVX1  _833_
timestamp 1727401709
transform -1 0 3630 0 -1 2870
box -12 -8 72 272
use NAND2X1  _834_
timestamp 1727424219
transform -1 0 3030 0 -1 2870
box -12 -8 92 272
use OAI21X1  _835_
timestamp 1727399082
transform -1 0 3290 0 -1 2870
box -12 -8 112 272
use INVX1  _836_
timestamp 1727401709
transform -1 0 3450 0 -1 1830
box -12 -8 72 272
use NAND2X1  _837_
timestamp 1727424219
transform 1 0 3310 0 1 1830
box -12 -8 92 272
use OAI21X1  _838_
timestamp 1727399082
transform -1 0 3350 0 -1 1830
box -12 -8 112 272
use INVX1  _839_
timestamp 1727401709
transform 1 0 4230 0 1 2350
box -12 -8 72 272
use NAND2X1  _840_
timestamp 1727424219
transform -1 0 4150 0 -1 2350
box -12 -8 92 272
use OAI21X1  _841_
timestamp 1727399082
transform -1 0 4210 0 1 2350
box -12 -8 112 272
use INVX1  _842_
timestamp 1727401709
transform -1 0 5370 0 1 2350
box -12 -8 72 272
use NAND2X1  _843_
timestamp 1727424219
transform 1 0 5450 0 -1 2870
box -12 -8 92 272
use OAI21X1  _844_
timestamp 1727399082
transform 1 0 5390 0 1 2350
box -12 -8 112 272
use INVX1  _845_
timestamp 1727401709
transform 1 0 5350 0 1 270
box -12 -8 72 272
use NAND2X1  _846_
timestamp 1727424219
transform 1 0 5430 0 1 790
box -12 -8 92 272
use OAI21X1  _847_
timestamp 1727399082
transform 1 0 5350 0 -1 790
box -12 -8 112 272
use INVX1  _848_
timestamp 1727401709
transform 1 0 5250 0 1 270
box -12 -8 72 272
use NAND2X1  _849_
timestamp 1727424219
transform -1 0 4610 0 1 270
box -12 -8 92 272
use OAI21X1  _850_
timestamp 1727399082
transform -1 0 5230 0 1 270
box -12 -8 112 272
use INVX1  _851_
timestamp 1727401709
transform -1 0 930 0 1 1830
box -12 -8 72 272
use NAND3X1  _852_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727401709
transform -1 0 1230 0 1 2350
box -12 -8 112 272
use OAI21X1  _853_
timestamp 1727399082
transform 1 0 990 0 -1 2350
box -12 -8 112 272
use INVX1  _854_
timestamp 1727401709
transform 1 0 530 0 -1 1830
box -12 -8 72 272
use NAND2X1  _855_
timestamp 1727424219
transform 1 0 1190 0 -1 2870
box -12 -8 92 272
use NAND2X1  _856_
timestamp 1727424219
transform 1 0 1410 0 1 2870
box -12 -8 92 272
use NOR2X1  _857_
timestamp 1727424219
transform -1 0 1170 0 -1 2870
box -12 -8 92 272
use INVX1  _858_
timestamp 1727401709
transform 1 0 790 0 1 2350
box -12 -8 72 272
use INVX1  _859_
timestamp 1727401709
transform 1 0 1690 0 -1 3390
box -12 -8 72 272
use INVX2  _860_
timestamp 1727401709
transform 1 0 3230 0 1 4430
box -12 -8 72 272
use OAI21X1  _861_
timestamp 1727399082
transform -1 0 1410 0 -1 2870
box -12 -8 112 272
use NAND3X1  _862_
timestamp 1727401709
transform -1 0 970 0 1 2350
box -12 -8 112 272
use OAI21X1  _863_
timestamp 1727399082
transform 1 0 630 0 1 1830
box -12 -8 112 272
use INVX1  _864_
timestamp 1727401709
transform -1 0 90 0 -1 1310
box -12 -8 72 272
use NAND2X1  _865_
timestamp 1727424219
transform 1 0 1290 0 1 2870
box -12 -8 92 272
use NAND2X1  _866_
timestamp 1727424219
transform 1 0 1190 0 -1 3390
box -12 -8 92 272
use NOR2X1  _867_
timestamp 1727424219
transform 1 0 1170 0 1 2870
box -12 -8 92 272
use AOI22X1  _868_
timestamp 1727401709
transform 1 0 1530 0 1 2870
box -14 -8 132 272
use OAI21X1  _869_
timestamp 1727399082
transform -1 0 1070 0 -1 2870
box -12 -8 112 272
use INVX1  _870_
timestamp 1727401709
transform -1 0 950 0 -1 2870
box -12 -8 72 272
use AND2X2  _871_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727424219
transform -1 0 1650 0 -1 3390
box -12 -8 112 273
use NAND3X1  _872_
timestamp 1727401709
transform -1 0 1410 0 -1 3390
box -12 -8 112 272
use INVX1  _873_
timestamp 1727401709
transform -1 0 1030 0 1 2870
box -12 -8 72 272
use NAND3X1  _874_
timestamp 1727401709
transform -1 0 730 0 -1 2870
box -12 -8 112 272
use NAND3X1  _875_
timestamp 1727401709
transform -1 0 750 0 1 2350
box -12 -8 112 272
use INVX1  _876_
timestamp 1727401709
transform -1 0 470 0 1 2350
box -12 -8 72 272
use AOI21X1  _877_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727401709
transform -1 0 610 0 1 2350
box -12 -8 112 272
use NOR2X1  _878_
timestamp 1727424219
transform -1 0 390 0 1 2350
box -12 -8 92 272
use NAND2X1  _879_
timestamp 1727424219
transform -1 0 410 0 1 1310
box -12 -8 92 272
use OAI21X1  _880_
timestamp 1727399082
transform 1 0 370 0 -1 1310
box -12 -8 112 272
use INVX1  _881_
timestamp 1727401709
transform -1 0 90 0 -1 270
box -12 -8 72 272
use NAND2X1  _882_
timestamp 1727424219
transform 1 0 1450 0 -1 3390
box -12 -8 92 272
use AOI21X1  _883_
timestamp 1727401709
transform -1 0 850 0 -1 2870
box -12 -8 112 272
use NAND2X1  _884_
timestamp 1727424219
transform 1 0 1330 0 1 3390
box -12 -8 92 272
use NAND2X1  _885_
timestamp 1727424219
transform -1 0 970 0 -1 3910
box -12 -8 92 272
use NOR2X1  _886_
timestamp 1727424219
transform -1 0 1150 0 -1 3390
box -12 -8 92 272
use AOI22X1  _887_
timestamp 1727401709
transform 1 0 1190 0 1 3910
box -14 -8 132 272
use OAI21X1  _888_
timestamp 1727399082
transform 1 0 790 0 1 3390
box -12 -8 112 272
use INVX1  _889_
timestamp 1727401709
transform 1 0 970 0 -1 3390
box -12 -8 72 272
use AND2X2  _890_
timestamp 1727424219
transform -1 0 870 0 -1 3910
box -12 -8 112 273
use NAND2X1  _891_
timestamp 1727424219
transform -1 0 1010 0 1 3390
box -12 -8 92 272
use INVX1  _892_
timestamp 1727401709
transform 1 0 870 0 -1 3390
box -12 -8 72 272
use NAND3X1  _893_
timestamp 1727401709
transform -1 0 710 0 -1 3390
box -12 -8 112 272
use NAND3X1  _894_
timestamp 1727401709
transform -1 0 650 0 1 2870
box -12 -8 112 272
use OAI21X1  _895_
timestamp 1727399082
transform -1 0 1150 0 1 2870
box -12 -8 112 272
use AOI21X1  _896_
timestamp 1727401709
transform -1 0 850 0 -1 3390
box -12 -8 112 272
use INVX2  _897_
timestamp 1727401709
transform 1 0 1330 0 1 3910
box -12 -8 72 272
use OAI21X1  _898_
timestamp 1727399082
transform -1 0 1290 0 1 3390
box -12 -8 112 272
use INVX2  _899_
timestamp 1727401709
transform -1 0 1970 0 -1 3910
box -12 -8 72 272
use INVX1  _900_
timestamp 1727401709
transform -1 0 3310 0 -1 4430
box -12 -8 72 272
use OAI21X1  _901_
timestamp 1727399082
transform -1 0 1890 0 1 3390
box -12 -8 112 272
use AOI21X1  _902_
timestamp 1727401709
transform -1 0 1150 0 1 3390
box -12 -8 112 272
use OAI21X1  _903_
timestamp 1727399082
transform 1 0 830 0 1 2870
box -12 -8 112 272
use NAND3X1  _904_
timestamp 1727401709
transform -1 0 510 0 1 2870
box -12 -8 112 272
use INVX1  _905_
timestamp 1727401709
transform -1 0 450 0 -1 3390
box -12 -8 72 272
use NAND3X1  _906_
timestamp 1727401709
transform -1 0 130 0 1 2870
box -12 -8 112 272
use OAI21X1  _907_
timestamp 1727399082
transform -1 0 790 0 1 2870
box -12 -8 112 272
use NAND3X1  _908_
timestamp 1727401709
transform -1 0 350 0 -1 2870
box -12 -8 112 272
use AOI21X1  _909_
timestamp 1727401709
transform -1 0 150 0 1 2350
box -12 -8 112 272
use NAND3X1  _910_
timestamp 1727401709
transform -1 0 290 0 1 2350
box -12 -8 112 272
use NAND2X1  _911_
timestamp 1727424219
transform -1 0 110 0 -1 2350
box -12 -8 92 272
use OAI22X1  _912_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727423652
transform -1 0 170 0 1 1310
box -12 -8 132 272
use INVX1  _913_
timestamp 1727401709
transform 1 0 1670 0 1 1830
box -12 -8 72 272
use INVX1  _914_
timestamp 1727401709
transform -1 0 210 0 -1 2350
box -12 -8 72 272
use AOI21X1  _915_
timestamp 1727401709
transform 1 0 150 0 1 2870
box -12 -8 112 272
use OAI21X1  _916_
timestamp 1727399082
transform -1 0 390 0 1 2870
box -12 -8 112 272
use OAI21X1  _917_
timestamp 1727399082
transform -1 0 770 0 1 3390
box -12 -8 112 272
use AND2X2  _918_
timestamp 1727424219
transform -1 0 950 0 -1 4950
box -12 -8 112 273
use NAND2X1  _919_
timestamp 1727424219
transform 1 0 810 0 1 3910
box -12 -8 92 272
use AOI22X1  _920_
timestamp 1727401709
transform 1 0 1030 0 1 3910
box -14 -8 132 272
use INVX1  _921_
timestamp 1727401709
transform 1 0 690 0 1 4430
box -12 -8 72 272
use NAND2X1  _922_
timestamp 1727424219
transform -1 0 1090 0 -1 4430
box -12 -8 92 272
use INVX1  _923_
timestamp 1727401709
transform -1 0 730 0 -1 4430
box -12 -8 72 272
use NAND3X1  _924_
timestamp 1727401709
transform 1 0 670 0 1 3910
box -12 -8 112 272
use NAND2X1  _925_
timestamp 1727424219
transform -1 0 1190 0 -1 4430
box -12 -8 92 272
use NOR2X1  _926_
timestamp 1727424219
transform -1 0 990 0 -1 4430
box -12 -8 92 272
use OAI21X1  _927_
timestamp 1727399082
transform 1 0 910 0 1 3910
box -12 -8 112 272
use AOI21X1  _928_
timestamp 1727401709
transform -1 0 610 0 -1 3910
box -12 -8 112 272
use AOI21X1  _929_
timestamp 1727401709
transform -1 0 570 0 -1 3390
box -12 -8 112 272
use NAND3X1  _930_
timestamp 1727401709
transform -1 0 490 0 1 3910
box -12 -8 112 272
use OAI21X1  _931_
timestamp 1727399082
transform -1 0 630 0 1 3910
box -12 -8 112 272
use AOI21X1  _932_
timestamp 1727401709
transform -1 0 370 0 -1 3910
box -12 -8 112 272
use NAND2X1  _933_
timestamp 1727424219
transform 1 0 1510 0 -1 3910
box -12 -8 92 272
use INVX2  _934_
timestamp 1727401709
transform 1 0 1750 0 -1 3910
box -12 -8 72 272
use NAND2X1  _935_
timestamp 1727424219
transform 1 0 1790 0 1 3910
box -12 -8 92 272
use OAI21X1  _936_
timestamp 1727399082
transform 1 0 1670 0 1 3390
box -12 -8 112 272
use OAI21X1  _937_
timestamp 1727399082
transform 1 0 1450 0 1 3390
box -12 -8 112 272
use OAI21X1  _938_
timestamp 1727399082
transform -1 0 510 0 1 3390
box -12 -8 112 272
use NAND3X1  _939_
timestamp 1727401709
transform -1 0 250 0 -1 3910
box -12 -8 112 272
use NAND3X1  _940_
timestamp 1727401709
transform -1 0 750 0 -1 3910
box -12 -8 112 272
use INVX1  _941_
timestamp 1727401709
transform -1 0 370 0 1 3390
box -12 -8 72 272
use NAND3X1  _942_
timestamp 1727401709
transform 1 0 190 0 1 3390
box -12 -8 112 272
use NAND3X1  _943_
timestamp 1727401709
transform 1 0 250 0 -1 3390
box -12 -8 112 272
use INVX1  _944_
timestamp 1727401709
transform -1 0 110 0 -1 2870
box -12 -8 72 272
use AOI21X1  _945_
timestamp 1727401709
transform -1 0 230 0 -1 2870
box -12 -8 112 272
use AOI21X1  _946_
timestamp 1727401709
transform -1 0 150 0 1 3390
box -12 -8 112 272
use INVX1  _947_
timestamp 1727401709
transform -1 0 230 0 -1 3390
box -12 -8 72 272
use OAI21X1  _948_
timestamp 1727399082
transform 1 0 30 0 -1 3390
box -12 -8 112 272
use AOI21X1  _949_
timestamp 1727401709
transform -1 0 350 0 -1 2350
box -12 -8 112 272
use NAND3X1  _950_
timestamp 1727401709
transform 1 0 370 0 -1 2350
box -12 -8 112 272
use NAND2X1  _951_
timestamp 1727424219
transform -1 0 970 0 -1 2350
box -12 -8 92 272
use OAI22X1  _952_
timestamp 1727423652
transform -1 0 1350 0 -1 2350
box -12 -8 132 272
use INVX1  _953_
timestamp 1727401709
transform 1 0 870 0 -1 1830
box -12 -8 72 272
use AND2X2  _954_
timestamp 1727424219
transform -1 0 2150 0 1 3910
box -12 -8 112 273
use NAND2X1  _955_
timestamp 1727424219
transform -1 0 470 0 -1 3910
box -12 -8 92 272
use INVX1  _956_
timestamp 1727401709
transform -1 0 350 0 1 3910
box -12 -8 72 272
use AOI21X1  _957_
timestamp 1727401709
transform -1 0 130 0 -1 3910
box -12 -8 112 272
use NAND2X1  _958_
timestamp 1727424219
transform 1 0 2410 0 1 3910
box -12 -8 92 272
use INVX1  _959_
timestamp 1727401709
transform -1 0 1830 0 -1 3390
box -12 -8 72 272
use AND2X2  _960_
timestamp 1727424219
transform 1 0 1130 0 -1 3910
box -12 -8 112 273
use OAI21X1  _961_
timestamp 1727399082
transform -1 0 1730 0 -1 3910
box -12 -8 112 272
use INVX2  _962_
timestamp 1727401709
transform 1 0 1830 0 -1 3910
box -12 -8 72 272
use OAI21X1  _963_
timestamp 1727399082
transform -1 0 2010 0 1 3910
box -12 -8 112 272
use NAND3X1  _964_
timestamp 1727401709
transform 1 0 1650 0 1 3910
box -12 -8 112 272
use INVX1  _965_
timestamp 1727401709
transform -1 0 1630 0 1 3910
box -12 -8 72 272
use NAND2X1  _966_
timestamp 1727424219
transform -1 0 1330 0 -1 3910
box -12 -8 92 272
use OAI21X1  _967_
timestamp 1727399082
transform 1 0 1370 0 -1 3910
box -12 -8 112 272
use NAND3X1  _968_
timestamp 1727401709
transform 1 0 1430 0 1 3910
box -12 -8 112 272
use NAND2X1  _969_
timestamp 1727424219
transform 1 0 890 0 1 4430
box -12 -8 92 272
use AOI21X1  _970_
timestamp 1727401709
transform -1 0 650 0 1 4430
box -12 -8 112 272
use NAND2X1  _971_
timestamp 1727424219
transform 1 0 850 0 1 4950
box -12 -8 92 272
use AND2X2  _972_
timestamp 1727424219
transform -1 0 1310 0 -1 5470
box -12 -8 112 273
use NAND2X1  _973_
timestamp 1727424219
transform 1 0 750 0 1 4950
box -12 -8 92 272
use NAND2X1  _974_
timestamp 1727424219
transform -1 0 1050 0 -1 5470
box -12 -8 92 272
use NAND2X1  _975_
timestamp 1727424219
transform -1 0 590 0 -1 5470
box -12 -8 92 272
use NAND3X1  _976_
timestamp 1727401709
transform 1 0 490 0 1 4950
box -12 -8 112 272
use INVX1  _977_
timestamp 1727401709
transform -1 0 350 0 -1 5470
box -12 -8 72 272
use NAND2X1  _978_
timestamp 1727424219
transform 1 0 730 0 -1 5470
box -12 -8 92 272
use OAI21X1  _979_
timestamp 1727399082
transform -1 0 1590 0 -1 4430
box -12 -8 112 272
use NAND3X1  _980_
timestamp 1727401709
transform -1 0 250 0 -1 5470
box -12 -8 112 272
use NAND3X1  _981_
timestamp 1727401709
transform -1 0 570 0 -1 4950
box -12 -8 112 272
use OAI21X1  _982_
timestamp 1727399082
transform -1 0 870 0 -1 4430
box -12 -8 112 272
use AOI21X1  _983_
timestamp 1727401709
transform -1 0 130 0 -1 5470
box -12 -8 112 272
use AOI21X1  _984_
timestamp 1727401709
transform -1 0 470 0 1 4950
box -12 -8 112 272
use OAI21X1  _985_
timestamp 1727399082
transform 1 0 230 0 1 4950
box -12 -8 112 272
use NAND3X1  _986_
timestamp 1727401709
transform -1 0 430 0 -1 4950
box -12 -8 112 272
use AND2X2  _987_
timestamp 1727424219
transform -1 0 870 0 1 4430
box -12 -8 112 273
use NAND3X1  _988_
timestamp 1727401709
transform 1 0 630 0 1 4950
box -12 -8 112 272
use OAI21X1  _989_
timestamp 1727399082
transform -1 0 130 0 1 4950
box -12 -8 112 272
use NAND3X1  _990_
timestamp 1727401709
transform -1 0 150 0 -1 4950
box -12 -8 112 272
use NAND3X1  _991_
timestamp 1727401709
transform -1 0 270 0 -1 4430
box -12 -8 112 272
use OAI21X1  _992_
timestamp 1727399082
transform 1 0 530 0 1 3390
box -12 -8 112 272
use NAND2X1  _993_
timestamp 1727424219
transform -1 0 130 0 1 4430
box -12 -8 92 272
use NAND2X1  _994_
timestamp 1727424219
transform -1 0 110 0 1 3910
box -12 -8 92 272
use NAND3X1  _995_
timestamp 1727401709
transform -1 0 250 0 1 3910
box -12 -8 112 272
use NAND3X1  _996_
timestamp 1727401709
transform 1 0 150 0 1 4430
box -12 -8 112 272
use NAND2X1  _997_
timestamp 1727424219
transform -1 0 130 0 -1 4430
box -12 -8 92 272
use NAND3X1  _998_
timestamp 1727401709
transform 1 0 310 0 -1 4430
box -12 -8 112 272
use NAND2X1  _999_
timestamp 1727424219
transform 1 0 530 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1000_
timestamp 1727424219
transform 1 0 490 0 -1 2350
box -12 -8 92 272
use OR2X2  _1001_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727424219
transform 1 0 610 0 -1 2350
box -12 -8 112 272
use AOI22X1  _1002_
timestamp 1727401709
transform -1 0 510 0 -1 2870
box -14 -8 132 272
use INVX1  _1003_
timestamp 1727401709
transform -1 0 1730 0 1 2870
box -12 -8 72 272
use NAND3X1  _1004_
timestamp 1727401709
transform -1 0 850 0 -1 2350
box -12 -8 112 272
use OAI21X1  _1005_
timestamp 1727399082
transform -1 0 850 0 1 1830
box -12 -8 112 272
use INVX1  _1006_
timestamp 1727401709
transform -1 0 1610 0 -1 1830
box -12 -8 72 272
use AOI21X1  _1007_
timestamp 1727401709
transform 1 0 270 0 1 4430
box -12 -8 112 272
use OAI21X1  _1008_
timestamp 1727399082
transform 1 0 410 0 1 4430
box -12 -8 112 272
use NAND2X1  _1009_
timestamp 1727424219
transform -1 0 1830 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1010_
timestamp 1727399082
transform -1 0 1710 0 -1 4430
box -12 -8 112 272
use INVX1  _1011_
timestamp 1727401709
transform 1 0 1670 0 1 4430
box -12 -8 72 272
use INVX1  _1012_
timestamp 1727401709
transform 1 0 150 0 1 4950
box -12 -8 72 272
use AOI21X1  _1013_
timestamp 1727401709
transform 1 0 190 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1014_
timestamp 1727424219
transform 1 0 2310 0 -1 4430
box -12 -8 92 272
use AND2X2  _1015_
timestamp 1727424219
transform -1 0 2750 0 1 3910
box -12 -8 112 273
use OAI21X1  _1016_
timestamp 1727399082
transform 1 0 2510 0 1 3910
box -12 -8 112 272
use AND2X2  _1017_
timestamp 1727424219
transform 1 0 2010 0 -1 3910
box -12 -8 112 273
use OAI21X1  _1018_
timestamp 1727399082
transform -1 0 2250 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1019_
timestamp 1727401709
transform -1 0 2370 0 1 3910
box -12 -8 112 272
use INVX1  _1020_
timestamp 1727401709
transform -1 0 2290 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1021_
timestamp 1727424219
transform 1 0 2170 0 1 3910
box -12 -8 92 272
use OAI21X1  _1022_
timestamp 1727399082
transform -1 0 1970 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1023_
timestamp 1727401709
transform 1 0 2090 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1024_
timestamp 1727424219
transform 1 0 2290 0 -1 4950
box -12 -8 92 272
use NOR2X1  _1025_
timestamp 1727424219
transform -1 0 710 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1026_
timestamp 1727401709
transform 1 0 370 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1027_
timestamp 1727424219
transform -1 0 2330 0 1 4430
box -12 -8 92 272
use AND2X2  _1028_
timestamp 1727424219
transform -1 0 3430 0 -1 4950
box -12 -8 112 273
use OAI21X1  _1029_
timestamp 1727399082
transform 1 0 2630 0 1 4430
box -12 -8 112 272
use NAND2X1  _1030_
timestamp 1727424219
transform -1 0 3110 0 1 4430
box -12 -8 92 272
use NAND3X1  _1031_
timestamp 1727401709
transform -1 0 3010 0 1 4430
box -12 -8 112 272
use NAND3X1  _1032_
timestamp 1727401709
transform -1 0 2590 0 1 4430
box -12 -8 112 272
use INVX1  _1033_
timestamp 1727401709
transform 1 0 2770 0 1 4950
box -12 -8 72 272
use AND2X2  _1034_
timestamp 1727424219
transform 1 0 3210 0 -1 4950
box -12 -8 112 273
use NAND2X1  _1035_
timestamp 1727424219
transform 1 0 3010 0 1 4950
box -12 -8 92 272
use OAI21X1  _1036_
timestamp 1727399082
transform 1 0 2770 0 1 4430
box -12 -8 112 272
use NAND3X1  _1037_
timestamp 1727401709
transform -1 0 2750 0 1 4950
box -12 -8 112 272
use NAND3X1  _1038_
timestamp 1727401709
transform -1 0 1450 0 -1 5470
box -12 -8 112 272
use AOI22X1  _1039_
timestamp 1727401709
transform 1 0 970 0 1 4950
box -14 -8 132 272
use OAI21X1  _1040_
timestamp 1727399082
transform -1 0 930 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1041_
timestamp 1727401709
transform -1 0 2630 0 1 4950
box -12 -8 112 272
use AOI21X1  _1042_
timestamp 1727401709
transform -1 0 2450 0 1 4430
box -12 -8 112 272
use OAI21X1  _1043_
timestamp 1727399082
transform -1 0 1490 0 1 4950
box -12 -8 112 272
use NAND3X1  _1044_
timestamp 1727401709
transform 1 0 1250 0 1 4950
box -12 -8 112 272
use AND2X2  _1045_
timestamp 1727424219
transform -1 0 2250 0 -1 4950
box -12 -8 112 273
use NAND3X1  _1046_
timestamp 1727401709
transform 1 0 1630 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1047_
timestamp 1727399082
transform -1 0 1610 0 1 4950
box -12 -8 112 272
use NAND3X1  _1048_
timestamp 1727401709
transform -1 0 1750 0 1 4950
box -12 -8 112 272
use NAND3X1  _1049_
timestamp 1727401709
transform -1 0 1450 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1050_
timestamp 1727401709
transform 1 0 610 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1051_
timestamp 1727399082
transform -1 0 830 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1052_
timestamp 1727401709
transform -1 0 1890 0 1 4950
box -12 -8 112 272
use AOI21X1  _1053_
timestamp 1727401709
transform -1 0 1230 0 1 4950
box -12 -8 112 272
use OAI21X1  _1054_
timestamp 1727399082
transform 1 0 1230 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1055_
timestamp 1727401709
transform -1 0 1250 0 1 4430
box -12 -8 112 272
use NAND3X1  _1056_
timestamp 1727401709
transform 1 0 1470 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1057_
timestamp 1727399082
transform -1 0 1210 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1058_
timestamp 1727401709
transform -1 0 1630 0 1 4430
box -12 -8 112 272
use NAND3X1  _1059_
timestamp 1727401709
transform -1 0 1110 0 1 4430
box -12 -8 112 272
use INVX1  _1060_
timestamp 1727401709
transform 1 0 430 0 -1 4430
box -12 -8 72 272
use AOI21X1  _1061_
timestamp 1727401709
transform 1 0 530 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1062_
timestamp 1727401709
transform -1 0 1510 0 1 4430
box -12 -8 112 272
use AOI21X1  _1063_
timestamp 1727401709
transform 1 0 1270 0 1 4430
box -12 -8 112 272
use OAI21X1  _1064_
timestamp 1727399082
transform -1 0 1450 0 -1 4430
box -12 -8 112 272
use AND2X2  _1065_
timestamp 1727424219
transform 1 0 1750 0 1 2870
box -12 -8 112 273
use NOR2X1  _1066_
timestamp 1727424219
transform 1 0 1450 0 -1 2870
box -12 -8 92 272
use INVX1  _1067_
timestamp 1727401709
transform 1 0 1550 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1068_
timestamp 1727399082
transform -1 0 1370 0 1 2350
box -12 -8 112 272
use OAI22X1  _1069_
timestamp 1727423652
transform -1 0 1530 0 1 2350
box -12 -8 132 272
use INVX1  _1070_
timestamp 1727401709
transform 1 0 1610 0 -1 2350
box -12 -8 72 272
use NAND3X1  _1071_
timestamp 1727401709
transform 1 0 2030 0 1 2870
box -12 -8 112 272
use AOI21X1  _1072_
timestamp 1727401709
transform 1 0 1590 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1073_
timestamp 1727399082
transform 1 0 1730 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1074_
timestamp 1727424219
transform -1 0 2210 0 1 4430
box -12 -8 92 272
use AOI21X1  _1075_
timestamp 1727401709
transform 1 0 1490 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1076_
timestamp 1727399082
transform 1 0 1770 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1077_
timestamp 1727424219
transform -1 0 2570 0 -1 4430
box -12 -8 92 272
use AND2X2  _1078_
timestamp 1727424219
transform -1 0 3230 0 1 3910
box -12 -8 112 273
use OAI21X1  _1079_
timestamp 1727399082
transform 1 0 2770 0 1 3910
box -12 -8 112 272
use AND2X2  _1080_
timestamp 1727424219
transform -1 0 2630 0 -1 3910
box -12 -8 112 273
use OAI21X1  _1081_
timestamp 1727399082
transform -1 0 2750 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1082_
timestamp 1727401709
transform 1 0 2710 0 -1 4430
box -12 -8 112 272
use INVX1  _1083_
timestamp 1727401709
transform -1 0 2670 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1084_
timestamp 1727424219
transform 1 0 2890 0 1 3910
box -12 -8 92 272
use NAND2X1  _1085_
timestamp 1727424219
transform -1 0 3350 0 1 3910
box -12 -8 92 272
use OAI21X1  _1086_
timestamp 1727399082
transform 1 0 2990 0 1 3910
box -12 -8 112 272
use NAND3X1  _1087_
timestamp 1727401709
transform -1 0 2950 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1088_
timestamp 1727424219
transform -1 0 2890 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1089_
timestamp 1727401709
transform -1 0 2990 0 1 4950
box -14 -8 132 272
use NAND2X1  _1090_
timestamp 1727424219
transform 1 0 4230 0 -1 5470
box -12 -8 92 272
use AND2X2  _1091_
timestamp 1727424219
transform 1 0 3450 0 -1 4950
box -12 -8 112 273
use OAI21X1  _1092_
timestamp 1727399082
transform 1 0 3430 0 1 4430
box -12 -8 112 272
use OAI21X1  _1093_
timestamp 1727399082
transform 1 0 3490 0 1 3910
box -12 -8 112 272
use NAND3X1  _1094_
timestamp 1727401709
transform 1 0 3490 0 1 4950
box -12 -8 112 272
use INVX1  _1095_
timestamp 1727401709
transform -1 0 4130 0 1 4950
box -12 -8 72 272
use NAND2X1  _1096_
timestamp 1727424219
transform -1 0 3710 0 1 4950
box -12 -8 92 272
use AOI22X1  _1097_
timestamp 1727401709
transform -1 0 3710 0 -1 4950
box -14 -8 132 272
use INVX1  _1098_
timestamp 1727401709
transform 1 0 3850 0 1 4950
box -12 -8 72 272
use NAND3X1  _1099_
timestamp 1727401709
transform -1 0 4050 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1100_
timestamp 1727401709
transform -1 0 3330 0 1 4950
box -12 -8 112 272
use AOI22X1  _1101_
timestamp 1727401709
transform -1 0 3170 0 -1 4950
box -14 -8 132 272
use OAI21X1  _1102_
timestamp 1727399082
transform 1 0 3110 0 1 4950
box -12 -8 112 272
use AOI21X1  _1103_
timestamp 1727401709
transform 1 0 4090 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1104_
timestamp 1727401709
transform -1 0 3450 0 1 4950
box -12 -8 112 272
use OAI21X1  _1105_
timestamp 1727399082
transform 1 0 3410 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1106_
timestamp 1727401709
transform -1 0 2630 0 -1 5470
box -12 -8 112 272
use AND2X2  _1107_
timestamp 1727424219
transform -1 0 3010 0 -1 4950
box -12 -8 112 273
use NAND3X1  _1108_
timestamp 1727401709
transform 1 0 3550 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1109_
timestamp 1727399082
transform -1 0 3370 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1110_
timestamp 1727401709
transform -1 0 2910 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1111_
timestamp 1727401709
transform 1 0 2390 0 -1 5470
box -12 -8 112 272
use INVX1  _1112_
timestamp 1727401709
transform 1 0 1910 0 -1 5470
box -12 -8 72 272
use AOI21X1  _1113_
timestamp 1727401709
transform 1 0 1930 0 1 4950
box -12 -8 112 272
use AOI21X1  _1114_
timestamp 1727401709
transform -1 0 3030 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1115_
timestamp 1727401709
transform -1 0 2770 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1116_
timestamp 1727399082
transform -1 0 2230 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1117_
timestamp 1727401709
transform -1 0 2510 0 -1 4950
box -12 -8 112 272
use INVX1  _1118_
timestamp 1727401709
transform -1 0 2490 0 1 4950
box -12 -8 72 272
use NAND3X1  _1119_
timestamp 1727401709
transform -1 0 2410 0 1 4950
box -12 -8 112 272
use OAI21X1  _1120_
timestamp 1727399082
transform -1 0 2110 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1121_
timestamp 1727401709
transform -1 0 2270 0 1 4950
box -12 -8 112 272
use AOI21X1  _1122_
timestamp 1727401709
transform -1 0 1970 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1123_
timestamp 1727401709
transform -1 0 2150 0 1 4950
box -12 -8 112 272
use NAND3X1  _1124_
timestamp 1727401709
transform -1 0 2650 0 -1 4950
box -12 -8 112 272
use AOI22X1  _1125_
timestamp 1727401709
transform 1 0 1750 0 1 4430
box -14 -8 132 272
use NOR2X1  _1126_
timestamp 1727424219
transform 1 0 1910 0 1 4430
box -12 -8 92 272
use AOI21X1  _1127_
timestamp 1727401709
transform -1 0 1990 0 1 2870
box -12 -8 112 272
use OAI21X1  _1128_
timestamp 1727399082
transform 1 0 1630 0 -1 2870
box -12 -8 112 272
use INVX1  _1129_
timestamp 1727401709
transform 1 0 2010 0 -1 4430
box -12 -8 72 272
use NAND3X1  _1130_
timestamp 1727401709
transform 1 0 2010 0 1 4430
box -12 -8 112 272
use NAND3X1  _1131_
timestamp 1727401709
transform 1 0 2010 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1132_
timestamp 1727424219
transform 1 0 2010 0 1 3390
box -12 -8 92 272
use NOR2X1  _1133_
timestamp 1727424219
transform 1 0 1910 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1134_
timestamp 1727399082
transform -1 0 1870 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1135_
timestamp 1727399082
transform -1 0 1650 0 1 2350
box -12 -8 112 272
use INVX1  _1136_
timestamp 1727401709
transform -1 0 3850 0 1 2350
box -12 -8 72 272
use NAND2X1  _1137_
timestamp 1727424219
transform -1 0 1990 0 1 3390
box -12 -8 92 272
use NAND2X1  _1138_
timestamp 1727424219
transform 1 0 2130 0 1 3390
box -12 -8 92 272
use OAI21X1  _1139_
timestamp 1727399082
transform 1 0 2150 0 1 2870
box -12 -8 112 272
use AOI21X1  _1140_
timestamp 1727401709
transform -1 0 2370 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1141_
timestamp 1727399082
transform 1 0 2690 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1142_
timestamp 1727424219
transform 1 0 2970 0 -1 4430
box -12 -8 92 272
use INVX1  _1143_
timestamp 1727401709
transform -1 0 4790 0 -1 4950
box -12 -8 72 272
use INVX1  _1144_
timestamp 1727401709
transform 1 0 3190 0 -1 5470
box -12 -8 72 272
use AOI21X1  _1145_
timestamp 1727401709
transform 1 0 3070 0 -1 5470
box -12 -8 112 272
use INVX2  _1146_
timestamp 1727401709
transform -1 0 3930 0 1 3910
box -12 -8 72 272
use NOR2X1  _1147_
timestamp 1727424219
transform 1 0 3570 0 -1 4430
box -12 -8 92 272
use AND2X2  _1148_
timestamp 1727424219
transform 1 0 3710 0 1 3390
box -12 -8 112 273
use NAND3X1  _1149_
timestamp 1727401709
transform 1 0 3750 0 1 3910
box -12 -8 112 272
use AOI22X1  _1150_
timestamp 1727401709
transform -1 0 3210 0 -1 4430
box -14 -8 132 272
use INVX1  _1151_
timestamp 1727401709
transform 1 0 3330 0 -1 4430
box -12 -8 72 272
use NAND3X1  _1152_
timestamp 1727401709
transform 1 0 3810 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1153_
timestamp 1727424219
transform -1 0 2850 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1154_
timestamp 1727424219
transform 1 0 3390 0 1 3910
box -12 -8 92 272
use OAI22X1  _1155_
timestamp 1727423652
transform -1 0 3530 0 -1 4430
box -12 -8 132 272
use NAND2X1  _1156_
timestamp 1727424219
transform 1 0 3890 0 -1 4950
box -12 -8 92 272
use AND2X2  _1157_
timestamp 1727424219
transform 1 0 3750 0 -1 4950
box -12 -8 112 273
use AOI22X1  _1158_
timestamp 1727401709
transform 1 0 3930 0 1 4950
box -14 -8 132 272
use NAND2X1  _1159_
timestamp 1727424219
transform 1 0 3730 0 1 4430
box -12 -8 92 272
use NAND2X1  _1160_
timestamp 1727424219
transform 1 0 3930 0 -1 4430
box -12 -8 92 272
use AOI22X1  _1161_
timestamp 1727401709
transform -1 0 3690 0 1 4430
box -14 -8 132 272
use INVX1  _1162_
timestamp 1727401709
transform -1 0 3890 0 1 4430
box -12 -8 72 272
use OAI21X1  _1163_
timestamp 1727399082
transform 1 0 3930 0 1 4430
box -12 -8 112 272
use NOR2X1  _1164_
timestamp 1727424219
transform -1 0 4350 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1165_
timestamp 1727399082
transform -1 0 3830 0 1 4950
box -12 -8 112 272
use INVX1  _1166_
timestamp 1727401709
transform -1 0 4130 0 1 4430
box -12 -8 72 272
use AOI21X1  _1167_
timestamp 1727401709
transform -1 0 4090 0 -1 4950
box -12 -8 112 272
use NOR2X1  _1168_
timestamp 1727424219
transform 1 0 4390 0 1 4950
box -12 -8 92 272
use OAI21X1  _1169_
timestamp 1727399082
transform 1 0 4730 0 1 4950
box -12 -8 112 272
use AND2X2  _1170_
timestamp 1727424219
transform 1 0 4130 0 -1 4950
box -12 -8 112 273
use NAND2X1  _1171_
timestamp 1727424219
transform -1 0 4250 0 1 4950
box -12 -8 92 272
use NAND2X1  _1172_
timestamp 1727424219
transform -1 0 4350 0 1 4950
box -12 -8 92 272
use NAND2X1  _1173_
timestamp 1727424219
transform -1 0 4550 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1174_
timestamp 1727424219
transform 1 0 4810 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1175_
timestamp 1727401709
transform 1 0 5190 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1176_
timestamp 1727401709
transform 1 0 3670 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1177_
timestamp 1727399082
transform 1 0 3810 0 -1 5470
box -12 -8 112 272
use NOR2X1  _1178_
timestamp 1727424219
transform -1 0 4790 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1179_
timestamp 1727401709
transform 1 0 4570 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1180_
timestamp 1727399082
transform 1 0 5050 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1181_
timestamp 1727401709
transform -1 0 5410 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1182_
timestamp 1727401709
transform -1 0 5250 0 1 4950
box -12 -8 112 272
use OAI21X1  _1183_
timestamp 1727399082
transform 1 0 4910 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1184_
timestamp 1727401709
transform -1 0 5010 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1185_
timestamp 1727401709
transform 1 0 5050 0 -1 4950
box -12 -8 112 272
use INVX1  _1186_
timestamp 1727401709
transform 1 0 4810 0 -1 4950
box -12 -8 72 272
use AOI21X1  _1187_
timestamp 1727401709
transform 1 0 4870 0 1 4950
box -12 -8 112 272
use AOI21X1  _1188_
timestamp 1727401709
transform 1 0 5430 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1189_
timestamp 1727399082
transform 1 0 5010 0 1 4950
box -12 -8 112 272
use NAND2X1  _1190_
timestamp 1727424219
transform -1 0 5190 0 -1 4430
box -12 -8 92 272
use INVX1  _1191_
timestamp 1727401709
transform 1 0 5210 0 1 2870
box -12 -8 72 272
use NOR2X1  _1192_
timestamp 1727424219
transform -1 0 5050 0 1 2870
box -12 -8 92 272
use INVX1  _1193_
timestamp 1727401709
transform -1 0 4910 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1194_
timestamp 1727399082
transform -1 0 4810 0 -1 2870
box -12 -8 112 272
use OAI22X1  _1195_
timestamp 1727423652
transform 1 0 4530 0 1 2350
box -12 -8 132 272
use INVX1  _1196_
timestamp 1727401709
transform 1 0 5210 0 1 1830
box -12 -8 72 272
use INVX8  _1197_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727424219
transform -1 0 4370 0 1 270
box -12 -8 133 272
use INVX1  _1198_
timestamp 1727401709
transform 1 0 5070 0 -1 3910
box -12 -8 72 272
use AOI21X1  _1199_
timestamp 1727401709
transform 1 0 5070 0 1 2870
box -12 -8 112 272
use AOI21X1  _1200_
timestamp 1727401709
transform 1 0 5290 0 1 4950
box -12 -8 112 272
use OAI21X1  _1201_
timestamp 1727399082
transform 1 0 5430 0 1 4950
box -12 -8 112 272
use AOI21X1  _1202_
timestamp 1727401709
transform 1 0 3670 0 -1 4430
box -12 -8 112 272
use INVX1  _1203_
timestamp 1727401709
transform -1 0 4810 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1204_
timestamp 1727424219
transform 1 0 4490 0 1 4950
box -12 -8 92 272
use OAI21X1  _1205_
timestamp 1727399082
transform -1 0 4710 0 1 4950
box -12 -8 112 272
use NOR2X1  _1206_
timestamp 1727424219
transform 1 0 3730 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1207_
timestamp 1727424219
transform -1 0 3690 0 1 3390
box -12 -8 92 272
use INVX1  _1208_
timestamp 1727401709
transform 1 0 3850 0 -1 3390
box -12 -8 72 272
use NAND2X1  _1209_
timestamp 1727424219
transform 1 0 3950 0 1 3390
box -12 -8 92 272
use OAI21X1  _1210_
timestamp 1727399082
transform -1 0 2990 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1211_
timestamp 1727401709
transform 1 0 3830 0 1 3390
box -12 -8 112 272
use NAND2X1  _1212_
timestamp 1727424219
transform -1 0 3210 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1213_
timestamp 1727399082
transform -1 0 3570 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1214_
timestamp 1727399082
transform -1 0 3710 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1215_
timestamp 1727424219
transform 1 0 4270 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1216_
timestamp 1727399082
transform 1 0 4150 0 1 4430
box -12 -8 112 272
use OAI21X1  _1217_
timestamp 1727399082
transform 1 0 4050 0 -1 4430
box -12 -8 112 272
use INVX1  _1218_
timestamp 1727401709
transform 1 0 4170 0 -1 4430
box -12 -8 72 272
use NAND3X1  _1219_
timestamp 1727401709
transform 1 0 4190 0 1 3910
box -12 -8 112 272
use NAND3X1  _1220_
timestamp 1727401709
transform -1 0 4370 0 1 4430
box -12 -8 112 272
use NAND2X1  _1221_
timestamp 1727424219
transform 1 0 4390 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1222_
timestamp 1727401709
transform 1 0 4510 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1223_
timestamp 1727401709
transform 1 0 4310 0 1 3910
box -12 -8 112 272
use INVX1  _1224_
timestamp 1727401709
transform -1 0 4450 0 -1 4430
box -12 -8 72 272
use OAI21X1  _1225_
timestamp 1727399082
transform 1 0 4610 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1226_
timestamp 1727401709
transform 1 0 4850 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1227_
timestamp 1727401709
transform 1 0 4390 0 1 4430
box -12 -8 112 272
use OAI21X1  _1228_
timestamp 1727399082
transform 1 0 4490 0 -1 4430
box -12 -8 112 272
use NAND3X1  _1229_
timestamp 1727401709
transform 1 0 4530 0 1 4430
box -12 -8 112 272
use AOI21X1  _1230_
timestamp 1727401709
transform 1 0 5430 0 1 4430
box -12 -8 112 272
use NAND3X1  _1231_
timestamp 1727401709
transform 1 0 4670 0 1 4430
box -12 -8 112 272
use NAND3X1  _1232_
timestamp 1727401709
transform 1 0 4790 0 1 4430
box -12 -8 112 272
use AOI22X1  _1233_
timestamp 1727401709
transform 1 0 4930 0 1 4430
box -14 -8 132 272
use NOR2X1  _1234_
timestamp 1727424219
transform -1 0 5150 0 1 4430
box -12 -8 92 272
use OR2X2  _1235_
timestamp 1727424219
transform 1 0 4810 0 1 2350
box -12 -8 112 272
use AOI21X1  _1236_
timestamp 1727401709
transform -1 0 4770 0 1 2350
box -12 -8 112 272
use AOI22X1  _1237_
timestamp 1727401709
transform -1 0 4990 0 -1 2350
box -14 -8 132 272
use INVX1  _1238_
timestamp 1727401709
transform -1 0 3830 0 -1 2870
box -12 -8 72 272
use NAND2X1  _1239_
timestamp 1727424219
transform -1 0 5390 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1240_
timestamp 1727401709
transform 1 0 5190 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1241_
timestamp 1727401709
transform -1 0 5510 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1242_
timestamp 1727424219
transform -1 0 5410 0 1 4430
box -12 -8 92 272
use NOR2X1  _1243_
timestamp 1727424219
transform -1 0 5290 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1244_
timestamp 1727399082
transform 1 0 5190 0 1 4430
box -12 -8 112 272
use AOI21X1  _1245_
timestamp 1727401709
transform 1 0 5050 0 1 3390
box -12 -8 112 272
use NAND2X1  _1246_
timestamp 1727424219
transform -1 0 5390 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1247_
timestamp 1727399082
transform 1 0 4370 0 -1 3910
box -12 -8 112 272
use INVX1  _1248_
timestamp 1727401709
transform -1 0 4910 0 1 3910
box -12 -8 72 272
use NAND2X1  _1249_
timestamp 1727424219
transform -1 0 4150 0 1 3910
box -12 -8 92 272
use NAND2X1  _1250_
timestamp 1727424219
transform -1 0 4030 0 1 3910
box -12 -8 92 272
use NAND2X1  _1251_
timestamp 1727424219
transform -1 0 3710 0 1 3910
box -12 -8 92 272
use OAI21X1  _1252_
timestamp 1727399082
transform 1 0 3250 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1253_
timestamp 1727424219
transform 1 0 4050 0 1 3390
box -12 -8 92 272
use OAI21X1  _1254_
timestamp 1727399082
transform -1 0 3990 0 -1 3910
box -12 -8 112 272
use OR2X2  _1255_
timestamp 1727424219
transform 1 0 4010 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1256_
timestamp 1727399082
transform 1 0 3750 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1257_
timestamp 1727424219
transform 1 0 4250 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1258_
timestamp 1727401709
transform 1 0 4450 0 1 3910
box -12 -8 112 272
use NAND3X1  _1259_
timestamp 1727401709
transform 1 0 4590 0 1 3910
box -12 -8 112 272
use INVX1  _1260_
timestamp 1727401709
transform -1 0 5130 0 1 3910
box -12 -8 72 272
use OAI21X1  _1261_
timestamp 1727399082
transform -1 0 5050 0 1 3910
box -12 -8 112 272
use INVX1  _1262_
timestamp 1727401709
transform 1 0 5150 0 1 3910
box -12 -8 72 272
use NAND3X1  _1263_
timestamp 1727401709
transform 1 0 5250 0 1 3910
box -12 -8 112 272
use NAND3X1  _1264_
timestamp 1727401709
transform -1 0 5470 0 1 3910
box -12 -8 112 272
use NAND2X1  _1265_
timestamp 1727424219
transform 1 0 5370 0 -1 270
box -12 -8 92 272
use NAND3X1  _1266_
timestamp 1727401709
transform 1 0 5430 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1267_
timestamp 1727424219
transform 1 0 5170 0 1 3390
box -12 -8 92 272
use NAND2X1  _1268_
timestamp 1727424219
transform 1 0 4990 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1269_
timestamp 1727401709
transform -1 0 1950 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1270_
timestamp 1727401709
transform -1 0 5090 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1271_
timestamp 1727401709
transform 1 0 3610 0 -1 3390
box -12 -8 112 272
use INVX1  _1272_
timestamp 1727401709
transform -1 0 4950 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1273_
timestamp 1727399082
transform 1 0 4750 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1274_
timestamp 1727401709
transform -1 0 4710 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1275_
timestamp 1727399082
transform 1 0 3810 0 1 2870
box -12 -8 112 272
use NAND2X1  _1276_
timestamp 1727424219
transform -1 0 4930 0 1 1310
box -12 -8 92 272
use AOI21X1  _1277_
timestamp 1727401709
transform -1 0 4830 0 1 3910
box -12 -8 112 272
use OAI21X1  _1278_
timestamp 1727399082
transform 1 0 4130 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1279_
timestamp 1727399082
transform 1 0 4170 0 1 3390
box -12 -8 112 272
use NOR2X1  _1280_
timestamp 1727424219
transform 1 0 3510 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1281_
timestamp 1727424219
transform -1 0 4030 0 -1 3390
box -12 -8 92 272
use AND2X2  _1282_
timestamp 1727424219
transform 1 0 4310 0 1 3390
box -12 -8 112 273
use OR2X2  _1283_
timestamp 1727424219
transform 1 0 4550 0 1 3390
box -12 -8 112 272
use NAND2X1  _1284_
timestamp 1727424219
transform -1 0 4530 0 1 3390
box -12 -8 92 272
use NAND2X1  _1285_
timestamp 1727424219
transform 1 0 4610 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1286_
timestamp 1727424219
transform -1 0 4810 0 -1 3910
box -12 -8 92 272
use AND2X2  _1287_
timestamp 1727424219
transform 1 0 4830 0 -1 3910
box -12 -8 112 273
use NOR2X1  _1288_
timestamp 1727424219
transform 1 0 5390 0 -1 3910
box -12 -8 92 272
use INVX1  _1289_
timestamp 1727401709
transform 1 0 5470 0 -1 3390
box -12 -8 72 272
use NAND3X1  _1290_
timestamp 1727401709
transform -1 0 5430 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1291_
timestamp 1727399082
transform 1 0 5110 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1292_
timestamp 1727424219
transform -1 0 5310 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1293_
timestamp 1727401709
transform 1 0 5310 0 1 2870
box -12 -8 112 272
use NAND2X1  _1294_
timestamp 1727424219
transform 1 0 5190 0 1 1310
box -12 -8 92 272
use INVX1  _1295_
timestamp 1727401709
transform -1 0 4430 0 -1 2870
box -12 -8 72 272
use NAND3X1  _1296_
timestamp 1727401709
transform -1 0 5390 0 1 3390
box -12 -8 112 272
use NOR2X1  _1297_
timestamp 1727424219
transform -1 0 4890 0 1 3390
box -12 -8 92 272
use INVX1  _1298_
timestamp 1727401709
transform -1 0 5030 0 -1 3910
box -12 -8 72 272
use NOR2X1  _1299_
timestamp 1727424219
transform 1 0 5270 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1300_
timestamp 1727424219
transform 1 0 5170 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1301_
timestamp 1727399082
transform 1 0 4910 0 1 3390
box -12 -8 112 272
use AOI21X1  _1302_
timestamp 1727401709
transform -1 0 4790 0 1 3390
box -12 -8 112 272
use INVX1  _1303_
timestamp 1727401709
transform -1 0 4350 0 -1 3390
box -12 -8 72 272
use NAND3X1  _1304_
timestamp 1727401709
transform 1 0 4150 0 -1 3390
box -12 -8 112 272
use INVX1  _1305_
timestamp 1727401709
transform -1 0 4130 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1306_
timestamp 1727399082
transform 1 0 4370 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1307_
timestamp 1727424219
transform 1 0 4530 0 1 2870
box -12 -8 92 272
use NAND2X1  _1308_
timestamp 1727424219
transform 1 0 4410 0 1 2870
box -12 -8 92 272
use INVX1  _1309_
timestamp 1727401709
transform -1 0 4390 0 1 2870
box -12 -8 72 272
use OAI21X1  _1310_
timestamp 1727399082
transform -1 0 4290 0 1 2870
box -12 -8 112 272
use OAI22X1  _1311_
timestamp 1727423652
transform -1 0 4330 0 -1 2870
box -12 -8 132 272
use INVX1  _1312_
timestamp 1727401709
transform 1 0 5350 0 -1 2870
box -12 -8 72 272
use OR2X2  _1313_
timestamp 1727424219
transform 1 0 4630 0 1 2870
box -12 -8 112 272
use INVX1  _1314_
timestamp 1727401709
transform 1 0 4770 0 1 2870
box -12 -8 72 272
use OAI21X1  _1315_
timestamp 1727399082
transform 1 0 4490 0 -1 3390
box -12 -8 112 272
use NOR2X1  _1316_
timestamp 1727424219
transform 1 0 4870 0 1 2870
box -12 -8 92 272
use AOI22X1  _1317_
timestamp 1727401709
transform -1 0 5070 0 -1 2870
box -14 -8 132 272
use NOR2X1  _1318_
timestamp 1727424219
transform -1 0 1010 0 1 790
box -12 -8 92 272
use INVX1  _1319_
timestamp 1727401709
transform 1 0 990 0 -1 790
box -12 -8 72 272
use NAND2X1  _1320_
timestamp 1727424219
transform -1 0 1110 0 1 790
box -12 -8 92 272
use NAND2X1  _1321_
timestamp 1727424219
transform -1 0 1170 0 -1 790
box -12 -8 92 272
use NAND2X1  _1322_
timestamp 1727424219
transform 1 0 2750 0 -1 790
box -12 -8 92 272
use OAI21X1  _1323_
timestamp 1727399082
transform 1 0 2390 0 -1 790
box -12 -8 112 272
use NOR2X1  _1324_
timestamp 1727424219
transform -1 0 510 0 1 1310
box -12 -8 92 272
use NOR2X1  _1325_
timestamp 1727424219
transform -1 0 290 0 1 1310
box -12 -8 92 272
use NOR2X1  _1326_
timestamp 1727424219
transform -1 0 670 0 1 790
box -12 -8 92 272
use NAND2X1  _1327_
timestamp 1727424219
transform -1 0 910 0 1 790
box -12 -8 92 272
use OAI21X1  _1328_
timestamp 1727399082
transform 1 0 710 0 1 790
box -12 -8 112 272
use NAND2X1  _1329_
timestamp 1727424219
transform 1 0 730 0 -1 790
box -12 -8 92 272
use NAND2X1  _1330_
timestamp 1727424219
transform 1 0 1390 0 1 270
box -12 -8 92 272
use OAI21X1  _1331_
timestamp 1727399082
transform 1 0 1010 0 1 270
box -12 -8 112 272
use OAI21X1  _1332_
timestamp 1727399082
transform 1 0 630 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1333_
timestamp 1727424219
transform -1 0 130 0 -1 790
box -12 -8 92 272
use NOR2X1  _1334_
timestamp 1727424219
transform -1 0 350 0 1 790
box -12 -8 92 272
use NOR2X1  _1335_
timestamp 1727424219
transform 1 0 170 0 -1 790
box -12 -8 92 272
use NAND2X1  _1336_
timestamp 1727424219
transform 1 0 530 0 -1 790
box -12 -8 92 272
use OR2X2  _1337_
timestamp 1727424219
transform 1 0 410 0 -1 790
box -12 -8 112 272
use NAND2X1  _1338_
timestamp 1727424219
transform 1 0 630 0 -1 790
box -12 -8 92 272
use NAND2X1  _1339_
timestamp 1727424219
transform 1 0 910 0 1 270
box -12 -8 92 272
use OAI21X1  _1340_
timestamp 1727399082
transform -1 0 950 0 -1 790
box -12 -8 112 272
use AOI21X1  _1341_
timestamp 1727401709
transform -1 0 370 0 -1 790
box -12 -8 112 272
use NOR2X1  _1342_
timestamp 1727424219
transform -1 0 210 0 -1 270
box -12 -8 92 272
use NOR2X1  _1343_
timestamp 1727424219
transform -1 0 410 0 -1 270
box -12 -8 92 272
use OAI21X1  _1344_
timestamp 1727399082
transform 1 0 450 0 -1 270
box -12 -8 112 272
use INVX1  _1345_
timestamp 1727401709
transform 1 0 890 0 -1 270
box -12 -8 72 272
use INVX1  _1346_
timestamp 1727401709
transform -1 0 750 0 -1 270
box -12 -8 72 272
use INVX1  _1347_
timestamp 1727401709
transform 1 0 590 0 -1 270
box -12 -8 72 272
use NAND3X1  _1348_
timestamp 1727401709
transform 1 0 970 0 -1 270
box -12 -8 112 272
use NAND2X1  _1349_
timestamp 1727424219
transform -1 0 1190 0 -1 270
box -12 -8 92 272
use NAND2X1  _1350_
timestamp 1727424219
transform 1 0 1730 0 1 270
box -12 -8 92 272
use OAI21X1  _1351_
timestamp 1727399082
transform 1 0 1330 0 -1 270
box -12 -8 112 272
use NAND2X1  _1352_
timestamp 1727424219
transform -1 0 2650 0 1 790
box -12 -8 92 272
use NOR2X1  _1353_
timestamp 1727424219
transform -1 0 2070 0 1 1830
box -12 -8 92 272
use NOR2X1  _1354_
timestamp 1727424219
transform -1 0 1850 0 1 1830
box -12 -8 92 272
use OAI21X1  _1355_
timestamp 1727399082
transform 1 0 770 0 -1 270
box -12 -8 112 272
use INVX1  _1356_
timestamp 1727401709
transform 1 0 2310 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1357_
timestamp 1727399082
transform 1 0 2170 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1358_
timestamp 1727424219
transform 1 0 2070 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1359_
timestamp 1727424219
transform 1 0 2210 0 1 790
box -12 -8 92 272
use NAND2X1  _1360_
timestamp 1727424219
transform 1 0 2330 0 1 790
box -12 -8 92 272
use OAI21X1  _1361_
timestamp 1727399082
transform 1 0 2450 0 1 790
box -12 -8 112 272
use INVX1  _1362_
timestamp 1727401709
transform -1 0 2410 0 1 270
box -12 -8 72 272
use AOI21X1  _1363_
timestamp 1727401709
transform -1 0 2190 0 1 790
box -12 -8 112 272
use NOR2X1  _1364_
timestamp 1727424219
transform -1 0 970 0 1 1310
box -12 -8 92 272
use NOR2X1  _1365_
timestamp 1727424219
transform 1 0 1110 0 1 1310
box -12 -8 92 272
use NOR2X1  _1366_
timestamp 1727424219
transform 1 0 990 0 1 1310
box -12 -8 92 272
use AND2X2  _1367_
timestamp 1727424219
transform -1 0 1990 0 -1 790
box -12 -8 112 273
use NOR2X1  _1368_
timestamp 1727424219
transform 1 0 2010 0 -1 790
box -12 -8 92 272
use OAI21X1  _1369_
timestamp 1727399082
transform 1 0 2130 0 -1 790
box -12 -8 112 272
use OAI21X1  _1370_
timestamp 1727399082
transform -1 0 2330 0 1 270
box -12 -8 112 272
use NAND2X1  _1371_
timestamp 1727424219
transform 1 0 1670 0 -1 790
box -12 -8 92 272
use NAND2X1  _1372_
timestamp 1727424219
transform -1 0 1430 0 1 1310
box -12 -8 92 272
use OAI21X1  _1373_
timestamp 1727399082
transform 1 0 1210 0 1 1310
box -12 -8 112 272
use AND2X2  _1374_
timestamp 1727424219
transform -1 0 2030 0 -1 1310
box -12 -8 112 273
use AOI21X1  _1375_
timestamp 1727401709
transform -1 0 1550 0 1 1310
box -12 -8 112 272
use NOR2X1  _1376_
timestamp 1727424219
transform 1 0 1650 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1377_
timestamp 1727424219
transform 1 0 1430 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1378_
timestamp 1727424219
transform 1 0 1750 0 -1 1830
box -12 -8 92 272
use INVX1  _1379_
timestamp 1727401709
transform -1 0 1590 0 1 790
box -12 -8 72 272
use AND2X2  _1380_
timestamp 1727424219
transform 1 0 1430 0 -1 790
box -12 -8 112 273
use OAI21X1  _1381_
timestamp 1727399082
transform -1 0 1490 0 1 790
box -12 -8 112 272
use OAI21X1  _1382_
timestamp 1727399082
transform 1 0 1550 0 -1 790
box -12 -8 112 272
use INVX1  _1383_
timestamp 1727401709
transform 1 0 1870 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1384_
timestamp 1727399082
transform 1 0 1790 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1385_
timestamp 1727424219
transform -1 0 1950 0 1 1830
box -12 -8 92 272
use NOR2X1  _1386_
timestamp 1727424219
transform -1 0 1790 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1387_
timestamp 1727424219
transform 1 0 1950 0 -1 1830
box -12 -8 92 272
use OR2X2  _1388_
timestamp 1727424219
transform 1 0 1950 0 1 790
box -12 -8 112 272
use NAND2X1  _1389_
timestamp 1727424219
transform 1 0 1710 0 1 790
box -12 -8 92 272
use NAND2X1  _1390_
timestamp 1727424219
transform 1 0 1830 0 1 790
box -12 -8 92 272
use NAND2X1  _1391_
timestamp 1727424219
transform 1 0 1970 0 1 270
box -12 -8 92 272
use OAI21X1  _1392_
timestamp 1727399082
transform -1 0 1930 0 1 270
box -12 -8 112 272
use NAND2X1  _1393_
timestamp 1727424219
transform -1 0 3430 0 -1 1310
box -12 -8 92 272
use INVX1  _1394_
timestamp 1727401709
transform 1 0 2190 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1395_
timestamp 1727399082
transform 1 0 2070 0 -1 1830
box -12 -8 112 272
use AND2X2  _1396_
timestamp 1727424219
transform 1 0 1570 0 1 1310
box -12 -8 112 273
use AOI21X1  _1397_
timestamp 1727401709
transform 1 0 1850 0 1 1310
box -12 -8 112 272
use NAND3X1  _1398_
timestamp 1727401709
transform 1 0 1710 0 1 1310
box -12 -8 112 272
use AND2X2  _1399_
timestamp 1727424219
transform 1 0 1970 0 1 1310
box -12 -8 112 273
use INVX1  _1400_
timestamp 1727401709
transform 1 0 3830 0 1 1310
box -12 -8 72 272
use NOR2X1  _1401_
timestamp 1727424219
transform 1 0 3670 0 1 2350
box -12 -8 92 272
use NOR2X1  _1402_
timestamp 1727424219
transform 1 0 3950 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1403_
timestamp 1727424219
transform 1 0 3990 0 1 1830
box -12 -8 92 272
use NOR2X1  _1404_
timestamp 1727424219
transform 1 0 3710 0 1 1310
box -12 -8 92 272
use INVX1  _1405_
timestamp 1727401709
transform -1 0 3670 0 1 1310
box -12 -8 72 272
use OAI21X1  _1406_
timestamp 1727399082
transform -1 0 3570 0 1 1310
box -12 -8 112 272
use OAI21X1  _1407_
timestamp 1727399082
transform -1 0 3570 0 -1 1310
box -12 -8 112 272
use AOI21X1  _1408_
timestamp 1727401709
transform 1 0 4210 0 1 1830
box -12 -8 112 272
use NOR2X1  _1409_
timestamp 1727424219
transform 1 0 5090 0 1 1830
box -12 -8 92 272
use NOR2X1  _1410_
timestamp 1727424219
transform 1 0 4710 0 1 1830
box -12 -8 92 272
use NOR2X1  _1411_
timestamp 1727424219
transform -1 0 5150 0 -1 1830
box -12 -8 92 272
use AND2X2  _1412_
timestamp 1727424219
transform -1 0 4570 0 1 1830
box -12 -8 112 273
use NOR2X1  _1413_
timestamp 1727424219
transform -1 0 4690 0 1 1830
box -12 -8 92 272
use OAI21X1  _1414_
timestamp 1727399082
transform -1 0 4450 0 1 1830
box -12 -8 112 272
use OAI21X1  _1415_
timestamp 1727399082
transform 1 0 4390 0 1 1310
box -12 -8 112 272
use NAND2X1  _1416_
timestamp 1727424219
transform 1 0 3710 0 -1 790
box -12 -8 92 272
use AND2X2  _1417_
timestamp 1727424219
transform 1 0 4450 0 -1 1830
box -12 -8 112 273
use OAI21X1  _1418_
timestamp 1727399082
transform -1 0 5050 0 1 1830
box -12 -8 112 272
use OAI21X1  _1419_
timestamp 1727399082
transform 1 0 4810 0 1 1830
box -12 -8 112 272
use AOI21X1  _1420_
timestamp 1727401709
transform 1 0 4690 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1421_
timestamp 1727424219
transform 1 0 3870 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1422_
timestamp 1727424219
transform 1 0 3650 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1423_
timestamp 1727424219
transform 1 0 4110 0 1 1830
box -12 -8 92 272
use INVX1  _1424_
timestamp 1727401709
transform 1 0 4170 0 -1 1830
box -12 -8 72 272
use AND2X2  _1425_
timestamp 1727424219
transform -1 0 4090 0 -1 1310
box -12 -8 112 273
use OAI21X1  _1426_
timestamp 1727399082
transform 1 0 4110 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1427_
timestamp 1727399082
transform -1 0 3950 0 -1 1310
box -12 -8 112 272
use INVX1  _1428_
timestamp 1727401709
transform -1 0 4030 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1429_
timestamp 1727399082
transform -1 0 4150 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1430_
timestamp 1727424219
transform 1 0 3370 0 1 1310
box -12 -8 92 272
use NAND2X1  _1431_
timestamp 1727424219
transform 1 0 3250 0 1 1310
box -12 -8 92 272
use INVX1  _1432_
timestamp 1727401709
transform -1 0 3230 0 1 1310
box -12 -8 72 272
use NOR2X1  _1433_
timestamp 1727424219
transform 1 0 3710 0 -1 1830
box -12 -8 92 272
use INVX1  _1434_
timestamp 1727401709
transform 1 0 4270 0 -1 1830
box -12 -8 72 272
use OR2X2  _1435_
timestamp 1727424219
transform -1 0 4130 0 1 790
box -12 -8 112 272
use AOI21X1  _1436_
timestamp 1727401709
transform -1 0 3990 0 1 790
box -12 -8 112 272
use AOI22X1  _1437_
timestamp 1727401709
transform 1 0 3830 0 -1 790
box -14 -8 132 272
use NAND2X1  _1438_
timestamp 1727424219
transform 1 0 4610 0 1 790
box -12 -8 92 272
use AOI21X1  _1439_
timestamp 1727401709
transform 1 0 3830 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1440_
timestamp 1727424219
transform 1 0 4350 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1441_
timestamp 1727424219
transform 1 0 4950 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1442_
timestamp 1727424219
transform 1 0 4830 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1443_
timestamp 1727424219
transform 1 0 4570 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1444_
timestamp 1727424219
transform -1 0 4610 0 1 1310
box -12 -8 92 272
use OR2X2  _1445_
timestamp 1727424219
transform 1 0 4730 0 1 1310
box -12 -8 112 272
use NOR2X1  _1446_
timestamp 1727424219
transform 1 0 4430 0 1 2350
box -12 -8 92 272
use NOR2X1  _1447_
timestamp 1727424219
transform 1 0 4310 0 1 2350
box -12 -8 92 272
use NOR2X1  _1448_
timestamp 1727424219
transform 1 0 4650 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1449_
timestamp 1727424219
transform 1 0 4770 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1450_
timestamp 1727424219
transform -1 0 4710 0 1 1310
box -12 -8 92 272
use INVX1  _1451_
timestamp 1727401709
transform 1 0 4890 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1452_
timestamp 1727399082
transform -1 0 4950 0 1 790
box -12 -8 112 272
use OAI21X1  _1453_
timestamp 1727399082
transform -1 0 4830 0 1 790
box -12 -8 112 272
use INVX1  _1454_
timestamp 1727401709
transform 1 0 4630 0 -1 4950
box -12 -8 72 272
use INVX1  _1455_
timestamp 1727401709
transform 1 0 4430 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1456_
timestamp 1727399082
transform -1 0 4610 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1457_
timestamp 1727424219
transform 1 0 5370 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1458_
timestamp 1727424219
transform -1 0 5270 0 1 2350
box -12 -8 92 272
use NOR2X1  _1459_
timestamp 1727424219
transform 1 0 5250 0 -1 2350
box -12 -8 92 272
use INVX1  _1460_
timestamp 1727401709
transform 1 0 5310 0 1 1310
box -12 -8 72 272
use OR2X2  _1461_
timestamp 1727424219
transform 1 0 4970 0 -1 790
box -12 -8 112 272
use AOI21X1  _1462_
timestamp 1727401709
transform -1 0 4950 0 -1 790
box -12 -8 112 272
use AOI22X1  _1463_
timestamp 1727401709
transform 1 0 4690 0 -1 790
box -14 -8 132 272
use NAND2X1  _1464_
timestamp 1727424219
transform -1 0 4390 0 -1 270
box -12 -8 92 272
use AOI21X1  _1465_
timestamp 1727401709
transform -1 0 5290 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1466_
timestamp 1727424219
transform 1 0 5230 0 1 790
box -12 -8 92 272
use INVX1  _1467_
timestamp 1727401709
transform 1 0 5350 0 1 790
box -12 -8 72 272
use OAI21X1  _1468_
timestamp 1727399082
transform -1 0 5210 0 1 790
box -12 -8 112 272
use NOR2X1  _1469_
timestamp 1727424219
transform -1 0 4870 0 -1 270
box -12 -8 92 272
use INVX1  _1470_
timestamp 1727401709
transform -1 0 5030 0 -1 1310
box -12 -8 72 272
use AOI21X1  _1471_
timestamp 1727401709
transform 1 0 4990 0 1 790
box -12 -8 112 272
use OAI21X1  _1472_
timestamp 1727399082
transform -1 0 4850 0 1 270
box -12 -8 112 272
use OAI21X1  _1473_
timestamp 1727399082
transform -1 0 4750 0 -1 270
box -12 -8 112 272
use NAND2X1  _1474_
timestamp 1727424219
transform 1 0 4190 0 -1 270
box -12 -8 92 272
use NAND3X1  _1475_
timestamp 1727401709
transform -1 0 4990 0 -1 270
box -12 -8 112 272
use OAI21X1  _1476_
timestamp 1727399082
transform 1 0 4990 0 1 270
box -12 -8 112 272
use NAND2X1  _1477_
timestamp 1727424219
transform 1 0 4870 0 1 270
box -12 -8 92 272
use OAI21X1  _1478_
timestamp 1727399082
transform -1 0 4230 0 1 270
box -12 -8 112 272
use INVX1  _1479_
timestamp 1727401709
transform 1 0 4170 0 1 790
box -12 -8 72 272
use NAND3X1  _1480_
timestamp 1727401709
transform 1 0 3330 0 -1 790
box -12 -8 112 272
use NAND2X1  _1481_
timestamp 1727424219
transform 1 0 3890 0 1 1830
box -12 -8 92 272
use OAI21X1  _1482_
timestamp 1727399082
transform -1 0 3850 0 1 1830
box -12 -8 112 272
use INVX1  _1483_
timestamp 1727401709
transform 1 0 5410 0 1 1310
box -12 -8 72 272
use NAND2X1  _1484_
timestamp 1727424219
transform -1 0 5370 0 1 1830
box -12 -8 92 272
use OAI21X1  _1485_
timestamp 1727399082
transform 1 0 5410 0 1 1830
box -12 -8 112 272
use INVX1  _1486_
timestamp 1727401709
transform 1 0 4650 0 1 270
box -12 -8 72 272
use NAND2X1  _1487_
timestamp 1727424219
transform -1 0 5270 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1488_
timestamp 1727399082
transform 1 0 5070 0 -1 1310
box -12 -8 112 272
use INVX1  _1489_
timestamp 1727401709
transform -1 0 3570 0 -1 270
box -12 -8 72 272
use NAND2X1  _1490_
timestamp 1727424219
transform 1 0 4110 0 -1 790
box -12 -8 92 272
use OAI21X1  _1491_
timestamp 1727399082
transform 1 0 3970 0 -1 790
box -12 -8 112 272
use NOR2X1  _1492_
timestamp 1727424219
transform -1 0 3190 0 -1 790
box -12 -8 92 272
use NOR2X1  _1493_
timestamp 1727424219
transform 1 0 3130 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1494_
timestamp 1727401709
transform -1 0 3090 0 -1 2350
box -12 -8 112 272
use NOR2X1  _1495_
timestamp 1727424219
transform -1 0 3330 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1496_
timestamp 1727401709
transform 1 0 3070 0 1 2350
box -12 -8 112 272
use NOR2X1  _1497_
timestamp 1727424219
transform 1 0 2970 0 1 2350
box -12 -8 92 272
use AOI21X1  _1498_
timestamp 1727401709
transform -1 0 2930 0 1 2350
box -12 -8 112 272
use NOR2X1  _1499_
timestamp 1727424219
transform -1 0 3510 0 1 1830
box -12 -8 92 272
use AOI21X1  _1500_
timestamp 1727401709
transform 1 0 3530 0 1 1830
box -12 -8 112 272
use INVX1  _1501_
timestamp 1727401709
transform 1 0 2910 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1502_
timestamp 1727399082
transform -1 0 3110 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1503_
timestamp 1727399082
transform 1 0 2950 0 1 1830
box -12 -8 112 272
use OAI21X1  _1504_
timestamp 1727399082
transform -1 0 2750 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1505_
timestamp 1727399082
transform -1 0 2870 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1506_
timestamp 1727399082
transform -1 0 2690 0 1 1310
box -12 -8 112 272
use OAI21X1  _1507_
timestamp 1727399082
transform 1 0 2450 0 1 1310
box -12 -8 112 272
use OAI21X1  _1508_
timestamp 1727399082
transform 1 0 2590 0 1 1830
box -12 -8 112 272
use OAI21X1  _1509_
timestamp 1727399082
transform -1 0 2830 0 1 1830
box -12 -8 112 272
use NOR2X1  _1510_
timestamp 1727424219
transform -1 0 2710 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1511_
timestamp 1727401709
transform -1 0 2850 0 -1 1310
box -12 -8 112 272
use NOR2X1  _1512_
timestamp 1727424219
transform -1 0 1970 0 1 2350
box -12 -8 92 272
use AOI21X1  _1513_
timestamp 1727401709
transform -1 0 2350 0 1 2350
box -12 -8 112 272
use NOR2X1  _1514_
timestamp 1727424219
transform -1 0 610 0 1 1310
box -12 -8 92 272
use AOI21X1  _1515_
timestamp 1727401709
transform -1 0 750 0 1 1310
box -12 -8 112 272
use NOR2X1  _1516_
timestamp 1727424219
transform -1 0 2170 0 -1 270
box -12 -8 92 272
use AOI21X1  _1517_
timestamp 1727401709
transform -1 0 2530 0 -1 270
box -12 -8 112 272
use NAND2X1  _1518_
timestamp 1727424219
transform 1 0 2150 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1519_
timestamp 1727399082
transform 1 0 2010 0 -1 2870
box -12 -8 112 272
use NAND2X1  _1520_
timestamp 1727424219
transform 1 0 1990 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1521_
timestamp 1727399082
transform 1 0 2090 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1522_
timestamp 1727424219
transform -1 0 2470 0 1 3390
box -12 -8 92 272
use OAI21X1  _1523_
timestamp 1727399082
transform 1 0 2510 0 1 3390
box -12 -8 112 272
use NAND2X1  _1524_
timestamp 1727424219
transform -1 0 2770 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1525_
timestamp 1727399082
transform 1 0 2570 0 -1 3390
box -12 -8 112 272
use DFFPOSX1  _1526_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727423275
transform 1 0 2950 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1527_
timestamp 1727423275
transform 1 0 2610 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1528_
timestamp 1727423275
transform 1 0 3090 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1529_
timestamp 1727423275
transform 1 0 3330 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1530_
timestamp 1727423275
transform -1 0 1410 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1531_
timestamp 1727423275
transform 1 0 10 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1532_
timestamp 1727423275
transform 1 0 10 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1533_
timestamp 1727423275
transform -1 0 490 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1534_
timestamp 1727423275
transform -1 0 2410 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1535_
timestamp 1727423275
transform -1 0 1390 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1536_
timestamp 1727423275
transform 1 0 930 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1537_
timestamp 1727423275
transform -1 0 2130 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1538_
timestamp 1727423275
transform 1 0 3410 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1539_
timestamp 1727423275
transform 1 0 4510 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1540_
timestamp 1727423275
transform 1 0 3290 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1541_
timestamp 1727423275
transform 1 0 2890 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1542_
timestamp 1727423275
transform 1 0 3950 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1543_
timestamp 1727423275
transform 1 0 4910 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1544_
timestamp 1727423275
transform -1 0 5310 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1545_
timestamp 1727423275
transform -1 0 5230 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1546_
timestamp 1727423275
transform -1 0 1170 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1547_
timestamp 1727423275
transform -1 0 590 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1548_
timestamp 1727423275
transform -1 0 330 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1549_
timestamp 1727423275
transform 1 0 10 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1550_
timestamp 1727423275
transform 1 0 1170 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1551_
timestamp 1727423275
transform 1 0 590 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1552_
timestamp 1727423275
transform 1 0 1410 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1553_
timestamp 1727423275
transform 1 0 1350 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1554_
timestamp 1727423275
transform -1 0 4090 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1555_
timestamp 1727423275
transform 1 0 4990 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1556_
timestamp 1727423275
transform 1 0 3530 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1557_
timestamp 1727423275
transform -1 0 5170 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1558_
timestamp 1727423275
transform -1 0 4670 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1559_
timestamp 1727423275
transform 1 0 5070 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1560_
timestamp 1727423275
transform 1 0 2490 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1561_
timestamp 1727423275
transform 1 0 1110 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1562_
timestamp 1727423275
transform 1 0 630 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1563_
timestamp 1727423275
transform 1 0 1430 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1564_
timestamp 1727423275
transform 1 0 2650 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1565_
timestamp 1727423275
transform 1 0 2410 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1566_
timestamp 1727423275
transform 1 0 1470 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1567_
timestamp 1727423275
transform 1 0 1670 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1568_
timestamp 1727423275
transform -1 0 3810 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1569_
timestamp 1727423275
transform 1 0 4130 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1570_
timestamp 1727423275
transform -1 0 3870 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1571_
timestamp 1727423275
transform 1 0 3510 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1572_
timestamp 1727423275
transform -1 0 4590 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1573_
timestamp 1727423275
transform -1 0 4670 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1574_
timestamp 1727423275
transform -1 0 4630 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1575_
timestamp 1727423275
transform -1 0 4150 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1576_
timestamp 1727423275
transform 1 0 3670 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1577_
timestamp 1727423275
transform -1 0 5530 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1578_
timestamp 1727423275
transform 1 0 5270 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1579_
timestamp 1727423275
transform 1 0 3850 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1580_
timestamp 1727423275
transform 1 0 2730 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1581_
timestamp 1727423275
transform 1 0 3170 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1582_
timestamp 1727423275
transform 1 0 2570 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1583_
timestamp 1727423275
transform -1 0 3690 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1584_
timestamp 1727423275
transform -1 0 3290 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1585_
timestamp 1727423275
transform -1 0 2610 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1586_
timestamp 1727423275
transform 1 0 2070 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1587_
timestamp 1727423275
transform -1 0 2730 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1588_
timestamp 1727423275
transform -1 0 2610 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1589_
timestamp 1727423275
transform -1 0 2210 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1590_
timestamp 1727423275
transform -1 0 970 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1591_
timestamp 1727423275
transform -1 0 2410 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1592_
timestamp 1727423275
transform 1 0 2230 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1593_
timestamp 1727423275
transform -1 0 2490 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1594_
timestamp 1727423275
transform 1 0 2590 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1595_
timestamp 1727423275
transform -1 0 2530 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1596_
timestamp 1727423275
transform 1 0 10 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1597_
timestamp 1727423275
transform 1 0 2530 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1598_
timestamp 1727423275
transform 1 0 2830 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1599_
timestamp 1727423275
transform -1 0 3670 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1600_
timestamp 1727423275
transform -1 0 3530 0 1 790
box -13 -8 253 272
use BUFX2  _1601_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727422626
transform 1 0 5430 0 1 270
box -12 -8 92 272
use BUFX2  _1602_
timestamp 1727422626
transform 1 0 5450 0 1 2870
box -12 -8 92 272
use BUFX2  _1603_
timestamp 1727422626
transform 1 0 5250 0 -1 270
box -12 -8 92 272
use BUFX2  _1604_
timestamp 1727422626
transform 1 0 5430 0 1 3390
box -12 -8 92 272
use BUFX2  _1605_
timestamp 1727422626
transform 1 0 4510 0 -1 3910
box -12 -8 92 272
use BUFX2  _1606_
timestamp 1727422626
transform 1 0 3410 0 -1 270
box -12 -8 92 272
use BUFX2  _1607_
timestamp 1727422626
transform 1 0 3310 0 -1 270
box -12 -8 92 272
use BUFX2  _1608_
timestamp 1727422626
transform -1 0 3130 0 -1 270
box -12 -8 92 272
use BUFX2  _1609_
timestamp 1727422626
transform -1 0 2890 0 -1 270
box -12 -8 92 272
use BUFX2  BUFX2_insert0
timestamp 1727422626
transform -1 0 3150 0 -1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert1
timestamp 1727422626
transform 1 0 4230 0 -1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert2
timestamp 1727422626
transform 1 0 4310 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert3
timestamp 1727422626
transform 1 0 3650 0 1 1830
box -12 -8 92 272
use BUFX2  BUFX2_insert4
timestamp 1727422626
transform -1 0 870 0 1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert5
timestamp 1727422626
transform -1 0 2390 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert6
timestamp 1727422626
transform -1 0 1070 0 -1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert7
timestamp 1727422626
transform -1 0 1210 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert16
timestamp 1727422626
transform -1 0 2350 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert17
timestamp 1727422626
transform -1 0 1850 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert18
timestamp 1727422626
transform 1 0 4410 0 1 270
box -12 -8 92 272
use BUFX2  BUFX2_insert19
timestamp 1727422626
transform 1 0 3090 0 1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert20
timestamp 1727422626
transform 1 0 4350 0 -1 790
box -12 -8 92 272
use BUFX2  BUFX2_insert21
timestamp 1727422626
transform -1 0 1170 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert22
timestamp 1727422626
transform -1 0 3390 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert23
timestamp 1727422626
transform -1 0 1090 0 -1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert24
timestamp 1727422626
transform -1 0 1650 0 1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert25
timestamp 1727422626
transform 1 0 1010 0 1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert26
timestamp 1727422626
transform -1 0 2910 0 1 270
box -12 -8 92 272
use BUFX2  BUFX2_insert27
timestamp 1727422626
transform 1 0 2510 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert28
timestamp 1727422626
transform 1 0 2870 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert29
timestamp 1727422626
transform 1 0 2810 0 1 1310
box -12 -8 92 272
use BUFX2  BUFX2_insert30
timestamp 1727422626
transform -1 0 1070 0 -1 4950
box -12 -8 92 272
use BUFX2  BUFX2_insert31
timestamp 1727422626
transform 1 0 3130 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert32
timestamp 1727422626
transform -1 0 1310 0 -1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert33
timestamp 1727422626
transform -1 0 4430 0 -1 5470
box -12 -8 92 272
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727396566
transform -1 0 3070 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1727396566
transform 1 0 3950 0 1 2870
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1727396566
transform -1 0 2690 0 -1 2870
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1727396566
transform 1 0 3110 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1727396566
transform 1 0 3930 0 1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert13
timestamp 1727396566
transform 1 0 2370 0 1 2350
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert14
timestamp 1727396566
transform -1 0 1750 0 -1 1310
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert15
timestamp 1727396566
transform -1 0 1870 0 1 2350
box -12 -8 212 272
use FILL  FILL81750x150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727399082
transform -1 0 5470 0 -1 270
box -12 -8 32 272
use FILL  FILL81750x7950
timestamp 1727399082
transform -1 0 5470 0 -1 790
box -12 -8 32 272
use FILL  FILL81750x31350
timestamp 1727399082
transform -1 0 5470 0 -1 2350
box -12 -8 32 272
use FILL  FILL82050x150
timestamp 1727399082
transform -1 0 5490 0 -1 270
box -12 -8 32 272
use FILL  FILL82050x7950
timestamp 1727399082
transform -1 0 5490 0 -1 790
box -12 -8 32 272
use FILL  FILL82050x19650
timestamp 1727399082
transform 1 0 5470 0 1 1310
box -12 -8 32 272
use FILL  FILL82050x31350
timestamp 1727399082
transform -1 0 5490 0 -1 2350
box -12 -8 32 272
use FILL  FILL82050x54750
timestamp 1727399082
transform -1 0 5490 0 -1 3910
box -12 -8 32 272
use FILL  FILL82050x58650
timestamp 1727399082
transform 1 0 5470 0 1 3910
box -12 -8 32 272
use FILL  FILL82350x150
timestamp 1727399082
transform -1 0 5510 0 -1 270
box -12 -8 32 272
use FILL  FILL82350x7950
timestamp 1727399082
transform -1 0 5510 0 -1 790
box -12 -8 32 272
use FILL  FILL82350x19650
timestamp 1727399082
transform 1 0 5490 0 1 1310
box -12 -8 32 272
use FILL  FILL82350x31350
timestamp 1727399082
transform -1 0 5510 0 -1 2350
box -12 -8 32 272
use FILL  FILL82350x35250
timestamp 1727399082
transform 1 0 5490 0 1 2350
box -12 -8 32 272
use FILL  FILL82350x54750
timestamp 1727399082
transform -1 0 5510 0 -1 3910
box -12 -8 32 272
use FILL  FILL82350x58650
timestamp 1727399082
transform 1 0 5490 0 1 3910
box -12 -8 32 272
use FILL  FILL82650x150
timestamp 1727399082
transform -1 0 5530 0 -1 270
box -12 -8 32 272
use FILL  FILL82650x4050
timestamp 1727399082
transform 1 0 5510 0 1 270
box -12 -8 32 272
use FILL  FILL82650x7950
timestamp 1727399082
transform -1 0 5530 0 -1 790
box -12 -8 32 272
use FILL  FILL82650x11850
timestamp 1727399082
transform 1 0 5510 0 1 790
box -12 -8 32 272
use FILL  FILL82650x15750
timestamp 1727399082
transform -1 0 5530 0 -1 1310
box -12 -8 32 272
use FILL  FILL82650x19650
timestamp 1727399082
transform 1 0 5510 0 1 1310
box -12 -8 32 272
use FILL  FILL82650x27450
timestamp 1727399082
transform 1 0 5510 0 1 1830
box -12 -8 32 272
use FILL  FILL82650x31350
timestamp 1727399082
transform -1 0 5530 0 -1 2350
box -12 -8 32 272
use FILL  FILL82650x35250
timestamp 1727399082
transform 1 0 5510 0 1 2350
box -12 -8 32 272
use FILL  FILL82650x50850
timestamp 1727399082
transform 1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL82650x54750
timestamp 1727399082
transform -1 0 5530 0 -1 3910
box -12 -8 32 272
use FILL  FILL82650x58650
timestamp 1727399082
transform 1 0 5510 0 1 3910
box -12 -8 32 272
use FILL  FILL82650x70350
timestamp 1727399082
transform -1 0 5530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__760_
timestamp 1727399082
transform 1 0 3530 0 1 790
box -12 -8 32 272
use FILL  FILL_0__761_
timestamp 1727399082
transform -1 0 3430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__762_
timestamp 1727399082
transform 1 0 2910 0 1 270
box -12 -8 32 272
use FILL  FILL_0__763_
timestamp 1727399082
transform -1 0 3210 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__764_
timestamp 1727399082
transform -1 0 2710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__765_
timestamp 1727399082
transform 1 0 3110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__766_
timestamp 1727399082
transform 1 0 2890 0 1 790
box -12 -8 32 272
use FILL  FILL_0__767_
timestamp 1727399082
transform -1 0 3190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__768_
timestamp 1727399082
transform 1 0 3030 0 1 270
box -12 -8 32 272
use FILL  FILL_0__769_
timestamp 1727399082
transform 1 0 4310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__770_
timestamp 1727399082
transform 1 0 4230 0 1 790
box -12 -8 32 272
use FILL  FILL_0__771_
timestamp 1727399082
transform 1 0 4190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__772_
timestamp 1727399082
transform -1 0 2670 0 1 270
box -12 -8 32 272
use FILL  FILL_0__773_
timestamp 1727399082
transform 1 0 3130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__774_
timestamp 1727399082
transform 1 0 3570 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__775_
timestamp 1727399082
transform -1 0 3290 0 1 270
box -12 -8 32 272
use FILL  FILL_0__776_
timestamp 1727399082
transform 1 0 2050 0 1 270
box -12 -8 32 272
use FILL  FILL_0__777_
timestamp 1727399082
transform -1 0 3150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__778_
timestamp 1727399082
transform 1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_0__779_
timestamp 1727399082
transform 1 0 3810 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__780_
timestamp 1727399082
transform -1 0 3690 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__781_
timestamp 1727399082
transform -1 0 1930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__782_
timestamp 1727399082
transform -1 0 2910 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__783_
timestamp 1727399082
transform 1 0 3450 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__784_
timestamp 1727399082
transform -1 0 3210 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__785_
timestamp 1727399082
transform 1 0 3310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__786_
timestamp 1727399082
transform -1 0 2410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__787_
timestamp 1727399082
transform -1 0 2270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__788_
timestamp 1727399082
transform -1 0 2390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__789_
timestamp 1727399082
transform -1 0 3010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__790_
timestamp 1727399082
transform -1 0 2790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__791_
timestamp 1727399082
transform -1 0 3230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__792_
timestamp 1727399082
transform -1 0 3370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__793_
timestamp 1727399082
transform -1 0 3010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__794_
timestamp 1727399082
transform 1 0 3350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__795_
timestamp 1727399082
transform 1 0 2690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__796_
timestamp 1727399082
transform -1 0 2810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__797_
timestamp 1727399082
transform 1 0 2190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__798_
timestamp 1727399082
transform -1 0 2230 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__799_
timestamp 1727399082
transform 1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__800_
timestamp 1727399082
transform -1 0 2990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__801_
timestamp 1727399082
transform 1 0 2870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__802_
timestamp 1727399082
transform -1 0 3110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__803_
timestamp 1727399082
transform -1 0 1130 0 1 790
box -12 -8 32 272
use FILL  FILL_0__804_
timestamp 1727399082
transform 1 0 1590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__805_
timestamp 1727399082
transform 1 0 1210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__806_
timestamp 1727399082
transform 1 0 390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__807_
timestamp 1727399082
transform 1 0 250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__808_
timestamp 1727399082
transform -1 0 270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__809_
timestamp 1727399082
transform 1 0 350 0 1 790
box -12 -8 32 272
use FILL  FILL_0__810_
timestamp 1727399082
transform 1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__811_
timestamp 1727399082
transform 1 0 430 0 1 790
box -12 -8 32 272
use FILL  FILL_0__812_
timestamp 1727399082
transform -1 0 230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__813_
timestamp 1727399082
transform 1 0 1190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__814_
timestamp 1727399082
transform 1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__815_
timestamp 1727399082
transform -1 0 2090 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__816_
timestamp 1727399082
transform 1 0 2830 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__817_
timestamp 1727399082
transform 1 0 2410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__818_
timestamp 1727399082
transform -1 0 1090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__819_
timestamp 1727399082
transform -1 0 2330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__820_
timestamp 1727399082
transform 1 0 1390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__821_
timestamp 1727399082
transform -1 0 1310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__822_
timestamp 1727399082
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__823_
timestamp 1727399082
transform 1 0 1170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__824_
timestamp 1727399082
transform -1 0 1810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__825_
timestamp 1727399082
transform 1 0 2390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__826_
timestamp 1727399082
transform -1 0 2150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__827_
timestamp 1727399082
transform -1 0 3610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__828_
timestamp 1727399082
transform -1 0 3350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__829_
timestamp 1727399082
transform -1 0 3470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__830_
timestamp 1727399082
transform 1 0 4750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__831_
timestamp 1727399082
transform -1 0 4170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__832_
timestamp 1727399082
transform -1 0 4410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__833_
timestamp 1727399082
transform -1 0 3550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__834_
timestamp 1727399082
transform -1 0 2950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__835_
timestamp 1727399082
transform -1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__836_
timestamp 1727399082
transform -1 0 3370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__837_
timestamp 1727399082
transform 1 0 3290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__838_
timestamp 1727399082
transform -1 0 3230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__839_
timestamp 1727399082
transform 1 0 4210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__840_
timestamp 1727399082
transform -1 0 4050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__841_
timestamp 1727399082
transform -1 0 4110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__842_
timestamp 1727399082
transform -1 0 5290 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__843_
timestamp 1727399082
transform 1 0 5410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__844_
timestamp 1727399082
transform 1 0 5370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__845_
timestamp 1727399082
transform 1 0 5310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__846_
timestamp 1727399082
transform 1 0 5410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__847_
timestamp 1727399082
transform 1 0 5310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__848_
timestamp 1727399082
transform 1 0 5230 0 1 270
box -12 -8 32 272
use FILL  FILL_0__849_
timestamp 1727399082
transform -1 0 4510 0 1 270
box -12 -8 32 272
use FILL  FILL_0__850_
timestamp 1727399082
transform -1 0 5110 0 1 270
box -12 -8 32 272
use FILL  FILL_0__851_
timestamp 1727399082
transform -1 0 870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__852_
timestamp 1727399082
transform -1 0 1110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__853_
timestamp 1727399082
transform 1 0 970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__854_
timestamp 1727399082
transform 1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__855_
timestamp 1727399082
transform 1 0 1170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__856_
timestamp 1727399082
transform 1 0 1370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__857_
timestamp 1727399082
transform -1 0 1090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__858_
timestamp 1727399082
transform 1 0 750 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__859_
timestamp 1727399082
transform 1 0 1650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__860_
timestamp 1727399082
transform 1 0 3210 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__861_
timestamp 1727399082
transform -1 0 1290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__862_
timestamp 1727399082
transform -1 0 870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__863_
timestamp 1727399082
transform 1 0 590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__864_
timestamp 1727399082
transform -1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__865_
timestamp 1727399082
transform 1 0 1250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__866_
timestamp 1727399082
transform 1 0 1150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__867_
timestamp 1727399082
transform 1 0 1150 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__868_
timestamp 1727399082
transform 1 0 1490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__869_
timestamp 1727399082
transform -1 0 970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__870_
timestamp 1727399082
transform -1 0 870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__871_
timestamp 1727399082
transform -1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__872_
timestamp 1727399082
transform -1 0 1290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__873_
timestamp 1727399082
transform -1 0 950 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__874_
timestamp 1727399082
transform -1 0 630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__875_
timestamp 1727399082
transform -1 0 630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__876_
timestamp 1727399082
transform -1 0 410 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__877_
timestamp 1727399082
transform -1 0 490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__878_
timestamp 1727399082
transform -1 0 310 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__879_
timestamp 1727399082
transform -1 0 310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__880_
timestamp 1727399082
transform 1 0 330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__881_
timestamp 1727399082
transform -1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__882_
timestamp 1727399082
transform 1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__883_
timestamp 1727399082
transform -1 0 750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__884_
timestamp 1727399082
transform 1 0 1290 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__885_
timestamp 1727399082
transform -1 0 890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__886_
timestamp 1727399082
transform -1 0 1050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__887_
timestamp 1727399082
transform 1 0 1150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__888_
timestamp 1727399082
transform 1 0 770 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__889_
timestamp 1727399082
transform 1 0 930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__890_
timestamp 1727399082
transform -1 0 770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__891_
timestamp 1727399082
transform -1 0 910 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__892_
timestamp 1727399082
transform 1 0 850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__893_
timestamp 1727399082
transform -1 0 590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__894_
timestamp 1727399082
transform -1 0 530 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__895_
timestamp 1727399082
transform -1 0 1050 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__896_
timestamp 1727399082
transform -1 0 730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__897_
timestamp 1727399082
transform 1 0 1310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__898_
timestamp 1727399082
transform -1 0 1170 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__899_
timestamp 1727399082
transform -1 0 1910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__900_
timestamp 1727399082
transform -1 0 3230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__901_
timestamp 1727399082
transform -1 0 1790 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__902_
timestamp 1727399082
transform -1 0 1030 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__903_
timestamp 1727399082
transform 1 0 790 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__904_
timestamp 1727399082
transform -1 0 410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__905_
timestamp 1727399082
transform -1 0 370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__906_
timestamp 1727399082
transform -1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__907_
timestamp 1727399082
transform -1 0 670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__908_
timestamp 1727399082
transform -1 0 250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__909_
timestamp 1727399082
transform -1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__910_
timestamp 1727399082
transform -1 0 170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__911_
timestamp 1727399082
transform -1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__912_
timestamp 1727399082
transform -1 0 30 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__913_
timestamp 1727399082
transform 1 0 1650 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__914_
timestamp 1727399082
transform -1 0 130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__915_
timestamp 1727399082
transform 1 0 130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__916_
timestamp 1727399082
transform -1 0 270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__917_
timestamp 1727399082
transform -1 0 650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__918_
timestamp 1727399082
transform -1 0 850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__919_
timestamp 1727399082
transform 1 0 770 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__920_
timestamp 1727399082
transform 1 0 1010 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__921_
timestamp 1727399082
transform 1 0 650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1727399082
transform -1 0 1010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1727399082
transform -1 0 650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1727399082
transform 1 0 630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1727399082
transform -1 0 1110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1727399082
transform -1 0 890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1727399082
transform 1 0 890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1727399082
transform -1 0 490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1727399082
transform -1 0 470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1727399082
transform -1 0 370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1727399082
transform -1 0 510 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1727399082
transform -1 0 270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1727399082
transform 1 0 1470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1727399082
transform 1 0 1730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1727399082
transform 1 0 1750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1727399082
transform 1 0 1650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1727399082
transform 1 0 1410 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1727399082
transform -1 0 390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1727399082
transform -1 0 150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1727399082
transform -1 0 630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1727399082
transform -1 0 310 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1727399082
transform 1 0 150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1727399082
transform 1 0 230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1727399082
transform -1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1727399082
transform -1 0 130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1727399082
transform -1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1727399082
transform -1 0 150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1727399082
transform 1 0 10 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1727399082
transform -1 0 230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1727399082
transform 1 0 350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1727399082
transform -1 0 870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1727399082
transform -1 0 1230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1727399082
transform 1 0 830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1727399082
transform -1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1727399082
transform -1 0 390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1727399082
transform -1 0 270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1727399082
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1727399082
transform 1 0 2370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1727399082
transform -1 0 1770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1727399082
transform 1 0 1090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1727399082
transform -1 0 1610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1727399082
transform 1 0 1810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1727399082
transform -1 0 1890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1727399082
transform 1 0 1630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1727399082
transform -1 0 1550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1727399082
transform -1 0 1250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1727399082
transform 1 0 1330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1727399082
transform 1 0 1390 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1727399082
transform 1 0 870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1727399082
transform -1 0 530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1727399082
transform 1 0 830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1727399082
transform -1 0 1190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1727399082
transform 1 0 730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1727399082
transform -1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1727399082
transform -1 0 490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1727399082
transform 1 0 470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1727399082
transform -1 0 270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1727399082
transform 1 0 710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1727399082
transform -1 0 1470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1727399082
transform -1 0 150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1727399082
transform -1 0 450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1727399082
transform -1 0 750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1727399082
transform -1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1727399082
transform -1 0 350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1727399082
transform 1 0 210 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1727399082
transform -1 0 310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1727399082
transform -1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1727399082
transform 1 0 590 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1727399082
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1727399082
transform -1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1727399082
transform -1 0 150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1727399082
transform 1 0 510 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1727399082
transform -1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1727399082
transform -1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1727399082
transform -1 0 130 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1727399082
transform 1 0 130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1727399082
transform -1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1727399082
transform 1 0 270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1727399082
transform 1 0 510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1727399082
transform 1 0 470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1727399082
transform 1 0 570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1727399082
transform -1 0 370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1727399082
transform -1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1727399082
transform -1 0 730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1727399082
transform -1 0 750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1727399082
transform -1 0 1530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1727399082
transform 1 0 250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1727399082
transform 1 0 370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1727399082
transform -1 0 1730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1727399082
transform -1 0 1610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1727399082
transform 1 0 1630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1727399082
transform 1 0 130 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1727399082
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1727399082
transform 1 0 2290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1727399082
transform -1 0 2630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1727399082
transform 1 0 2490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1727399082
transform 1 0 1970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1727399082
transform -1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1727399082
transform -1 0 2270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1727399082
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1727399082
transform 1 0 2150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1727399082
transform -1 0 1850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1727399082
transform 1 0 2070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1727399082
transform 1 0 2250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1727399082
transform -1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1727399082
transform 1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1727399082
transform -1 0 2230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1727399082
transform -1 0 3330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1727399082
transform 1 0 2590 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1727399082
transform -1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1727399082
transform -1 0 2890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1727399082
transform -1 0 2470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1727399082
transform 1 0 2750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1727399082
transform 1 0 3170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1727399082
transform 1 0 2990 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1727399082
transform 1 0 2730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1727399082
transform -1 0 2650 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1727399082
transform -1 0 1330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1727399082
transform 1 0 930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1727399082
transform -1 0 830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1727399082
transform -1 0 2510 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1727399082
transform -1 0 2350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1727399082
transform -1 0 1370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1727399082
transform 1 0 1230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1727399082
transform -1 0 2130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1727399082
transform 1 0 1590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1727399082
transform -1 0 1510 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1727399082
transform -1 0 1630 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1727399082
transform -1 0 1350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1727399082
transform 1 0 570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1727399082
transform -1 0 730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1727399082
transform -1 0 1770 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1727399082
transform -1 0 1110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1727399082
transform 1 0 1210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1727399082
transform -1 0 1130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1727399082
transform 1 0 1450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1727399082
transform -1 0 1090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1727399082
transform -1 0 1530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1727399082
transform -1 0 990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1727399082
transform 1 0 410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1727399082
transform 1 0 490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1727399082
transform -1 0 1390 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1727399082
transform 1 0 1250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1727399082
transform -1 0 1330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1727399082
transform 1 0 1730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1727399082
transform 1 0 1410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1727399082
transform 1 0 1530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1727399082
transform -1 0 1250 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1727399082
transform -1 0 1390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1727399082
transform 1 0 1590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1727399082
transform 1 0 1990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1727399082
transform 1 0 1570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1727399082
transform 1 0 1690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1727399082
transform -1 0 2130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1727399082
transform 1 0 1450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1727399082
transform 1 0 1730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1727399082
transform -1 0 2490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1727399082
transform -1 0 3110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1727399082
transform 1 0 2750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1727399082
transform -1 0 2510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1727399082
transform -1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1727399082
transform 1 0 2670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1727399082
transform -1 0 2590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1727399082
transform 1 0 2870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1727399082
transform -1 0 3250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1727399082
transform 1 0 2970 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1727399082
transform -1 0 2830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1727399082
transform -1 0 2810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1727399082
transform -1 0 2850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1727399082
transform 1 0 4190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1727399082
transform 1 0 3430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1727399082
transform 1 0 3390 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1727399082
transform 1 0 3470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1727399082
transform 1 0 3450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1727399082
transform -1 0 4070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1727399082
transform -1 0 3610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1727399082
transform -1 0 3570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1727399082
transform 1 0 3830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1727399082
transform -1 0 3930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1727399082
transform -1 0 3230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1727399082
transform -1 0 3030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1727399082
transform 1 0 3090 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1727399082
transform 1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1727399082
transform -1 0 3350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1727399082
transform 1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1727399082
transform -1 0 2510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1727399082
transform -1 0 2910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1727399082
transform 1 0 3510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1727399082
transform -1 0 3270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1727399082
transform -1 0 2790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1727399082
transform 1 0 2370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1727399082
transform 1 0 1870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1727399082
transform 1 0 1890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1727399082
transform -1 0 2930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1727399082
transform -1 0 2650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1727399082
transform -1 0 2130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1727399082
transform -1 0 2390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1727399082
transform -1 0 2430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1727399082
transform -1 0 2290 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1727399082
transform -1 0 1990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1727399082
transform -1 0 2170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1727399082
transform -1 0 1850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1727399082
transform -1 0 2050 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1727399082
transform -1 0 2530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1727399082
transform 1 0 1730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1727399082
transform 1 0 1870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1727399082
transform -1 0 1870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1727399082
transform 1 0 1610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1727399082
transform 1 0 1970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1727399082
transform 1 0 1990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1727399082
transform 1 0 1970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1727399082
transform 1 0 1990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1727399082
transform 1 0 1870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1727399082
transform -1 0 1750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1727399082
transform -1 0 1550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1727399082
transform -1 0 3770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1727399082
transform -1 0 1910 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1727399082
transform 1 0 2090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1727399082
transform 1 0 2130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1727399082
transform -1 0 2250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1727399082
transform 1 0 2650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1727399082
transform 1 0 2950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1727399082
transform -1 0 4710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1727399082
transform 1 0 3170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1727399082
transform 1 0 3030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1727399082
transform -1 0 3870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1727399082
transform 1 0 3530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1727399082
transform 1 0 3690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1727399082
transform 1 0 3710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1727399082
transform -1 0 3070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1727399082
transform 1 0 3310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1727399082
transform 1 0 3770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1727399082
transform -1 0 2770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1727399082
transform 1 0 3350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1727399082
transform -1 0 3410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1727399082
transform 1 0 3850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1727399082
transform 1 0 3710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1727399082
transform 1 0 3910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1727399082
transform 1 0 3690 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1727399082
transform 1 0 3910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1727399082
transform -1 0 3550 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1727399082
transform -1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1727399082
transform 1 0 3890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1727399082
transform -1 0 4250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1727399082
transform -1 0 3730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1727399082
transform -1 0 4050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1727399082
transform -1 0 3990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1727399082
transform 1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1727399082
transform 1 0 4710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1727399082
transform 1 0 4090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1727399082
transform -1 0 4150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1727399082
transform -1 0 4270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1727399082
transform -1 0 4450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1727399082
transform 1 0 4790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1727399082
transform 1 0 5150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1727399082
transform 1 0 3650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1727399082
transform 1 0 3770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1727399082
transform -1 0 4690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1727399082
transform 1 0 4550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1727399082
transform 1 0 5010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1727399082
transform -1 0 5310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1727399082
transform -1 0 5130 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1727399082
transform 1 0 4890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1727399082
transform -1 0 4890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1727399082
transform 1 0 5010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1727399082
transform 1 0 4790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1727399082
transform 1 0 4830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1727399082
transform 1 0 5410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1727399082
transform 1 0 4970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1727399082
transform -1 0 5110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1727399082
transform 1 0 5170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1727399082
transform -1 0 4970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1727399082
transform -1 0 4830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1727399082
transform -1 0 4690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1727399082
transform 1 0 4510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1727399082
transform 1 0 5170 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1727399082
transform -1 0 4250 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1727399082
transform 1 0 5030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1727399082
transform 1 0 5050 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1727399082
transform 1 0 5250 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1727399082
transform 1 0 5390 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1727399082
transform 1 0 3650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1727399082
transform -1 0 4730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1727399082
transform 1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1727399082
transform -1 0 4590 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1727399082
transform 1 0 3710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1727399082
transform -1 0 3590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1727399082
transform 1 0 3810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1727399082
transform 1 0 3930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1727399082
transform -1 0 2870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1727399082
transform 1 0 3810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1727399082
transform -1 0 3110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1727399082
transform -1 0 3470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1727399082
transform -1 0 3590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1727399082
transform 1 0 4230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1727399082
transform 1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1727399082
transform 1 0 4010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1727399082
transform 1 0 4150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1727399082
transform 1 0 4150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1727399082
transform -1 0 4270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1727399082
transform 1 0 4350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1727399082
transform 1 0 4470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1727399082
transform 1 0 4290 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1727399082
transform -1 0 4370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1727399082
transform 1 0 4590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1727399082
transform 1 0 4810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1727399082
transform 1 0 4370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1727399082
transform 1 0 4450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1727399082
transform 1 0 4490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1727399082
transform 1 0 5410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1727399082
transform 1 0 4630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1727399082
transform 1 0 4770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1727399082
transform 1 0 4890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1727399082
transform -1 0 5070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1727399082
transform 1 0 4770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1727399082
transform -1 0 4670 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1727399082
transform -1 0 4850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1727399082
transform -1 0 3750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1727399082
transform -1 0 5310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1727399082
transform 1 0 5150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1727399082
transform -1 0 5410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1727399082
transform -1 0 5310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1727399082
transform -1 0 5210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1727399082
transform 1 0 5150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1727399082
transform 1 0 5010 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1727399082
transform -1 0 5310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1727399082
transform 1 0 4330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1727399082
transform -1 0 4850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1727399082
transform -1 0 4050 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1727399082
transform -1 0 3950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1727399082
transform -1 0 3610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1727399082
transform 1 0 3210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1727399082
transform 1 0 4030 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1727399082
transform -1 0 3870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1727399082
transform 1 0 3990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1727399082
transform 1 0 3710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1727399082
transform 1 0 4230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1727399082
transform 1 0 4410 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1727399082
transform 1 0 4550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1727399082
transform -1 0 5070 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1727399082
transform -1 0 4930 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1727399082
transform 1 0 5130 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1727399082
transform 1 0 5210 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1727399082
transform -1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1727399082
transform 1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1727399082
transform 1 0 5390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1727399082
transform 1 0 5150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1727399082
transform 1 0 4950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1727399082
transform -1 0 1850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1727399082
transform -1 0 4970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1727399082
transform 1 0 3590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1727399082
transform -1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1727399082
transform 1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1727399082
transform -1 0 4610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1727399082
transform 1 0 3770 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1727399082
transform -1 0 4850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1727399082
transform -1 0 4710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1727399082
transform 1 0 4110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1727399082
transform 1 0 4130 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1727399082
transform 1 0 3490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1727399082
transform -1 0 3930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1727399082
transform 1 0 4270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1727399082
transform 1 0 4530 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1727399082
transform -1 0 4430 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1727399082
transform 1 0 4590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1727399082
transform -1 0 4710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1727399082
transform 1 0 4810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1727399082
transform 1 0 5350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1727399082
transform 1 0 5430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1727399082
transform -1 0 5330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1727399082
transform 1 0 5070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1727399082
transform -1 0 5230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1727399082
transform 1 0 5270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1727399082
transform 1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1727399082
transform -1 0 4350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1727399082
transform -1 0 5270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1727399082
transform -1 0 4810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1727399082
transform -1 0 4950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1727399082
transform 1 0 5250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1727399082
transform 1 0 5130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1727399082
transform 1 0 4890 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1727399082
transform -1 0 4670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1727399082
transform -1 0 4270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1727399082
transform 1 0 4130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1727399082
transform -1 0 4050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1727399082
transform 1 0 4350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1727399082
transform 1 0 4490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1727399082
transform 1 0 4390 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1727399082
transform -1 0 4310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1727399082
transform -1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1727399082
transform -1 0 4210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1727399082
transform 1 0 5310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1727399082
transform 1 0 4610 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1727399082
transform 1 0 4730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1727399082
transform 1 0 4470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1727399082
transform 1 0 4830 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1727399082
transform -1 0 4930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1727399082
transform -1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1727399082
transform 1 0 950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1727399082
transform -1 0 1030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1727399082
transform -1 0 1070 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1727399082
transform 1 0 2730 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1727399082
transform 1 0 2350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1727399082
transform -1 0 430 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1727399082
transform -1 0 190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1727399082
transform -1 0 570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1727399082
transform -1 0 830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1727399082
transform 1 0 670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1727399082
transform 1 0 710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1727399082
transform 1 0 1350 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1727399082
transform 1 0 990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1727399082
transform 1 0 590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1727399082
transform -1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1727399082
transform -1 0 270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1727399082
transform 1 0 130 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1727399082
transform 1 0 510 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1727399082
transform 1 0 370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1727399082
transform 1 0 610 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1727399082
transform 1 0 870 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1727399082
transform -1 0 830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1727399082
transform -1 0 270 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1727399082
transform -1 0 110 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1727399082
transform -1 0 330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1727399082
transform 1 0 410 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1727399082
transform 1 0 870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1727399082
transform -1 0 670 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1727399082
transform 1 0 550 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1727399082
transform 1 0 950 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1727399082
transform -1 0 1090 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1727399082
transform 1 0 1710 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1727399082
transform 1 0 1290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1727399082
transform -1 0 2570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1727399082
transform -1 0 1970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1727399082
transform -1 0 1750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1727399082
transform 1 0 750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1727399082
transform 1 0 2270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1727399082
transform 1 0 2150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1727399082
transform 1 0 2030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1727399082
transform 1 0 2190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1727399082
transform 1 0 2290 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1727399082
transform 1 0 2410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1727399082
transform -1 0 2350 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1727399082
transform -1 0 2070 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1727399082
transform -1 0 890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1727399082
transform 1 0 1070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1727399082
transform 1 0 970 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1727399082
transform -1 0 1870 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1727399082
transform 1 0 1990 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1727399082
transform 1 0 2090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1727399082
transform -1 0 2210 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1727399082
transform 1 0 1650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1727399082
transform -1 0 1330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1727399082
transform 1 0 1190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1727399082
transform -1 0 1910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1727399082
transform -1 0 1450 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1727399082
transform 1 0 1610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1727399082
transform 1 0 1390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1727399082
transform 1 0 1730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1727399082
transform -1 0 1510 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1727399082
transform 1 0 1410 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1727399082
transform -1 0 1370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1727399082
transform 1 0 1530 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1727399082
transform 1 0 1830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1727399082
transform 1 0 1750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1727399082
transform -1 0 1870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1727399082
transform -1 0 1690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1727399082
transform 1 0 1930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1727399082
transform 1 0 1910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1727399082
transform 1 0 1690 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1727399082
transform 1 0 1790 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1727399082
transform 1 0 1930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1727399082
transform -1 0 1830 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1727399082
transform -1 0 3330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1727399082
transform 1 0 2170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1727399082
transform 1 0 2030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1727399082
transform 1 0 1550 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1727399082
transform 1 0 1810 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1727399082
transform 1 0 1670 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1727399082
transform 1 0 1950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1727399082
transform 1 0 3790 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1727399082
transform 1 0 3650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1727399082
transform 1 0 3910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1727399082
transform 1 0 3970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1727399082
transform 1 0 3670 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1727399082
transform -1 0 3590 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1727399082
transform -1 0 3470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1727399082
transform -1 0 3450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1727399082
transform 1 0 4190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1727399082
transform 1 0 5050 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1727399082
transform 1 0 4690 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1727399082
transform -1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1727399082
transform -1 0 4470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1727399082
transform -1 0 4590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1727399082
transform -1 0 4330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1727399082
transform 1 0 4370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1727399082
transform 1 0 3670 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1727399082
transform 1 0 4430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1727399082
transform -1 0 4930 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1727399082
transform 1 0 4790 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1727399082
transform 1 0 4650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1727399082
transform 1 0 3830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1727399082
transform 1 0 3630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1727399082
transform 1 0 4070 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1727399082
transform 1 0 4150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1727399082
transform -1 0 3970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1727399082
transform 1 0 4090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1727399082
transform -1 0 3830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1727399082
transform -1 0 3950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1727399082
transform -1 0 4050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1727399082
transform 1 0 3330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1727399082
transform 1 0 3230 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1727399082
transform -1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1727399082
transform 1 0 3690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1727399082
transform 1 0 4230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1727399082
transform -1 0 4010 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1727399082
transform -1 0 3890 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1727399082
transform 1 0 3790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1727399082
transform 1 0 4590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1727399082
transform 1 0 3790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1727399082
transform 1 0 4330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1727399082
transform 1 0 4910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1727399082
transform 1 0 4790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1727399082
transform 1 0 4550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1727399082
transform -1 0 4510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1727399082
transform 1 0 4710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1727399082
transform 1 0 4390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1727399082
transform 1 0 4290 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1727399082
transform 1 0 4610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1727399082
transform 1 0 4730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1727399082
transform -1 0 4630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1727399082
transform 1 0 4850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1452_
timestamp 1727399082
transform -1 0 4850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1453_
timestamp 1727399082
transform -1 0 4710 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1454_
timestamp 1727399082
transform 1 0 4610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1455_
timestamp 1727399082
transform 1 0 4390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1456_
timestamp 1727399082
transform -1 0 4510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1457_
timestamp 1727399082
transform 1 0 5330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1458_
timestamp 1727399082
transform -1 0 5170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1459_
timestamp 1727399082
transform 1 0 5230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1460_
timestamp 1727399082
transform 1 0 5270 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1461_
timestamp 1727399082
transform 1 0 4950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1462_
timestamp 1727399082
transform -1 0 4830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1463_
timestamp 1727399082
transform 1 0 4670 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1464_
timestamp 1727399082
transform -1 0 4290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1465_
timestamp 1727399082
transform -1 0 5170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1466_
timestamp 1727399082
transform 1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1467_
timestamp 1727399082
transform 1 0 5310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1468_
timestamp 1727399082
transform -1 0 5110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1469_
timestamp 1727399082
transform -1 0 4770 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1470_
timestamp 1727399082
transform -1 0 4970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1471_
timestamp 1727399082
transform 1 0 4950 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1472_
timestamp 1727399082
transform -1 0 4730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1473_
timestamp 1727399082
transform -1 0 4650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1474_
timestamp 1727399082
transform 1 0 4150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1475_
timestamp 1727399082
transform -1 0 4890 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1476_
timestamp 1727399082
transform 1 0 4950 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1477_
timestamp 1727399082
transform 1 0 4850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1478_
timestamp 1727399082
transform -1 0 4110 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1479_
timestamp 1727399082
transform 1 0 4130 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1480_
timestamp 1727399082
transform 1 0 3310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1481_
timestamp 1727399082
transform 1 0 3850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1482_
timestamp 1727399082
transform -1 0 3750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1483_
timestamp 1727399082
transform 1 0 5370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1484_
timestamp 1727399082
transform -1 0 5290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1485_
timestamp 1727399082
transform 1 0 5370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1486_
timestamp 1727399082
transform 1 0 4610 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1487_
timestamp 1727399082
transform -1 0 5190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1488_
timestamp 1727399082
transform 1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1489_
timestamp 1727399082
transform -1 0 3510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1490_
timestamp 1727399082
transform 1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1491_
timestamp 1727399082
transform 1 0 3950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1492_
timestamp 1727399082
transform -1 0 3090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1493_
timestamp 1727399082
transform 1 0 3090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1494_
timestamp 1727399082
transform -1 0 2990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1495_
timestamp 1727399082
transform -1 0 3230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1496_
timestamp 1727399082
transform 1 0 3050 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1497_
timestamp 1727399082
transform 1 0 2930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1498_
timestamp 1727399082
transform -1 0 2830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1499_
timestamp 1727399082
transform -1 0 3410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1500_
timestamp 1727399082
transform 1 0 3510 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1501_
timestamp 1727399082
transform 1 0 2870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1502_
timestamp 1727399082
transform -1 0 2990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1503_
timestamp 1727399082
transform 1 0 2930 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1504_
timestamp 1727399082
transform -1 0 2630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1505_
timestamp 1727399082
transform -1 0 2770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1506_
timestamp 1727399082
transform -1 0 2570 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1507_
timestamp 1727399082
transform 1 0 2430 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1508_
timestamp 1727399082
transform 1 0 2550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1509_
timestamp 1727399082
transform -1 0 2710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1510_
timestamp 1727399082
transform -1 0 2630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1511_
timestamp 1727399082
transform -1 0 2730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1512_
timestamp 1727399082
transform -1 0 1890 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1513_
timestamp 1727399082
transform -1 0 2230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1514_
timestamp 1727399082
transform -1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1515_
timestamp 1727399082
transform -1 0 630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1516_
timestamp 1727399082
transform -1 0 2070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1517_
timestamp 1727399082
transform -1 0 2430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1518_
timestamp 1727399082
transform 1 0 2110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1519_
timestamp 1727399082
transform 1 0 1990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1520_
timestamp 1727399082
transform 1 0 1950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1521_
timestamp 1727399082
transform 1 0 2070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1522_
timestamp 1727399082
transform -1 0 2370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1523_
timestamp 1727399082
transform 1 0 2470 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1524_
timestamp 1727399082
transform -1 0 2690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1525_
timestamp 1727399082
transform 1 0 2530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1601_
timestamp 1727399082
transform 1 0 5410 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1602_
timestamp 1727399082
transform 1 0 5410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1603_
timestamp 1727399082
transform 1 0 5230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1604_
timestamp 1727399082
transform 1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1605_
timestamp 1727399082
transform 1 0 4470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1606_
timestamp 1727399082
transform 1 0 3390 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1607_
timestamp 1727399082
transform 1 0 3270 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1608_
timestamp 1727399082
transform -1 0 3050 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1609_
timestamp 1727399082
transform -1 0 2790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1727399082
transform -1 0 3050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1727399082
transform 1 0 4210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1727399082
transform 1 0 4270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1727399082
transform 1 0 3630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1727399082
transform -1 0 770 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1727399082
transform -1 0 2290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1727399082
transform -1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1727399082
transform -1 0 1110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1727399082
transform -1 0 2250 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1727399082
transform -1 0 1770 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1727399082
transform 1 0 4370 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1727399082
transform 1 0 3050 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1727399082
transform 1 0 4330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1727399082
transform -1 0 1070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1727399082
transform -1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1727399082
transform -1 0 990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1727399082
transform -1 0 1570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1727399082
transform 1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1727399082
transform -1 0 2810 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1727399082
transform 1 0 2490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1727399082
transform 1 0 2830 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1727399082
transform 1 0 2790 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1727399082
transform -1 0 970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1727399082
transform 1 0 3110 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1727399082
transform -1 0 1210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1727399082
transform -1 0 4330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1727399082
transform -1 0 2870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1727399082
transform 1 0 3910 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1727399082
transform -1 0 2490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1727399082
transform 1 0 3070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1727399082
transform 1 0 3890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert13
timestamp 1727399082
transform 1 0 2350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert14
timestamp 1727399082
transform -1 0 1530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert15
timestamp 1727399082
transform -1 0 1670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__761_
timestamp 1727399082
transform -1 0 3450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__762_
timestamp 1727399082
transform 1 0 2930 0 1 270
box -12 -8 32 272
use FILL  FILL_1__764_
timestamp 1727399082
transform -1 0 2730 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__766_
timestamp 1727399082
transform 1 0 2910 0 1 790
box -12 -8 32 272
use FILL  FILL_1__768_
timestamp 1727399082
transform 1 0 3050 0 1 270
box -12 -8 32 272
use FILL  FILL_1__770_
timestamp 1727399082
transform 1 0 4250 0 1 790
box -12 -8 32 272
use FILL  FILL_1__771_
timestamp 1727399082
transform 1 0 4210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__773_
timestamp 1727399082
transform 1 0 3150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__775_
timestamp 1727399082
transform -1 0 3310 0 1 270
box -12 -8 32 272
use FILL  FILL_1__777_
timestamp 1727399082
transform -1 0 3170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__778_
timestamp 1727399082
transform 1 0 3770 0 1 270
box -12 -8 32 272
use FILL  FILL_1__780_
timestamp 1727399082
transform -1 0 3710 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__782_
timestamp 1727399082
transform -1 0 2930 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__784_
timestamp 1727399082
transform -1 0 3230 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__785_
timestamp 1727399082
transform 1 0 3330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__787_
timestamp 1727399082
transform -1 0 2290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__789_
timestamp 1727399082
transform -1 0 3030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__791_
timestamp 1727399082
transform -1 0 3250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__792_
timestamp 1727399082
transform -1 0 3390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__794_
timestamp 1727399082
transform 1 0 3370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__796_
timestamp 1727399082
transform -1 0 2830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__798_
timestamp 1727399082
transform -1 0 2250 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__799_
timestamp 1727399082
transform 1 0 2870 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__801_
timestamp 1727399082
transform 1 0 2890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__803_
timestamp 1727399082
transform -1 0 1150 0 1 790
box -12 -8 32 272
use FILL  FILL_1__805_
timestamp 1727399082
transform 1 0 1230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__806_
timestamp 1727399082
transform 1 0 410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__808_
timestamp 1727399082
transform -1 0 290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__810_
timestamp 1727399082
transform 1 0 490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__812_
timestamp 1727399082
transform -1 0 250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__814_
timestamp 1727399082
transform 1 0 510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__815_
timestamp 1727399082
transform -1 0 2110 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__817_
timestamp 1727399082
transform 1 0 2430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__819_
timestamp 1727399082
transform -1 0 2350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__821_
timestamp 1727399082
transform -1 0 1330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__822_
timestamp 1727399082
transform 1 0 2270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__824_
timestamp 1727399082
transform -1 0 1830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__826_
timestamp 1727399082
transform -1 0 2170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__828_
timestamp 1727399082
transform -1 0 3370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__829_
timestamp 1727399082
transform -1 0 3490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__831_
timestamp 1727399082
transform -1 0 4190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__833_
timestamp 1727399082
transform -1 0 3570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__835_
timestamp 1727399082
transform -1 0 3190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__836_
timestamp 1727399082
transform -1 0 3390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__838_
timestamp 1727399082
transform -1 0 3250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__840_
timestamp 1727399082
transform -1 0 4070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__842_
timestamp 1727399082
transform -1 0 5310 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__843_
timestamp 1727399082
transform 1 0 5430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__845_
timestamp 1727399082
transform 1 0 5330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__847_
timestamp 1727399082
transform 1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__849_
timestamp 1727399082
transform -1 0 4530 0 1 270
box -12 -8 32 272
use FILL  FILL_1__850_
timestamp 1727399082
transform -1 0 5130 0 1 270
box -12 -8 32 272
use FILL  FILL_1__852_
timestamp 1727399082
transform -1 0 1130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__854_
timestamp 1727399082
transform 1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__856_
timestamp 1727399082
transform 1 0 1390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__858_
timestamp 1727399082
transform 1 0 770 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__859_
timestamp 1727399082
transform 1 0 1670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__861_
timestamp 1727399082
transform -1 0 1310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__863_
timestamp 1727399082
transform 1 0 610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__865_
timestamp 1727399082
transform 1 0 1270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__866_
timestamp 1727399082
transform 1 0 1170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__868_
timestamp 1727399082
transform 1 0 1510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__870_
timestamp 1727399082
transform -1 0 890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__872_
timestamp 1727399082
transform -1 0 1310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__873_
timestamp 1727399082
transform -1 0 970 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__875_
timestamp 1727399082
transform -1 0 650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__877_
timestamp 1727399082
transform -1 0 510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__879_
timestamp 1727399082
transform -1 0 330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__880_
timestamp 1727399082
transform 1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__882_
timestamp 1727399082
transform 1 0 1430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__884_
timestamp 1727399082
transform 1 0 1310 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__886_
timestamp 1727399082
transform -1 0 1070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__887_
timestamp 1727399082
transform 1 0 1170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__889_
timestamp 1727399082
transform 1 0 950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__891_
timestamp 1727399082
transform -1 0 930 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__893_
timestamp 1727399082
transform -1 0 610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__894_
timestamp 1727399082
transform -1 0 550 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__896_
timestamp 1727399082
transform -1 0 750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__898_
timestamp 1727399082
transform -1 0 1190 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__900_
timestamp 1727399082
transform -1 0 3250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__902_
timestamp 1727399082
transform -1 0 1050 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__903_
timestamp 1727399082
transform 1 0 810 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__905_
timestamp 1727399082
transform -1 0 390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__907_
timestamp 1727399082
transform -1 0 690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__909_
timestamp 1727399082
transform -1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__910_
timestamp 1727399082
transform -1 0 190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__912_
timestamp 1727399082
transform -1 0 50 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__914_
timestamp 1727399082
transform -1 0 150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__916_
timestamp 1727399082
transform -1 0 290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__917_
timestamp 1727399082
transform -1 0 670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__919_
timestamp 1727399082
transform 1 0 790 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__921_
timestamp 1727399082
transform 1 0 670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1727399082
transform -1 0 670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1727399082
transform 1 0 650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1727399082
transform -1 0 910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1727399082
transform -1 0 510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1727399082
transform -1 0 390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1727399082
transform -1 0 530 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1727399082
transform 1 0 1490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1727399082
transform 1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1727399082
transform 1 0 1430 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1727399082
transform -1 0 410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1727399082
transform -1 0 650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1727399082
transform 1 0 170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1727399082
transform -1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1727399082
transform -1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1727399082
transform -1 0 170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1727399082
transform -1 0 250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1727399082
transform -1 0 890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1727399082
transform 1 0 850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1727399082
transform -1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1727399082
transform -1 0 290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1727399082
transform 1 0 2390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1727399082
transform 1 0 1110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1727399082
transform -1 0 1630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1727399082
transform -1 0 1910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1727399082
transform -1 0 1570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1727399082
transform 1 0 1350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1727399082
transform 1 0 1410 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1727399082
transform -1 0 550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1727399082
transform -1 0 1210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1727399082
transform -1 0 970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1727399082
transform -1 0 510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1727399082
transform -1 0 290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1727399082
transform -1 0 1490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1727399082
transform -1 0 470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1727399082
transform -1 0 770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1727399082
transform -1 0 370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1727399082
transform -1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1727399082
transform 1 0 610 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1727399082
transform -1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1727399082
transform -1 0 170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1727399082
transform -1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1727399082
transform -1 0 150 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1727399082
transform -1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1727399082
transform 1 0 290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1727399082
transform 1 0 590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1727399082
transform -1 0 390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1727399082
transform -1 0 750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1727399082
transform -1 0 1550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1727399082
transform 1 0 390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1727399082
transform -1 0 1750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1727399082
transform 1 0 1650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1727399082
transform 1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1727399082
transform -1 0 2650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1727399082
transform 1 0 1990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1727399082
transform -1 0 2150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1727399082
transform -1 0 2230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1727399082
transform -1 0 1870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1727399082
transform 1 0 2270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1727399082
transform -1 0 630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1727399082
transform -1 0 2250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1727399082
transform 1 0 2610 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1727399082
transform -1 0 2910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1727399082
transform -1 0 2490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1727399082
transform 1 0 3190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1727399082
transform 1 0 2750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1727399082
transform -1 0 1350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1727399082
transform 1 0 950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1727399082
transform -1 0 2530 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1727399082
transform -1 0 1390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1727399082
transform -1 0 2150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1727399082
transform 1 0 1610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1727399082
transform -1 0 1650 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1727399082
transform 1 0 590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1727399082
transform -1 0 1790 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1727399082
transform -1 0 1130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1727399082
transform -1 0 1150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1727399082
transform -1 0 1110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1727399082
transform -1 0 1010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1727399082
transform 1 0 510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1727399082
transform -1 0 1410 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1727399082
transform -1 0 1350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1727399082
transform 1 0 1430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1727399082
transform -1 0 1270 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1727399082
transform -1 0 1410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1727399082
transform 1 0 2010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1727399082
transform 1 0 1710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1727399082
transform 1 0 1470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1727399082
transform 1 0 1750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1727399082
transform -1 0 3130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1727399082
transform -1 0 2530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1727399082
transform 1 0 2690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1727399082
transform -1 0 2610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1727399082
transform -1 0 3270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1727399082
transform -1 0 2850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1727399082
transform -1 0 2870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1727399082
transform 1 0 4210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1727399082
transform 1 0 3410 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1727399082
transform 1 0 3470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1727399082
transform -1 0 3630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1727399082
transform -1 0 3590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1727399082
transform -1 0 3950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1727399082
transform -1 0 3050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1727399082
transform 1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1727399082
transform 1 0 3390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1727399082
transform -1 0 2530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1727399082
transform 1 0 3530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1727399082
transform -1 0 2810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1727399082
transform 1 0 1890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1727399082
transform 1 0 1910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1727399082
transform -1 0 2670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1727399082
transform -1 0 2410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1727399082
transform -1 0 2310 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1727399082
transform -1 0 2010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1727399082
transform -1 0 1870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1727399082
transform -1 0 2550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1727399082
transform 1 0 1890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1727399082
transform -1 0 1890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1727399082
transform 1 0 1990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1727399082
transform 1 0 1990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1727399082
transform 1 0 1890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1727399082
transform -1 0 1770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1727399082
transform -1 0 3790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1727399082
transform 1 0 2110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1727399082
transform -1 0 2270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1727399082
transform 1 0 2670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1727399082
transform -1 0 4730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1727399082
transform 1 0 3050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1727399082
transform 1 0 3550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1727399082
transform 1 0 3730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1727399082
transform -1 0 3090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1727399082
transform 1 0 3790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1727399082
transform 1 0 3370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1727399082
transform 1 0 3870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1727399082
transform 1 0 3730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1727399082
transform 1 0 3710 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1727399082
transform -1 0 3570 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1727399082
transform 1 0 3910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1727399082
transform -1 0 4270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1727399082
transform -1 0 4070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1727399082
transform 1 0 4370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1727399082
transform 1 0 4110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1727399082
transform -1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1727399082
transform -1 0 4470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1727399082
transform 1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1727399082
transform 1 0 3790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1727399082
transform -1 0 4710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1727399082
transform 1 0 5030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1727399082
transform -1 0 5150 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1727399082
transform -1 0 4910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1727399082
transform 1 0 5030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1727399082
transform 1 0 4850 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1727399082
transform 1 0 4990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1727399082
transform 1 0 5190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1727399082
transform -1 0 4850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1727399082
transform -1 0 4710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1727399082
transform 1 0 5190 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1727399082
transform 1 0 5050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1727399082
transform 1 0 5270 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1727399082
transform 1 0 5410 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1727399082
transform -1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1727399082
transform -1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1727399082
transform -1 0 3610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1727399082
transform 1 0 3830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1727399082
transform -1 0 2890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1727399082
transform -1 0 3130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1727399082
transform -1 0 3610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1727399082
transform 1 0 4250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1727399082
transform 1 0 4030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1727399082
transform 1 0 4170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1727399082
transform 1 0 4370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1727399082
transform 1 0 4490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1727399082
transform -1 0 4390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1727399082
transform 1 0 4830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1727399082
transform 1 0 4470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1727399082
transform 1 0 4510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1727399082
transform 1 0 4650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1727399082
transform 1 0 4910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1727399082
transform 1 0 4790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1727399082
transform -1 0 4870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1727399082
transform -1 0 3770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1727399082
transform 1 0 5170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1727399082
transform -1 0 5330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1727399082
transform 1 0 5170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1727399082
transform 1 0 5030 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1727399082
transform 1 0 4350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1727399082
transform -1 0 4070 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1727399082
transform -1 0 3630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1727399082
transform 1 0 3230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1727399082
transform -1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1727399082
transform 1 0 3730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1727399082
transform 1 0 4430 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1727399082
transform 1 0 4570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1727399082
transform -1 0 4950 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1727399082
transform 1 0 5230 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1727399082
transform 1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1727399082
transform 1 0 5410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1727399082
transform 1 0 4970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1727399082
transform -1 0 4990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1727399082
transform -1 0 4890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1727399082
transform 1 0 4730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1727399082
transform 1 0 3790 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1727399082
transform -1 0 4730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1727399082
transform 1 0 4150 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1727399082
transform -1 0 3950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1727399082
transform 1 0 4290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1727399082
transform -1 0 4450 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1727399082
transform -1 0 4730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1727399082
transform 1 0 5370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1727399082
transform 1 0 5450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1727399082
transform 1 0 5090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1727399082
transform 1 0 5290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1727399082
transform -1 0 4370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1727399082
transform -1 0 5290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1727399082
transform -1 0 4970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1727399082
transform 1 0 5150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1727399082
transform -1 0 4690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1727399082
transform -1 0 4290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1727399082
transform -1 0 4070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1727399082
transform 1 0 4510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1727399082
transform -1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1727399082
transform -1 0 4190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1727399082
transform 1 0 5330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1727399082
transform 1 0 4750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1727399082
transform 1 0 4850 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1727399082
transform -1 0 4950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1727399082
transform 1 0 970 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1727399082
transform -1 0 1090 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1727399082
transform 1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1727399082
transform -1 0 210 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1727399082
transform -1 0 590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1727399082
transform 1 0 690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1727399082
transform 1 0 1370 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1727399082
transform 1 0 610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1727399082
transform -1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1727399082
transform 1 0 150 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1727399082
transform 1 0 390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1727399082
transform 1 0 890 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1727399082
transform -1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1727399082
transform -1 0 130 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1727399082
transform 1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1727399082
transform -1 0 690 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1727399082
transform 1 0 570 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1727399082
transform -1 0 1110 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1727399082
transform 1 0 1310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1727399082
transform -1 0 1990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1727399082
transform -1 0 1770 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1727399082
transform 1 0 2290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1727399082
transform 1 0 2050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1727399082
transform 1 0 2310 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1727399082
transform 1 0 2430 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1727399082
transform -1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1727399082
transform 1 0 1090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1727399082
transform -1 0 1890 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1727399082
transform 1 0 2110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1727399082
transform -1 0 2230 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1727399082
transform -1 0 1350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1727399082
transform -1 0 1930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1727399082
transform 1 0 1630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1727399082
transform 1 0 1410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1727399082
transform -1 0 1530 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1727399082
transform -1 0 1390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1727399082
transform 1 0 1850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1727399082
transform 1 0 1770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1727399082
transform -1 0 1710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1727399082
transform 1 0 1930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1727399082
transform 1 0 1810 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1727399082
transform 1 0 1950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1727399082
transform -1 0 3350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1727399082
transform 1 0 2050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1727399082
transform 1 0 1830 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1727399082
transform 1 0 1690 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1727399082
transform 1 0 3810 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1727399082
transform 1 0 3930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1727399082
transform 1 0 3690 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1727399082
transform -1 0 3610 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1727399082
transform -1 0 3470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1727399082
transform 1 0 5070 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1727399082
transform -1 0 5070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1727399082
transform -1 0 4610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1727399082
transform -1 0 4350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1727399082
transform 1 0 3690 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1727399082
transform -1 0 4950 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1727399082
transform 1 0 4670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1727399082
transform 1 0 3850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1727399082
transform 1 0 4090 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1727399082
transform -1 0 3990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1727399082
transform -1 0 3850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1727399082
transform -1 0 3970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1727399082
transform 1 0 3350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1727399082
transform -1 0 3170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1727399082
transform 1 0 4250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1727399082
transform -1 0 4030 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1727399082
transform 1 0 3810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1727399082
transform 1 0 3810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1727399082
transform 1 0 4930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1727399082
transform 1 0 4810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1727399082
transform -1 0 4530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1727399082
transform 1 0 4410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1727399082
transform 1 0 4630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1727399082
transform 1 0 4750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1727399082
transform 1 0 4870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1453_
timestamp 1727399082
transform -1 0 4730 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1455_
timestamp 1727399082
transform 1 0 4410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1457_
timestamp 1727399082
transform 1 0 5350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1458_
timestamp 1727399082
transform -1 0 5190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1460_
timestamp 1727399082
transform 1 0 5290 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1462_
timestamp 1727399082
transform -1 0 4850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1464_
timestamp 1727399082
transform -1 0 4310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1465_
timestamp 1727399082
transform -1 0 5190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1467_
timestamp 1727399082
transform 1 0 5330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1469_
timestamp 1727399082
transform -1 0 4790 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1471_
timestamp 1727399082
transform 1 0 4970 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1472_
timestamp 1727399082
transform -1 0 4750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1474_
timestamp 1727399082
transform 1 0 4170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1476_
timestamp 1727399082
transform 1 0 4970 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1478_
timestamp 1727399082
transform -1 0 4130 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1479_
timestamp 1727399082
transform 1 0 4150 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1481_
timestamp 1727399082
transform 1 0 3870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1483_
timestamp 1727399082
transform 1 0 5390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1485_
timestamp 1727399082
transform 1 0 5390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1486_
timestamp 1727399082
transform 1 0 4630 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1488_
timestamp 1727399082
transform 1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1490_
timestamp 1727399082
transform 1 0 4090 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1492_
timestamp 1727399082
transform -1 0 3110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1493_
timestamp 1727399082
transform 1 0 3110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1495_
timestamp 1727399082
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1497_
timestamp 1727399082
transform 1 0 2950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1499_
timestamp 1727399082
transform -1 0 3430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1501_
timestamp 1727399082
transform 1 0 2890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1502_
timestamp 1727399082
transform -1 0 3010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1504_
timestamp 1727399082
transform -1 0 2650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1506_
timestamp 1727399082
transform -1 0 2590 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1508_
timestamp 1727399082
transform 1 0 2570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1509_
timestamp 1727399082
transform -1 0 2730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1511_
timestamp 1727399082
transform -1 0 2750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1513_
timestamp 1727399082
transform -1 0 2250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1515_
timestamp 1727399082
transform -1 0 650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1516_
timestamp 1727399082
transform -1 0 2090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1518_
timestamp 1727399082
transform 1 0 2130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1520_
timestamp 1727399082
transform 1 0 1970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1522_
timestamp 1727399082
transform -1 0 2390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1523_
timestamp 1727399082
transform 1 0 2490 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1525_
timestamp 1727399082
transform 1 0 2550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1602_
timestamp 1727399082
transform 1 0 5430 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1604_
timestamp 1727399082
transform 1 0 5410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1605_
timestamp 1727399082
transform 1 0 4490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1607_
timestamp 1727399082
transform 1 0 3290 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1609_
timestamp 1727399082
transform -1 0 2810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1727399082
transform -1 0 3070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1727399082
transform 1 0 4290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1727399082
transform -1 0 790 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1727399082
transform -1 0 2310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1727399082
transform -1 0 1130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1727399082
transform -1 0 2270 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1727399082
transform 1 0 4390 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1727399082
transform 1 0 3070 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1727399082
transform -1 0 1090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1727399082
transform -1 0 1010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1727399082
transform 1 0 990 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1727399082
transform -1 0 2830 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1727399082
transform 1 0 2850 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1727399082
transform -1 0 990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1727399082
transform -1 0 1230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1727399082
transform -1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1727399082
transform 1 0 3930 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1727399082
transform 1 0 3090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1727399082
transform 1 0 3910 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert14
timestamp 1727399082
transform -1 0 1550 0 -1 1310
box -12 -8 32 272
<< labels >>
flabel metal1 s 5543 2 5603 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 2537 5517 2543 5523 3 FreeSans 16 90 0 0 Cin[5]
port 2 nsew
flabel metal2 s 3117 5517 3123 5523 3 FreeSans 16 90 0 0 Cin[4]
port 3 nsew
flabel metal2 s 3217 5517 3223 5523 3 FreeSans 16 90 0 0 Cin[3]
port 4 nsew
flabel metal2 s 4257 5517 4263 5523 3 FreeSans 16 90 0 0 Cin[2]
port 5 nsew
flabel metal2 s 4377 5517 4383 5523 3 FreeSans 16 90 0 0 Cin[1]
port 6 nsew
flabel metal2 s 4417 5517 4423 5523 3 FreeSans 16 90 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 1956 -16 1964 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal3 s 5576 396 5584 404 3 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal3 s -24 3556 -16 3564 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 3256 -16 3264 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2736 -16 2744 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal3 s 5576 3776 5584 3784 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal3 s 5576 3516 5584 3524 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal3 s 5576 3036 5584 3044 3 FreeSans 16 0 0 0 Xout[1]
port 16 nsew
flabel metal3 s 5576 2996 5584 3004 3 FreeSans 16 0 0 0 Xout[0]
port 17 nsew
flabel metal2 s 3537 -23 3543 -17 7 FreeSans 16 270 0 0 Yin[3]
port 18 nsew
flabel metal2 s 4677 -23 4683 -17 7 FreeSans 16 270 0 0 Yin[2]
port 19 nsew
flabel metal2 s 5397 -23 5403 -17 7 FreeSans 16 270 0 0 Yin[1]
port 20 nsew
flabel metal2 s 5437 -23 5443 -17 7 FreeSans 16 270 0 0 Yin[0]
port 21 nsew
flabel metal2 s 2837 -23 2843 -17 7 FreeSans 16 270 0 0 Yout[3]
port 22 nsew
flabel metal2 s 3077 -23 3083 -17 7 FreeSans 16 270 0 0 Yout[2]
port 23 nsew
flabel metal2 s 3337 -23 3343 -17 7 FreeSans 16 270 0 0 Yout[1]
port 24 nsew
flabel metal2 s 3437 -23 3443 -17 7 FreeSans 16 270 0 0 Yout[0]
port 25 nsew
flabel metal2 s 4457 5517 4463 5523 3 FreeSans 16 90 0 0 clk
port 26 nsew
<< properties >>
string FIXED_BBOX -40 -40 5580 5520
<< end >>
