magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -120 -120 2520 5180
<< metal1 >>
rect 352 4520 2048 4580
rect 394 2960 2006 3020
rect 0 0 80 1560
rect 2300 1460 2400 1560
rect 100 1400 2400 1460
rect 2300 0 2400 1400
<< metal2 >>
rect 516 4680 1884 5060
rect 0 0 80 1560
rect 264 141 372 1380
rect 394 180 494 4500
rect 516 141 624 4680
rect 646 180 746 4500
rect 768 141 876 4680
rect 898 180 998 4500
rect 1020 141 1128 4680
rect 1150 180 1250 4500
rect 1272 141 1380 4680
rect 1402 180 1502 4500
rect 1524 141 1632 4680
rect 1654 180 1754 4500
rect 1776 141 1884 4680
rect 1906 180 2006 4500
rect 2028 141 2136 1380
rect 264 0 2136 141
rect 2300 0 2400 1560
use VIA2  VIA2_0
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 568 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_1
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 1578 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_2
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 1326 0 1 4260
box -8 -8 8 8
use VIA2  VIA2_3
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 1328 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_4
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 1074 0 1 4260
box -8 -8 8 8
use VIA2  VIA2_5
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 1581 0 1 4260
box -8 -8 8 8
use VIA2  VIA2_6
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 569 0 1 4260
box -8 -8 8 8
use VIA2  VIA2_7
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 1829 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_8
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 823 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_9
array 0 0 0 0 41 36
timestamp 1537935238
transform 1 0 1075 0 1 2304
box -8 -8 8 8
use VIA2  VIA2_10
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 822 0 1 4260
box -8 -8 8 8
use VIA2  VIA2_11
array 0 0 0 0 6 36
timestamp 1537935238
transform 1 0 1833 0 1 4260
box -8 -8 8 8
<< end >>
