magic
tech scmos
magscale 1 3
timestamp 1756367991
<< checkpaint >>
rect -430 18085 14990 18900
rect -430 15010 18085 18085
rect -430 3960 18470 15010
rect -430 915 18085 3960
rect -430 760 15180 915
rect -430 20 14990 760
use MY_LOGO1  MY_LOGO1_0
timestamp 1756365015
transform 1 0 15364 0 1 1490
box 6 0 2466 2172
use MY_LOGO2  MY_LOGO2_0
timestamp 1756367800
transform 1 0 15214 0 1 15140
box 6 0 2466 2172
<< end >>
