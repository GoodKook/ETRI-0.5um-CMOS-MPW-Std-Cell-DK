magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 44
rect 42 14 46 54
rect 62 14 66 54
<< ptransistor >>
rect 20 186 24 246
rect 42 166 46 246
rect 62 166 66 246
<< ndiffusion >>
rect 18 14 20 44
rect 24 14 28 44
rect 40 14 42 54
rect 46 14 48 54
rect 60 14 62 54
rect 66 14 68 54
<< pdiffusion >>
rect 18 186 20 246
rect 24 186 28 246
rect 40 168 42 246
rect 28 166 42 168
rect 46 168 48 246
rect 60 168 62 246
rect 46 166 62 168
rect 66 166 68 246
<< ndcontact >>
rect 6 14 18 44
rect 28 14 40 54
rect 48 14 60 54
rect 68 14 80 54
<< pdcontact >>
rect 6 186 18 246
rect 28 168 40 246
rect 48 168 60 246
rect 68 166 80 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 42 246 46 250
rect 62 246 66 250
rect 20 129 24 186
rect 42 162 46 166
rect 62 162 66 166
rect 47 156 66 162
rect 16 117 24 129
rect 20 44 24 117
rect 47 60 66 66
rect 42 54 46 60
rect 62 54 66 60
rect 20 10 24 14
rect 42 10 46 14
rect 62 10 66 14
<< polycontact >>
rect 35 150 47 162
rect 4 117 16 129
rect 35 60 47 72
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 28 246 40 252
rect 68 246 80 252
rect 6 162 14 186
rect 6 156 35 162
rect 35 72 43 150
rect 53 117 60 168
rect 53 103 63 117
rect 6 60 35 66
rect 6 44 14 60
rect 53 54 60 103
rect 28 8 40 14
rect 68 8 80 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 103 17 117
rect 63 103 77 117
<< metal2 >>
rect 63 117 77 137
rect 3 83 17 103
<< m2p >>
rect 63 123 77 137
rect 3 83 17 97
<< labels >>
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 63 123 77 137 0 Y
port 1 nsew signal output
rlabel metal1 -6 252 106 268 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
