magic
tech scmos
magscale 1 6
timestamp 1555589239
<< checkpaint >>
rect -127 -120 147 5132
<< nwell >>
rect -7 4201 27 4571
rect -7 2241 27 3839
<< metal3 >>
rect 0 4680 20 5012
rect 0 4220 20 4552
rect 0 2260 20 3820
rect 0 0 20 1560
<< end >>
