VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU8_Mult
  CLASS BLOCK ;
  FOREIGN ALU8_Mult ;
  ORIGIN 6.000 6.000 ;
  SIZE 885.000 BY 879.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 873.300 830.700 882.300 866.700 ;
        RECT 0.600 828.300 882.300 830.700 ;
        RECT 873.300 758.700 882.300 828.300 ;
        RECT 0.600 756.300 882.300 758.700 ;
        RECT 873.300 686.700 882.300 756.300 ;
        RECT 0.600 684.300 882.300 686.700 ;
        RECT 873.300 614.700 882.300 684.300 ;
        RECT 0.600 612.300 882.300 614.700 ;
        RECT 873.300 542.700 882.300 612.300 ;
        RECT 0.600 540.300 882.300 542.700 ;
        RECT 873.300 470.700 882.300 540.300 ;
        RECT 0.600 468.300 882.300 470.700 ;
        RECT 873.300 398.700 882.300 468.300 ;
        RECT 0.600 396.300 882.300 398.700 ;
        RECT 873.300 326.700 882.300 396.300 ;
        RECT 0.600 324.300 882.300 326.700 ;
        RECT 873.300 254.700 882.300 324.300 ;
        RECT 0.600 252.300 882.300 254.700 ;
        RECT 873.300 182.700 882.300 252.300 ;
        RECT 0.600 180.300 882.300 182.700 ;
        RECT 873.300 110.700 882.300 180.300 ;
        RECT 0.600 108.300 882.300 110.700 ;
        RECT 873.300 38.700 882.300 108.300 ;
        RECT 0.600 36.300 882.300 38.700 ;
        RECT 873.300 0.300 882.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 864.300 872.400 866.700 ;
        RECT -9.300 794.700 -0.300 864.300 ;
        RECT -9.300 792.300 872.400 794.700 ;
        RECT -9.300 722.700 -0.300 792.300 ;
        RECT -9.300 720.300 872.400 722.700 ;
        RECT -9.300 650.700 -0.300 720.300 ;
        RECT -9.300 648.300 872.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT -9.300 576.300 872.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT -9.300 504.300 872.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT -9.300 432.300 872.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT 655.950 430.950 658.050 432.300 ;
        RECT -9.300 360.300 872.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT 379.950 358.950 382.050 360.300 ;
        RECT 652.950 358.950 655.050 360.300 ;
        RECT 673.950 358.950 676.050 360.300 ;
        RECT -9.300 288.300 872.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT 397.950 286.950 400.050 288.300 ;
        RECT 415.950 286.950 418.050 288.300 ;
        RECT -9.300 216.300 872.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT 319.950 214.950 322.050 216.300 ;
        RECT 484.950 214.950 487.050 216.300 ;
        RECT -9.300 144.300 872.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT -9.300 72.300 872.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT -9.300 0.300 872.400 2.700 ;
      LAYER metal2 ;
        RECT 655.950 430.950 658.050 433.050 ;
        RECT 656.400 382.050 657.450 430.950 ;
        RECT 655.950 379.950 658.050 382.050 ;
        RECT 676.950 381.450 679.050 382.050 ;
        RECT 674.400 380.400 679.050 381.450 ;
        RECT 674.400 361.050 675.450 380.400 ;
        RECT 676.950 379.950 679.050 380.400 ;
        RECT 379.950 358.950 382.050 361.050 ;
        RECT 652.950 358.950 655.050 361.050 ;
        RECT 673.950 358.950 676.050 361.050 ;
        RECT 380.400 343.050 381.450 358.950 ;
        RECT 653.400 343.050 654.450 358.950 ;
        RECT 367.950 340.950 370.050 343.050 ;
        RECT 379.950 340.950 382.050 343.050 ;
        RECT 640.950 340.950 643.050 343.050 ;
        RECT 652.950 340.950 655.050 343.050 ;
        RECT 409.950 309.450 412.050 310.050 ;
        RECT 409.950 308.400 414.450 309.450 ;
        RECT 409.950 307.950 412.050 308.400 ;
        RECT 397.950 286.950 400.050 289.050 ;
        RECT 413.400 288.450 414.450 308.400 ;
        RECT 415.950 288.450 418.050 289.050 ;
        RECT 413.400 287.400 418.050 288.450 ;
        RECT 415.950 286.950 418.050 287.400 ;
        RECT 398.400 271.050 399.450 286.950 ;
        RECT 385.950 268.950 388.050 271.050 ;
        RECT 397.950 268.950 400.050 271.050 ;
        RECT 322.950 237.450 325.050 238.050 ;
        RECT 320.400 236.400 325.050 237.450 ;
        RECT 320.400 217.050 321.450 236.400 ;
        RECT 322.950 235.950 325.050 236.400 ;
        RECT 466.950 235.950 469.050 238.050 ;
        RECT 484.950 235.950 487.050 238.050 ;
        RECT 485.400 217.050 486.450 235.950 ;
        RECT 319.950 214.950 322.050 217.050 ;
        RECT 484.950 214.950 487.050 217.050 ;
      LAYER metal3 ;
        RECT 367.950 342.600 370.050 343.050 ;
        RECT 379.950 342.600 382.050 343.050 ;
        RECT 367.950 341.400 382.050 342.600 ;
        RECT 367.950 340.950 370.050 341.400 ;
        RECT 379.950 340.950 382.050 341.400 ;
        RECT 640.950 342.600 643.050 343.050 ;
        RECT 652.950 342.600 655.050 343.050 ;
        RECT 640.950 341.400 655.050 342.600 ;
        RECT 640.950 340.950 643.050 341.400 ;
        RECT 652.950 340.950 655.050 341.400 ;
        RECT 385.950 270.600 388.050 271.050 ;
        RECT 397.950 270.600 400.050 271.050 ;
        RECT 385.950 269.400 400.050 270.600 ;
        RECT 385.950 268.950 388.050 269.400 ;
        RECT 397.950 268.950 400.050 269.400 ;
        RECT 466.950 237.600 469.050 238.050 ;
        RECT 484.950 237.600 487.050 238.050 ;
        RECT 466.950 236.400 487.050 237.600 ;
        RECT 466.950 235.950 469.050 236.400 ;
        RECT 484.950 235.950 487.050 236.400 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal2 ;
        RECT 860.400 832.050 861.450 873.450 ;
        RECT 850.950 829.950 853.050 832.050 ;
        RECT 859.950 829.950 862.050 832.050 ;
        RECT 851.400 811.050 852.450 829.950 ;
        RECT 844.950 808.950 847.050 811.050 ;
        RECT 850.950 808.950 853.050 811.050 ;
        RECT 851.400 781.050 852.450 808.950 ;
        RECT 835.950 778.950 838.050 781.050 ;
        RECT 850.950 778.950 853.050 781.050 ;
        RECT 836.400 745.050 837.450 778.950 ;
        RECT 835.950 744.450 838.050 745.050 ;
        RECT 833.400 743.400 838.050 744.450 ;
        RECT 829.950 738.450 832.050 739.050 ;
        RECT 833.400 738.450 834.450 743.400 ;
        RECT 835.950 742.950 838.050 743.400 ;
        RECT 829.950 737.400 834.450 738.450 ;
        RECT 829.950 736.950 832.050 737.400 ;
        RECT 859.950 736.950 862.050 739.050 ;
      LAYER metal3 ;
        RECT 850.950 831.600 853.050 832.050 ;
        RECT 859.950 831.600 862.050 832.050 ;
        RECT 850.950 830.400 862.050 831.600 ;
        RECT 850.950 829.950 853.050 830.400 ;
        RECT 859.950 829.950 862.050 830.400 ;
        RECT 844.950 810.600 847.050 811.050 ;
        RECT 850.950 810.600 853.050 811.050 ;
        RECT 844.950 809.400 853.050 810.600 ;
        RECT 844.950 808.950 847.050 809.400 ;
        RECT 850.950 808.950 853.050 809.400 ;
        RECT 835.950 780.600 838.050 781.050 ;
        RECT 850.950 780.600 853.050 781.050 ;
        RECT 835.950 779.400 853.050 780.600 ;
        RECT 835.950 778.950 838.050 779.400 ;
        RECT 850.950 778.950 853.050 779.400 ;
        RECT 835.950 744.600 838.050 745.050 ;
        RECT 835.950 743.400 861.600 744.600 ;
        RECT 835.950 742.950 838.050 743.400 ;
        RECT 860.400 739.050 861.600 743.400 ;
        RECT 859.950 736.950 862.050 739.050 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal2 ;
        RECT 854.400 810.450 855.450 873.450 ;
        RECT 856.950 810.450 859.050 811.050 ;
        RECT 854.400 809.400 859.050 810.450 ;
        RECT 854.400 778.050 855.450 809.400 ;
        RECT 856.950 808.950 859.050 809.400 ;
        RECT 853.950 777.450 856.050 778.050 ;
        RECT 851.400 776.400 856.050 777.450 ;
        RECT 851.400 739.050 852.450 776.400 ;
        RECT 853.950 775.950 856.050 776.400 ;
        RECT 844.950 736.950 847.050 739.050 ;
        RECT 850.950 736.950 853.050 739.050 ;
      LAYER metal3 ;
        RECT 844.950 738.600 847.050 739.050 ;
        RECT 850.950 738.600 853.050 739.050 ;
        RECT 844.950 737.400 853.050 738.600 ;
        RECT 844.950 736.950 847.050 737.400 ;
        RECT 850.950 736.950 853.050 737.400 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal2 ;
        RECT 845.400 853.050 846.450 873.450 ;
        RECT 769.950 850.950 772.050 853.050 ;
        RECT 775.950 850.950 778.050 853.050 ;
        RECT 844.950 850.950 847.050 853.050 ;
        RECT 766.950 849.450 769.050 850.050 ;
        RECT 770.400 849.450 771.450 850.950 ;
        RECT 776.400 850.050 777.450 850.950 ;
        RECT 766.950 848.400 771.450 849.450 ;
        RECT 766.950 847.950 769.050 848.400 ;
        RECT 770.400 844.050 771.450 848.400 ;
        RECT 775.950 847.950 778.050 850.050 ;
        RECT 769.950 841.950 772.050 844.050 ;
        RECT 781.950 841.950 784.050 844.050 ;
        RECT 782.400 799.050 783.450 841.950 ;
        RECT 781.950 796.950 784.050 799.050 ;
        RECT 838.950 796.950 841.050 799.050 ;
        RECT 839.400 778.050 840.450 796.950 ;
        RECT 838.950 775.950 841.050 778.050 ;
      LAYER metal3 ;
        RECT 769.950 852.600 772.050 853.050 ;
        RECT 775.950 852.600 778.050 853.050 ;
        RECT 844.950 852.600 847.050 853.050 ;
        RECT 769.950 851.400 847.050 852.600 ;
        RECT 769.950 850.950 772.050 851.400 ;
        RECT 775.950 850.950 778.050 851.400 ;
        RECT 844.950 850.950 847.050 851.400 ;
        RECT 769.950 843.600 772.050 844.050 ;
        RECT 781.950 843.600 784.050 844.050 ;
        RECT 769.950 842.400 784.050 843.600 ;
        RECT 769.950 841.950 772.050 842.400 ;
        RECT 781.950 841.950 784.050 842.400 ;
        RECT 781.950 798.600 784.050 799.050 ;
        RECT 838.950 798.600 841.050 799.050 ;
        RECT 781.950 797.400 841.050 798.600 ;
        RECT 781.950 796.950 784.050 797.400 ;
        RECT 838.950 796.950 841.050 797.400 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal2 ;
        RECT 839.400 868.050 840.450 873.450 ;
        RECT 808.950 865.950 811.050 868.050 ;
        RECT 838.950 865.950 841.050 868.050 ;
        RECT 766.950 703.950 769.050 706.050 ;
        RECT 772.950 703.950 775.050 706.050 ;
        RECT 767.400 700.050 768.450 703.950 ;
        RECT 766.950 697.950 769.050 700.050 ;
        RECT 796.950 697.950 799.050 700.050 ;
        RECT 797.400 691.050 798.450 697.950 ;
        RECT 809.400 691.050 810.450 865.950 ;
        RECT 796.950 688.950 799.050 691.050 ;
        RECT 808.950 688.950 811.050 691.050 ;
        RECT 797.400 627.450 798.450 688.950 ;
        RECT 794.400 626.400 798.450 627.450 ;
        RECT 794.400 610.050 795.450 626.400 ;
        RECT 784.950 607.950 787.050 610.050 ;
        RECT 793.950 607.950 796.050 610.050 ;
        RECT 785.400 562.050 786.450 607.950 ;
        RECT 757.950 559.950 760.050 562.050 ;
        RECT 784.950 559.950 787.050 562.050 ;
        RECT 823.950 559.950 826.050 562.050 ;
        RECT 824.400 523.050 825.450 559.950 ;
        RECT 823.950 520.950 826.050 523.050 ;
        RECT 829.950 520.950 832.050 523.050 ;
      LAYER metal3 ;
        RECT 808.950 867.600 811.050 868.050 ;
        RECT 838.950 867.600 841.050 868.050 ;
        RECT 808.950 866.400 841.050 867.600 ;
        RECT 808.950 865.950 811.050 866.400 ;
        RECT 838.950 865.950 841.050 866.400 ;
        RECT 766.950 705.600 769.050 706.050 ;
        RECT 772.950 705.600 775.050 706.050 ;
        RECT 766.950 704.400 775.050 705.600 ;
        RECT 766.950 703.950 769.050 704.400 ;
        RECT 772.950 703.950 775.050 704.400 ;
        RECT 766.950 699.600 769.050 700.050 ;
        RECT 796.950 699.600 799.050 700.050 ;
        RECT 766.950 698.400 799.050 699.600 ;
        RECT 766.950 697.950 769.050 698.400 ;
        RECT 796.950 697.950 799.050 698.400 ;
        RECT 796.950 690.600 799.050 691.050 ;
        RECT 808.950 690.600 811.050 691.050 ;
        RECT 796.950 689.400 811.050 690.600 ;
        RECT 796.950 688.950 799.050 689.400 ;
        RECT 808.950 688.950 811.050 689.400 ;
        RECT 784.950 609.600 787.050 610.050 ;
        RECT 793.950 609.600 796.050 610.050 ;
        RECT 784.950 608.400 796.050 609.600 ;
        RECT 784.950 607.950 787.050 608.400 ;
        RECT 793.950 607.950 796.050 608.400 ;
        RECT 757.950 561.600 760.050 562.050 ;
        RECT 784.950 561.600 787.050 562.050 ;
        RECT 823.950 561.600 826.050 562.050 ;
        RECT 757.950 560.400 826.050 561.600 ;
        RECT 757.950 559.950 760.050 560.400 ;
        RECT 784.950 559.950 787.050 560.400 ;
        RECT 823.950 559.950 826.050 560.400 ;
        RECT 823.950 522.600 826.050 523.050 ;
        RECT 829.950 522.600 832.050 523.050 ;
        RECT 823.950 521.400 832.050 522.600 ;
        RECT 823.950 520.950 826.050 521.400 ;
        RECT 829.950 520.950 832.050 521.400 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal2 ;
        RECT 833.400 865.050 834.450 873.450 ;
        RECT 772.950 862.950 775.050 865.050 ;
        RECT 832.950 862.950 835.050 865.050 ;
        RECT 773.400 813.450 774.450 862.950 ;
        RECT 770.400 812.400 774.450 813.450 ;
        RECT 770.400 766.050 771.450 812.400 ;
        RECT 739.950 763.950 742.050 766.050 ;
        RECT 769.950 763.950 772.050 766.050 ;
        RECT 740.400 694.050 741.450 763.950 ;
        RECT 721.950 691.950 724.050 694.050 ;
        RECT 739.950 691.950 742.050 694.050 ;
        RECT 722.400 622.050 723.450 691.950 ;
        RECT 721.950 619.950 724.050 622.050 ;
        RECT 748.950 619.950 751.050 622.050 ;
        RECT 749.400 523.050 750.450 619.950 ;
        RECT 667.950 520.950 670.050 523.050 ;
        RECT 676.950 520.950 679.050 523.050 ;
        RECT 733.950 520.950 736.050 523.050 ;
        RECT 748.950 520.950 751.050 523.050 ;
      LAYER metal3 ;
        RECT 772.950 864.600 775.050 865.050 ;
        RECT 832.950 864.600 835.050 865.050 ;
        RECT 772.950 863.400 835.050 864.600 ;
        RECT 772.950 862.950 775.050 863.400 ;
        RECT 832.950 862.950 835.050 863.400 ;
        RECT 739.950 765.600 742.050 766.050 ;
        RECT 769.950 765.600 772.050 766.050 ;
        RECT 739.950 764.400 772.050 765.600 ;
        RECT 739.950 763.950 742.050 764.400 ;
        RECT 769.950 763.950 772.050 764.400 ;
        RECT 721.950 693.600 724.050 694.050 ;
        RECT 739.950 693.600 742.050 694.050 ;
        RECT 721.950 692.400 742.050 693.600 ;
        RECT 721.950 691.950 724.050 692.400 ;
        RECT 739.950 691.950 742.050 692.400 ;
        RECT 721.950 621.600 724.050 622.050 ;
        RECT 748.950 621.600 751.050 622.050 ;
        RECT 721.950 620.400 751.050 621.600 ;
        RECT 721.950 619.950 724.050 620.400 ;
        RECT 748.950 619.950 751.050 620.400 ;
        RECT 667.950 522.600 670.050 523.050 ;
        RECT 676.950 522.600 679.050 523.050 ;
        RECT 733.950 522.600 736.050 523.050 ;
        RECT 748.950 522.600 751.050 523.050 ;
        RECT 667.950 521.400 751.050 522.600 ;
        RECT 667.950 520.950 670.050 521.400 ;
        RECT 676.950 520.950 679.050 521.400 ;
        RECT 733.950 520.950 736.050 521.400 ;
        RECT 748.950 520.950 751.050 521.400 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal2 ;
        RECT 736.950 448.950 739.050 451.050 ;
        RECT 745.950 448.950 748.050 451.050 ;
        RECT 737.400 448.050 738.450 448.950 ;
        RECT 746.400 448.050 747.450 448.950 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 776.400 418.050 777.450 445.950 ;
        RECT 775.950 415.950 778.050 418.050 ;
      LAYER metal3 ;
        RECT 736.950 447.600 739.050 448.050 ;
        RECT 745.950 447.600 748.050 448.050 ;
        RECT 775.950 447.600 778.050 448.050 ;
        RECT 736.950 446.400 778.050 447.600 ;
        RECT 736.950 445.950 739.050 446.400 ;
        RECT 745.950 445.950 748.050 446.400 ;
        RECT 775.950 445.950 778.050 446.400 ;
        RECT 775.950 417.600 778.050 418.050 ;
        RECT 775.950 416.400 879.600 417.600 ;
        RECT 775.950 415.950 778.050 416.400 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal2 ;
        RECT 835.950 847.950 838.050 850.050 ;
        RECT 844.950 847.950 847.050 850.050 ;
        RECT 845.400 822.450 846.450 847.950 ;
        RECT 845.400 821.400 849.450 822.450 ;
        RECT 848.400 711.450 849.450 821.400 ;
        RECT 845.400 710.400 849.450 711.450 ;
        RECT 845.400 532.050 846.450 710.400 ;
        RECT 805.950 529.950 808.050 532.050 ;
        RECT 844.950 529.950 847.050 532.050 ;
        RECT 806.400 523.050 807.450 529.950 ;
        RECT 772.950 520.950 775.050 523.050 ;
        RECT 805.950 520.950 808.050 523.050 ;
        RECT 773.400 490.050 774.450 520.950 ;
        RECT 739.950 487.950 742.050 490.050 ;
        RECT 772.950 487.950 775.050 490.050 ;
      LAYER metal3 ;
        RECT 835.950 849.600 838.050 850.050 ;
        RECT 844.950 849.600 847.050 850.050 ;
        RECT 835.950 848.400 879.600 849.600 ;
        RECT 835.950 847.950 838.050 848.400 ;
        RECT 844.950 847.950 847.050 848.400 ;
        RECT 878.400 845.400 879.600 848.400 ;
        RECT 805.950 531.600 808.050 532.050 ;
        RECT 844.950 531.600 847.050 532.050 ;
        RECT 805.950 530.400 847.050 531.600 ;
        RECT 805.950 529.950 808.050 530.400 ;
        RECT 844.950 529.950 847.050 530.400 ;
        RECT 772.950 522.600 775.050 523.050 ;
        RECT 805.950 522.600 808.050 523.050 ;
        RECT 772.950 521.400 808.050 522.600 ;
        RECT 772.950 520.950 775.050 521.400 ;
        RECT 805.950 520.950 808.050 521.400 ;
        RECT 739.950 489.600 742.050 490.050 ;
        RECT 772.950 489.600 775.050 490.050 ;
        RECT 739.950 488.400 775.050 489.600 ;
        RECT 739.950 487.950 742.050 488.400 ;
        RECT 772.950 487.950 775.050 488.400 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal2 ;
        RECT 871.950 850.950 874.050 853.050 ;
        RECT 872.400 592.050 873.450 850.950 ;
        RECT 862.950 589.950 865.050 592.050 ;
        RECT 871.950 589.950 874.050 592.050 ;
        RECT 863.400 562.050 864.450 589.950 ;
        RECT 841.950 559.950 844.050 562.050 ;
        RECT 862.950 559.950 865.050 562.050 ;
        RECT 842.400 490.050 843.450 559.950 ;
        RECT 793.950 487.950 796.050 490.050 ;
        RECT 841.950 487.950 844.050 490.050 ;
        RECT 853.950 487.950 856.050 490.050 ;
      LAYER metal3 ;
        RECT 871.950 852.600 874.050 853.050 ;
        RECT 871.950 851.400 879.600 852.600 ;
        RECT 871.950 850.950 874.050 851.400 ;
        RECT 862.950 591.600 865.050 592.050 ;
        RECT 871.950 591.600 874.050 592.050 ;
        RECT 862.950 590.400 874.050 591.600 ;
        RECT 862.950 589.950 865.050 590.400 ;
        RECT 871.950 589.950 874.050 590.400 ;
        RECT 841.950 561.600 844.050 562.050 ;
        RECT 862.950 561.600 865.050 562.050 ;
        RECT 841.950 560.400 865.050 561.600 ;
        RECT 841.950 559.950 844.050 560.400 ;
        RECT 862.950 559.950 865.050 560.400 ;
        RECT 793.950 489.600 796.050 490.050 ;
        RECT 841.950 489.600 844.050 490.050 ;
        RECT 853.950 489.600 856.050 490.050 ;
        RECT 793.950 488.400 856.050 489.600 ;
        RECT 793.950 487.950 796.050 488.400 ;
        RECT 841.950 487.950 844.050 488.400 ;
        RECT 853.950 487.950 856.050 488.400 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal2 ;
        RECT 583.950 24.450 586.050 25.050 ;
        RECT 583.950 23.400 588.450 24.450 ;
        RECT 583.950 22.950 586.050 23.400 ;
        RECT 587.400 -2.550 588.450 23.400 ;
        RECT 584.400 -3.600 588.450 -2.550 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal1 ;
        RECT 568.950 169.950 571.050 172.050 ;
        RECT 569.550 160.050 570.450 169.950 ;
        RECT 568.950 157.950 571.050 160.050 ;
        RECT 577.950 132.450 580.050 133.050 ;
        RECT 572.550 131.550 580.050 132.450 ;
        RECT 568.950 117.450 571.050 118.050 ;
        RECT 572.550 117.450 573.450 131.550 ;
        RECT 577.950 130.950 580.050 131.550 ;
        RECT 568.950 116.550 573.450 117.450 ;
        RECT 568.950 115.950 571.050 116.550 ;
        RECT 580.950 99.450 583.050 100.050 ;
        RECT 578.550 98.550 583.050 99.450 ;
        RECT 578.550 94.050 579.450 98.550 ;
        RECT 580.950 97.950 583.050 98.550 ;
        RECT 577.950 91.950 580.050 94.050 ;
      LAYER metal2 ;
        RECT 574.950 238.950 577.050 241.050 ;
        RECT 580.950 238.950 583.050 241.050 ;
        RECT 575.400 216.450 576.450 238.950 ;
        RECT 575.400 215.400 579.450 216.450 ;
        RECT 578.400 178.050 579.450 215.400 ;
        RECT 568.950 175.950 571.050 178.050 ;
        RECT 577.950 175.950 580.050 178.050 ;
        RECT 569.400 172.050 570.450 175.950 ;
        RECT 568.950 169.950 571.050 172.050 ;
        RECT 568.950 157.950 571.050 160.050 ;
        RECT 569.400 142.050 570.450 157.950 ;
        RECT 568.950 139.950 571.050 142.050 ;
        RECT 577.950 139.950 580.050 142.050 ;
        RECT 578.400 133.050 579.450 139.950 ;
        RECT 577.950 130.950 580.050 133.050 ;
        RECT 568.950 115.950 571.050 118.050 ;
        RECT 569.400 109.050 570.450 115.950 ;
        RECT 568.950 106.950 571.050 109.050 ;
        RECT 583.950 106.950 586.050 109.050 ;
        RECT 580.950 99.450 583.050 100.050 ;
        RECT 584.400 99.450 585.450 106.950 ;
        RECT 580.950 98.400 585.450 99.450 ;
        RECT 580.950 97.950 583.050 98.400 ;
        RECT 577.950 91.950 580.050 94.050 ;
        RECT 578.400 64.050 579.450 91.950 ;
        RECT 577.950 61.950 580.050 64.050 ;
        RECT 583.950 61.950 586.050 64.050 ;
        RECT 584.400 27.450 585.450 61.950 ;
        RECT 581.400 26.400 585.450 27.450 ;
        RECT 581.400 -2.550 582.450 26.400 ;
        RECT 578.400 -3.600 582.450 -2.550 ;
      LAYER metal3 ;
        RECT 574.950 240.600 577.050 241.050 ;
        RECT 580.950 240.600 583.050 241.050 ;
        RECT 574.950 239.400 583.050 240.600 ;
        RECT 574.950 238.950 577.050 239.400 ;
        RECT 580.950 238.950 583.050 239.400 ;
        RECT 568.950 177.600 571.050 178.050 ;
        RECT 577.950 177.600 580.050 178.050 ;
        RECT 568.950 176.400 580.050 177.600 ;
        RECT 568.950 175.950 571.050 176.400 ;
        RECT 577.950 175.950 580.050 176.400 ;
        RECT 568.950 141.600 571.050 142.050 ;
        RECT 577.950 141.600 580.050 142.050 ;
        RECT 568.950 140.400 580.050 141.600 ;
        RECT 568.950 139.950 571.050 140.400 ;
        RECT 577.950 139.950 580.050 140.400 ;
        RECT 568.950 108.600 571.050 109.050 ;
        RECT 583.950 108.600 586.050 109.050 ;
        RECT 568.950 107.400 586.050 108.600 ;
        RECT 568.950 106.950 571.050 107.400 ;
        RECT 583.950 106.950 586.050 107.400 ;
        RECT 577.950 63.600 580.050 64.050 ;
        RECT 583.950 63.600 586.050 64.050 ;
        RECT 577.950 62.400 586.050 63.600 ;
        RECT 577.950 61.950 580.050 62.400 ;
        RECT 583.950 61.950 586.050 62.400 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal2 ;
        RECT 562.950 24.450 565.050 25.050 ;
        RECT 562.950 23.400 567.450 24.450 ;
        RECT 562.950 22.950 565.050 23.400 ;
        RECT 566.400 -2.550 567.450 23.400 ;
        RECT 563.400 -3.600 567.450 -2.550 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal2 ;
        RECT 523.950 193.950 526.050 196.050 ;
        RECT 524.400 184.050 525.450 193.950 ;
        RECT 511.950 181.950 514.050 184.050 ;
        RECT 523.950 181.950 526.050 184.050 ;
        RECT 512.400 127.050 513.450 181.950 ;
        RECT 511.950 124.950 514.050 127.050 ;
        RECT 520.950 124.950 523.050 127.050 ;
        RECT 521.400 -2.550 522.450 124.950 ;
        RECT 521.400 -3.600 525.450 -2.550 ;
      LAYER metal3 ;
        RECT 511.950 183.600 514.050 184.050 ;
        RECT 523.950 183.600 526.050 184.050 ;
        RECT 511.950 182.400 526.050 183.600 ;
        RECT 511.950 181.950 514.050 182.400 ;
        RECT 523.950 181.950 526.050 182.400 ;
        RECT 511.950 126.600 514.050 127.050 ;
        RECT 520.950 126.600 523.050 127.050 ;
        RECT 511.950 125.400 523.050 126.600 ;
        RECT 511.950 124.950 514.050 125.400 ;
        RECT 520.950 124.950 523.050 125.400 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal2 ;
        RECT 337.950 24.450 340.050 25.050 ;
        RECT 337.950 23.400 342.450 24.450 ;
        RECT 337.950 22.950 340.050 23.400 ;
        RECT 341.400 7.050 342.450 23.400 ;
        RECT 340.950 4.950 343.050 7.050 ;
        RECT 400.950 4.950 403.050 7.050 ;
        RECT 401.400 -3.600 402.450 4.950 ;
      LAYER metal3 ;
        RECT 340.950 6.600 343.050 7.050 ;
        RECT 400.950 6.600 403.050 7.050 ;
        RECT 340.950 5.400 403.050 6.600 ;
        RECT 340.950 4.950 343.050 5.400 ;
        RECT 400.950 4.950 403.050 5.400 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal2 ;
        RECT 13.950 340.950 16.050 343.050 ;
        RECT 14.400 313.050 15.450 340.950 ;
        RECT 13.950 310.950 16.050 313.050 ;
      LAYER metal3 ;
        RECT -3.600 342.600 -2.400 345.600 ;
        RECT 13.950 342.600 16.050 343.050 ;
        RECT -3.600 341.400 16.050 342.600 ;
        RECT 13.950 340.950 16.050 341.400 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal2 ;
        RECT 10.950 337.950 13.050 340.050 ;
      LAYER metal3 ;
        RECT 10.950 339.600 13.050 340.050 ;
        RECT -3.600 338.400 13.050 339.600 ;
        RECT 10.950 337.950 13.050 338.400 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal2 ;
        RECT 211.950 240.450 214.050 241.050 ;
        RECT 209.400 239.400 214.050 240.450 ;
        RECT 1.950 232.950 4.050 235.050 ;
        RECT 2.400 226.050 3.450 232.950 ;
        RECT 209.400 226.050 210.450 239.400 ;
        RECT 211.950 238.950 214.050 239.400 ;
        RECT 1.950 223.950 4.050 226.050 ;
        RECT 208.950 223.950 211.050 226.050 ;
      LAYER metal3 ;
        RECT 1.950 234.600 4.050 235.050 ;
        RECT -3.600 233.400 4.050 234.600 ;
        RECT 1.950 232.950 4.050 233.400 ;
        RECT 1.950 225.600 4.050 226.050 ;
        RECT 208.950 225.600 211.050 226.050 ;
        RECT 1.950 224.400 211.050 225.600 ;
        RECT 1.950 223.950 4.050 224.400 ;
        RECT 208.950 223.950 211.050 224.400 ;
    END
  END ACC_o[0]
  PIN Flag_i
    PORT
      LAYER metal2 ;
        RECT 481.950 310.950 484.050 313.050 ;
        RECT 487.950 310.950 490.050 313.050 ;
        RECT 482.400 271.050 483.450 310.950 ;
        RECT 481.950 268.950 484.050 271.050 ;
        RECT 442.950 265.950 445.050 268.050 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 406.950 196.950 409.050 199.050 ;
        RECT 406.950 190.950 409.050 193.050 ;
        RECT 407.400 178.050 408.450 190.950 ;
        RECT 443.400 178.050 444.450 265.950 ;
        RECT 481.950 193.950 484.050 196.050 ;
        RECT 482.400 178.050 483.450 193.950 ;
        RECT 406.950 175.950 409.050 178.050 ;
        RECT 421.950 175.950 424.050 178.050 ;
        RECT 442.950 175.950 445.050 178.050 ;
        RECT 448.950 175.950 451.050 178.050 ;
        RECT 481.950 175.950 484.050 178.050 ;
        RECT 407.400 172.050 408.450 175.950 ;
        RECT 406.950 169.950 409.050 172.050 ;
        RECT 422.400 169.050 423.450 175.950 ;
        RECT 421.950 166.950 424.050 169.050 ;
        RECT 449.400 121.050 450.450 175.950 ;
        RECT 482.400 169.050 483.450 175.950 ;
        RECT 481.950 166.950 484.050 169.050 ;
        RECT 442.950 118.950 445.050 121.050 ;
        RECT 448.950 118.950 451.050 121.050 ;
        RECT 443.400 4.050 444.450 118.950 ;
        RECT 394.950 1.950 397.050 4.050 ;
        RECT 442.950 1.950 445.050 4.050 ;
        RECT 395.400 -3.600 396.450 1.950 ;
      LAYER metal3 ;
        RECT 481.950 312.600 484.050 313.050 ;
        RECT 487.950 312.600 490.050 313.050 ;
        RECT 481.950 311.400 490.050 312.600 ;
        RECT 481.950 310.950 484.050 311.400 ;
        RECT 487.950 310.950 490.050 311.400 ;
        RECT 481.950 268.950 484.050 271.050 ;
        RECT 442.950 267.600 445.050 268.050 ;
        RECT 463.950 267.600 466.050 268.050 ;
        RECT 482.400 267.600 483.600 268.950 ;
        RECT 442.950 266.400 483.600 267.600 ;
        RECT 442.950 265.950 445.050 266.400 ;
        RECT 463.950 265.950 466.050 266.400 ;
        RECT 406.950 196.950 409.050 199.050 ;
        RECT 407.400 193.050 408.600 196.950 ;
        RECT 406.950 190.950 409.050 193.050 ;
        RECT 406.950 177.600 409.050 178.050 ;
        RECT 421.950 177.600 424.050 178.050 ;
        RECT 442.950 177.600 445.050 178.050 ;
        RECT 448.950 177.600 451.050 178.050 ;
        RECT 481.950 177.600 484.050 178.050 ;
        RECT 406.950 176.400 484.050 177.600 ;
        RECT 406.950 175.950 409.050 176.400 ;
        RECT 421.950 175.950 424.050 176.400 ;
        RECT 442.950 175.950 445.050 176.400 ;
        RECT 448.950 175.950 451.050 176.400 ;
        RECT 481.950 175.950 484.050 176.400 ;
        RECT 442.950 120.600 445.050 121.050 ;
        RECT 448.950 120.600 451.050 121.050 ;
        RECT 442.950 119.400 451.050 120.600 ;
        RECT 442.950 118.950 445.050 119.400 ;
        RECT 448.950 118.950 451.050 119.400 ;
        RECT 394.950 3.600 397.050 4.050 ;
        RECT 442.950 3.600 445.050 4.050 ;
        RECT 394.950 2.400 445.050 3.600 ;
        RECT 394.950 1.950 397.050 2.400 ;
        RECT 442.950 1.950 445.050 2.400 ;
    END
  END Flag_i
  PIN LoadA_i
    PORT
      LAYER metal2 ;
        RECT 779.400 872.400 783.450 873.450 ;
        RECT 782.400 850.050 783.450 872.400 ;
        RECT 781.950 849.450 784.050 850.050 ;
        RECT 781.950 848.400 786.450 849.450 ;
        RECT 781.950 847.950 784.050 848.400 ;
        RECT 676.950 841.950 679.050 844.050 ;
        RECT 677.400 835.050 678.450 841.950 ;
        RECT 785.400 835.050 786.450 848.400 ;
        RECT 676.950 832.950 679.050 835.050 ;
        RECT 784.950 832.950 787.050 835.050 ;
        RECT 785.400 823.050 786.450 832.950 ;
        RECT 784.950 820.950 787.050 823.050 ;
        RECT 814.950 820.950 817.050 823.050 ;
        RECT 785.400 811.050 786.450 820.950 ;
        RECT 815.400 817.050 816.450 820.950 ;
        RECT 814.950 814.950 817.050 817.050 ;
        RECT 772.950 808.950 775.050 811.050 ;
        RECT 784.950 808.950 787.050 811.050 ;
        RECT 862.950 808.950 865.050 811.050 ;
        RECT 773.400 745.050 774.450 808.950 ;
        RECT 785.400 808.050 786.450 808.950 ;
        RECT 863.400 808.050 864.450 808.950 ;
        RECT 784.950 805.950 787.050 808.050 ;
        RECT 862.950 805.950 865.050 808.050 ;
        RECT 757.950 742.950 760.050 745.050 ;
        RECT 763.950 742.950 766.050 745.050 ;
        RECT 772.950 742.950 775.050 745.050 ;
        RECT 758.400 733.050 759.450 742.950 ;
        RECT 823.950 736.950 826.050 739.050 ;
        RECT 824.400 733.050 825.450 736.950 ;
        RECT 757.950 730.950 760.050 733.050 ;
        RECT 823.950 730.950 826.050 733.050 ;
        RECT 758.400 709.050 759.450 730.950 ;
        RECT 742.950 706.950 745.050 709.050 ;
        RECT 757.950 706.950 760.050 709.050 ;
        RECT 778.950 706.950 781.050 709.050 ;
        RECT 743.400 700.050 744.450 706.950 ;
        RECT 779.400 706.050 780.450 706.950 ;
        RECT 778.950 703.950 781.050 706.050 ;
        RECT 742.950 697.950 745.050 700.050 ;
        RECT 751.950 697.950 754.050 700.050 ;
        RECT 637.950 529.950 640.050 532.050 ;
        RECT 685.950 529.950 688.050 532.050 ;
        RECT 638.400 529.050 639.450 529.950 ;
        RECT 637.950 526.950 640.050 529.050 ;
        RECT 682.950 522.450 685.050 523.050 ;
        RECT 686.400 522.450 687.450 529.950 ;
        RECT 682.950 521.400 687.450 522.450 ;
        RECT 682.950 520.950 685.050 521.400 ;
        RECT 683.400 493.050 684.450 520.950 ;
        RECT 743.400 493.050 744.450 697.950 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 706.950 490.950 709.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 787.950 490.950 790.050 493.050 ;
        RECT 631.950 481.950 634.050 484.050 ;
        RECT 632.400 481.050 633.450 481.950 ;
        RECT 686.400 481.050 687.450 490.950 ;
        RECT 707.400 483.450 708.450 490.950 ;
        RECT 709.950 483.450 712.050 484.050 ;
        RECT 707.400 482.400 712.050 483.450 ;
        RECT 709.950 481.950 712.050 482.400 ;
        RECT 631.950 478.950 634.050 481.050 ;
        RECT 685.950 478.950 688.050 481.050 ;
        RECT 686.400 457.050 687.450 478.950 ;
        RECT 685.950 454.950 688.050 457.050 ;
        RECT 722.400 451.050 723.450 490.950 ;
        RECT 734.400 490.050 735.450 490.950 ;
        RECT 788.400 490.050 789.450 490.950 ;
        RECT 733.950 487.950 736.050 490.050 ;
        RECT 787.950 487.950 790.050 490.050 ;
        RECT 721.950 448.950 724.050 451.050 ;
        RECT 730.950 448.950 733.050 451.050 ;
      LAYER metal3 ;
        RECT 676.950 834.600 679.050 835.050 ;
        RECT 784.950 834.600 787.050 835.050 ;
        RECT 676.950 833.400 787.050 834.600 ;
        RECT 676.950 832.950 679.050 833.400 ;
        RECT 784.950 832.950 787.050 833.400 ;
        RECT 784.950 822.600 787.050 823.050 ;
        RECT 814.950 822.600 817.050 823.050 ;
        RECT 784.950 821.400 817.050 822.600 ;
        RECT 784.950 820.950 787.050 821.400 ;
        RECT 814.950 820.950 817.050 821.400 ;
        RECT 772.950 810.600 775.050 811.050 ;
        RECT 784.950 810.600 787.050 811.050 ;
        RECT 772.950 809.400 787.050 810.600 ;
        RECT 772.950 808.950 775.050 809.400 ;
        RECT 784.950 808.950 787.050 809.400 ;
        RECT 784.950 807.600 787.050 808.050 ;
        RECT 862.950 807.600 865.050 808.050 ;
        RECT 784.950 806.400 865.050 807.600 ;
        RECT 784.950 805.950 787.050 806.400 ;
        RECT 862.950 805.950 865.050 806.400 ;
        RECT 757.950 744.600 760.050 745.050 ;
        RECT 763.950 744.600 766.050 745.050 ;
        RECT 772.950 744.600 775.050 745.050 ;
        RECT 757.950 743.400 775.050 744.600 ;
        RECT 757.950 742.950 760.050 743.400 ;
        RECT 763.950 742.950 766.050 743.400 ;
        RECT 772.950 742.950 775.050 743.400 ;
        RECT 757.950 732.600 760.050 733.050 ;
        RECT 823.950 732.600 826.050 733.050 ;
        RECT 757.950 731.400 826.050 732.600 ;
        RECT 757.950 730.950 760.050 731.400 ;
        RECT 823.950 730.950 826.050 731.400 ;
        RECT 742.950 708.600 745.050 709.050 ;
        RECT 757.950 708.600 760.050 709.050 ;
        RECT 778.950 708.600 781.050 709.050 ;
        RECT 742.950 707.400 781.050 708.600 ;
        RECT 742.950 706.950 745.050 707.400 ;
        RECT 757.950 706.950 760.050 707.400 ;
        RECT 778.950 706.950 781.050 707.400 ;
        RECT 742.950 699.600 745.050 700.050 ;
        RECT 751.950 699.600 754.050 700.050 ;
        RECT 742.950 698.400 754.050 699.600 ;
        RECT 742.950 697.950 745.050 698.400 ;
        RECT 751.950 697.950 754.050 698.400 ;
        RECT 637.950 531.600 640.050 532.050 ;
        RECT 685.950 531.600 688.050 532.050 ;
        RECT 637.950 530.400 688.050 531.600 ;
        RECT 637.950 529.950 640.050 530.400 ;
        RECT 685.950 529.950 688.050 530.400 ;
        RECT 682.950 492.600 685.050 493.050 ;
        RECT 685.950 492.600 688.050 493.050 ;
        RECT 706.950 492.600 709.050 493.050 ;
        RECT 721.950 492.600 724.050 493.050 ;
        RECT 733.950 492.600 736.050 493.050 ;
        RECT 742.950 492.600 745.050 493.050 ;
        RECT 787.950 492.600 790.050 493.050 ;
        RECT 682.950 491.400 790.050 492.600 ;
        RECT 682.950 490.950 685.050 491.400 ;
        RECT 685.950 490.950 688.050 491.400 ;
        RECT 706.950 490.950 709.050 491.400 ;
        RECT 721.950 490.950 724.050 491.400 ;
        RECT 733.950 490.950 736.050 491.400 ;
        RECT 742.950 490.950 745.050 491.400 ;
        RECT 787.950 490.950 790.050 491.400 ;
        RECT 631.950 480.600 634.050 481.050 ;
        RECT 685.950 480.600 688.050 481.050 ;
        RECT 631.950 479.400 688.050 480.600 ;
        RECT 631.950 478.950 634.050 479.400 ;
        RECT 685.950 478.950 688.050 479.400 ;
        RECT 721.950 450.600 724.050 451.050 ;
        RECT 730.950 450.600 733.050 451.050 ;
        RECT 721.950 449.400 733.050 450.600 ;
        RECT 721.950 448.950 724.050 449.400 ;
        RECT 730.950 448.950 733.050 449.400 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal2 ;
        RECT 785.400 868.050 786.450 873.450 ;
        RECT 760.950 865.950 763.050 868.050 ;
        RECT 784.950 865.950 787.050 868.050 ;
        RECT 761.400 850.050 762.450 865.950 ;
        RECT 760.950 849.450 763.050 850.050 ;
        RECT 758.400 848.400 763.050 849.450 ;
        RECT 758.400 844.050 759.450 848.400 ;
        RECT 760.950 847.950 763.050 848.400 ;
        RECT 748.950 841.950 751.050 844.050 ;
        RECT 757.950 841.950 760.050 844.050 ;
        RECT 749.400 840.450 750.450 841.950 ;
        RECT 746.400 839.400 750.450 840.450 ;
        RECT 746.400 739.050 747.450 839.400 ;
        RECT 859.950 777.450 862.050 778.050 ;
        RECT 859.950 776.400 864.450 777.450 ;
        RECT 859.950 775.950 862.050 776.400 ;
        RECT 863.400 772.050 864.450 776.400 ;
        RECT 814.950 769.950 817.050 772.050 ;
        RECT 856.950 769.950 859.050 772.050 ;
        RECT 862.950 769.950 865.050 772.050 ;
        RECT 815.400 739.050 816.450 769.950 ;
        RECT 745.950 736.950 748.050 739.050 ;
        RECT 769.950 736.950 772.050 739.050 ;
        RECT 814.950 736.950 817.050 739.050 ;
        RECT 770.400 682.050 771.450 736.950 ;
        RECT 815.400 736.050 816.450 736.950 ;
        RECT 857.400 736.050 858.450 769.950 ;
        RECT 865.950 736.950 868.050 739.050 ;
        RECT 866.400 736.050 867.450 736.950 ;
        RECT 814.950 733.950 817.050 736.050 ;
        RECT 856.950 733.950 859.050 736.050 ;
        RECT 865.950 733.950 868.050 736.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 794.400 679.050 795.450 679.950 ;
        RECT 793.950 676.950 796.050 679.050 ;
        RECT 802.950 676.950 805.050 679.050 ;
        RECT 794.400 637.050 795.450 676.950 ;
        RECT 803.400 673.050 804.450 676.950 ;
        RECT 802.950 670.950 805.050 673.050 ;
        RECT 793.950 634.950 796.050 637.050 ;
        RECT 850.950 628.950 853.050 631.050 ;
        RECT 851.400 600.450 852.450 628.950 ;
        RECT 853.950 600.450 856.050 601.050 ;
        RECT 851.400 599.400 856.050 600.450 ;
        RECT 851.400 589.050 852.450 599.400 ;
        RECT 853.950 598.950 856.050 599.400 ;
        RECT 850.950 586.950 853.050 589.050 ;
        RECT 856.950 586.950 859.050 589.050 ;
        RECT 857.400 565.050 858.450 586.950 ;
        RECT 751.950 562.950 754.050 565.050 ;
        RECT 772.950 562.950 775.050 565.050 ;
        RECT 856.950 562.950 859.050 565.050 ;
        RECT 752.400 562.050 753.450 562.950 ;
        RECT 751.950 559.950 754.050 562.050 ;
        RECT 773.400 556.050 774.450 562.950 ;
        RECT 857.400 562.050 858.450 562.950 ;
        RECT 856.950 559.950 859.050 562.050 ;
        RECT 709.950 553.950 712.050 556.050 ;
        RECT 772.950 553.950 775.050 556.050 ;
        RECT 773.400 529.050 774.450 553.950 ;
        RECT 760.950 526.950 763.050 529.050 ;
        RECT 769.950 526.950 772.050 529.050 ;
        RECT 772.950 526.950 775.050 529.050 ;
        RECT 661.950 520.950 664.050 523.050 ;
        RECT 662.400 504.450 663.450 520.950 ;
        RECT 770.400 520.050 771.450 526.950 ;
        RECT 778.950 520.950 781.050 523.050 ;
        RECT 779.400 520.050 780.450 520.950 ;
        RECT 766.950 517.950 769.050 520.050 ;
        RECT 769.950 517.950 772.050 520.050 ;
        RECT 778.950 517.950 781.050 520.050 ;
        RECT 662.400 503.400 666.450 504.450 ;
        RECT 652.950 481.950 655.050 484.050 ;
        RECT 653.400 466.050 654.450 481.950 ;
        RECT 665.400 466.050 666.450 503.400 ;
        RECT 652.950 463.950 655.050 466.050 ;
        RECT 664.950 463.950 667.050 466.050 ;
        RECT 706.950 463.950 709.050 466.050 ;
        RECT 707.400 460.050 708.450 463.950 ;
        RECT 767.400 460.050 768.450 517.950 ;
        RECT 706.950 457.950 709.050 460.050 ;
        RECT 766.950 457.950 769.050 460.050 ;
        RECT 707.400 457.050 708.450 457.950 ;
        RECT 706.950 454.950 709.050 457.050 ;
        RECT 767.400 451.050 768.450 457.950 ;
        RECT 751.950 448.950 754.050 451.050 ;
        RECT 766.950 448.950 769.050 451.050 ;
      LAYER metal3 ;
        RECT 760.950 867.600 763.050 868.050 ;
        RECT 784.950 867.600 787.050 868.050 ;
        RECT 760.950 866.400 787.050 867.600 ;
        RECT 760.950 865.950 763.050 866.400 ;
        RECT 784.950 865.950 787.050 866.400 ;
        RECT 748.950 843.600 751.050 844.050 ;
        RECT 757.950 843.600 760.050 844.050 ;
        RECT 748.950 842.400 760.050 843.600 ;
        RECT 748.950 841.950 751.050 842.400 ;
        RECT 757.950 841.950 760.050 842.400 ;
        RECT 856.950 771.600 859.050 772.050 ;
        RECT 862.950 771.600 865.050 772.050 ;
        RECT 856.950 770.400 865.050 771.600 ;
        RECT 856.950 769.950 859.050 770.400 ;
        RECT 862.950 769.950 865.050 770.400 ;
        RECT 745.950 738.600 748.050 739.050 ;
        RECT 769.950 738.600 772.050 739.050 ;
        RECT 814.950 738.600 817.050 739.050 ;
        RECT 745.950 737.400 817.050 738.600 ;
        RECT 745.950 736.950 748.050 737.400 ;
        RECT 769.950 736.950 772.050 737.400 ;
        RECT 814.950 736.950 817.050 737.400 ;
        RECT 814.950 735.600 817.050 736.050 ;
        RECT 856.950 735.600 859.050 736.050 ;
        RECT 865.950 735.600 868.050 736.050 ;
        RECT 814.950 734.400 868.050 735.600 ;
        RECT 814.950 733.950 817.050 734.400 ;
        RECT 856.950 733.950 859.050 734.400 ;
        RECT 865.950 733.950 868.050 734.400 ;
        RECT 769.950 681.600 772.050 682.050 ;
        RECT 793.950 681.600 796.050 682.050 ;
        RECT 769.950 680.400 796.050 681.600 ;
        RECT 769.950 679.950 772.050 680.400 ;
        RECT 793.950 679.950 796.050 680.400 ;
        RECT 793.950 678.600 796.050 679.050 ;
        RECT 802.950 678.600 805.050 679.050 ;
        RECT 793.950 677.400 805.050 678.600 ;
        RECT 793.950 676.950 796.050 677.400 ;
        RECT 802.950 676.950 805.050 677.400 ;
        RECT 793.950 636.600 796.050 637.050 ;
        RECT 793.950 635.400 828.600 636.600 ;
        RECT 793.950 634.950 796.050 635.400 ;
        RECT 827.400 630.600 828.600 635.400 ;
        RECT 850.950 630.600 853.050 631.050 ;
        RECT 827.400 629.400 853.050 630.600 ;
        RECT 850.950 628.950 853.050 629.400 ;
        RECT 850.950 588.600 853.050 589.050 ;
        RECT 856.950 588.600 859.050 589.050 ;
        RECT 850.950 587.400 859.050 588.600 ;
        RECT 850.950 586.950 853.050 587.400 ;
        RECT 856.950 586.950 859.050 587.400 ;
        RECT 751.950 564.600 754.050 565.050 ;
        RECT 772.950 564.600 775.050 565.050 ;
        RECT 856.950 564.600 859.050 565.050 ;
        RECT 751.950 563.400 859.050 564.600 ;
        RECT 751.950 562.950 754.050 563.400 ;
        RECT 772.950 562.950 775.050 563.400 ;
        RECT 856.950 562.950 859.050 563.400 ;
        RECT 709.950 555.600 712.050 556.050 ;
        RECT 772.950 555.600 775.050 556.050 ;
        RECT 709.950 554.400 775.050 555.600 ;
        RECT 709.950 553.950 712.050 554.400 ;
        RECT 772.950 553.950 775.050 554.400 ;
        RECT 760.950 528.600 763.050 529.050 ;
        RECT 769.950 528.600 772.050 529.050 ;
        RECT 772.950 528.600 775.050 529.050 ;
        RECT 760.950 527.400 775.050 528.600 ;
        RECT 760.950 526.950 763.050 527.400 ;
        RECT 769.950 526.950 772.050 527.400 ;
        RECT 772.950 526.950 775.050 527.400 ;
        RECT 766.950 519.600 769.050 520.050 ;
        RECT 769.950 519.600 772.050 520.050 ;
        RECT 778.950 519.600 781.050 520.050 ;
        RECT 766.950 518.400 781.050 519.600 ;
        RECT 766.950 517.950 769.050 518.400 ;
        RECT 769.950 517.950 772.050 518.400 ;
        RECT 778.950 517.950 781.050 518.400 ;
        RECT 652.950 465.600 655.050 466.050 ;
        RECT 664.950 465.600 667.050 466.050 ;
        RECT 706.950 465.600 709.050 466.050 ;
        RECT 652.950 464.400 709.050 465.600 ;
        RECT 652.950 463.950 655.050 464.400 ;
        RECT 664.950 463.950 667.050 464.400 ;
        RECT 706.950 463.950 709.050 464.400 ;
        RECT 706.950 459.600 709.050 460.050 ;
        RECT 766.950 459.600 769.050 460.050 ;
        RECT 706.950 458.400 769.050 459.600 ;
        RECT 706.950 457.950 709.050 458.400 ;
        RECT 766.950 457.950 769.050 458.400 ;
        RECT 751.950 450.600 754.050 451.050 ;
        RECT 766.950 450.600 769.050 451.050 ;
        RECT 751.950 449.400 769.050 450.600 ;
        RECT 751.950 448.950 754.050 449.400 ;
        RECT 766.950 448.950 769.050 449.400 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal2 ;
        RECT 827.400 849.450 828.450 873.450 ;
        RECT 829.950 849.450 832.050 850.050 ;
        RECT 827.400 848.400 832.050 849.450 ;
        RECT 827.400 844.050 828.450 848.400 ;
        RECT 829.950 847.950 832.050 848.400 ;
        RECT 826.950 841.950 829.050 844.050 ;
        RECT 835.950 841.950 838.050 844.050 ;
        RECT 836.400 805.050 837.450 841.950 ;
        RECT 838.950 808.950 841.050 811.050 ;
        RECT 839.400 805.050 840.450 808.950 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 844.950 802.950 847.050 805.050 ;
        RECT 845.400 778.050 846.450 802.950 ;
        RECT 760.950 775.950 763.050 778.050 ;
        RECT 844.950 775.950 847.050 778.050 ;
        RECT 761.400 769.050 762.450 775.950 ;
        RECT 778.950 769.950 781.050 772.050 ;
        RECT 779.400 769.050 780.450 769.950 ;
        RECT 760.950 766.950 763.050 769.050 ;
        RECT 778.950 766.950 781.050 769.050 ;
        RECT 761.400 721.050 762.450 766.950 ;
        RECT 838.950 736.950 841.050 739.050 ;
        RECT 839.400 735.450 840.450 736.950 ;
        RECT 839.400 734.400 843.450 735.450 ;
        RECT 842.400 721.050 843.450 734.400 ;
        RECT 760.950 718.950 763.050 721.050 ;
        RECT 841.950 718.950 844.050 721.050 ;
        RECT 865.950 718.950 868.050 721.050 ;
        RECT 866.400 700.050 867.450 718.950 ;
        RECT 859.950 697.950 862.050 700.050 ;
        RECT 865.950 697.950 868.050 700.050 ;
        RECT 856.950 672.450 859.050 673.050 ;
        RECT 860.400 672.450 861.450 697.950 ;
        RECT 856.950 671.400 861.450 672.450 ;
        RECT 856.950 670.950 859.050 671.400 ;
        RECT 860.400 664.050 861.450 671.400 ;
        RECT 835.950 661.950 838.050 664.050 ;
        RECT 859.950 661.950 862.050 664.050 ;
        RECT 836.400 628.050 837.450 661.950 ;
        RECT 820.950 625.950 823.050 628.050 ;
        RECT 835.950 625.950 838.050 628.050 ;
        RECT 836.400 529.050 837.450 625.950 ;
        RECT 835.950 526.950 838.050 529.050 ;
        RECT 838.950 526.950 841.050 529.050 ;
        RECT 844.950 526.950 847.050 529.050 ;
        RECT 739.950 520.950 742.050 523.050 ;
        RECT 835.950 522.450 838.050 523.050 ;
        RECT 839.400 522.450 840.450 526.950 ;
        RECT 835.950 521.400 840.450 522.450 ;
        RECT 835.950 520.950 838.050 521.400 ;
        RECT 740.400 505.050 741.450 520.950 ;
        RECT 836.400 517.050 837.450 520.950 ;
        RECT 835.950 514.950 838.050 517.050 ;
        RECT 847.950 514.950 850.050 517.050 ;
        RECT 739.950 502.950 742.050 505.050 ;
        RECT 745.950 502.950 748.050 505.050 ;
        RECT 746.400 484.050 747.450 502.950 ;
        RECT 848.400 490.050 849.450 514.950 ;
        RECT 847.950 489.450 850.050 490.050 ;
        RECT 845.400 488.400 850.050 489.450 ;
        RECT 845.400 484.050 846.450 488.400 ;
        RECT 847.950 487.950 850.050 488.400 ;
        RECT 742.950 481.950 745.050 484.050 ;
        RECT 745.950 481.950 748.050 484.050 ;
        RECT 760.950 481.950 763.050 484.050 ;
        RECT 820.950 481.950 823.050 484.050 ;
        RECT 844.950 481.950 847.050 484.050 ;
        RECT 743.400 418.050 744.450 481.950 ;
        RECT 742.950 415.950 745.050 418.050 ;
        RECT 769.950 415.950 772.050 418.050 ;
        RECT 743.400 412.050 744.450 415.950 ;
        RECT 742.950 409.950 745.050 412.050 ;
        RECT 748.950 409.950 751.050 412.050 ;
        RECT 841.950 409.950 844.050 412.050 ;
        RECT 749.400 409.050 750.450 409.950 ;
        RECT 842.400 409.050 843.450 409.950 ;
        RECT 748.950 406.950 751.050 409.050 ;
        RECT 841.950 406.950 844.050 409.050 ;
      LAYER metal3 ;
        RECT 826.950 843.600 829.050 844.050 ;
        RECT 835.950 843.600 838.050 844.050 ;
        RECT 826.950 842.400 838.050 843.600 ;
        RECT 826.950 841.950 829.050 842.400 ;
        RECT 835.950 841.950 838.050 842.400 ;
        RECT 835.950 804.600 838.050 805.050 ;
        RECT 838.950 804.600 841.050 805.050 ;
        RECT 844.950 804.600 847.050 805.050 ;
        RECT 835.950 803.400 847.050 804.600 ;
        RECT 835.950 802.950 838.050 803.400 ;
        RECT 838.950 802.950 841.050 803.400 ;
        RECT 844.950 802.950 847.050 803.400 ;
        RECT 760.950 777.600 763.050 778.050 ;
        RECT 844.950 777.600 847.050 778.050 ;
        RECT 760.950 776.400 847.050 777.600 ;
        RECT 760.950 775.950 763.050 776.400 ;
        RECT 844.950 775.950 847.050 776.400 ;
        RECT 760.950 768.600 763.050 769.050 ;
        RECT 778.950 768.600 781.050 769.050 ;
        RECT 760.950 767.400 781.050 768.600 ;
        RECT 760.950 766.950 763.050 767.400 ;
        RECT 778.950 766.950 781.050 767.400 ;
        RECT 760.950 720.600 763.050 721.050 ;
        RECT 841.950 720.600 844.050 721.050 ;
        RECT 865.950 720.600 868.050 721.050 ;
        RECT 760.950 719.400 868.050 720.600 ;
        RECT 760.950 718.950 763.050 719.400 ;
        RECT 841.950 718.950 844.050 719.400 ;
        RECT 865.950 718.950 868.050 719.400 ;
        RECT 859.950 699.600 862.050 700.050 ;
        RECT 865.950 699.600 868.050 700.050 ;
        RECT 859.950 698.400 868.050 699.600 ;
        RECT 859.950 697.950 862.050 698.400 ;
        RECT 865.950 697.950 868.050 698.400 ;
        RECT 835.950 663.600 838.050 664.050 ;
        RECT 859.950 663.600 862.050 664.050 ;
        RECT 835.950 662.400 862.050 663.600 ;
        RECT 835.950 661.950 838.050 662.400 ;
        RECT 859.950 661.950 862.050 662.400 ;
        RECT 820.950 627.600 823.050 628.050 ;
        RECT 835.950 627.600 838.050 628.050 ;
        RECT 820.950 626.400 838.050 627.600 ;
        RECT 820.950 625.950 823.050 626.400 ;
        RECT 835.950 625.950 838.050 626.400 ;
        RECT 835.950 528.600 838.050 529.050 ;
        RECT 838.950 528.600 841.050 529.050 ;
        RECT 844.950 528.600 847.050 529.050 ;
        RECT 835.950 527.400 847.050 528.600 ;
        RECT 835.950 526.950 838.050 527.400 ;
        RECT 838.950 526.950 841.050 527.400 ;
        RECT 844.950 526.950 847.050 527.400 ;
        RECT 835.950 516.600 838.050 517.050 ;
        RECT 847.950 516.600 850.050 517.050 ;
        RECT 835.950 515.400 850.050 516.600 ;
        RECT 835.950 514.950 838.050 515.400 ;
        RECT 847.950 514.950 850.050 515.400 ;
        RECT 739.950 504.600 742.050 505.050 ;
        RECT 745.950 504.600 748.050 505.050 ;
        RECT 739.950 503.400 748.050 504.600 ;
        RECT 739.950 502.950 742.050 503.400 ;
        RECT 745.950 502.950 748.050 503.400 ;
        RECT 742.950 483.600 745.050 484.050 ;
        RECT 745.950 483.600 748.050 484.050 ;
        RECT 760.950 483.600 763.050 484.050 ;
        RECT 820.950 483.600 823.050 484.050 ;
        RECT 844.950 483.600 847.050 484.050 ;
        RECT 742.950 482.400 847.050 483.600 ;
        RECT 742.950 481.950 745.050 482.400 ;
        RECT 745.950 481.950 748.050 482.400 ;
        RECT 760.950 481.950 763.050 482.400 ;
        RECT 820.950 481.950 823.050 482.400 ;
        RECT 844.950 481.950 847.050 482.400 ;
        RECT 742.950 417.600 745.050 418.050 ;
        RECT 769.950 417.600 772.050 418.050 ;
        RECT 742.950 416.400 772.050 417.600 ;
        RECT 742.950 415.950 745.050 416.400 ;
        RECT 769.950 415.950 772.050 416.400 ;
        RECT 742.950 411.600 745.050 412.050 ;
        RECT 748.950 411.600 751.050 412.050 ;
        RECT 742.950 410.400 751.050 411.600 ;
        RECT 742.950 409.950 745.050 410.400 ;
        RECT 748.950 409.950 751.050 410.400 ;
        RECT 748.950 408.600 751.050 409.050 ;
        RECT 841.950 408.600 844.050 409.050 ;
        RECT 748.950 407.400 844.050 408.600 ;
        RECT 748.950 406.950 751.050 407.400 ;
        RECT 841.950 406.950 844.050 407.400 ;
    END
  END LoadCmd_i
  PIN MulH_i
    PORT
      LAYER metal1 ;
        RECT 559.950 387.450 562.050 388.050 ;
        RECT 557.550 386.550 562.050 387.450 ;
        RECT 557.550 382.050 558.450 386.550 ;
        RECT 559.950 385.950 562.050 386.550 ;
        RECT 556.950 379.950 559.050 382.050 ;
      LAYER metal2 ;
        RECT 508.950 556.950 511.050 559.050 ;
        RECT 509.400 538.050 510.450 556.950 ;
        RECT 496.950 535.950 499.050 538.050 ;
        RECT 508.950 535.950 511.050 538.050 ;
        RECT 382.950 511.950 385.050 514.050 ;
        RECT 436.950 511.950 439.050 514.050 ;
        RECT 383.400 505.050 384.450 511.950 ;
        RECT 437.400 508.050 438.450 511.950 ;
        RECT 497.400 511.050 498.450 535.950 ;
        RECT 496.950 508.950 499.050 511.050 ;
        RECT 538.950 508.950 541.050 511.050 ;
        RECT 436.950 505.950 439.050 508.050 ;
        RECT 154.950 502.950 157.050 505.050 ;
        RECT 382.950 502.950 385.050 505.050 ;
        RECT 155.400 472.050 156.450 502.950 ;
        RECT 539.400 495.450 540.450 508.950 ;
        RECT 536.400 494.400 540.450 495.450 ;
        RECT 536.400 472.050 537.450 494.400 ;
        RECT 1.950 469.950 4.050 472.050 ;
        RECT 154.950 469.950 157.050 472.050 ;
        RECT 535.950 469.950 538.050 472.050 ;
        RECT 541.950 469.950 544.050 472.050 ;
        RECT 2.400 454.050 3.450 469.950 ;
        RECT 155.400 454.050 156.450 469.950 ;
        RECT 1.950 451.950 4.050 454.050 ;
        RECT 145.950 451.950 148.050 454.050 ;
        RECT 154.950 451.950 157.050 454.050 ;
        RECT 542.400 412.050 543.450 469.950 ;
        RECT 550.950 412.950 553.050 415.050 ;
        RECT 551.400 412.050 552.450 412.950 ;
        RECT 541.950 409.950 544.050 412.050 ;
        RECT 550.950 409.950 553.050 412.050 ;
        RECT 559.950 409.950 562.050 412.050 ;
        RECT 560.400 388.050 561.450 409.950 ;
        RECT 559.950 385.950 562.050 388.050 ;
        RECT 556.950 379.950 559.050 382.050 ;
        RECT 557.400 367.050 558.450 379.950 ;
        RECT 511.950 364.950 514.050 367.050 ;
        RECT 556.950 364.950 559.050 367.050 ;
        RECT 512.400 343.050 513.450 364.950 ;
        RECT 487.950 340.950 490.050 343.050 ;
        RECT 493.950 340.950 496.050 343.050 ;
        RECT 511.950 340.950 514.050 343.050 ;
        RECT 488.400 328.050 489.450 340.950 ;
        RECT 487.950 325.950 490.050 328.050 ;
        RECT 499.950 325.950 502.050 328.050 ;
        RECT 500.400 307.050 501.450 325.950 ;
        RECT 532.950 307.950 535.050 310.050 ;
        RECT 556.950 307.950 559.050 310.050 ;
        RECT 533.400 307.050 534.450 307.950 ;
        RECT 499.950 304.950 502.050 307.050 ;
        RECT 532.950 304.950 535.050 307.050 ;
      LAYER metal3 ;
        RECT 496.950 537.600 499.050 538.050 ;
        RECT 508.950 537.600 511.050 538.050 ;
        RECT 496.950 536.400 511.050 537.600 ;
        RECT 496.950 535.950 499.050 536.400 ;
        RECT 508.950 535.950 511.050 536.400 ;
        RECT 382.950 513.600 385.050 514.050 ;
        RECT 436.950 513.600 439.050 514.050 ;
        RECT 382.950 512.400 439.050 513.600 ;
        RECT 382.950 511.950 385.050 512.400 ;
        RECT 436.950 511.950 439.050 512.400 ;
        RECT 496.950 510.600 499.050 511.050 ;
        RECT 538.950 510.600 541.050 511.050 ;
        RECT 485.400 509.400 541.050 510.600 ;
        RECT 436.950 507.600 439.050 508.050 ;
        RECT 485.400 507.600 486.600 509.400 ;
        RECT 496.950 508.950 499.050 509.400 ;
        RECT 538.950 508.950 541.050 509.400 ;
        RECT 436.950 506.400 486.600 507.600 ;
        RECT 436.950 505.950 439.050 506.400 ;
        RECT 154.950 504.600 157.050 505.050 ;
        RECT 382.950 504.600 385.050 505.050 ;
        RECT 154.950 503.400 385.050 504.600 ;
        RECT 154.950 502.950 157.050 503.400 ;
        RECT 382.950 502.950 385.050 503.400 ;
        RECT 1.950 471.600 4.050 472.050 ;
        RECT 154.950 471.600 157.050 472.050 ;
        RECT 1.950 470.400 157.050 471.600 ;
        RECT 1.950 469.950 4.050 470.400 ;
        RECT 154.950 469.950 157.050 470.400 ;
        RECT 535.950 471.600 538.050 472.050 ;
        RECT 541.950 471.600 544.050 472.050 ;
        RECT 535.950 470.400 544.050 471.600 ;
        RECT 535.950 469.950 538.050 470.400 ;
        RECT 541.950 469.950 544.050 470.400 ;
        RECT 1.950 453.600 4.050 454.050 ;
        RECT -3.600 452.400 4.050 453.600 ;
        RECT 1.950 451.950 4.050 452.400 ;
        RECT 145.950 453.600 148.050 454.050 ;
        RECT 154.950 453.600 157.050 454.050 ;
        RECT 145.950 452.400 157.050 453.600 ;
        RECT 145.950 451.950 148.050 452.400 ;
        RECT 154.950 451.950 157.050 452.400 ;
        RECT 541.950 411.600 544.050 412.050 ;
        RECT 550.950 411.600 553.050 412.050 ;
        RECT 559.950 411.600 562.050 412.050 ;
        RECT 541.950 410.400 562.050 411.600 ;
        RECT 541.950 409.950 544.050 410.400 ;
        RECT 550.950 409.950 553.050 410.400 ;
        RECT 559.950 409.950 562.050 410.400 ;
        RECT 511.950 366.600 514.050 367.050 ;
        RECT 556.950 366.600 559.050 367.050 ;
        RECT 511.950 365.400 559.050 366.600 ;
        RECT 511.950 364.950 514.050 365.400 ;
        RECT 556.950 364.950 559.050 365.400 ;
        RECT 487.950 342.600 490.050 343.050 ;
        RECT 493.950 342.600 496.050 343.050 ;
        RECT 511.950 342.600 514.050 343.050 ;
        RECT 487.950 341.400 514.050 342.600 ;
        RECT 487.950 340.950 490.050 341.400 ;
        RECT 493.950 340.950 496.050 341.400 ;
        RECT 511.950 340.950 514.050 341.400 ;
        RECT 487.950 327.600 490.050 328.050 ;
        RECT 499.950 327.600 502.050 328.050 ;
        RECT 487.950 326.400 502.050 327.600 ;
        RECT 487.950 325.950 490.050 326.400 ;
        RECT 499.950 325.950 502.050 326.400 ;
        RECT 532.950 309.600 535.050 310.050 ;
        RECT 556.950 309.600 559.050 310.050 ;
        RECT 532.950 308.400 559.050 309.600 ;
        RECT 532.950 307.950 535.050 308.400 ;
        RECT 556.950 307.950 559.050 308.400 ;
        RECT 499.950 306.600 502.050 307.050 ;
        RECT 532.950 306.600 535.050 307.050 ;
        RECT 499.950 305.400 535.050 306.600 ;
        RECT 499.950 304.950 502.050 305.400 ;
        RECT 532.950 304.950 535.050 305.400 ;
    END
  END MulH_i
  PIN MulL_i
    PORT
      LAYER metal2 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 85.950 525.450 88.050 526.050 ;
        RECT 83.400 524.400 88.050 525.450 ;
        RECT 83.400 523.050 84.450 524.400 ;
        RECT 85.950 523.950 88.050 524.400 ;
        RECT 82.950 520.950 85.050 523.050 ;
        RECT 83.400 517.050 84.450 520.950 ;
        RECT 82.950 514.950 85.050 517.050 ;
        RECT 88.950 514.950 91.050 517.050 ;
        RECT 89.400 442.050 90.450 514.950 ;
        RECT 103.950 453.450 106.050 454.050 ;
        RECT 103.950 452.400 108.450 453.450 ;
        RECT 103.950 451.950 106.050 452.400 ;
        RECT 107.400 442.050 108.450 452.400 ;
        RECT 88.950 439.950 91.050 442.050 ;
        RECT 106.950 439.950 109.050 442.050 ;
        RECT 172.950 439.950 175.050 442.050 ;
        RECT 173.400 427.050 174.450 439.950 ;
        RECT 172.950 424.950 175.050 427.050 ;
        RECT 442.950 424.950 445.050 427.050 ;
        RECT 490.950 424.950 493.050 427.050 ;
        RECT 173.400 378.450 174.450 424.950 ;
        RECT 439.950 414.450 442.050 415.050 ;
        RECT 443.400 414.450 444.450 424.950 ;
        RECT 439.950 413.400 444.450 414.450 ;
        RECT 491.400 414.450 492.450 424.950 ;
        RECT 493.950 414.450 496.050 415.050 ;
        RECT 491.400 413.400 496.050 414.450 ;
        RECT 439.950 412.950 442.050 413.400 ;
        RECT 170.400 377.400 174.450 378.450 ;
        RECT 170.400 343.050 171.450 377.400 ;
        RECT 169.950 340.950 172.050 343.050 ;
        RECT 443.400 319.050 444.450 413.400 ;
        RECT 493.950 412.950 496.050 413.400 ;
        RECT 442.950 316.950 445.050 319.050 ;
        RECT 493.950 316.950 496.050 319.050 ;
        RECT 443.400 301.050 444.450 316.950 ;
        RECT 494.400 313.050 495.450 316.950 ;
        RECT 493.950 310.950 496.050 313.050 ;
        RECT 442.950 298.950 445.050 301.050 ;
        RECT 454.950 298.950 457.050 301.050 ;
        RECT 455.400 274.050 456.450 298.950 ;
        RECT 430.950 271.950 433.050 274.050 ;
        RECT 454.950 271.950 457.050 274.050 ;
      LAYER metal3 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 11.400 522.600 12.600 523.950 ;
        RECT 82.950 522.600 85.050 523.050 ;
        RECT -3.600 521.400 85.050 522.600 ;
        RECT 82.950 520.950 85.050 521.400 ;
        RECT 82.950 516.600 85.050 517.050 ;
        RECT 88.950 516.600 91.050 517.050 ;
        RECT 82.950 515.400 91.050 516.600 ;
        RECT 82.950 514.950 85.050 515.400 ;
        RECT 88.950 514.950 91.050 515.400 ;
        RECT 88.950 441.600 91.050 442.050 ;
        RECT 106.950 441.600 109.050 442.050 ;
        RECT 172.950 441.600 175.050 442.050 ;
        RECT 88.950 440.400 175.050 441.600 ;
        RECT 88.950 439.950 91.050 440.400 ;
        RECT 106.950 439.950 109.050 440.400 ;
        RECT 172.950 439.950 175.050 440.400 ;
        RECT 172.950 426.600 175.050 427.050 ;
        RECT 442.950 426.600 445.050 427.050 ;
        RECT 490.950 426.600 493.050 427.050 ;
        RECT 172.950 425.400 493.050 426.600 ;
        RECT 172.950 424.950 175.050 425.400 ;
        RECT 442.950 424.950 445.050 425.400 ;
        RECT 490.950 424.950 493.050 425.400 ;
        RECT 442.950 318.600 445.050 319.050 ;
        RECT 493.950 318.600 496.050 319.050 ;
        RECT 442.950 317.400 496.050 318.600 ;
        RECT 442.950 316.950 445.050 317.400 ;
        RECT 493.950 316.950 496.050 317.400 ;
        RECT 442.950 300.600 445.050 301.050 ;
        RECT 454.950 300.600 457.050 301.050 ;
        RECT 442.950 299.400 457.050 300.600 ;
        RECT 442.950 298.950 445.050 299.400 ;
        RECT 454.950 298.950 457.050 299.400 ;
        RECT 430.950 273.600 433.050 274.050 ;
        RECT 454.950 273.600 457.050 274.050 ;
        RECT 430.950 272.400 457.050 273.600 ;
        RECT 430.950 271.950 433.050 272.400 ;
        RECT 454.950 271.950 457.050 272.400 ;
    END
  END MulL_i
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 707.400 850.050 708.450 873.450 ;
        RECT 706.950 847.950 709.050 850.050 ;
        RECT 709.950 847.950 712.050 850.050 ;
        RECT 730.950 847.950 733.050 850.050 ;
        RECT 710.400 847.050 711.450 847.950 ;
        RECT 709.950 844.950 712.050 847.050 ;
        RECT 731.400 802.050 732.450 847.950 ;
        RECT 730.950 799.950 733.050 802.050 ;
        RECT 775.950 799.950 778.050 802.050 ;
        RECT 776.400 727.050 777.450 799.950 ;
        RECT 775.950 724.950 778.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 785.400 666.450 786.450 724.950 ;
        RECT 782.400 665.400 786.450 666.450 ;
        RECT 782.400 622.050 783.450 665.400 ;
        RECT 781.950 619.950 784.050 622.050 ;
        RECT 805.950 619.950 808.050 622.050 ;
        RECT 806.400 559.050 807.450 619.950 ;
        RECT 805.950 558.450 808.050 559.050 ;
        RECT 803.400 557.400 808.050 558.450 ;
        RECT 803.400 544.050 804.450 557.400 ;
        RECT 805.950 556.950 808.050 557.400 ;
        RECT 802.950 541.950 805.050 544.050 ;
        RECT 817.950 541.950 820.050 544.050 ;
        RECT 818.400 439.050 819.450 541.950 ;
        RECT 823.950 451.950 826.050 454.050 ;
        RECT 824.400 439.050 825.450 451.950 ;
        RECT 817.950 436.950 820.050 439.050 ;
        RECT 823.950 436.950 826.050 439.050 ;
        RECT 818.400 382.050 819.450 436.950 ;
        RECT 805.950 379.950 808.050 382.050 ;
        RECT 817.950 379.950 820.050 382.050 ;
        RECT 823.950 379.950 826.050 382.050 ;
      LAYER metal3 ;
        RECT 706.950 849.600 709.050 850.050 ;
        RECT 709.950 849.600 712.050 850.050 ;
        RECT 730.950 849.600 733.050 850.050 ;
        RECT 706.950 848.400 733.050 849.600 ;
        RECT 706.950 847.950 709.050 848.400 ;
        RECT 709.950 847.950 712.050 848.400 ;
        RECT 730.950 847.950 733.050 848.400 ;
        RECT 730.950 801.600 733.050 802.050 ;
        RECT 775.950 801.600 778.050 802.050 ;
        RECT 730.950 800.400 778.050 801.600 ;
        RECT 730.950 799.950 733.050 800.400 ;
        RECT 775.950 799.950 778.050 800.400 ;
        RECT 775.950 726.600 778.050 727.050 ;
        RECT 784.950 726.600 787.050 727.050 ;
        RECT 775.950 725.400 787.050 726.600 ;
        RECT 775.950 724.950 778.050 725.400 ;
        RECT 784.950 724.950 787.050 725.400 ;
        RECT 781.950 621.600 784.050 622.050 ;
        RECT 805.950 621.600 808.050 622.050 ;
        RECT 781.950 620.400 808.050 621.600 ;
        RECT 781.950 619.950 784.050 620.400 ;
        RECT 805.950 619.950 808.050 620.400 ;
        RECT 802.950 543.600 805.050 544.050 ;
        RECT 817.950 543.600 820.050 544.050 ;
        RECT 802.950 542.400 820.050 543.600 ;
        RECT 802.950 541.950 805.050 542.400 ;
        RECT 817.950 541.950 820.050 542.400 ;
        RECT 817.950 438.600 820.050 439.050 ;
        RECT 823.950 438.600 826.050 439.050 ;
        RECT 817.950 437.400 826.050 438.600 ;
        RECT 817.950 436.950 820.050 437.400 ;
        RECT 823.950 436.950 826.050 437.400 ;
        RECT 805.950 381.600 808.050 382.050 ;
        RECT 817.950 381.600 820.050 382.050 ;
        RECT 823.950 381.600 826.050 382.050 ;
        RECT 805.950 380.400 826.050 381.600 ;
        RECT 805.950 379.950 808.050 380.400 ;
        RECT 817.950 379.950 820.050 380.400 ;
        RECT 823.950 379.950 826.050 380.400 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal2 ;
        RECT 847.950 268.950 850.050 271.050 ;
      LAYER metal3 ;
        RECT 847.950 270.600 850.050 271.050 ;
        RECT 847.950 269.400 879.600 270.600 ;
        RECT 847.950 268.950 850.050 269.400 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 11.400 857.400 13.200 863.250 ;
        RECT 14.700 851.400 16.500 863.250 ;
        RECT 18.900 851.400 20.700 863.250 ;
        RECT 30.300 851.400 32.100 863.250 ;
        RECT 34.500 851.400 36.300 863.250 ;
        RECT 37.800 857.400 39.600 863.250 ;
        RECT 55.650 851.400 57.450 863.250 ;
        RECT 58.650 852.300 60.450 863.250 ;
        RECT 61.650 853.200 63.450 863.250 ;
        RECT 64.650 852.300 66.450 863.250 ;
        RECT 74.550 857.400 76.350 863.250 ;
        RECT 77.550 857.400 79.350 863.250 ;
        RECT 80.550 858.000 82.350 863.250 ;
        RECT 77.700 857.100 79.350 857.400 ;
        RECT 83.550 857.400 85.350 863.250 ;
        RECT 98.400 857.400 100.200 863.250 ;
        RECT 83.550 857.100 84.750 857.400 ;
        RECT 77.700 856.200 84.750 857.100 ;
        RECT 58.650 851.400 66.450 852.300 ;
        RECT 77.100 852.150 78.900 853.950 ;
        RECT 11.250 849.150 13.050 850.950 ;
        RECT 10.950 847.050 13.050 849.150 ;
        RECT 14.850 846.150 16.050 851.400 ;
        RECT 20.100 846.150 21.900 847.950 ;
        RECT 29.100 846.150 30.900 847.950 ;
        RECT 34.950 846.150 36.150 851.400 ;
        RECT 37.950 849.150 39.750 850.950 ;
        RECT 37.950 847.050 40.050 849.150 ;
        RECT 56.100 846.150 57.300 851.400 ;
        RECT 74.100 849.150 75.900 850.950 ;
        RECT 76.950 850.050 79.050 852.150 ;
        RECT 80.250 849.150 82.050 850.950 ;
        RECT 73.950 847.050 76.050 849.150 ;
        RECT 79.950 847.050 82.050 849.150 ;
        RECT 83.700 847.950 84.750 856.200 ;
        RECT 101.700 851.400 103.500 863.250 ;
        RECT 105.900 851.400 107.700 863.250 ;
        RECT 118.650 857.400 120.450 863.250 ;
        RECT 121.650 857.400 123.450 863.250 ;
        RECT 124.650 857.400 126.450 863.250 ;
        RECT 98.250 849.150 100.050 850.950 ;
        RECT 13.950 844.050 16.050 846.150 ;
        RECT 13.950 840.750 15.150 844.050 ;
        RECT 16.950 842.850 19.050 844.950 ;
        RECT 19.950 844.050 22.050 846.150 ;
        RECT 28.950 844.050 31.050 846.150 ;
        RECT 31.950 842.850 34.050 844.950 ;
        RECT 34.950 844.050 37.050 846.150 ;
        RECT 55.950 844.050 58.050 846.150 ;
        RECT 82.950 845.850 85.050 847.950 ;
        RECT 97.950 847.050 100.050 849.150 ;
        RECT 101.850 846.150 103.050 851.400 ;
        RECT 122.250 849.150 123.450 857.400 ;
        RECT 136.650 851.400 138.450 863.250 ;
        RECT 139.650 852.300 141.450 863.250 ;
        RECT 142.650 853.200 144.450 863.250 ;
        RECT 145.650 852.300 147.450 863.250 ;
        RECT 139.650 851.400 147.450 852.300 ;
        RECT 158.550 851.400 160.350 863.250 ;
        RECT 162.750 851.400 164.550 863.250 ;
        RECT 183.150 852.900 184.950 863.250 ;
        RECT 107.100 846.150 108.900 847.950 ;
        RECT 17.100 841.050 18.900 842.850 ;
        RECT 32.100 841.050 33.900 842.850 ;
        RECT 35.850 840.750 37.050 844.050 ;
        RECT 11.250 839.700 15.000 840.750 ;
        RECT 36.000 839.700 39.750 840.750 ;
        RECT 11.250 837.600 12.450 839.700 ;
        RECT 10.650 831.750 12.450 837.600 ;
        RECT 13.650 836.700 21.450 838.050 ;
        RECT 13.650 831.750 15.450 836.700 ;
        RECT 16.650 831.750 18.450 835.800 ;
        RECT 19.650 831.750 21.450 836.700 ;
        RECT 29.550 836.700 37.350 838.050 ;
        RECT 29.550 831.750 31.350 836.700 ;
        RECT 32.550 831.750 34.350 835.800 ;
        RECT 35.550 831.750 37.350 836.700 ;
        RECT 38.550 837.600 39.750 839.700 ;
        RECT 56.100 837.600 57.300 844.050 ;
        RECT 58.950 842.850 61.050 844.950 ;
        RECT 62.100 843.150 63.900 844.950 ;
        RECT 59.100 841.050 60.900 842.850 ;
        RECT 61.950 841.050 64.050 843.150 ;
        RECT 64.950 842.850 67.050 844.950 ;
        RECT 65.100 841.050 66.900 842.850 ;
        RECT 83.400 841.650 84.600 845.850 ;
        RECT 38.550 831.750 40.350 837.600 ;
        RECT 56.100 835.950 61.800 837.600 ;
        RECT 56.700 831.750 58.500 834.600 ;
        RECT 60.000 831.750 61.800 835.950 ;
        RECT 64.200 831.750 66.000 837.600 ;
        RECT 74.700 831.750 76.500 840.600 ;
        RECT 80.100 840.000 84.600 841.650 ;
        RECT 100.950 844.050 103.050 846.150 ;
        RECT 100.950 840.750 102.150 844.050 ;
        RECT 103.950 842.850 106.050 844.950 ;
        RECT 106.950 844.050 109.050 846.150 ;
        RECT 118.950 845.850 121.050 847.950 ;
        RECT 121.950 847.050 124.050 849.150 ;
        RECT 119.100 844.050 120.900 845.850 ;
        RECT 104.100 841.050 105.900 842.850 ;
        RECT 80.100 831.750 81.900 840.000 ;
        RECT 98.250 839.700 102.000 840.750 ;
        RECT 122.250 839.700 123.450 847.050 ;
        RECT 124.950 845.850 127.050 847.950 ;
        RECT 137.100 846.150 138.300 851.400 ;
        RECT 162.000 850.350 164.550 851.400 ;
        RECT 182.550 851.550 184.950 852.900 ;
        RECT 186.150 851.550 187.950 863.250 ;
        RECT 158.100 846.150 159.900 847.950 ;
        RECT 125.100 844.050 126.900 845.850 ;
        RECT 136.950 844.050 139.050 846.150 ;
        RECT 98.250 837.600 99.450 839.700 ;
        RECT 119.850 838.800 123.450 839.700 ;
        RECT 97.650 831.750 99.450 837.600 ;
        RECT 100.650 836.700 108.450 838.050 ;
        RECT 100.650 831.750 102.450 836.700 ;
        RECT 103.650 831.750 105.450 835.800 ;
        RECT 106.650 831.750 108.450 836.700 ;
        RECT 119.850 831.750 121.650 838.800 ;
        RECT 137.100 837.600 138.300 844.050 ;
        RECT 139.950 842.850 142.050 844.950 ;
        RECT 143.100 843.150 144.900 844.950 ;
        RECT 140.100 841.050 141.900 842.850 ;
        RECT 142.950 841.050 145.050 843.150 ;
        RECT 145.950 842.850 148.050 844.950 ;
        RECT 157.950 844.050 160.050 846.150 ;
        RECT 162.000 843.150 163.050 850.350 ;
        RECT 164.100 846.150 165.900 847.950 ;
        RECT 163.950 844.050 166.050 846.150 ;
        RECT 182.550 844.950 183.900 851.550 ;
        RECT 190.650 851.400 192.450 863.250 ;
        RECT 202.050 851.400 203.850 863.250 ;
        RECT 205.050 851.400 206.850 863.250 ;
        RECT 208.650 857.400 210.450 863.250 ;
        RECT 211.650 857.400 213.450 863.250 ;
        RECT 223.650 857.400 225.450 863.250 ;
        RECT 226.650 858.000 228.450 863.250 ;
        RECT 185.250 850.200 187.050 850.650 ;
        RECT 191.250 850.200 192.450 851.400 ;
        RECT 185.250 849.000 192.450 850.200 ;
        RECT 185.250 848.850 187.050 849.000 ;
        RECT 146.100 841.050 147.900 842.850 ;
        RECT 160.950 841.050 163.050 843.150 ;
        RECT 124.350 831.750 126.150 837.600 ;
        RECT 137.100 835.950 142.800 837.600 ;
        RECT 137.700 831.750 139.500 834.600 ;
        RECT 141.000 831.750 142.800 835.950 ;
        RECT 145.200 831.750 147.000 837.600 ;
        RECT 162.000 834.600 163.050 841.050 ;
        RECT 181.950 842.850 184.050 844.950 ;
        RECT 181.950 837.600 183.000 842.850 ;
        RECT 185.400 840.600 186.300 848.850 ;
        RECT 188.100 846.150 189.900 847.950 ;
        RECT 202.650 846.150 203.850 851.400 ;
        RECT 187.950 844.050 190.050 846.150 ;
        RECT 191.100 843.150 192.900 844.950 ;
        RECT 202.650 844.050 205.050 846.150 ;
        RECT 205.950 845.850 208.050 847.950 ;
        RECT 206.100 844.050 207.900 845.850 ;
        RECT 190.950 841.050 193.050 843.150 ;
        RECT 185.250 839.700 187.050 840.600 ;
        RECT 185.250 838.800 188.550 839.700 ;
        RECT 158.550 831.750 160.350 834.600 ;
        RECT 161.550 831.750 163.350 834.600 ;
        RECT 164.550 831.750 166.350 834.600 ;
        RECT 181.650 831.750 183.450 837.600 ;
        RECT 187.650 834.600 188.550 838.800 ;
        RECT 202.650 837.600 203.850 844.050 ;
        RECT 209.100 840.300 210.300 857.400 ;
        RECT 224.250 857.100 225.450 857.400 ;
        RECT 229.650 857.400 231.450 863.250 ;
        RECT 232.650 857.400 234.450 863.250 ;
        RECT 229.650 857.100 231.300 857.400 ;
        RECT 224.250 856.200 231.300 857.100 ;
        RECT 224.250 847.950 225.300 856.200 ;
        RECT 230.100 852.150 231.900 853.950 ;
        RECT 226.950 849.150 228.750 850.950 ;
        RECT 229.950 850.050 232.050 852.150 ;
        RECT 247.650 851.400 249.450 863.250 ;
        RECT 250.650 852.300 252.450 863.250 ;
        RECT 253.650 853.200 255.450 863.250 ;
        RECT 256.650 852.300 258.450 863.250 ;
        RECT 268.650 857.400 270.450 863.250 ;
        RECT 271.650 858.000 273.450 863.250 ;
        RECT 250.650 851.400 258.450 852.300 ;
        RECT 269.250 857.100 270.450 857.400 ;
        RECT 274.650 857.400 276.450 863.250 ;
        RECT 277.650 857.400 279.450 863.250 ;
        RECT 287.550 857.400 289.350 863.250 ;
        RECT 290.550 857.400 292.350 863.250 ;
        RECT 305.400 857.400 307.200 863.250 ;
        RECT 274.650 857.100 276.300 857.400 ;
        RECT 269.250 856.200 276.300 857.100 ;
        RECT 233.100 849.150 234.900 850.950 ;
        RECT 212.100 846.150 213.900 847.950 ;
        RECT 211.950 844.050 214.050 846.150 ;
        RECT 223.950 845.850 226.050 847.950 ;
        RECT 226.950 847.050 229.050 849.150 ;
        RECT 232.950 847.050 235.050 849.150 ;
        RECT 248.100 846.150 249.300 851.400 ;
        RECT 269.250 847.950 270.300 856.200 ;
        RECT 275.100 852.150 276.900 853.950 ;
        RECT 271.950 849.150 273.750 850.950 ;
        RECT 274.950 850.050 277.050 852.150 ;
        RECT 278.100 849.150 279.900 850.950 ;
        RECT 224.400 841.650 225.600 845.850 ;
        RECT 247.950 844.050 250.050 846.150 ;
        RECT 268.950 845.850 271.050 847.950 ;
        RECT 271.950 847.050 274.050 849.150 ;
        RECT 277.950 847.050 280.050 849.150 ;
        RECT 205.950 839.100 213.450 840.300 ;
        RECT 224.400 840.000 228.900 841.650 ;
        RECT 205.950 838.500 207.750 839.100 ;
        RECT 202.650 836.100 205.950 837.600 ;
        RECT 184.650 831.750 186.450 834.600 ;
        RECT 187.650 831.750 189.450 834.600 ;
        RECT 190.650 831.750 192.450 834.600 ;
        RECT 204.150 831.750 205.950 836.100 ;
        RECT 207.150 831.750 208.950 837.600 ;
        RECT 211.650 831.750 213.450 839.100 ;
        RECT 227.100 831.750 228.900 840.000 ;
        RECT 232.500 831.750 234.300 840.600 ;
        RECT 248.100 837.600 249.300 844.050 ;
        RECT 250.950 842.850 253.050 844.950 ;
        RECT 254.100 843.150 255.900 844.950 ;
        RECT 251.100 841.050 252.900 842.850 ;
        RECT 253.950 841.050 256.050 843.150 ;
        RECT 256.950 842.850 259.050 844.950 ;
        RECT 257.100 841.050 258.900 842.850 ;
        RECT 269.400 841.650 270.600 845.850 ;
        RECT 290.400 844.950 291.600 857.400 ;
        RECT 308.700 851.400 310.500 863.250 ;
        RECT 312.900 851.400 314.700 863.250 ;
        RECT 324.300 851.400 326.100 863.250 ;
        RECT 328.500 851.400 330.300 863.250 ;
        RECT 331.800 857.400 333.600 863.250 ;
        RECT 344.550 852.300 346.350 863.250 ;
        RECT 347.550 853.200 349.350 863.250 ;
        RECT 350.550 852.300 352.350 863.250 ;
        RECT 344.550 851.400 352.350 852.300 ;
        RECT 353.550 851.400 355.350 863.250 ;
        RECT 367.650 857.400 369.450 863.250 ;
        RECT 370.650 857.400 372.450 863.250 ;
        RECT 373.650 857.400 375.450 863.250 ;
        RECT 385.650 857.400 387.450 863.250 ;
        RECT 388.650 858.000 390.450 863.250 ;
        RECT 305.250 849.150 307.050 850.950 ;
        RECT 304.950 847.050 307.050 849.150 ;
        RECT 308.850 846.150 310.050 851.400 ;
        RECT 314.100 846.150 315.900 847.950 ;
        RECT 323.100 846.150 324.900 847.950 ;
        RECT 328.950 846.150 330.150 851.400 ;
        RECT 331.950 849.150 333.750 850.950 ;
        RECT 331.950 847.050 334.050 849.150 ;
        RECT 353.700 846.150 354.900 851.400 ;
        RECT 371.250 849.150 372.450 857.400 ;
        RECT 386.250 857.100 387.450 857.400 ;
        RECT 391.650 857.400 393.450 863.250 ;
        RECT 394.650 857.400 396.450 863.250 ;
        RECT 406.650 857.400 408.450 863.250 ;
        RECT 409.650 858.000 411.450 863.250 ;
        RECT 391.650 857.100 393.300 857.400 ;
        RECT 386.250 856.200 393.300 857.100 ;
        RECT 407.250 857.100 408.450 857.400 ;
        RECT 412.650 857.400 414.450 863.250 ;
        RECT 415.650 857.400 417.450 863.250 ;
        RECT 425.550 857.400 427.350 863.250 ;
        RECT 428.550 857.400 430.350 863.250 ;
        RECT 431.550 857.400 433.350 863.250 ;
        RECT 445.650 857.400 447.450 863.250 ;
        RECT 448.650 857.400 450.450 863.250 ;
        RECT 461.400 857.400 463.200 863.250 ;
        RECT 412.650 857.100 414.300 857.400 ;
        RECT 407.250 856.200 414.300 857.100 ;
        RECT 287.100 843.150 288.900 844.950 ;
        RECT 269.400 840.000 273.900 841.650 ;
        RECT 286.950 841.050 289.050 843.150 ;
        RECT 289.950 842.850 292.050 844.950 ;
        RECT 307.950 844.050 310.050 846.150 ;
        RECT 248.100 835.950 253.800 837.600 ;
        RECT 248.700 831.750 250.500 834.600 ;
        RECT 252.000 831.750 253.800 835.950 ;
        RECT 256.200 831.750 258.000 837.600 ;
        RECT 272.100 831.750 273.900 840.000 ;
        RECT 277.500 831.750 279.300 840.600 ;
        RECT 290.400 834.600 291.600 842.850 ;
        RECT 307.950 840.750 309.150 844.050 ;
        RECT 310.950 842.850 313.050 844.950 ;
        RECT 313.950 844.050 316.050 846.150 ;
        RECT 322.950 844.050 325.050 846.150 ;
        RECT 325.950 842.850 328.050 844.950 ;
        RECT 328.950 844.050 331.050 846.150 ;
        RECT 311.100 841.050 312.900 842.850 ;
        RECT 326.100 841.050 327.900 842.850 ;
        RECT 329.850 840.750 331.050 844.050 ;
        RECT 343.950 842.850 346.050 844.950 ;
        RECT 347.100 843.150 348.900 844.950 ;
        RECT 344.100 841.050 345.900 842.850 ;
        RECT 346.950 841.050 349.050 843.150 ;
        RECT 349.950 842.850 352.050 844.950 ;
        RECT 352.950 844.050 355.050 846.150 ;
        RECT 367.950 845.850 370.050 847.950 ;
        RECT 370.950 847.050 373.050 849.150 ;
        RECT 386.250 847.950 387.300 856.200 ;
        RECT 392.100 852.150 393.900 853.950 ;
        RECT 388.950 849.150 390.750 850.950 ;
        RECT 391.950 850.050 394.050 852.150 ;
        RECT 395.100 849.150 396.900 850.950 ;
        RECT 368.100 844.050 369.900 845.850 ;
        RECT 350.100 841.050 351.900 842.850 ;
        RECT 305.250 839.700 309.000 840.750 ;
        RECT 330.000 839.700 333.750 840.750 ;
        RECT 305.250 837.600 306.450 839.700 ;
        RECT 287.550 831.750 289.350 834.600 ;
        RECT 290.550 831.750 292.350 834.600 ;
        RECT 304.650 831.750 306.450 837.600 ;
        RECT 307.650 836.700 315.450 838.050 ;
        RECT 307.650 831.750 309.450 836.700 ;
        RECT 310.650 831.750 312.450 835.800 ;
        RECT 313.650 831.750 315.450 836.700 ;
        RECT 323.550 836.700 331.350 838.050 ;
        RECT 323.550 831.750 325.350 836.700 ;
        RECT 326.550 831.750 328.350 835.800 ;
        RECT 329.550 831.750 331.350 836.700 ;
        RECT 332.550 837.600 333.750 839.700 ;
        RECT 353.700 837.600 354.900 844.050 ;
        RECT 371.250 839.700 372.450 847.050 ;
        RECT 373.950 845.850 376.050 847.950 ;
        RECT 385.950 845.850 388.050 847.950 ;
        RECT 388.950 847.050 391.050 849.150 ;
        RECT 394.950 847.050 397.050 849.150 ;
        RECT 407.250 847.950 408.300 856.200 ;
        RECT 413.100 852.150 414.900 853.950 ;
        RECT 409.950 849.150 411.750 850.950 ;
        RECT 412.950 850.050 415.050 852.150 ;
        RECT 416.100 849.150 417.900 850.950 ;
        RECT 428.550 849.150 429.750 857.400 ;
        RECT 406.950 845.850 409.050 847.950 ;
        RECT 409.950 847.050 412.050 849.150 ;
        RECT 415.950 847.050 418.050 849.150 ;
        RECT 424.950 845.850 427.050 847.950 ;
        RECT 427.950 847.050 430.050 849.150 ;
        RECT 374.100 844.050 375.900 845.850 ;
        RECT 386.400 841.650 387.600 845.850 ;
        RECT 407.400 841.650 408.600 845.850 ;
        RECT 425.100 844.050 426.900 845.850 ;
        RECT 386.400 840.000 390.900 841.650 ;
        RECT 332.550 831.750 334.350 837.600 ;
        RECT 345.000 831.750 346.800 837.600 ;
        RECT 349.200 835.950 354.900 837.600 ;
        RECT 368.850 838.800 372.450 839.700 ;
        RECT 349.200 831.750 351.000 835.950 ;
        RECT 352.500 831.750 354.300 834.600 ;
        RECT 368.850 831.750 370.650 838.800 ;
        RECT 373.350 831.750 375.150 837.600 ;
        RECT 389.100 831.750 390.900 840.000 ;
        RECT 394.500 831.750 396.300 840.600 ;
        RECT 407.400 840.000 411.900 841.650 ;
        RECT 410.100 831.750 411.900 840.000 ;
        RECT 415.500 831.750 417.300 840.600 ;
        RECT 428.550 839.700 429.750 847.050 ;
        RECT 430.950 845.850 433.050 847.950 ;
        RECT 431.100 844.050 432.900 845.850 ;
        RECT 446.400 844.950 447.600 857.400 ;
        RECT 464.700 851.400 466.500 863.250 ;
        RECT 468.900 851.400 470.700 863.250 ;
        RECT 484.050 851.400 485.850 863.250 ;
        RECT 487.050 851.400 488.850 863.250 ;
        RECT 490.650 857.400 492.450 863.250 ;
        RECT 493.650 857.400 495.450 863.250 ;
        RECT 461.250 849.150 463.050 850.950 ;
        RECT 460.950 847.050 463.050 849.150 ;
        RECT 464.850 846.150 466.050 851.400 ;
        RECT 470.100 846.150 471.900 847.950 ;
        RECT 484.650 846.150 485.850 851.400 ;
        RECT 445.950 842.850 448.050 844.950 ;
        RECT 449.100 843.150 450.900 844.950 ;
        RECT 463.950 844.050 466.050 846.150 ;
        RECT 428.550 838.800 432.150 839.700 ;
        RECT 425.850 831.750 427.650 837.600 ;
        RECT 430.350 831.750 432.150 838.800 ;
        RECT 446.400 834.600 447.600 842.850 ;
        RECT 448.950 841.050 451.050 843.150 ;
        RECT 463.950 840.750 465.150 844.050 ;
        RECT 466.950 842.850 469.050 844.950 ;
        RECT 469.950 844.050 472.050 846.150 ;
        RECT 484.650 844.050 487.050 846.150 ;
        RECT 487.950 845.850 490.050 847.950 ;
        RECT 488.100 844.050 489.900 845.850 ;
        RECT 467.100 841.050 468.900 842.850 ;
        RECT 461.250 839.700 465.000 840.750 ;
        RECT 461.250 837.600 462.450 839.700 ;
        RECT 445.650 831.750 447.450 834.600 ;
        RECT 448.650 831.750 450.450 834.600 ;
        RECT 460.650 831.750 462.450 837.600 ;
        RECT 463.650 836.700 471.450 838.050 ;
        RECT 463.650 831.750 465.450 836.700 ;
        RECT 466.650 831.750 468.450 835.800 ;
        RECT 469.650 831.750 471.450 836.700 ;
        RECT 484.650 837.600 485.850 844.050 ;
        RECT 491.100 840.300 492.300 857.400 ;
        RECT 507.450 851.400 509.250 863.250 ;
        RECT 511.650 851.400 513.450 863.250 ;
        RECT 523.650 857.400 525.450 863.250 ;
        RECT 526.650 858.000 528.450 863.250 ;
        RECT 524.250 857.100 525.450 857.400 ;
        RECT 529.650 857.400 531.450 863.250 ;
        RECT 532.650 857.400 534.450 863.250 ;
        RECT 547.650 857.400 549.450 863.250 ;
        RECT 550.650 857.400 552.450 863.250 ;
        RECT 562.650 857.400 564.450 863.250 ;
        RECT 565.650 857.400 567.450 863.250 ;
        RECT 575.550 857.400 577.350 863.250 ;
        RECT 578.550 857.400 580.350 863.250 ;
        RECT 529.650 857.100 531.300 857.400 ;
        RECT 524.250 856.200 531.300 857.100 ;
        RECT 507.450 850.350 510.000 851.400 ;
        RECT 494.100 846.150 495.900 847.950 ;
        RECT 506.100 846.150 507.900 847.950 ;
        RECT 493.950 844.050 496.050 846.150 ;
        RECT 505.950 844.050 508.050 846.150 ;
        RECT 508.950 843.150 510.000 850.350 ;
        RECT 524.250 847.950 525.300 856.200 ;
        RECT 530.100 852.150 531.900 853.950 ;
        RECT 526.950 849.150 528.750 850.950 ;
        RECT 529.950 850.050 532.050 852.150 ;
        RECT 533.100 849.150 534.900 850.950 ;
        RECT 512.100 846.150 513.900 847.950 ;
        RECT 511.950 844.050 514.050 846.150 ;
        RECT 523.950 845.850 526.050 847.950 ;
        RECT 526.950 847.050 529.050 849.150 ;
        RECT 532.950 847.050 535.050 849.150 ;
        RECT 508.950 841.050 511.050 843.150 ;
        RECT 524.400 841.650 525.600 845.850 ;
        RECT 548.400 844.950 549.600 857.400 ;
        RECT 563.400 844.950 564.600 857.400 ;
        RECT 578.400 844.950 579.600 857.400 ;
        RECT 591.300 851.400 593.100 863.250 ;
        RECT 595.500 851.400 597.300 863.250 ;
        RECT 598.800 857.400 600.600 863.250 ;
        RECT 611.550 857.400 613.350 863.250 ;
        RECT 614.550 857.400 616.350 863.250 ;
        RECT 590.100 846.150 591.900 847.950 ;
        RECT 595.950 846.150 597.150 851.400 ;
        RECT 598.950 849.150 600.750 850.950 ;
        RECT 598.950 847.050 601.050 849.150 ;
        RECT 547.950 842.850 550.050 844.950 ;
        RECT 551.100 843.150 552.900 844.950 ;
        RECT 487.950 839.100 495.450 840.300 ;
        RECT 487.950 838.500 489.750 839.100 ;
        RECT 484.650 836.100 487.950 837.600 ;
        RECT 486.150 831.750 487.950 836.100 ;
        RECT 489.150 831.750 490.950 837.600 ;
        RECT 493.650 831.750 495.450 839.100 ;
        RECT 508.950 834.600 510.000 841.050 ;
        RECT 524.400 840.000 528.900 841.650 ;
        RECT 505.650 831.750 507.450 834.600 ;
        RECT 508.650 831.750 510.450 834.600 ;
        RECT 511.650 831.750 513.450 834.600 ;
        RECT 527.100 831.750 528.900 840.000 ;
        RECT 532.500 831.750 534.300 840.600 ;
        RECT 548.400 834.600 549.600 842.850 ;
        RECT 550.950 841.050 553.050 843.150 ;
        RECT 562.950 842.850 565.050 844.950 ;
        RECT 566.100 843.150 567.900 844.950 ;
        RECT 575.100 843.150 576.900 844.950 ;
        RECT 563.400 834.600 564.600 842.850 ;
        RECT 565.950 841.050 568.050 843.150 ;
        RECT 574.950 841.050 577.050 843.150 ;
        RECT 577.950 842.850 580.050 844.950 ;
        RECT 589.950 844.050 592.050 846.150 ;
        RECT 592.950 842.850 595.050 844.950 ;
        RECT 595.950 844.050 598.050 846.150 ;
        RECT 614.400 844.950 615.600 857.400 ;
        RECT 620.550 851.400 622.350 863.250 ;
        RECT 623.550 860.400 625.350 863.250 ;
        RECT 628.050 857.400 629.850 863.250 ;
        RECT 632.250 857.400 634.050 863.250 ;
        RECT 625.950 855.300 629.850 857.400 ;
        RECT 636.150 856.500 637.950 863.250 ;
        RECT 639.150 857.400 640.950 863.250 ;
        RECT 643.950 857.400 645.750 863.250 ;
        RECT 649.050 857.400 650.850 863.250 ;
        RECT 644.250 856.500 645.450 857.400 ;
        RECT 634.950 854.700 641.850 856.500 ;
        RECT 644.250 854.400 649.050 856.500 ;
        RECT 627.150 852.600 629.850 854.400 ;
        RECT 630.750 853.800 632.550 854.400 ;
        RECT 630.750 852.900 637.050 853.800 ;
        RECT 644.250 853.500 645.450 854.400 ;
        RECT 630.750 852.600 632.550 852.900 ;
        RECT 628.950 851.700 629.850 852.600 ;
        RECT 578.400 834.600 579.600 842.850 ;
        RECT 593.100 841.050 594.900 842.850 ;
        RECT 596.850 840.750 598.050 844.050 ;
        RECT 611.100 843.150 612.900 844.950 ;
        RECT 610.950 841.050 613.050 843.150 ;
        RECT 613.950 842.850 616.050 844.950 ;
        RECT 597.000 839.700 600.750 840.750 ;
        RECT 590.550 836.700 598.350 838.050 ;
        RECT 547.650 831.750 549.450 834.600 ;
        RECT 550.650 831.750 552.450 834.600 ;
        RECT 562.650 831.750 564.450 834.600 ;
        RECT 565.650 831.750 567.450 834.600 ;
        RECT 575.550 831.750 577.350 834.600 ;
        RECT 578.550 831.750 580.350 834.600 ;
        RECT 590.550 831.750 592.350 836.700 ;
        RECT 593.550 831.750 595.350 835.800 ;
        RECT 596.550 831.750 598.350 836.700 ;
        RECT 599.550 837.600 600.750 839.700 ;
        RECT 599.550 831.750 601.350 837.600 ;
        RECT 614.400 834.600 615.600 842.850 ;
        RECT 620.550 841.950 621.750 851.400 ;
        RECT 625.950 850.800 628.050 851.700 ;
        RECT 628.950 850.800 634.950 851.700 ;
        RECT 623.850 849.600 628.050 850.800 ;
        RECT 622.950 847.800 624.750 849.600 ;
        RECT 634.050 846.150 634.950 850.800 ;
        RECT 636.150 850.800 637.050 852.900 ;
        RECT 637.950 852.300 645.450 853.500 ;
        RECT 637.950 851.700 639.750 852.300 ;
        RECT 652.050 851.400 653.850 863.250 ;
        RECT 668.400 857.400 670.200 863.250 ;
        RECT 671.700 851.400 673.500 863.250 ;
        RECT 675.900 851.400 677.700 863.250 ;
        RECT 688.650 851.400 690.450 863.250 ;
        RECT 642.750 850.800 653.850 851.400 ;
        RECT 636.150 850.200 653.850 850.800 ;
        RECT 636.150 849.900 644.550 850.200 ;
        RECT 642.750 849.600 644.550 849.900 ;
        RECT 634.050 844.050 637.050 846.150 ;
        RECT 640.950 845.100 643.050 846.150 ;
        RECT 640.950 844.050 648.900 845.100 ;
        RECT 622.950 843.750 625.050 844.050 ;
        RECT 622.950 841.950 626.850 843.750 ;
        RECT 620.550 839.850 625.050 841.950 ;
        RECT 634.050 840.000 634.950 844.050 ;
        RECT 647.100 843.300 648.900 844.050 ;
        RECT 650.100 843.150 651.900 844.950 ;
        RECT 644.100 842.400 645.900 843.000 ;
        RECT 650.100 842.400 651.000 843.150 ;
        RECT 644.100 841.200 651.000 842.400 ;
        RECT 644.100 840.000 645.150 841.200 ;
        RECT 620.550 837.600 621.750 839.850 ;
        RECT 634.050 839.100 645.150 840.000 ;
        RECT 634.050 838.800 634.950 839.100 ;
        RECT 611.550 831.750 613.350 834.600 ;
        RECT 614.550 831.750 616.350 834.600 ;
        RECT 620.550 831.750 622.350 837.600 ;
        RECT 625.950 836.700 628.050 837.600 ;
        RECT 633.150 837.000 634.950 838.800 ;
        RECT 644.100 838.200 645.150 839.100 ;
        RECT 640.350 837.450 642.150 838.200 ;
        RECT 625.950 835.500 629.700 836.700 ;
        RECT 628.650 834.600 629.700 835.500 ;
        RECT 637.200 836.400 642.150 837.450 ;
        RECT 643.650 836.400 645.450 838.200 ;
        RECT 652.950 837.600 653.850 850.200 ;
        RECT 668.250 849.150 670.050 850.950 ;
        RECT 667.950 847.050 670.050 849.150 ;
        RECT 671.850 846.150 673.050 851.400 ;
        RECT 691.650 850.500 693.450 863.250 ;
        RECT 694.650 851.400 696.450 863.250 ;
        RECT 697.650 850.500 699.450 863.250 ;
        RECT 700.650 851.400 702.450 863.250 ;
        RECT 703.650 850.500 705.450 863.250 ;
        RECT 706.650 851.400 708.450 863.250 ;
        RECT 709.650 850.500 711.450 863.250 ;
        RECT 712.650 851.400 714.450 863.250 ;
        RECT 724.650 857.400 726.450 863.250 ;
        RECT 727.650 857.400 729.450 863.250 ;
        RECT 740.400 857.400 742.200 863.250 ;
        RECT 690.750 849.300 693.450 850.500 ;
        RECT 695.700 849.300 699.450 850.500 ;
        RECT 701.700 849.300 705.450 850.500 ;
        RECT 707.550 849.300 711.450 850.500 ;
        RECT 677.100 846.150 678.900 847.950 ;
        RECT 670.950 844.050 673.050 846.150 ;
        RECT 670.950 840.750 672.150 844.050 ;
        RECT 673.950 842.850 676.050 844.950 ;
        RECT 676.950 844.050 679.050 846.150 ;
        RECT 690.750 844.950 691.800 849.300 ;
        RECT 688.950 842.850 691.800 844.950 ;
        RECT 674.100 841.050 675.900 842.850 ;
        RECT 668.250 839.700 672.000 840.750 ;
        RECT 690.750 839.700 691.800 842.850 ;
        RECT 695.700 842.400 696.900 849.300 ;
        RECT 701.700 842.400 702.900 849.300 ;
        RECT 707.550 842.400 708.750 849.300 ;
        RECT 725.400 844.950 726.600 857.400 ;
        RECT 743.700 851.400 745.500 863.250 ;
        RECT 747.900 851.400 749.700 863.250 ;
        RECT 760.650 857.400 762.450 863.250 ;
        RECT 763.650 857.400 765.450 863.250 ;
        RECT 766.650 857.400 768.450 863.250 ;
        RECT 776.550 857.400 778.350 863.250 ;
        RECT 779.550 857.400 781.350 863.250 ;
        RECT 782.550 857.400 784.350 863.250 ;
        RECT 740.250 849.150 742.050 850.950 ;
        RECT 739.950 847.050 742.050 849.150 ;
        RECT 743.850 846.150 745.050 851.400 ;
        RECT 764.250 849.150 765.450 857.400 ;
        RECT 779.550 849.150 780.750 857.400 ;
        RECT 795.300 851.400 797.100 863.250 ;
        RECT 799.500 851.400 801.300 863.250 ;
        RECT 802.800 857.400 804.600 863.250 ;
        RECT 815.550 857.400 817.350 863.250 ;
        RECT 818.550 857.400 820.350 863.250 ;
        RECT 830.550 857.400 832.350 863.250 ;
        RECT 833.550 857.400 835.350 863.250 ;
        RECT 836.550 857.400 838.350 863.250 ;
        RECT 848.550 857.400 850.350 863.250 ;
        RECT 851.550 857.400 853.350 863.250 ;
        RECT 749.100 846.150 750.900 847.950 ;
        RECT 709.950 842.850 712.050 844.950 ;
        RECT 724.950 842.850 727.050 844.950 ;
        RECT 728.100 843.150 729.900 844.950 ;
        RECT 742.950 844.050 745.050 846.150 ;
        RECT 692.700 840.600 696.900 842.400 ;
        RECT 698.700 840.600 702.900 842.400 ;
        RECT 704.700 840.600 708.750 842.400 ;
        RECT 710.100 841.050 711.900 842.850 ;
        RECT 695.700 839.700 696.900 840.600 ;
        RECT 701.700 839.700 702.900 840.600 ;
        RECT 707.550 839.700 708.750 840.600 ;
        RECT 668.250 837.600 669.450 839.700 ;
        RECT 690.750 838.650 693.600 839.700 ;
        RECT 690.900 838.500 693.600 838.650 ;
        RECT 695.700 838.500 699.600 839.700 ;
        RECT 701.700 838.500 705.450 839.700 ;
        RECT 707.550 838.500 711.600 839.700 ;
        RECT 637.200 834.600 638.250 836.400 ;
        RECT 646.950 835.500 649.050 837.600 ;
        RECT 646.950 834.600 648.000 835.500 ;
        RECT 623.850 831.750 625.650 834.600 ;
        RECT 628.350 831.750 630.150 834.600 ;
        RECT 632.550 831.750 634.350 834.600 ;
        RECT 636.450 831.750 638.250 834.600 ;
        RECT 639.750 831.750 641.550 834.600 ;
        RECT 644.250 833.700 648.000 834.600 ;
        RECT 644.250 831.750 646.050 833.700 ;
        RECT 649.050 831.750 650.850 834.600 ;
        RECT 652.050 831.750 653.850 837.600 ;
        RECT 667.650 831.750 669.450 837.600 ;
        RECT 670.650 836.700 678.450 838.050 ;
        RECT 691.800 837.600 693.600 838.500 ;
        RECT 697.800 837.600 699.600 838.500 ;
        RECT 670.650 831.750 672.450 836.700 ;
        RECT 673.650 831.750 675.450 835.800 ;
        RECT 676.650 831.750 678.450 836.700 ;
        RECT 688.650 831.750 690.450 837.600 ;
        RECT 691.650 831.750 693.450 837.600 ;
        RECT 694.650 831.750 696.450 837.600 ;
        RECT 697.650 831.750 699.450 837.600 ;
        RECT 700.650 831.750 702.450 837.600 ;
        RECT 703.650 831.750 705.450 838.500 ;
        RECT 709.800 837.600 711.600 838.500 ;
        RECT 706.650 831.750 708.450 837.600 ;
        RECT 709.650 831.750 711.450 837.600 ;
        RECT 712.650 831.750 714.450 837.600 ;
        RECT 725.400 834.600 726.600 842.850 ;
        RECT 727.950 841.050 730.050 843.150 ;
        RECT 742.950 840.750 744.150 844.050 ;
        RECT 745.950 842.850 748.050 844.950 ;
        RECT 748.950 844.050 751.050 846.150 ;
        RECT 760.950 845.850 763.050 847.950 ;
        RECT 763.950 847.050 766.050 849.150 ;
        RECT 761.100 844.050 762.900 845.850 ;
        RECT 746.100 841.050 747.900 842.850 ;
        RECT 740.250 839.700 744.000 840.750 ;
        RECT 764.250 839.700 765.450 847.050 ;
        RECT 766.950 845.850 769.050 847.950 ;
        RECT 775.950 845.850 778.050 847.950 ;
        RECT 778.950 847.050 781.050 849.150 ;
        RECT 767.100 844.050 768.900 845.850 ;
        RECT 776.100 844.050 777.900 845.850 ;
        RECT 740.250 837.600 741.450 839.700 ;
        RECT 761.850 838.800 765.450 839.700 ;
        RECT 779.550 839.700 780.750 847.050 ;
        RECT 781.950 845.850 784.050 847.950 ;
        RECT 794.100 846.150 795.900 847.950 ;
        RECT 799.950 846.150 801.150 851.400 ;
        RECT 802.950 849.150 804.750 850.950 ;
        RECT 802.950 847.050 805.050 849.150 ;
        RECT 782.100 844.050 783.900 845.850 ;
        RECT 793.950 844.050 796.050 846.150 ;
        RECT 796.950 842.850 799.050 844.950 ;
        RECT 799.950 844.050 802.050 846.150 ;
        RECT 818.400 844.950 819.600 857.400 ;
        RECT 833.550 849.150 834.750 857.400 ;
        RECT 829.950 845.850 832.050 847.950 ;
        RECT 832.950 847.050 835.050 849.150 ;
        RECT 797.100 841.050 798.900 842.850 ;
        RECT 800.850 840.750 802.050 844.050 ;
        RECT 815.100 843.150 816.900 844.950 ;
        RECT 814.950 841.050 817.050 843.150 ;
        RECT 817.950 842.850 820.050 844.950 ;
        RECT 830.100 844.050 831.900 845.850 ;
        RECT 801.000 839.700 804.750 840.750 ;
        RECT 779.550 838.800 783.150 839.700 ;
        RECT 724.650 831.750 726.450 834.600 ;
        RECT 727.650 831.750 729.450 834.600 ;
        RECT 739.650 831.750 741.450 837.600 ;
        RECT 742.650 836.700 750.450 838.050 ;
        RECT 742.650 831.750 744.450 836.700 ;
        RECT 745.650 831.750 747.450 835.800 ;
        RECT 748.650 831.750 750.450 836.700 ;
        RECT 761.850 831.750 763.650 838.800 ;
        RECT 766.350 831.750 768.150 837.600 ;
        RECT 776.850 831.750 778.650 837.600 ;
        RECT 781.350 831.750 783.150 838.800 ;
        RECT 794.550 836.700 802.350 838.050 ;
        RECT 794.550 831.750 796.350 836.700 ;
        RECT 797.550 831.750 799.350 835.800 ;
        RECT 800.550 831.750 802.350 836.700 ;
        RECT 803.550 837.600 804.750 839.700 ;
        RECT 803.550 831.750 805.350 837.600 ;
        RECT 818.400 834.600 819.600 842.850 ;
        RECT 833.550 839.700 834.750 847.050 ;
        RECT 835.950 845.850 838.050 847.950 ;
        RECT 836.100 844.050 837.900 845.850 ;
        RECT 851.400 844.950 852.600 857.400 ;
        RECT 848.100 843.150 849.900 844.950 ;
        RECT 847.950 841.050 850.050 843.150 ;
        RECT 850.950 842.850 853.050 844.950 ;
        RECT 833.550 838.800 837.150 839.700 ;
        RECT 815.550 831.750 817.350 834.600 ;
        RECT 818.550 831.750 820.350 834.600 ;
        RECT 830.850 831.750 832.650 837.600 ;
        RECT 835.350 831.750 837.150 838.800 ;
        RECT 851.400 834.600 852.600 842.850 ;
        RECT 848.550 831.750 850.350 834.600 ;
        RECT 851.550 831.750 853.350 834.600 ;
        RECT 10.650 821.400 12.450 827.250 ;
        RECT 11.250 819.300 12.450 821.400 ;
        RECT 13.650 822.300 15.450 827.250 ;
        RECT 16.650 823.200 18.450 827.250 ;
        RECT 19.650 822.300 21.450 827.250 ;
        RECT 13.650 820.950 21.450 822.300 ;
        RECT 11.250 818.250 15.000 819.300 ;
        RECT 38.100 819.000 39.900 827.250 ;
        RECT 13.950 814.950 15.150 818.250 ;
        RECT 17.100 816.150 18.900 817.950 ;
        RECT 35.400 817.350 39.900 819.000 ;
        RECT 43.500 818.400 45.300 827.250 ;
        RECT 59.100 819.000 60.900 827.250 ;
        RECT 56.400 817.350 60.900 819.000 ;
        RECT 64.500 818.400 66.300 827.250 ;
        RECT 80.100 819.000 81.900 827.250 ;
        RECT 77.400 817.350 81.900 819.000 ;
        RECT 85.500 818.400 87.300 827.250 ;
        RECT 98.700 818.400 100.500 827.250 ;
        RECT 104.100 819.000 105.900 827.250 ;
        RECT 119.550 822.300 121.350 827.250 ;
        RECT 122.550 823.200 124.350 827.250 ;
        RECT 125.550 822.300 127.350 827.250 ;
        RECT 119.550 820.950 127.350 822.300 ;
        RECT 128.550 821.400 130.350 827.250 ;
        RECT 128.550 819.300 129.750 821.400 ;
        RECT 104.100 817.350 108.600 819.000 ;
        RECT 126.000 818.250 129.750 819.300 ;
        RECT 140.700 818.400 142.500 827.250 ;
        RECT 146.100 819.000 147.900 827.250 ;
        RECT 164.700 824.400 166.500 827.250 ;
        RECT 168.000 823.050 169.800 827.250 ;
        RECT 164.100 821.400 169.800 823.050 ;
        RECT 172.200 821.400 174.000 827.250 ;
        RECT 13.950 812.850 16.050 814.950 ;
        RECT 16.950 814.050 19.050 816.150 ;
        RECT 19.950 812.850 22.050 814.950 ;
        RECT 35.400 813.150 36.600 817.350 ;
        RECT 56.400 813.150 57.600 817.350 ;
        RECT 77.400 813.150 78.600 817.350 ;
        RECT 107.400 813.150 108.600 817.350 ;
        RECT 122.100 816.150 123.900 817.950 ;
        RECT 10.950 809.850 13.050 811.950 ;
        RECT 11.250 808.050 13.050 809.850 ;
        RECT 14.850 807.600 16.050 812.850 ;
        RECT 20.100 811.050 21.900 812.850 ;
        RECT 34.950 811.050 37.050 813.150 ;
        RECT 11.400 795.750 13.200 801.600 ;
        RECT 14.700 795.750 16.500 807.600 ;
        RECT 18.900 795.750 20.700 807.600 ;
        RECT 35.250 802.800 36.300 811.050 ;
        RECT 37.950 809.850 40.050 811.950 ;
        RECT 43.950 809.850 46.050 811.950 ;
        RECT 55.950 811.050 58.050 813.150 ;
        RECT 37.950 808.050 39.750 809.850 ;
        RECT 40.950 806.850 43.050 808.950 ;
        RECT 44.100 808.050 45.900 809.850 ;
        RECT 41.100 805.050 42.900 806.850 ;
        RECT 56.250 802.800 57.300 811.050 ;
        RECT 58.950 809.850 61.050 811.950 ;
        RECT 64.950 809.850 67.050 811.950 ;
        RECT 76.950 811.050 79.050 813.150 ;
        RECT 58.950 808.050 60.750 809.850 ;
        RECT 61.950 806.850 64.050 808.950 ;
        RECT 65.100 808.050 66.900 809.850 ;
        RECT 62.100 805.050 63.900 806.850 ;
        RECT 77.250 802.800 78.300 811.050 ;
        RECT 79.950 809.850 82.050 811.950 ;
        RECT 85.950 809.850 88.050 811.950 ;
        RECT 97.950 809.850 100.050 811.950 ;
        RECT 103.950 809.850 106.050 811.950 ;
        RECT 106.950 811.050 109.050 813.150 ;
        RECT 118.950 812.850 121.050 814.950 ;
        RECT 121.950 814.050 124.050 816.150 ;
        RECT 125.850 814.950 127.050 818.250 ;
        RECT 146.100 817.350 150.600 819.000 ;
        RECT 124.950 812.850 127.050 814.950 ;
        RECT 149.400 813.150 150.600 817.350 ;
        RECT 164.100 814.950 165.300 821.400 ;
        RECT 182.700 818.400 184.500 827.250 ;
        RECT 188.100 819.000 189.900 827.250 ;
        RECT 206.550 824.400 208.350 827.250 ;
        RECT 209.550 824.400 211.350 827.250 ;
        RECT 212.550 824.400 214.350 827.250 ;
        RECT 167.100 816.150 168.900 817.950 ;
        RECT 119.100 811.050 120.900 812.850 ;
        RECT 79.950 808.050 81.750 809.850 ;
        RECT 82.950 806.850 85.050 808.950 ;
        RECT 86.100 808.050 87.900 809.850 ;
        RECT 98.100 808.050 99.900 809.850 ;
        RECT 100.950 806.850 103.050 808.950 ;
        RECT 104.250 808.050 106.050 809.850 ;
        RECT 83.100 805.050 84.900 806.850 ;
        RECT 101.100 805.050 102.900 806.850 ;
        RECT 107.700 802.800 108.750 811.050 ;
        RECT 124.950 807.600 126.150 812.850 ;
        RECT 127.950 809.850 130.050 811.950 ;
        RECT 139.950 809.850 142.050 811.950 ;
        RECT 145.950 809.850 148.050 811.950 ;
        RECT 148.950 811.050 151.050 813.150 ;
        RECT 163.950 812.850 166.050 814.950 ;
        RECT 166.950 814.050 169.050 816.150 ;
        RECT 169.950 815.850 172.050 817.950 ;
        RECT 173.100 816.150 174.900 817.950 ;
        RECT 188.100 817.350 192.600 819.000 ;
        RECT 210.000 817.950 211.050 824.400 ;
        RECT 230.100 819.000 231.900 827.250 ;
        RECT 170.100 814.050 171.900 815.850 ;
        RECT 172.950 814.050 175.050 816.150 ;
        RECT 191.400 813.150 192.600 817.350 ;
        RECT 208.950 815.850 211.050 817.950 ;
        RECT 127.950 808.050 129.750 809.850 ;
        RECT 140.100 808.050 141.900 809.850 ;
        RECT 35.250 801.900 42.300 802.800 ;
        RECT 35.250 801.600 36.450 801.900 ;
        RECT 34.650 795.750 36.450 801.600 ;
        RECT 40.650 801.600 42.300 801.900 ;
        RECT 56.250 801.900 63.300 802.800 ;
        RECT 56.250 801.600 57.450 801.900 ;
        RECT 37.650 795.750 39.450 801.000 ;
        RECT 40.650 795.750 42.450 801.600 ;
        RECT 43.650 795.750 45.450 801.600 ;
        RECT 55.650 795.750 57.450 801.600 ;
        RECT 61.650 801.600 63.300 801.900 ;
        RECT 77.250 801.900 84.300 802.800 ;
        RECT 77.250 801.600 78.450 801.900 ;
        RECT 58.650 795.750 60.450 801.000 ;
        RECT 61.650 795.750 63.450 801.600 ;
        RECT 64.650 795.750 66.450 801.600 ;
        RECT 76.650 795.750 78.450 801.600 ;
        RECT 82.650 801.600 84.300 801.900 ;
        RECT 101.700 801.900 108.750 802.800 ;
        RECT 101.700 801.600 103.350 801.900 ;
        RECT 79.650 795.750 81.450 801.000 ;
        RECT 82.650 795.750 84.450 801.600 ;
        RECT 85.650 795.750 87.450 801.600 ;
        RECT 98.550 795.750 100.350 801.600 ;
        RECT 101.550 795.750 103.350 801.600 ;
        RECT 107.550 801.600 108.750 801.900 ;
        RECT 104.550 795.750 106.350 801.000 ;
        RECT 107.550 795.750 109.350 801.600 ;
        RECT 120.300 795.750 122.100 807.600 ;
        RECT 124.500 795.750 126.300 807.600 ;
        RECT 142.950 806.850 145.050 808.950 ;
        RECT 146.250 808.050 148.050 809.850 ;
        RECT 143.100 805.050 144.900 806.850 ;
        RECT 149.700 802.800 150.750 811.050 ;
        RECT 164.100 807.600 165.300 812.850 ;
        RECT 166.950 810.450 169.050 811.050 ;
        RECT 178.950 810.450 181.050 811.050 ;
        RECT 166.950 809.550 181.050 810.450 ;
        RECT 181.950 809.850 184.050 811.950 ;
        RECT 187.950 809.850 190.050 811.950 ;
        RECT 190.950 811.050 193.050 813.150 ;
        RECT 205.950 812.850 208.050 814.950 ;
        RECT 206.100 811.050 207.900 812.850 ;
        RECT 166.950 808.950 169.050 809.550 ;
        RECT 178.950 808.950 181.050 809.550 ;
        RECT 182.100 808.050 183.900 809.850 ;
        RECT 143.700 801.900 150.750 802.800 ;
        RECT 143.700 801.600 145.350 801.900 ;
        RECT 127.800 795.750 129.600 801.600 ;
        RECT 140.550 795.750 142.350 801.600 ;
        RECT 143.550 795.750 145.350 801.600 ;
        RECT 149.550 801.600 150.750 801.900 ;
        RECT 146.550 795.750 148.350 801.000 ;
        RECT 149.550 795.750 151.350 801.600 ;
        RECT 163.650 795.750 165.450 807.600 ;
        RECT 166.650 806.700 174.450 807.600 ;
        RECT 184.950 806.850 187.050 808.950 ;
        RECT 188.250 808.050 190.050 809.850 ;
        RECT 166.650 795.750 168.450 806.700 ;
        RECT 169.650 795.750 171.450 805.800 ;
        RECT 172.650 795.750 174.450 806.700 ;
        RECT 185.100 805.050 186.900 806.850 ;
        RECT 191.700 802.800 192.750 811.050 ;
        RECT 210.000 808.650 211.050 815.850 ;
        RECT 227.400 817.350 231.900 819.000 ;
        RECT 235.500 818.400 237.300 827.250 ;
        RECT 245.550 822.300 247.350 827.250 ;
        RECT 248.550 823.200 250.350 827.250 ;
        RECT 251.550 822.300 253.350 827.250 ;
        RECT 245.550 820.950 253.350 822.300 ;
        RECT 254.550 821.400 256.350 827.250 ;
        RECT 254.550 819.300 255.750 821.400 ;
        RECT 252.000 818.250 255.750 819.300 ;
        RECT 272.100 819.000 273.900 827.250 ;
        RECT 211.950 812.850 214.050 814.950 ;
        RECT 227.400 813.150 228.600 817.350 ;
        RECT 248.100 816.150 249.900 817.950 ;
        RECT 212.100 811.050 213.900 812.850 ;
        RECT 226.950 811.050 229.050 813.150 ;
        RECT 244.950 812.850 247.050 814.950 ;
        RECT 247.950 814.050 250.050 816.150 ;
        RECT 251.850 814.950 253.050 818.250 ;
        RECT 250.950 812.850 253.050 814.950 ;
        RECT 269.400 817.350 273.900 819.000 ;
        RECT 277.500 818.400 279.300 827.250 ;
        RECT 293.100 819.000 294.900 827.250 ;
        RECT 290.400 817.350 294.900 819.000 ;
        RECT 298.500 818.400 300.300 827.250 ;
        RECT 308.850 821.400 310.650 827.250 ;
        RECT 313.350 820.200 315.150 827.250 ;
        RECT 331.650 824.400 333.450 827.250 ;
        RECT 334.650 824.400 336.450 827.250 ;
        RECT 311.550 819.300 315.150 820.200 ;
        RECT 269.400 813.150 270.600 817.350 ;
        RECT 290.400 813.150 291.600 817.350 ;
        RECT 308.100 813.150 309.900 814.950 ;
        RECT 210.000 807.600 212.550 808.650 ;
        RECT 185.700 801.900 192.750 802.800 ;
        RECT 185.700 801.600 187.350 801.900 ;
        RECT 182.550 795.750 184.350 801.600 ;
        RECT 185.550 795.750 187.350 801.600 ;
        RECT 191.550 801.600 192.750 801.900 ;
        RECT 188.550 795.750 190.350 801.000 ;
        RECT 191.550 795.750 193.350 801.600 ;
        RECT 206.550 795.750 208.350 807.600 ;
        RECT 210.750 795.750 212.550 807.600 ;
        RECT 227.250 802.800 228.300 811.050 ;
        RECT 229.950 809.850 232.050 811.950 ;
        RECT 235.950 809.850 238.050 811.950 ;
        RECT 245.100 811.050 246.900 812.850 ;
        RECT 229.950 808.050 231.750 809.850 ;
        RECT 232.950 806.850 235.050 808.950 ;
        RECT 236.100 808.050 237.900 809.850 ;
        RECT 250.950 807.600 252.150 812.850 ;
        RECT 253.950 809.850 256.050 811.950 ;
        RECT 268.950 811.050 271.050 813.150 ;
        RECT 253.950 808.050 255.750 809.850 ;
        RECT 233.100 805.050 234.900 806.850 ;
        RECT 227.250 801.900 234.300 802.800 ;
        RECT 227.250 801.600 228.450 801.900 ;
        RECT 226.650 795.750 228.450 801.600 ;
        RECT 232.650 801.600 234.300 801.900 ;
        RECT 229.650 795.750 231.450 801.000 ;
        RECT 232.650 795.750 234.450 801.600 ;
        RECT 235.650 795.750 237.450 801.600 ;
        RECT 246.300 795.750 248.100 807.600 ;
        RECT 250.500 795.750 252.300 807.600 ;
        RECT 269.250 802.800 270.300 811.050 ;
        RECT 271.950 809.850 274.050 811.950 ;
        RECT 277.950 809.850 280.050 811.950 ;
        RECT 289.950 811.050 292.050 813.150 ;
        RECT 271.950 808.050 273.750 809.850 ;
        RECT 274.950 806.850 277.050 808.950 ;
        RECT 278.100 808.050 279.900 809.850 ;
        RECT 275.100 805.050 276.900 806.850 ;
        RECT 290.250 802.800 291.300 811.050 ;
        RECT 292.950 809.850 295.050 811.950 ;
        RECT 298.950 809.850 301.050 811.950 ;
        RECT 307.950 811.050 310.050 813.150 ;
        RECT 311.550 811.950 312.750 819.300 ;
        RECT 332.400 816.150 333.600 824.400 ;
        RECT 348.150 822.900 349.950 827.250 ;
        RECT 346.650 821.400 349.950 822.900 ;
        RECT 351.150 821.400 352.950 827.250 ;
        RECT 314.100 813.150 315.900 814.950 ;
        RECT 331.950 814.050 334.050 816.150 ;
        RECT 334.950 815.850 337.050 817.950 ;
        RECT 335.100 814.050 336.900 815.850 ;
        RECT 346.650 814.950 347.850 821.400 ;
        RECT 349.950 819.900 351.750 820.500 ;
        RECT 355.650 819.900 357.450 827.250 ;
        RECT 365.550 822.300 367.350 827.250 ;
        RECT 368.550 823.200 370.350 827.250 ;
        RECT 371.550 822.300 373.350 827.250 ;
        RECT 365.550 820.950 373.350 822.300 ;
        RECT 374.550 821.400 376.350 827.250 ;
        RECT 349.950 818.700 357.450 819.900 ;
        RECT 374.550 819.300 375.750 821.400 ;
        RECT 310.950 809.850 313.050 811.950 ;
        RECT 313.950 811.050 316.050 813.150 ;
        RECT 292.950 808.050 294.750 809.850 ;
        RECT 295.950 806.850 298.050 808.950 ;
        RECT 299.100 808.050 300.900 809.850 ;
        RECT 296.100 805.050 297.900 806.850 ;
        RECT 269.250 801.900 276.300 802.800 ;
        RECT 269.250 801.600 270.450 801.900 ;
        RECT 253.800 795.750 255.600 801.600 ;
        RECT 268.650 795.750 270.450 801.600 ;
        RECT 274.650 801.600 276.300 801.900 ;
        RECT 290.250 801.900 297.300 802.800 ;
        RECT 290.250 801.600 291.450 801.900 ;
        RECT 271.650 795.750 273.450 801.000 ;
        RECT 274.650 795.750 276.450 801.600 ;
        RECT 277.650 795.750 279.450 801.600 ;
        RECT 289.650 795.750 291.450 801.600 ;
        RECT 295.650 801.600 297.300 801.900 ;
        RECT 311.550 801.600 312.750 809.850 ;
        RECT 332.400 801.600 333.600 814.050 ;
        RECT 346.650 812.850 349.050 814.950 ;
        RECT 350.100 813.150 351.900 814.950 ;
        RECT 346.650 807.600 347.850 812.850 ;
        RECT 349.950 811.050 352.050 813.150 ;
        RECT 292.650 795.750 294.450 801.000 ;
        RECT 295.650 795.750 297.450 801.600 ;
        RECT 298.650 795.750 300.450 801.600 ;
        RECT 308.550 795.750 310.350 801.600 ;
        RECT 311.550 795.750 313.350 801.600 ;
        RECT 314.550 795.750 316.350 801.600 ;
        RECT 331.650 795.750 333.450 801.600 ;
        RECT 334.650 795.750 336.450 801.600 ;
        RECT 346.050 795.750 347.850 807.600 ;
        RECT 349.050 795.750 350.850 807.600 ;
        RECT 353.100 801.600 354.300 818.700 ;
        RECT 372.000 818.250 375.750 819.300 ;
        RECT 395.100 819.000 396.900 827.250 ;
        RECT 368.100 816.150 369.900 817.950 ;
        RECT 355.950 812.850 358.050 814.950 ;
        RECT 364.950 812.850 367.050 814.950 ;
        RECT 367.950 814.050 370.050 816.150 ;
        RECT 371.850 814.950 373.050 818.250 ;
        RECT 370.950 812.850 373.050 814.950 ;
        RECT 392.400 817.350 396.900 819.000 ;
        RECT 400.500 818.400 402.300 827.250 ;
        RECT 416.100 819.000 417.900 827.250 ;
        RECT 413.400 817.350 417.900 819.000 ;
        RECT 421.500 818.400 423.300 827.250 ;
        RECT 431.550 822.300 433.350 827.250 ;
        RECT 434.550 823.200 436.350 827.250 ;
        RECT 437.550 822.300 439.350 827.250 ;
        RECT 431.550 820.950 439.350 822.300 ;
        RECT 440.550 821.400 442.350 827.250 ;
        RECT 452.550 824.400 454.350 827.250 ;
        RECT 455.550 824.400 457.350 827.250 ;
        RECT 440.550 819.300 441.750 821.400 ;
        RECT 438.000 818.250 441.750 819.300 ;
        RECT 392.400 813.150 393.600 817.350 ;
        RECT 413.400 813.150 414.600 817.350 ;
        RECT 434.100 816.150 435.900 817.950 ;
        RECT 356.100 811.050 357.900 812.850 ;
        RECT 365.100 811.050 366.900 812.850 ;
        RECT 370.950 807.600 372.150 812.850 ;
        RECT 373.950 809.850 376.050 811.950 ;
        RECT 391.950 811.050 394.050 813.150 ;
        RECT 373.950 808.050 375.750 809.850 ;
        RECT 352.650 795.750 354.450 801.600 ;
        RECT 355.650 795.750 357.450 801.600 ;
        RECT 366.300 795.750 368.100 807.600 ;
        RECT 370.500 795.750 372.300 807.600 ;
        RECT 392.250 802.800 393.300 811.050 ;
        RECT 394.950 809.850 397.050 811.950 ;
        RECT 400.950 809.850 403.050 811.950 ;
        RECT 412.950 811.050 415.050 813.150 ;
        RECT 430.950 812.850 433.050 814.950 ;
        RECT 433.950 814.050 436.050 816.150 ;
        RECT 437.850 814.950 439.050 818.250 ;
        RECT 451.950 815.850 454.050 817.950 ;
        RECT 455.400 816.150 456.600 824.400 ;
        RECT 467.850 821.400 469.650 827.250 ;
        RECT 472.350 820.200 474.150 827.250 ;
        RECT 470.550 819.300 474.150 820.200 ;
        RECT 436.950 812.850 439.050 814.950 ;
        RECT 452.100 814.050 453.900 815.850 ;
        RECT 454.950 814.050 457.050 816.150 ;
        RECT 394.950 808.050 396.750 809.850 ;
        RECT 397.950 806.850 400.050 808.950 ;
        RECT 401.100 808.050 402.900 809.850 ;
        RECT 398.100 805.050 399.900 806.850 ;
        RECT 413.250 802.800 414.300 811.050 ;
        RECT 415.950 809.850 418.050 811.950 ;
        RECT 421.950 809.850 424.050 811.950 ;
        RECT 431.100 811.050 432.900 812.850 ;
        RECT 415.950 808.050 417.750 809.850 ;
        RECT 418.950 806.850 421.050 808.950 ;
        RECT 422.100 808.050 423.900 809.850 ;
        RECT 436.950 807.600 438.150 812.850 ;
        RECT 439.950 809.850 442.050 811.950 ;
        RECT 439.950 808.050 441.750 809.850 ;
        RECT 419.100 805.050 420.900 806.850 ;
        RECT 392.250 801.900 399.300 802.800 ;
        RECT 392.250 801.600 393.450 801.900 ;
        RECT 373.800 795.750 375.600 801.600 ;
        RECT 391.650 795.750 393.450 801.600 ;
        RECT 397.650 801.600 399.300 801.900 ;
        RECT 413.250 801.900 420.300 802.800 ;
        RECT 413.250 801.600 414.450 801.900 ;
        RECT 394.650 795.750 396.450 801.000 ;
        RECT 397.650 795.750 399.450 801.600 ;
        RECT 400.650 795.750 402.450 801.600 ;
        RECT 412.650 795.750 414.450 801.600 ;
        RECT 418.650 801.600 420.300 801.900 ;
        RECT 415.650 795.750 417.450 801.000 ;
        RECT 418.650 795.750 420.450 801.600 ;
        RECT 421.650 795.750 423.450 801.600 ;
        RECT 432.300 795.750 434.100 807.600 ;
        RECT 436.500 795.750 438.300 807.600 ;
        RECT 455.400 801.600 456.600 814.050 ;
        RECT 467.100 813.150 468.900 814.950 ;
        RECT 466.950 811.050 469.050 813.150 ;
        RECT 470.550 811.950 471.750 819.300 ;
        RECT 488.700 818.400 490.500 827.250 ;
        RECT 494.100 819.000 495.900 827.250 ;
        RECT 509.850 821.400 511.650 827.250 ;
        RECT 514.350 820.200 516.150 827.250 ;
        RECT 527.550 824.400 529.350 827.250 ;
        RECT 530.550 824.400 532.350 827.250 ;
        RECT 533.550 824.400 535.350 827.250 ;
        RECT 512.550 819.300 516.150 820.200 ;
        RECT 531.450 820.200 532.350 824.400 ;
        RECT 536.550 821.400 538.350 827.250 ;
        RECT 531.450 819.300 534.750 820.200 ;
        RECT 494.100 817.350 498.600 819.000 ;
        RECT 473.100 813.150 474.900 814.950 ;
        RECT 497.400 813.150 498.600 817.350 ;
        RECT 509.100 813.150 510.900 814.950 ;
        RECT 469.950 809.850 472.050 811.950 ;
        RECT 472.950 811.050 475.050 813.150 ;
        RECT 487.950 809.850 490.050 811.950 ;
        RECT 493.950 809.850 496.050 811.950 ;
        RECT 496.950 811.050 499.050 813.150 ;
        RECT 508.950 811.050 511.050 813.150 ;
        RECT 512.550 811.950 513.750 819.300 ;
        RECT 532.950 818.400 534.750 819.300 ;
        RECT 526.950 815.850 529.050 817.950 ;
        RECT 515.100 813.150 516.900 814.950 ;
        RECT 527.100 814.050 528.900 815.850 ;
        RECT 470.550 801.600 471.750 809.850 ;
        RECT 488.100 808.050 489.900 809.850 ;
        RECT 490.950 806.850 493.050 808.950 ;
        RECT 494.250 808.050 496.050 809.850 ;
        RECT 491.100 805.050 492.900 806.850 ;
        RECT 497.700 802.800 498.750 811.050 ;
        RECT 511.950 809.850 514.050 811.950 ;
        RECT 514.950 811.050 517.050 813.150 ;
        RECT 529.950 812.850 532.050 814.950 ;
        RECT 530.100 811.050 531.900 812.850 ;
        RECT 533.700 810.150 534.600 818.400 ;
        RECT 537.000 816.150 538.050 821.400 ;
        RECT 554.100 819.000 555.900 827.250 ;
        RECT 535.950 814.050 538.050 816.150 ;
        RECT 551.400 817.350 555.900 819.000 ;
        RECT 559.500 818.400 561.300 827.250 ;
        RECT 572.700 824.400 574.500 827.250 ;
        RECT 576.000 823.050 577.800 827.250 ;
        RECT 572.100 821.400 577.800 823.050 ;
        RECT 580.200 821.400 582.000 827.250 ;
        RECT 590.850 821.400 592.650 827.250 ;
        RECT 532.950 810.000 534.750 810.150 ;
        RECT 491.700 801.900 498.750 802.800 ;
        RECT 491.700 801.600 493.350 801.900 ;
        RECT 439.800 795.750 441.600 801.600 ;
        RECT 452.550 795.750 454.350 801.600 ;
        RECT 455.550 795.750 457.350 801.600 ;
        RECT 467.550 795.750 469.350 801.600 ;
        RECT 470.550 795.750 472.350 801.600 ;
        RECT 473.550 795.750 475.350 801.600 ;
        RECT 488.550 795.750 490.350 801.600 ;
        RECT 491.550 795.750 493.350 801.600 ;
        RECT 497.550 801.600 498.750 801.900 ;
        RECT 512.550 801.600 513.750 809.850 ;
        RECT 527.550 808.800 534.750 810.000 ;
        RECT 527.550 807.600 528.750 808.800 ;
        RECT 532.950 808.350 534.750 808.800 ;
        RECT 494.550 795.750 496.350 801.000 ;
        RECT 497.550 795.750 499.350 801.600 ;
        RECT 509.550 795.750 511.350 801.600 ;
        RECT 512.550 795.750 514.350 801.600 ;
        RECT 515.550 795.750 517.350 801.600 ;
        RECT 527.550 795.750 529.350 807.600 ;
        RECT 536.100 807.450 537.450 814.050 ;
        RECT 551.400 813.150 552.600 817.350 ;
        RECT 572.100 814.950 573.300 821.400 ;
        RECT 595.350 820.200 597.150 827.250 ;
        RECT 610.650 821.400 612.450 827.250 ;
        RECT 593.550 819.300 597.150 820.200 ;
        RECT 611.250 819.300 612.450 821.400 ;
        RECT 613.650 822.300 615.450 827.250 ;
        RECT 616.650 823.200 618.450 827.250 ;
        RECT 619.650 822.300 621.450 827.250 ;
        RECT 613.650 820.950 621.450 822.300 ;
        RECT 632.850 820.200 634.650 827.250 ;
        RECT 637.350 821.400 639.150 827.250 ;
        RECT 632.850 819.300 636.450 820.200 ;
        RECT 575.100 816.150 576.900 817.950 ;
        RECT 550.950 811.050 553.050 813.150 ;
        RECT 571.950 812.850 574.050 814.950 ;
        RECT 574.950 814.050 577.050 816.150 ;
        RECT 577.950 815.850 580.050 817.950 ;
        RECT 581.100 816.150 582.900 817.950 ;
        RECT 578.100 814.050 579.900 815.850 ;
        RECT 580.950 814.050 583.050 816.150 ;
        RECT 590.100 813.150 591.900 814.950 ;
        RECT 532.050 795.750 533.850 807.450 ;
        RECT 535.050 806.100 537.450 807.450 ;
        RECT 535.050 795.750 536.850 806.100 ;
        RECT 551.250 802.800 552.300 811.050 ;
        RECT 553.950 809.850 556.050 811.950 ;
        RECT 559.950 809.850 562.050 811.950 ;
        RECT 553.950 808.050 555.750 809.850 ;
        RECT 556.950 806.850 559.050 808.950 ;
        RECT 560.100 808.050 561.900 809.850 ;
        RECT 572.100 807.600 573.300 812.850 ;
        RECT 589.950 811.050 592.050 813.150 ;
        RECT 593.550 811.950 594.750 819.300 ;
        RECT 611.250 818.250 615.000 819.300 ;
        RECT 613.950 814.950 615.150 818.250 ;
        RECT 617.100 816.150 618.900 817.950 ;
        RECT 596.100 813.150 597.900 814.950 ;
        RECT 592.950 809.850 595.050 811.950 ;
        RECT 595.950 811.050 598.050 813.150 ;
        RECT 613.950 812.850 616.050 814.950 ;
        RECT 616.950 814.050 619.050 816.150 ;
        RECT 619.950 812.850 622.050 814.950 ;
        RECT 632.100 813.150 633.900 814.950 ;
        RECT 610.950 809.850 613.050 811.950 ;
        RECT 557.100 805.050 558.900 806.850 ;
        RECT 551.250 801.900 558.300 802.800 ;
        RECT 551.250 801.600 552.450 801.900 ;
        RECT 550.650 795.750 552.450 801.600 ;
        RECT 556.650 801.600 558.300 801.900 ;
        RECT 553.650 795.750 555.450 801.000 ;
        RECT 556.650 795.750 558.450 801.600 ;
        RECT 559.650 795.750 561.450 801.600 ;
        RECT 571.650 795.750 573.450 807.600 ;
        RECT 574.650 806.700 582.450 807.600 ;
        RECT 574.650 795.750 576.450 806.700 ;
        RECT 577.650 795.750 579.450 805.800 ;
        RECT 580.650 795.750 582.450 806.700 ;
        RECT 593.550 801.600 594.750 809.850 ;
        RECT 611.250 808.050 613.050 809.850 ;
        RECT 614.850 807.600 616.050 812.850 ;
        RECT 620.100 811.050 621.900 812.850 ;
        RECT 631.950 811.050 634.050 813.150 ;
        RECT 635.250 811.950 636.450 819.300 ;
        RECT 653.100 819.000 654.900 827.250 ;
        RECT 650.400 817.350 654.900 819.000 ;
        RECT 658.500 818.400 660.300 827.250 ;
        RECT 672.000 821.400 673.800 827.250 ;
        RECT 676.200 823.050 678.000 827.250 ;
        RECT 679.500 824.400 681.300 827.250 ;
        RECT 692.550 824.400 694.350 827.250 ;
        RECT 695.550 824.400 697.350 827.250 ;
        RECT 676.200 821.400 681.900 823.050 ;
        RECT 638.100 813.150 639.900 814.950 ;
        RECT 650.400 813.150 651.600 817.350 ;
        RECT 671.100 816.150 672.900 817.950 ;
        RECT 670.950 814.050 673.050 816.150 ;
        RECT 673.950 815.850 676.050 817.950 ;
        RECT 677.100 816.150 678.900 817.950 ;
        RECT 674.100 814.050 675.900 815.850 ;
        RECT 676.950 814.050 679.050 816.150 ;
        RECT 680.700 814.950 681.900 821.400 ;
        RECT 691.950 815.850 694.050 817.950 ;
        RECT 695.400 816.150 696.600 824.400 ;
        RECT 707.550 822.300 709.350 827.250 ;
        RECT 710.550 823.200 712.350 827.250 ;
        RECT 713.550 822.300 715.350 827.250 ;
        RECT 707.550 820.950 715.350 822.300 ;
        RECT 716.550 821.400 718.350 827.250 ;
        RECT 722.550 821.400 724.350 827.250 ;
        RECT 725.850 824.400 727.650 827.250 ;
        RECT 730.350 824.400 732.150 827.250 ;
        RECT 734.550 824.400 736.350 827.250 ;
        RECT 738.450 824.400 740.250 827.250 ;
        RECT 741.750 824.400 743.550 827.250 ;
        RECT 746.250 825.300 748.050 827.250 ;
        RECT 746.250 824.400 750.000 825.300 ;
        RECT 751.050 824.400 752.850 827.250 ;
        RECT 730.650 823.500 731.700 824.400 ;
        RECT 727.950 822.300 731.700 823.500 ;
        RECT 739.200 822.600 740.250 824.400 ;
        RECT 748.950 823.500 750.000 824.400 ;
        RECT 727.950 821.400 730.050 822.300 ;
        RECT 716.550 819.300 717.750 821.400 ;
        RECT 714.000 818.250 717.750 819.300 ;
        RECT 722.550 819.150 723.750 821.400 ;
        RECT 735.150 820.200 736.950 822.000 ;
        RECT 739.200 821.550 744.150 822.600 ;
        RECT 742.350 820.800 744.150 821.550 ;
        RECT 745.650 820.800 747.450 822.600 ;
        RECT 748.950 821.400 751.050 823.500 ;
        RECT 754.050 821.400 755.850 827.250 ;
        RECT 764.550 824.400 766.350 827.250 ;
        RECT 767.550 824.400 769.350 827.250 ;
        RECT 736.050 819.900 736.950 820.200 ;
        RECT 746.100 819.900 747.150 820.800 ;
        RECT 710.100 816.150 711.900 817.950 ;
        RECT 634.950 809.850 637.050 811.950 ;
        RECT 637.950 811.050 640.050 813.150 ;
        RECT 649.950 811.050 652.050 813.150 ;
        RECT 679.950 812.850 682.050 814.950 ;
        RECT 692.100 814.050 693.900 815.850 ;
        RECT 694.950 814.050 697.050 816.150 ;
        RECT 590.550 795.750 592.350 801.600 ;
        RECT 593.550 795.750 595.350 801.600 ;
        RECT 596.550 795.750 598.350 801.600 ;
        RECT 611.400 795.750 613.200 801.600 ;
        RECT 614.700 795.750 616.500 807.600 ;
        RECT 618.900 795.750 620.700 807.600 ;
        RECT 635.250 801.600 636.450 809.850 ;
        RECT 650.250 802.800 651.300 811.050 ;
        RECT 652.950 809.850 655.050 811.950 ;
        RECT 658.950 809.850 661.050 811.950 ;
        RECT 652.950 808.050 654.750 809.850 ;
        RECT 655.950 806.850 658.050 808.950 ;
        RECT 659.100 808.050 660.900 809.850 ;
        RECT 680.700 807.600 681.900 812.850 ;
        RECT 656.100 805.050 657.900 806.850 ;
        RECT 671.550 806.700 679.350 807.600 ;
        RECT 650.250 801.900 657.300 802.800 ;
        RECT 650.250 801.600 651.450 801.900 ;
        RECT 631.650 795.750 633.450 801.600 ;
        RECT 634.650 795.750 636.450 801.600 ;
        RECT 637.650 795.750 639.450 801.600 ;
        RECT 649.650 795.750 651.450 801.600 ;
        RECT 655.650 801.600 657.300 801.900 ;
        RECT 652.650 795.750 654.450 801.000 ;
        RECT 655.650 795.750 657.450 801.600 ;
        RECT 658.650 795.750 660.450 801.600 ;
        RECT 671.550 795.750 673.350 806.700 ;
        RECT 674.550 795.750 676.350 805.800 ;
        RECT 677.550 795.750 679.350 806.700 ;
        RECT 680.550 795.750 682.350 807.600 ;
        RECT 695.400 801.600 696.600 814.050 ;
        RECT 706.950 812.850 709.050 814.950 ;
        RECT 709.950 814.050 712.050 816.150 ;
        RECT 713.850 814.950 715.050 818.250 ;
        RECT 712.950 812.850 715.050 814.950 ;
        RECT 722.550 817.050 727.050 819.150 ;
        RECT 736.050 819.000 747.150 819.900 ;
        RECT 707.100 811.050 708.900 812.850 ;
        RECT 712.950 807.600 714.150 812.850 ;
        RECT 715.950 809.850 718.050 811.950 ;
        RECT 715.950 808.050 717.750 809.850 ;
        RECT 722.550 807.600 723.750 817.050 ;
        RECT 724.950 815.250 728.850 817.050 ;
        RECT 724.950 814.950 727.050 815.250 ;
        RECT 736.050 814.950 736.950 819.000 ;
        RECT 746.100 817.800 747.150 819.000 ;
        RECT 746.100 816.600 753.000 817.800 ;
        RECT 746.100 816.000 747.900 816.600 ;
        RECT 752.100 815.850 753.000 816.600 ;
        RECT 749.100 814.950 750.900 815.700 ;
        RECT 736.050 812.850 739.050 814.950 ;
        RECT 742.950 813.900 750.900 814.950 ;
        RECT 752.100 814.050 753.900 815.850 ;
        RECT 742.950 812.850 745.050 813.900 ;
        RECT 724.950 809.400 726.750 811.200 ;
        RECT 725.850 808.200 730.050 809.400 ;
        RECT 736.050 808.200 736.950 812.850 ;
        RECT 744.750 809.100 746.550 809.400 ;
        RECT 692.550 795.750 694.350 801.600 ;
        RECT 695.550 795.750 697.350 801.600 ;
        RECT 708.300 795.750 710.100 807.600 ;
        RECT 712.500 795.750 714.300 807.600 ;
        RECT 715.800 795.750 717.600 801.600 ;
        RECT 722.550 795.750 724.350 807.600 ;
        RECT 727.950 807.300 730.050 808.200 ;
        RECT 730.950 807.300 736.950 808.200 ;
        RECT 738.150 808.800 746.550 809.100 ;
        RECT 754.950 808.800 755.850 821.400 ;
        RECT 763.950 815.850 766.050 817.950 ;
        RECT 767.400 816.150 768.600 824.400 ;
        RECT 773.550 821.400 775.350 827.250 ;
        RECT 776.850 824.400 778.650 827.250 ;
        RECT 781.350 824.400 783.150 827.250 ;
        RECT 785.550 824.400 787.350 827.250 ;
        RECT 789.450 824.400 791.250 827.250 ;
        RECT 792.750 824.400 794.550 827.250 ;
        RECT 797.250 825.300 799.050 827.250 ;
        RECT 797.250 824.400 801.000 825.300 ;
        RECT 802.050 824.400 803.850 827.250 ;
        RECT 781.650 823.500 782.700 824.400 ;
        RECT 778.950 822.300 782.700 823.500 ;
        RECT 790.200 822.600 791.250 824.400 ;
        RECT 799.950 823.500 801.000 824.400 ;
        RECT 778.950 821.400 781.050 822.300 ;
        RECT 773.550 819.150 774.750 821.400 ;
        RECT 786.150 820.200 787.950 822.000 ;
        RECT 790.200 821.550 795.150 822.600 ;
        RECT 793.350 820.800 795.150 821.550 ;
        RECT 796.650 820.800 798.450 822.600 ;
        RECT 799.950 821.400 802.050 823.500 ;
        RECT 805.050 821.400 806.850 827.250 ;
        RECT 787.050 819.900 787.950 820.200 ;
        RECT 797.100 819.900 798.150 820.800 ;
        RECT 773.550 817.050 778.050 819.150 ;
        RECT 787.050 819.000 798.150 819.900 ;
        RECT 764.100 814.050 765.900 815.850 ;
        RECT 766.950 814.050 769.050 816.150 ;
        RECT 738.150 808.200 755.850 808.800 ;
        RECT 730.950 806.400 731.850 807.300 ;
        RECT 729.150 804.600 731.850 806.400 ;
        RECT 732.750 806.100 734.550 806.400 ;
        RECT 738.150 806.100 739.050 808.200 ;
        RECT 744.750 807.600 755.850 808.200 ;
        RECT 732.750 805.200 739.050 806.100 ;
        RECT 739.950 806.700 741.750 807.300 ;
        RECT 739.950 805.500 747.450 806.700 ;
        RECT 732.750 804.600 734.550 805.200 ;
        RECT 746.250 804.600 747.450 805.500 ;
        RECT 727.950 801.600 731.850 803.700 ;
        RECT 736.950 802.500 743.850 804.300 ;
        RECT 746.250 802.500 751.050 804.600 ;
        RECT 725.550 795.750 727.350 798.600 ;
        RECT 730.050 795.750 731.850 801.600 ;
        RECT 734.250 795.750 736.050 801.600 ;
        RECT 738.150 795.750 739.950 802.500 ;
        RECT 746.250 801.600 747.450 802.500 ;
        RECT 741.150 795.750 742.950 801.600 ;
        RECT 745.950 795.750 747.750 801.600 ;
        RECT 751.050 795.750 752.850 801.600 ;
        RECT 754.050 795.750 755.850 807.600 ;
        RECT 767.400 801.600 768.600 814.050 ;
        RECT 773.550 807.600 774.750 817.050 ;
        RECT 775.950 815.250 779.850 817.050 ;
        RECT 775.950 814.950 778.050 815.250 ;
        RECT 787.050 814.950 787.950 819.000 ;
        RECT 797.100 817.800 798.150 819.000 ;
        RECT 797.100 816.600 804.000 817.800 ;
        RECT 797.100 816.000 798.900 816.600 ;
        RECT 803.100 815.850 804.000 816.600 ;
        RECT 800.100 814.950 801.900 815.700 ;
        RECT 787.050 812.850 790.050 814.950 ;
        RECT 793.950 813.900 801.900 814.950 ;
        RECT 803.100 814.050 804.900 815.850 ;
        RECT 793.950 812.850 796.050 813.900 ;
        RECT 775.950 809.400 777.750 811.200 ;
        RECT 776.850 808.200 781.050 809.400 ;
        RECT 787.050 808.200 787.950 812.850 ;
        RECT 795.750 809.100 797.550 809.400 ;
        RECT 764.550 795.750 766.350 801.600 ;
        RECT 767.550 795.750 769.350 801.600 ;
        RECT 773.550 795.750 775.350 807.600 ;
        RECT 778.950 807.300 781.050 808.200 ;
        RECT 781.950 807.300 787.950 808.200 ;
        RECT 789.150 808.800 797.550 809.100 ;
        RECT 805.950 808.800 806.850 821.400 ;
        RECT 815.550 822.300 817.350 827.250 ;
        RECT 818.550 823.200 820.350 827.250 ;
        RECT 821.550 822.300 823.350 827.250 ;
        RECT 815.550 820.950 823.350 822.300 ;
        RECT 824.550 821.400 826.350 827.250 ;
        RECT 839.850 821.400 841.650 827.250 ;
        RECT 824.550 819.300 825.750 821.400 ;
        RECT 844.350 820.200 846.150 827.250 ;
        RECT 857.850 821.400 859.650 827.250 ;
        RECT 862.350 820.200 864.150 827.250 ;
        RECT 822.000 818.250 825.750 819.300 ;
        RECT 842.550 819.300 846.150 820.200 ;
        RECT 856.950 819.450 859.050 820.050 ;
        RECT 818.100 816.150 819.900 817.950 ;
        RECT 814.950 812.850 817.050 814.950 ;
        RECT 817.950 814.050 820.050 816.150 ;
        RECT 821.850 814.950 823.050 818.250 ;
        RECT 820.950 812.850 823.050 814.950 ;
        RECT 839.100 813.150 840.900 814.950 ;
        RECT 815.100 811.050 816.900 812.850 ;
        RECT 789.150 808.200 806.850 808.800 ;
        RECT 781.950 806.400 782.850 807.300 ;
        RECT 780.150 804.600 782.850 806.400 ;
        RECT 783.750 806.100 785.550 806.400 ;
        RECT 789.150 806.100 790.050 808.200 ;
        RECT 795.750 807.600 806.850 808.200 ;
        RECT 820.950 807.600 822.150 812.850 ;
        RECT 823.950 809.850 826.050 811.950 ;
        RECT 838.950 811.050 841.050 813.150 ;
        RECT 842.550 811.950 843.750 819.300 ;
        RECT 854.550 818.550 859.050 819.450 ;
        RECT 845.100 813.150 846.900 814.950 ;
        RECT 841.950 809.850 844.050 811.950 ;
        RECT 844.950 811.050 847.050 813.150 ;
        RECT 823.950 808.050 825.750 809.850 ;
        RECT 783.750 805.200 790.050 806.100 ;
        RECT 790.950 806.700 792.750 807.300 ;
        RECT 790.950 805.500 798.450 806.700 ;
        RECT 783.750 804.600 785.550 805.200 ;
        RECT 797.250 804.600 798.450 805.500 ;
        RECT 778.950 801.600 782.850 803.700 ;
        RECT 787.950 802.500 794.850 804.300 ;
        RECT 797.250 802.500 802.050 804.600 ;
        RECT 776.550 795.750 778.350 798.600 ;
        RECT 781.050 795.750 782.850 801.600 ;
        RECT 785.250 795.750 787.050 801.600 ;
        RECT 789.150 795.750 790.950 802.500 ;
        RECT 797.250 801.600 798.450 802.500 ;
        RECT 792.150 795.750 793.950 801.600 ;
        RECT 796.950 795.750 798.750 801.600 ;
        RECT 802.050 795.750 803.850 801.600 ;
        RECT 805.050 795.750 806.850 807.600 ;
        RECT 816.300 795.750 818.100 807.600 ;
        RECT 820.500 795.750 822.300 807.600 ;
        RECT 842.550 801.600 843.750 809.850 ;
        RECT 854.550 807.450 855.450 818.550 ;
        RECT 856.950 817.950 859.050 818.550 ;
        RECT 860.550 819.300 864.150 820.200 ;
        RECT 857.100 813.150 858.900 814.950 ;
        RECT 856.950 811.050 859.050 813.150 ;
        RECT 860.550 811.950 861.750 819.300 ;
        RECT 863.100 813.150 864.900 814.950 ;
        RECT 859.950 809.850 862.050 811.950 ;
        RECT 862.950 811.050 865.050 813.150 ;
        RECT 856.950 807.450 859.050 808.050 ;
        RECT 854.550 806.550 859.050 807.450 ;
        RECT 856.950 805.950 859.050 806.550 ;
        RECT 860.550 801.600 861.750 809.850 ;
        RECT 823.800 795.750 825.600 801.600 ;
        RECT 839.550 795.750 841.350 801.600 ;
        RECT 842.550 795.750 844.350 801.600 ;
        RECT 845.550 795.750 847.350 801.600 ;
        RECT 857.550 795.750 859.350 801.600 ;
        RECT 860.550 795.750 862.350 801.600 ;
        RECT 863.550 795.750 865.350 801.600 ;
        RECT 10.650 785.400 12.450 791.250 ;
        RECT 13.650 786.000 15.450 791.250 ;
        RECT 11.250 785.100 12.450 785.400 ;
        RECT 16.650 785.400 18.450 791.250 ;
        RECT 19.650 785.400 21.450 791.250 ;
        RECT 16.650 785.100 18.300 785.400 ;
        RECT 11.250 784.200 18.300 785.100 ;
        RECT 11.250 775.950 12.300 784.200 ;
        RECT 17.100 780.150 18.900 781.950 ;
        RECT 29.550 780.300 31.350 791.250 ;
        RECT 32.550 781.200 34.350 791.250 ;
        RECT 35.550 780.300 37.350 791.250 ;
        RECT 13.950 777.150 15.750 778.950 ;
        RECT 16.950 778.050 19.050 780.150 ;
        RECT 29.550 779.400 37.350 780.300 ;
        RECT 38.550 779.400 40.350 791.250 ;
        RECT 50.550 785.400 52.350 791.250 ;
        RECT 53.550 785.400 55.350 791.250 ;
        RECT 67.650 785.400 69.450 791.250 ;
        RECT 70.650 786.000 72.450 791.250 ;
        RECT 20.100 777.150 21.900 778.950 ;
        RECT 10.950 773.850 13.050 775.950 ;
        RECT 13.950 775.050 16.050 777.150 ;
        RECT 19.950 775.050 22.050 777.150 ;
        RECT 38.700 774.150 39.900 779.400 ;
        RECT 11.400 769.650 12.600 773.850 ;
        RECT 28.950 770.850 31.050 772.950 ;
        RECT 32.100 771.150 33.900 772.950 ;
        RECT 11.400 768.000 15.900 769.650 ;
        RECT 29.100 769.050 30.900 770.850 ;
        RECT 31.950 769.050 34.050 771.150 ;
        RECT 34.950 770.850 37.050 772.950 ;
        RECT 37.950 772.050 40.050 774.150 ;
        RECT 53.400 772.950 54.600 785.400 ;
        RECT 68.250 785.100 69.450 785.400 ;
        RECT 73.650 785.400 75.450 791.250 ;
        RECT 76.650 785.400 78.450 791.250 ;
        RECT 73.650 785.100 75.300 785.400 ;
        RECT 68.250 784.200 75.300 785.100 ;
        RECT 68.250 775.950 69.300 784.200 ;
        RECT 74.100 780.150 75.900 781.950 ;
        RECT 86.550 780.300 88.350 791.250 ;
        RECT 89.550 781.200 91.350 791.250 ;
        RECT 92.550 780.300 94.350 791.250 ;
        RECT 70.950 777.150 72.750 778.950 ;
        RECT 73.950 778.050 76.050 780.150 ;
        RECT 86.550 779.400 94.350 780.300 ;
        RECT 95.550 779.400 97.350 791.250 ;
        RECT 109.650 779.400 111.450 791.250 ;
        RECT 112.650 780.300 114.450 791.250 ;
        RECT 115.650 781.200 117.450 791.250 ;
        RECT 118.650 780.300 120.450 791.250 ;
        RECT 128.550 785.400 130.350 791.250 ;
        RECT 131.550 785.400 133.350 791.250 ;
        RECT 134.550 786.000 136.350 791.250 ;
        RECT 131.700 785.100 133.350 785.400 ;
        RECT 137.550 785.400 139.350 791.250 ;
        RECT 151.650 785.400 153.450 791.250 ;
        RECT 154.650 786.000 156.450 791.250 ;
        RECT 137.550 785.100 138.750 785.400 ;
        RECT 131.700 784.200 138.750 785.100 ;
        RECT 112.650 779.400 120.450 780.300 ;
        RECT 131.100 780.150 132.900 781.950 ;
        RECT 77.100 777.150 78.900 778.950 ;
        RECT 67.950 773.850 70.050 775.950 ;
        RECT 70.950 775.050 73.050 777.150 ;
        RECT 76.950 775.050 79.050 777.150 ;
        RECT 95.700 774.150 96.900 779.400 ;
        RECT 110.100 774.150 111.300 779.400 ;
        RECT 128.100 777.150 129.900 778.950 ;
        RECT 130.950 778.050 133.050 780.150 ;
        RECT 134.250 777.150 136.050 778.950 ;
        RECT 127.950 775.050 130.050 777.150 ;
        RECT 133.950 775.050 136.050 777.150 ;
        RECT 137.700 775.950 138.750 784.200 ;
        RECT 152.250 785.100 153.450 785.400 ;
        RECT 157.650 785.400 159.450 791.250 ;
        RECT 160.650 785.400 162.450 791.250 ;
        RECT 170.550 785.400 172.350 791.250 ;
        RECT 173.550 785.400 175.350 791.250 ;
        RECT 187.650 785.400 189.450 791.250 ;
        RECT 190.650 786.000 192.450 791.250 ;
        RECT 157.650 785.100 159.300 785.400 ;
        RECT 152.250 784.200 159.300 785.100 ;
        RECT 152.250 775.950 153.300 784.200 ;
        RECT 158.100 780.150 159.900 781.950 ;
        RECT 154.950 777.150 156.750 778.950 ;
        RECT 157.950 778.050 160.050 780.150 ;
        RECT 161.100 777.150 162.900 778.950 ;
        RECT 35.100 769.050 36.900 770.850 ;
        RECT 14.100 759.750 15.900 768.000 ;
        RECT 19.500 759.750 21.300 768.600 ;
        RECT 38.700 765.600 39.900 772.050 ;
        RECT 50.100 771.150 51.900 772.950 ;
        RECT 49.950 769.050 52.050 771.150 ;
        RECT 52.950 770.850 55.050 772.950 ;
        RECT 30.000 759.750 31.800 765.600 ;
        RECT 34.200 763.950 39.900 765.600 ;
        RECT 34.200 759.750 36.000 763.950 ;
        RECT 53.400 762.600 54.600 770.850 ;
        RECT 68.400 769.650 69.600 773.850 ;
        RECT 85.950 770.850 88.050 772.950 ;
        RECT 89.100 771.150 90.900 772.950 ;
        RECT 68.400 768.000 72.900 769.650 ;
        RECT 86.100 769.050 87.900 770.850 ;
        RECT 88.950 769.050 91.050 771.150 ;
        RECT 91.950 770.850 94.050 772.950 ;
        RECT 94.950 772.050 97.050 774.150 ;
        RECT 109.950 772.050 112.050 774.150 ;
        RECT 136.950 773.850 139.050 775.950 ;
        RECT 151.950 773.850 154.050 775.950 ;
        RECT 154.950 775.050 157.050 777.150 ;
        RECT 160.950 775.050 163.050 777.150 ;
        RECT 92.100 769.050 93.900 770.850 ;
        RECT 37.500 759.750 39.300 762.600 ;
        RECT 50.550 759.750 52.350 762.600 ;
        RECT 53.550 759.750 55.350 762.600 ;
        RECT 71.100 759.750 72.900 768.000 ;
        RECT 76.500 759.750 78.300 768.600 ;
        RECT 95.700 765.600 96.900 772.050 ;
        RECT 87.000 759.750 88.800 765.600 ;
        RECT 91.200 763.950 96.900 765.600 ;
        RECT 110.100 765.600 111.300 772.050 ;
        RECT 112.950 770.850 115.050 772.950 ;
        RECT 116.100 771.150 117.900 772.950 ;
        RECT 113.100 769.050 114.900 770.850 ;
        RECT 115.950 769.050 118.050 771.150 ;
        RECT 118.950 770.850 121.050 772.950 ;
        RECT 119.100 769.050 120.900 770.850 ;
        RECT 137.400 769.650 138.600 773.850 ;
        RECT 110.100 763.950 115.800 765.600 ;
        RECT 91.200 759.750 93.000 763.950 ;
        RECT 94.500 759.750 96.300 762.600 ;
        RECT 110.700 759.750 112.500 762.600 ;
        RECT 114.000 759.750 115.800 763.950 ;
        RECT 118.200 759.750 120.000 765.600 ;
        RECT 128.700 759.750 130.500 768.600 ;
        RECT 134.100 768.000 138.600 769.650 ;
        RECT 152.400 769.650 153.600 773.850 ;
        RECT 173.400 772.950 174.600 785.400 ;
        RECT 188.250 785.100 189.450 785.400 ;
        RECT 193.650 785.400 195.450 791.250 ;
        RECT 196.650 785.400 198.450 791.250 ;
        RECT 212.400 785.400 214.200 791.250 ;
        RECT 193.650 785.100 195.300 785.400 ;
        RECT 188.250 784.200 195.300 785.100 ;
        RECT 188.250 775.950 189.300 784.200 ;
        RECT 194.100 780.150 195.900 781.950 ;
        RECT 190.950 777.150 192.750 778.950 ;
        RECT 193.950 778.050 196.050 780.150 ;
        RECT 215.700 779.400 217.500 791.250 ;
        RECT 219.900 779.400 221.700 791.250 ;
        RECT 232.650 785.400 234.450 791.250 ;
        RECT 235.650 785.400 237.450 791.250 ;
        RECT 248.400 785.400 250.200 791.250 ;
        RECT 197.100 777.150 198.900 778.950 ;
        RECT 212.250 777.150 214.050 778.950 ;
        RECT 187.950 773.850 190.050 775.950 ;
        RECT 190.950 775.050 193.050 777.150 ;
        RECT 196.950 775.050 199.050 777.150 ;
        RECT 211.950 775.050 214.050 777.150 ;
        RECT 215.850 774.150 217.050 779.400 ;
        RECT 221.100 774.150 222.900 775.950 ;
        RECT 170.100 771.150 171.900 772.950 ;
        RECT 152.400 768.000 156.900 769.650 ;
        RECT 169.950 769.050 172.050 771.150 ;
        RECT 172.950 770.850 175.050 772.950 ;
        RECT 134.100 759.750 135.900 768.000 ;
        RECT 155.100 759.750 156.900 768.000 ;
        RECT 160.500 759.750 162.300 768.600 ;
        RECT 173.400 762.600 174.600 770.850 ;
        RECT 188.400 769.650 189.600 773.850 ;
        RECT 214.950 772.050 217.050 774.150 ;
        RECT 188.400 768.000 192.900 769.650 ;
        RECT 214.950 768.750 216.150 772.050 ;
        RECT 217.950 770.850 220.050 772.950 ;
        RECT 220.950 772.050 223.050 774.150 ;
        RECT 233.400 772.950 234.600 785.400 ;
        RECT 251.700 779.400 253.500 791.250 ;
        RECT 255.900 779.400 257.700 791.250 ;
        RECT 271.050 790.500 278.850 791.250 ;
        RECT 271.050 781.200 272.850 790.500 ;
        RECT 274.050 781.800 275.850 789.600 ;
        RECT 274.650 779.400 275.850 781.800 ;
        RECT 277.050 781.800 278.850 790.500 ;
        RECT 280.650 790.500 288.450 791.250 ;
        RECT 280.650 782.700 282.450 790.500 ;
        RECT 283.650 781.800 285.450 789.600 ;
        RECT 277.050 780.900 285.450 781.800 ;
        RECT 286.650 781.500 288.450 790.500 ;
        RECT 289.650 782.400 291.450 791.250 ;
        RECT 292.650 781.500 294.450 791.250 ;
        RECT 286.650 780.600 294.450 781.500 ;
        RECT 304.650 790.500 312.450 791.250 ;
        RECT 304.650 779.400 306.450 790.500 ;
        RECT 307.650 779.400 309.450 789.600 ;
        RECT 310.650 780.600 312.450 790.500 ;
        RECT 313.650 781.500 315.450 791.250 ;
        RECT 316.650 780.600 318.450 791.250 ;
        RECT 326.550 785.400 328.350 791.250 ;
        RECT 329.550 785.400 331.350 791.250 ;
        RECT 332.550 785.400 334.350 791.250 ;
        RECT 346.650 785.400 348.450 791.250 ;
        RECT 349.650 786.000 351.450 791.250 ;
        RECT 310.650 779.700 318.450 780.600 ;
        RECT 248.250 777.150 250.050 778.950 ;
        RECT 247.950 775.050 250.050 777.150 ;
        RECT 251.850 774.150 253.050 779.400 ;
        RECT 274.650 778.200 278.100 779.400 ;
        RECT 257.100 774.150 258.900 775.950 ;
        RECT 232.950 770.850 235.050 772.950 ;
        RECT 236.100 771.150 237.900 772.950 ;
        RECT 250.950 772.050 253.050 774.150 ;
        RECT 218.100 769.050 219.900 770.850 ;
        RECT 170.550 759.750 172.350 762.600 ;
        RECT 173.550 759.750 175.350 762.600 ;
        RECT 191.100 759.750 192.900 768.000 ;
        RECT 196.500 759.750 198.300 768.600 ;
        RECT 212.250 767.700 216.000 768.750 ;
        RECT 212.250 765.600 213.450 767.700 ;
        RECT 211.650 759.750 213.450 765.600 ;
        RECT 214.650 764.700 222.450 766.050 ;
        RECT 214.650 759.750 216.450 764.700 ;
        RECT 217.650 759.750 219.450 763.800 ;
        RECT 220.650 759.750 222.450 764.700 ;
        RECT 233.400 762.600 234.600 770.850 ;
        RECT 235.950 769.050 238.050 771.150 ;
        RECT 250.950 768.750 252.150 772.050 ;
        RECT 253.950 770.850 256.050 772.950 ;
        RECT 256.950 772.050 259.050 774.150 ;
        RECT 276.900 772.950 278.100 778.200 ;
        RECT 307.800 778.500 309.600 779.400 ;
        RECT 307.800 777.600 311.850 778.500 ;
        RECT 281.100 774.150 282.900 775.950 ;
        RECT 290.100 774.150 291.900 775.950 ;
        RECT 305.100 774.150 306.900 775.950 ;
        RECT 310.950 774.150 311.850 777.600 ;
        RECT 329.550 777.150 330.750 785.400 ;
        RECT 347.250 785.100 348.450 785.400 ;
        RECT 352.650 785.400 354.450 791.250 ;
        RECT 355.650 785.400 357.450 791.250 ;
        RECT 352.650 785.100 354.300 785.400 ;
        RECT 347.250 784.200 354.300 785.100 ;
        RECT 316.950 774.150 318.750 775.950 ;
        RECT 274.950 770.850 278.100 772.950 ;
        RECT 280.950 772.050 283.050 774.150 ;
        RECT 283.950 770.850 286.050 772.950 ;
        RECT 289.950 772.050 292.050 774.150 ;
        RECT 304.950 772.050 307.050 774.150 ;
        RECT 307.950 770.850 310.050 772.950 ;
        RECT 310.950 772.050 313.050 774.150 ;
        RECT 254.100 769.050 255.900 770.850 ;
        RECT 248.250 767.700 252.000 768.750 ;
        RECT 235.950 765.450 238.050 766.050 ;
        RECT 241.950 765.450 244.050 766.050 ;
        RECT 248.250 765.600 249.450 767.700 ;
        RECT 235.950 764.550 244.050 765.450 ;
        RECT 235.950 763.950 238.050 764.550 ;
        RECT 241.950 763.950 244.050 764.550 ;
        RECT 232.650 759.750 234.450 762.600 ;
        RECT 235.650 759.750 237.450 762.600 ;
        RECT 247.650 759.750 249.450 765.600 ;
        RECT 250.650 764.700 258.450 766.050 ;
        RECT 250.650 759.750 252.450 764.700 ;
        RECT 253.650 759.750 255.450 763.800 ;
        RECT 256.650 759.750 258.450 764.700 ;
        RECT 276.900 764.400 278.100 770.850 ;
        RECT 284.100 769.050 285.900 770.850 ;
        RECT 308.250 769.050 310.050 770.850 ;
        RECT 312.000 765.600 313.050 772.050 ;
        RECT 313.950 770.850 316.050 772.950 ;
        RECT 316.950 772.050 319.050 774.150 ;
        RECT 325.950 773.850 328.050 775.950 ;
        RECT 328.950 775.050 331.050 777.150 ;
        RECT 347.250 775.950 348.300 784.200 ;
        RECT 353.100 780.150 354.900 781.950 ;
        RECT 349.950 777.150 351.750 778.950 ;
        RECT 352.950 778.050 355.050 780.150 ;
        RECT 367.650 779.400 369.450 791.250 ;
        RECT 370.650 780.300 372.450 791.250 ;
        RECT 373.650 781.200 375.450 791.250 ;
        RECT 376.650 780.300 378.450 791.250 ;
        RECT 388.650 785.400 390.450 791.250 ;
        RECT 391.650 785.400 393.450 791.250 ;
        RECT 404.400 785.400 406.200 791.250 ;
        RECT 370.650 779.400 378.450 780.300 ;
        RECT 356.100 777.150 357.900 778.950 ;
        RECT 326.100 772.050 327.900 773.850 ;
        RECT 313.950 769.050 315.750 770.850 ;
        RECT 329.550 767.700 330.750 775.050 ;
        RECT 331.950 773.850 334.050 775.950 ;
        RECT 346.950 773.850 349.050 775.950 ;
        RECT 349.950 775.050 352.050 777.150 ;
        RECT 355.950 775.050 358.050 777.150 ;
        RECT 368.100 774.150 369.300 779.400 ;
        RECT 332.100 772.050 333.900 773.850 ;
        RECT 347.400 769.650 348.600 773.850 ;
        RECT 367.950 772.050 370.050 774.150 ;
        RECT 389.400 772.950 390.600 785.400 ;
        RECT 407.700 779.400 409.500 791.250 ;
        RECT 411.900 779.400 413.700 791.250 ;
        RECT 428.400 785.400 430.200 791.250 ;
        RECT 431.700 779.400 433.500 791.250 ;
        RECT 435.900 779.400 437.700 791.250 ;
        RECT 448.050 779.400 449.850 791.250 ;
        RECT 451.050 779.400 452.850 791.250 ;
        RECT 454.650 785.400 456.450 791.250 ;
        RECT 457.650 785.400 459.450 791.250 ;
        RECT 404.250 777.150 406.050 778.950 ;
        RECT 403.950 775.050 406.050 777.150 ;
        RECT 407.850 774.150 409.050 779.400 ;
        RECT 428.250 777.150 430.050 778.950 ;
        RECT 413.100 774.150 414.900 775.950 ;
        RECT 427.950 775.050 430.050 777.150 ;
        RECT 431.850 774.150 433.050 779.400 ;
        RECT 437.100 774.150 438.900 775.950 ;
        RECT 448.650 774.150 449.850 779.400 ;
        RECT 347.400 768.000 351.900 769.650 ;
        RECT 329.550 766.800 333.150 767.700 ;
        RECT 276.900 763.500 287.700 764.400 ;
        RECT 280.650 762.600 281.700 763.500 ;
        RECT 286.650 762.600 287.700 763.500 ;
        RECT 280.650 759.750 282.450 762.600 ;
        RECT 283.650 759.750 285.450 762.600 ;
        RECT 286.650 759.750 288.450 762.600 ;
        RECT 289.650 759.750 291.750 762.600 ;
        RECT 307.800 759.750 309.600 765.600 ;
        RECT 312.000 759.750 313.800 765.600 ;
        RECT 316.200 759.750 318.000 765.600 ;
        RECT 326.850 759.750 328.650 765.600 ;
        RECT 331.350 759.750 333.150 766.800 ;
        RECT 350.100 759.750 351.900 768.000 ;
        RECT 355.500 759.750 357.300 768.600 ;
        RECT 368.100 765.600 369.300 772.050 ;
        RECT 370.950 770.850 373.050 772.950 ;
        RECT 374.100 771.150 375.900 772.950 ;
        RECT 371.100 769.050 372.900 770.850 ;
        RECT 373.950 769.050 376.050 771.150 ;
        RECT 376.950 770.850 379.050 772.950 ;
        RECT 388.950 770.850 391.050 772.950 ;
        RECT 392.100 771.150 393.900 772.950 ;
        RECT 406.950 772.050 409.050 774.150 ;
        RECT 377.100 769.050 378.900 770.850 ;
        RECT 368.100 763.950 373.800 765.600 ;
        RECT 368.700 759.750 370.500 762.600 ;
        RECT 372.000 759.750 373.800 763.950 ;
        RECT 376.200 759.750 378.000 765.600 ;
        RECT 389.400 762.600 390.600 770.850 ;
        RECT 391.950 769.050 394.050 771.150 ;
        RECT 406.950 768.750 408.150 772.050 ;
        RECT 409.950 770.850 412.050 772.950 ;
        RECT 412.950 772.050 415.050 774.150 ;
        RECT 430.950 772.050 433.050 774.150 ;
        RECT 410.100 769.050 411.900 770.850 ;
        RECT 430.950 768.750 432.150 772.050 ;
        RECT 433.950 770.850 436.050 772.950 ;
        RECT 436.950 772.050 439.050 774.150 ;
        RECT 448.650 772.050 451.050 774.150 ;
        RECT 451.950 773.850 454.050 775.950 ;
        RECT 452.100 772.050 453.900 773.850 ;
        RECT 434.100 769.050 435.900 770.850 ;
        RECT 404.250 767.700 408.000 768.750 ;
        RECT 428.250 767.700 432.000 768.750 ;
        RECT 404.250 765.600 405.450 767.700 ;
        RECT 388.650 759.750 390.450 762.600 ;
        RECT 391.650 759.750 393.450 762.600 ;
        RECT 403.650 759.750 405.450 765.600 ;
        RECT 406.650 764.700 414.450 766.050 ;
        RECT 428.250 765.600 429.450 767.700 ;
        RECT 406.650 759.750 408.450 764.700 ;
        RECT 409.650 759.750 411.450 763.800 ;
        RECT 412.650 759.750 414.450 764.700 ;
        RECT 427.650 759.750 429.450 765.600 ;
        RECT 430.650 764.700 438.450 766.050 ;
        RECT 430.650 759.750 432.450 764.700 ;
        RECT 433.650 759.750 435.450 763.800 ;
        RECT 436.650 759.750 438.450 764.700 ;
        RECT 448.650 765.600 449.850 772.050 ;
        RECT 455.100 768.300 456.300 785.400 ;
        RECT 467.550 779.400 469.350 791.250 ;
        RECT 471.750 779.400 473.550 791.250 ;
        RECT 490.650 785.400 492.450 791.250 ;
        RECT 493.650 785.400 495.450 791.250 ;
        RECT 471.000 778.350 473.550 779.400 ;
        RECT 458.100 774.150 459.900 775.950 ;
        RECT 467.100 774.150 468.900 775.950 ;
        RECT 457.950 772.050 460.050 774.150 ;
        RECT 466.950 772.050 469.050 774.150 ;
        RECT 471.000 771.150 472.050 778.350 ;
        RECT 473.100 774.150 474.900 775.950 ;
        RECT 472.950 772.050 475.050 774.150 ;
        RECT 491.400 772.950 492.600 785.400 ;
        RECT 507.450 779.400 509.250 791.250 ;
        RECT 511.650 779.400 513.450 791.250 ;
        RECT 527.400 785.400 529.200 791.250 ;
        RECT 530.700 779.400 532.500 791.250 ;
        RECT 534.900 779.400 536.700 791.250 ;
        RECT 545.550 785.400 547.350 791.250 ;
        RECT 548.550 785.400 550.350 791.250 ;
        RECT 551.550 785.400 553.350 791.250 ;
        RECT 565.650 785.400 567.450 791.250 ;
        RECT 568.650 785.400 570.450 791.250 ;
        RECT 571.650 785.400 573.450 791.250 ;
        RECT 586.650 785.400 588.450 791.250 ;
        RECT 589.650 785.400 591.450 791.250 ;
        RECT 592.650 785.400 594.450 791.250 ;
        RECT 602.550 785.400 604.350 791.250 ;
        RECT 605.550 785.400 607.350 791.250 ;
        RECT 608.550 786.000 610.350 791.250 ;
        RECT 507.450 778.350 510.000 779.400 ;
        RECT 506.100 774.150 507.900 775.950 ;
        RECT 469.950 769.050 472.050 771.150 ;
        RECT 490.950 770.850 493.050 772.950 ;
        RECT 494.100 771.150 495.900 772.950 ;
        RECT 505.950 772.050 508.050 774.150 ;
        RECT 508.950 771.150 510.000 778.350 ;
        RECT 527.250 777.150 529.050 778.950 ;
        RECT 512.100 774.150 513.900 775.950 ;
        RECT 526.950 775.050 529.050 777.150 ;
        RECT 530.850 774.150 532.050 779.400 ;
        RECT 548.550 777.150 549.750 785.400 ;
        RECT 569.250 777.150 570.450 785.400 ;
        RECT 590.250 777.150 591.450 785.400 ;
        RECT 605.700 785.100 607.350 785.400 ;
        RECT 611.550 785.400 613.350 791.250 ;
        RECT 626.400 785.400 628.200 791.250 ;
        RECT 611.550 785.100 612.750 785.400 ;
        RECT 605.700 784.200 612.750 785.100 ;
        RECT 592.950 780.450 595.050 781.050 ;
        RECT 592.950 779.550 597.450 780.450 ;
        RECT 605.100 780.150 606.900 781.950 ;
        RECT 592.950 778.950 595.050 779.550 ;
        RECT 536.100 774.150 537.900 775.950 ;
        RECT 511.950 772.050 514.050 774.150 ;
        RECT 529.950 772.050 532.050 774.150 ;
        RECT 451.950 767.100 459.450 768.300 ;
        RECT 451.950 766.500 453.750 767.100 ;
        RECT 448.650 764.100 451.950 765.600 ;
        RECT 450.150 759.750 451.950 764.100 ;
        RECT 453.150 759.750 454.950 765.600 ;
        RECT 457.650 759.750 459.450 767.100 ;
        RECT 471.000 762.600 472.050 769.050 ;
        RECT 491.400 762.600 492.600 770.850 ;
        RECT 493.950 769.050 496.050 771.150 ;
        RECT 508.950 769.050 511.050 771.150 ;
        RECT 508.950 762.600 510.000 769.050 ;
        RECT 529.950 768.750 531.150 772.050 ;
        RECT 532.950 770.850 535.050 772.950 ;
        RECT 535.950 772.050 538.050 774.150 ;
        RECT 544.950 773.850 547.050 775.950 ;
        RECT 547.950 775.050 550.050 777.150 ;
        RECT 545.100 772.050 546.900 773.850 ;
        RECT 533.100 769.050 534.900 770.850 ;
        RECT 527.250 767.700 531.000 768.750 ;
        RECT 548.550 767.700 549.750 775.050 ;
        RECT 550.950 773.850 553.050 775.950 ;
        RECT 565.950 773.850 568.050 775.950 ;
        RECT 568.950 775.050 571.050 777.150 ;
        RECT 551.100 772.050 552.900 773.850 ;
        RECT 566.100 772.050 567.900 773.850 ;
        RECT 569.250 767.700 570.450 775.050 ;
        RECT 571.950 773.850 574.050 775.950 ;
        RECT 586.950 773.850 589.050 775.950 ;
        RECT 589.950 775.050 592.050 777.150 ;
        RECT 572.100 772.050 573.900 773.850 ;
        RECT 587.100 772.050 588.900 773.850 ;
        RECT 590.250 767.700 591.450 775.050 ;
        RECT 592.950 773.850 595.050 775.950 ;
        RECT 593.100 772.050 594.900 773.850 ;
        RECT 596.550 771.450 597.450 779.550 ;
        RECT 602.100 777.150 603.900 778.950 ;
        RECT 604.950 778.050 607.050 780.150 ;
        RECT 608.250 777.150 610.050 778.950 ;
        RECT 601.950 775.050 604.050 777.150 ;
        RECT 607.950 775.050 610.050 777.150 ;
        RECT 611.700 775.950 612.750 784.200 ;
        RECT 629.700 779.400 631.500 791.250 ;
        RECT 633.900 779.400 635.700 791.250 ;
        RECT 648.300 779.400 650.100 791.250 ;
        RECT 652.500 779.400 654.300 791.250 ;
        RECT 655.800 785.400 657.600 791.250 ;
        RECT 668.550 785.400 670.350 791.250 ;
        RECT 671.550 785.400 673.350 791.250 ;
        RECT 685.650 785.400 687.450 791.250 ;
        RECT 688.650 786.000 690.450 791.250 ;
        RECT 626.250 777.150 628.050 778.950 ;
        RECT 610.950 773.850 613.050 775.950 ;
        RECT 625.950 775.050 628.050 777.150 ;
        RECT 629.850 774.150 631.050 779.400 ;
        RECT 635.100 774.150 636.900 775.950 ;
        RECT 647.100 774.150 648.900 775.950 ;
        RECT 652.950 774.150 654.150 779.400 ;
        RECT 655.950 777.150 657.750 778.950 ;
        RECT 655.950 775.050 658.050 777.150 ;
        RECT 601.950 771.450 604.050 772.050 ;
        RECT 596.550 770.550 604.050 771.450 ;
        RECT 601.950 769.950 604.050 770.550 ;
        RECT 611.400 769.650 612.600 773.850 ;
        RECT 527.250 765.600 528.450 767.700 ;
        RECT 548.550 766.800 552.150 767.700 ;
        RECT 467.550 759.750 469.350 762.600 ;
        RECT 470.550 759.750 472.350 762.600 ;
        RECT 473.550 759.750 475.350 762.600 ;
        RECT 490.650 759.750 492.450 762.600 ;
        RECT 493.650 759.750 495.450 762.600 ;
        RECT 505.650 759.750 507.450 762.600 ;
        RECT 508.650 759.750 510.450 762.600 ;
        RECT 511.650 759.750 513.450 762.600 ;
        RECT 526.650 759.750 528.450 765.600 ;
        RECT 529.650 764.700 537.450 766.050 ;
        RECT 529.650 759.750 531.450 764.700 ;
        RECT 532.650 759.750 534.450 763.800 ;
        RECT 535.650 759.750 537.450 764.700 ;
        RECT 545.850 759.750 547.650 765.600 ;
        RECT 550.350 759.750 552.150 766.800 ;
        RECT 566.850 766.800 570.450 767.700 ;
        RECT 587.850 766.800 591.450 767.700 ;
        RECT 566.850 759.750 568.650 766.800 ;
        RECT 571.350 759.750 573.150 765.600 ;
        RECT 587.850 759.750 589.650 766.800 ;
        RECT 592.350 759.750 594.150 765.600 ;
        RECT 602.700 759.750 604.500 768.600 ;
        RECT 608.100 768.000 612.600 769.650 ;
        RECT 628.950 772.050 631.050 774.150 ;
        RECT 628.950 768.750 630.150 772.050 ;
        RECT 631.950 770.850 634.050 772.950 ;
        RECT 634.950 772.050 637.050 774.150 ;
        RECT 646.950 772.050 649.050 774.150 ;
        RECT 649.950 770.850 652.050 772.950 ;
        RECT 652.950 772.050 655.050 774.150 ;
        RECT 671.400 772.950 672.600 785.400 ;
        RECT 686.250 785.100 687.450 785.400 ;
        RECT 691.650 785.400 693.450 791.250 ;
        RECT 694.650 785.400 696.450 791.250 ;
        RECT 691.650 785.100 693.300 785.400 ;
        RECT 686.250 784.200 693.300 785.100 ;
        RECT 686.250 775.950 687.300 784.200 ;
        RECT 692.100 780.150 693.900 781.950 ;
        RECT 704.550 780.300 706.350 791.250 ;
        RECT 707.550 781.200 709.350 791.250 ;
        RECT 710.550 780.300 712.350 791.250 ;
        RECT 688.950 777.150 690.750 778.950 ;
        RECT 691.950 778.050 694.050 780.150 ;
        RECT 704.550 779.400 712.350 780.300 ;
        RECT 713.550 779.400 715.350 791.250 ;
        RECT 725.550 779.400 727.350 791.250 ;
        RECT 729.750 779.400 731.550 791.250 ;
        RECT 695.100 777.150 696.900 778.950 ;
        RECT 685.950 773.850 688.050 775.950 ;
        RECT 688.950 775.050 691.050 777.150 ;
        RECT 694.950 775.050 697.050 777.150 ;
        RECT 713.700 774.150 714.900 779.400 ;
        RECT 729.000 778.350 731.550 779.400 ;
        RECT 737.550 779.400 739.350 791.250 ;
        RECT 740.550 788.400 742.350 791.250 ;
        RECT 745.050 785.400 746.850 791.250 ;
        RECT 749.250 785.400 751.050 791.250 ;
        RECT 742.950 783.300 746.850 785.400 ;
        RECT 753.150 784.500 754.950 791.250 ;
        RECT 756.150 785.400 757.950 791.250 ;
        RECT 760.950 785.400 762.750 791.250 ;
        RECT 766.050 785.400 767.850 791.250 ;
        RECT 761.250 784.500 762.450 785.400 ;
        RECT 751.950 782.700 758.850 784.500 ;
        RECT 761.250 782.400 766.050 784.500 ;
        RECT 744.150 780.600 746.850 782.400 ;
        RECT 747.750 781.800 749.550 782.400 ;
        RECT 747.750 780.900 754.050 781.800 ;
        RECT 761.250 781.500 762.450 782.400 ;
        RECT 747.750 780.600 749.550 780.900 ;
        RECT 745.950 779.700 746.850 780.600 ;
        RECT 725.100 774.150 726.900 775.950 ;
        RECT 632.100 769.050 633.900 770.850 ;
        RECT 650.100 769.050 651.900 770.850 ;
        RECT 653.850 768.750 655.050 772.050 ;
        RECT 668.100 771.150 669.900 772.950 ;
        RECT 667.950 769.050 670.050 771.150 ;
        RECT 670.950 770.850 673.050 772.950 ;
        RECT 608.100 759.750 609.900 768.000 ;
        RECT 626.250 767.700 630.000 768.750 ;
        RECT 654.000 767.700 657.750 768.750 ;
        RECT 626.250 765.600 627.450 767.700 ;
        RECT 625.650 759.750 627.450 765.600 ;
        RECT 628.650 764.700 636.450 766.050 ;
        RECT 628.650 759.750 630.450 764.700 ;
        RECT 631.650 759.750 633.450 763.800 ;
        RECT 634.650 759.750 636.450 764.700 ;
        RECT 647.550 764.700 655.350 766.050 ;
        RECT 647.550 759.750 649.350 764.700 ;
        RECT 650.550 759.750 652.350 763.800 ;
        RECT 653.550 759.750 655.350 764.700 ;
        RECT 656.550 765.600 657.750 767.700 ;
        RECT 656.550 759.750 658.350 765.600 ;
        RECT 671.400 762.600 672.600 770.850 ;
        RECT 686.400 769.650 687.600 773.850 ;
        RECT 703.950 770.850 706.050 772.950 ;
        RECT 707.100 771.150 708.900 772.950 ;
        RECT 686.400 768.000 690.900 769.650 ;
        RECT 704.100 769.050 705.900 770.850 ;
        RECT 706.950 769.050 709.050 771.150 ;
        RECT 709.950 770.850 712.050 772.950 ;
        RECT 712.950 772.050 715.050 774.150 ;
        RECT 724.950 772.050 727.050 774.150 ;
        RECT 710.100 769.050 711.900 770.850 ;
        RECT 668.550 759.750 670.350 762.600 ;
        RECT 671.550 759.750 673.350 762.600 ;
        RECT 689.100 759.750 690.900 768.000 ;
        RECT 694.500 759.750 696.300 768.600 ;
        RECT 713.700 765.600 714.900 772.050 ;
        RECT 729.000 771.150 730.050 778.350 ;
        RECT 731.100 774.150 732.900 775.950 ;
        RECT 730.950 772.050 733.050 774.150 ;
        RECT 727.950 769.050 730.050 771.150 ;
        RECT 705.000 759.750 706.800 765.600 ;
        RECT 709.200 763.950 714.900 765.600 ;
        RECT 709.200 759.750 711.000 763.950 ;
        RECT 729.000 762.600 730.050 769.050 ;
        RECT 737.550 769.950 738.750 779.400 ;
        RECT 742.950 778.800 745.050 779.700 ;
        RECT 745.950 778.800 751.950 779.700 ;
        RECT 740.850 777.600 745.050 778.800 ;
        RECT 739.950 775.800 741.750 777.600 ;
        RECT 751.050 774.150 751.950 778.800 ;
        RECT 753.150 778.800 754.050 780.900 ;
        RECT 754.950 780.300 762.450 781.500 ;
        RECT 754.950 779.700 756.750 780.300 ;
        RECT 769.050 779.400 770.850 791.250 ;
        RECT 780.300 779.400 782.100 791.250 ;
        RECT 784.500 779.400 786.300 791.250 ;
        RECT 787.800 785.400 789.600 791.250 ;
        RECT 800.550 785.400 802.350 791.250 ;
        RECT 803.550 785.400 805.350 791.250 ;
        RECT 759.750 778.800 770.850 779.400 ;
        RECT 753.150 778.200 770.850 778.800 ;
        RECT 753.150 777.900 761.550 778.200 ;
        RECT 759.750 777.600 761.550 777.900 ;
        RECT 751.050 772.050 754.050 774.150 ;
        RECT 757.950 773.100 760.050 774.150 ;
        RECT 757.950 772.050 765.900 773.100 ;
        RECT 739.950 771.750 742.050 772.050 ;
        RECT 739.950 769.950 743.850 771.750 ;
        RECT 737.550 767.850 742.050 769.950 ;
        RECT 751.050 768.000 751.950 772.050 ;
        RECT 764.100 771.300 765.900 772.050 ;
        RECT 767.100 771.150 768.900 772.950 ;
        RECT 761.100 770.400 762.900 771.000 ;
        RECT 767.100 770.400 768.000 771.150 ;
        RECT 761.100 769.200 768.000 770.400 ;
        RECT 761.100 768.000 762.150 769.200 ;
        RECT 737.550 765.600 738.750 767.850 ;
        RECT 751.050 767.100 762.150 768.000 ;
        RECT 751.050 766.800 751.950 767.100 ;
        RECT 712.500 759.750 714.300 762.600 ;
        RECT 725.550 759.750 727.350 762.600 ;
        RECT 728.550 759.750 730.350 762.600 ;
        RECT 731.550 759.750 733.350 762.600 ;
        RECT 737.550 759.750 739.350 765.600 ;
        RECT 742.950 764.700 745.050 765.600 ;
        RECT 750.150 765.000 751.950 766.800 ;
        RECT 761.100 766.200 762.150 767.100 ;
        RECT 757.350 765.450 759.150 766.200 ;
        RECT 742.950 763.500 746.700 764.700 ;
        RECT 745.650 762.600 746.700 763.500 ;
        RECT 754.200 764.400 759.150 765.450 ;
        RECT 760.650 764.400 762.450 766.200 ;
        RECT 769.950 765.600 770.850 778.200 ;
        RECT 779.100 774.150 780.900 775.950 ;
        RECT 784.950 774.150 786.150 779.400 ;
        RECT 787.950 777.150 789.750 778.950 ;
        RECT 787.950 775.050 790.050 777.150 ;
        RECT 778.950 772.050 781.050 774.150 ;
        RECT 781.950 770.850 784.050 772.950 ;
        RECT 784.950 772.050 787.050 774.150 ;
        RECT 803.400 772.950 804.600 785.400 ;
        RECT 816.300 779.400 818.100 791.250 ;
        RECT 820.500 779.400 822.300 791.250 ;
        RECT 823.800 785.400 825.600 791.250 ;
        RECT 838.650 785.400 840.450 791.250 ;
        RECT 841.650 785.400 843.450 791.250 ;
        RECT 844.650 785.400 846.450 791.250 ;
        RECT 854.550 785.400 856.350 791.250 ;
        RECT 857.550 785.400 859.350 791.250 ;
        RECT 860.550 785.400 862.350 791.250 ;
        RECT 815.100 774.150 816.900 775.950 ;
        RECT 820.950 774.150 822.150 779.400 ;
        RECT 823.950 777.150 825.750 778.950 ;
        RECT 842.250 777.150 843.450 785.400 ;
        RECT 857.550 777.150 858.750 785.400 ;
        RECT 862.950 778.950 865.050 781.050 ;
        RECT 823.950 775.050 826.050 777.150 ;
        RECT 782.100 769.050 783.900 770.850 ;
        RECT 785.850 768.750 787.050 772.050 ;
        RECT 800.100 771.150 801.900 772.950 ;
        RECT 799.950 769.050 802.050 771.150 ;
        RECT 802.950 770.850 805.050 772.950 ;
        RECT 814.950 772.050 817.050 774.150 ;
        RECT 817.950 770.850 820.050 772.950 ;
        RECT 820.950 772.050 823.050 774.150 ;
        RECT 838.950 773.850 841.050 775.950 ;
        RECT 841.950 775.050 844.050 777.150 ;
        RECT 839.100 772.050 840.900 773.850 ;
        RECT 786.000 767.700 789.750 768.750 ;
        RECT 754.200 762.600 755.250 764.400 ;
        RECT 763.950 763.500 766.050 765.600 ;
        RECT 763.950 762.600 765.000 763.500 ;
        RECT 740.850 759.750 742.650 762.600 ;
        RECT 745.350 759.750 747.150 762.600 ;
        RECT 749.550 759.750 751.350 762.600 ;
        RECT 753.450 759.750 755.250 762.600 ;
        RECT 756.750 759.750 758.550 762.600 ;
        RECT 761.250 761.700 765.000 762.600 ;
        RECT 761.250 759.750 763.050 761.700 ;
        RECT 766.050 759.750 767.850 762.600 ;
        RECT 769.050 759.750 770.850 765.600 ;
        RECT 779.550 764.700 787.350 766.050 ;
        RECT 779.550 759.750 781.350 764.700 ;
        RECT 782.550 759.750 784.350 763.800 ;
        RECT 785.550 759.750 787.350 764.700 ;
        RECT 788.550 765.600 789.750 767.700 ;
        RECT 788.550 759.750 790.350 765.600 ;
        RECT 803.400 762.600 804.600 770.850 ;
        RECT 818.100 769.050 819.900 770.850 ;
        RECT 821.850 768.750 823.050 772.050 ;
        RECT 822.000 767.700 825.750 768.750 ;
        RECT 842.250 767.700 843.450 775.050 ;
        RECT 844.950 773.850 847.050 775.950 ;
        RECT 853.950 773.850 856.050 775.950 ;
        RECT 856.950 775.050 859.050 777.150 ;
        RECT 845.100 772.050 846.900 773.850 ;
        RECT 854.100 772.050 855.900 773.850 ;
        RECT 815.550 764.700 823.350 766.050 ;
        RECT 800.550 759.750 802.350 762.600 ;
        RECT 803.550 759.750 805.350 762.600 ;
        RECT 815.550 759.750 817.350 764.700 ;
        RECT 818.550 759.750 820.350 763.800 ;
        RECT 821.550 759.750 823.350 764.700 ;
        RECT 824.550 765.600 825.750 767.700 ;
        RECT 839.850 766.800 843.450 767.700 ;
        RECT 857.550 767.700 858.750 775.050 ;
        RECT 859.950 773.850 862.050 775.950 ;
        RECT 860.100 772.050 861.900 773.850 ;
        RECT 863.550 769.050 864.450 778.950 ;
        RECT 857.550 766.800 861.150 767.700 ;
        RECT 862.950 766.950 865.050 769.050 ;
        RECT 824.550 759.750 826.350 765.600 ;
        RECT 839.850 759.750 841.650 766.800 ;
        RECT 844.350 759.750 846.150 765.600 ;
        RECT 854.850 759.750 856.650 765.600 ;
        RECT 859.350 759.750 861.150 766.800 ;
        RECT 10.650 749.400 12.450 755.250 ;
        RECT 11.250 747.300 12.450 749.400 ;
        RECT 13.650 750.300 15.450 755.250 ;
        RECT 16.650 751.200 18.450 755.250 ;
        RECT 19.650 750.300 21.450 755.250 ;
        RECT 13.650 748.950 21.450 750.300 ;
        RECT 11.250 746.250 15.000 747.300 ;
        RECT 35.100 747.000 36.900 755.250 ;
        RECT 13.950 742.950 15.150 746.250 ;
        RECT 17.100 744.150 18.900 745.950 ;
        RECT 32.400 745.350 36.900 747.000 ;
        RECT 40.500 746.400 42.300 755.250 ;
        RECT 50.700 746.400 52.500 755.250 ;
        RECT 56.100 747.000 57.900 755.250 ;
        RECT 71.550 750.300 73.350 755.250 ;
        RECT 74.550 751.200 76.350 755.250 ;
        RECT 77.550 750.300 79.350 755.250 ;
        RECT 71.550 748.950 79.350 750.300 ;
        RECT 80.550 749.400 82.350 755.250 ;
        RECT 80.550 747.300 81.750 749.400 ;
        RECT 95.850 748.200 97.650 755.250 ;
        RECT 100.350 749.400 102.150 755.250 ;
        RECT 112.650 749.400 114.450 755.250 ;
        RECT 95.850 747.300 99.450 748.200 ;
        RECT 56.100 745.350 60.600 747.000 ;
        RECT 78.000 746.250 81.750 747.300 ;
        RECT 13.950 740.850 16.050 742.950 ;
        RECT 16.950 742.050 19.050 744.150 ;
        RECT 19.950 740.850 22.050 742.950 ;
        RECT 32.400 741.150 33.600 745.350 ;
        RECT 59.400 741.150 60.600 745.350 ;
        RECT 74.100 744.150 75.900 745.950 ;
        RECT 10.950 737.850 13.050 739.950 ;
        RECT 11.250 736.050 13.050 737.850 ;
        RECT 14.850 735.600 16.050 740.850 ;
        RECT 20.100 739.050 21.900 740.850 ;
        RECT 31.950 739.050 34.050 741.150 ;
        RECT 11.400 723.750 13.200 729.600 ;
        RECT 14.700 723.750 16.500 735.600 ;
        RECT 18.900 723.750 20.700 735.600 ;
        RECT 32.250 730.800 33.300 739.050 ;
        RECT 34.950 737.850 37.050 739.950 ;
        RECT 40.950 737.850 43.050 739.950 ;
        RECT 49.950 737.850 52.050 739.950 ;
        RECT 55.950 737.850 58.050 739.950 ;
        RECT 58.950 739.050 61.050 741.150 ;
        RECT 70.950 740.850 73.050 742.950 ;
        RECT 73.950 742.050 76.050 744.150 ;
        RECT 77.850 742.950 79.050 746.250 ;
        RECT 76.950 740.850 79.050 742.950 ;
        RECT 95.100 741.150 96.900 742.950 ;
        RECT 71.100 739.050 72.900 740.850 ;
        RECT 34.950 736.050 36.750 737.850 ;
        RECT 37.950 734.850 40.050 736.950 ;
        RECT 41.100 736.050 42.900 737.850 ;
        RECT 50.100 736.050 51.900 737.850 ;
        RECT 52.950 734.850 55.050 736.950 ;
        RECT 56.250 736.050 58.050 737.850 ;
        RECT 38.100 733.050 39.900 734.850 ;
        RECT 53.100 733.050 54.900 734.850 ;
        RECT 59.700 730.800 60.750 739.050 ;
        RECT 76.950 735.600 78.150 740.850 ;
        RECT 79.950 737.850 82.050 739.950 ;
        RECT 94.950 739.050 97.050 741.150 ;
        RECT 98.250 739.950 99.450 747.300 ;
        RECT 113.250 747.300 114.450 749.400 ;
        RECT 115.650 750.300 117.450 755.250 ;
        RECT 118.650 751.200 120.450 755.250 ;
        RECT 121.650 750.300 123.450 755.250 ;
        RECT 115.650 748.950 123.450 750.300 ;
        RECT 133.650 749.400 135.450 755.250 ;
        RECT 134.250 747.300 135.450 749.400 ;
        RECT 136.650 750.300 138.450 755.250 ;
        RECT 139.650 751.200 141.450 755.250 ;
        RECT 142.650 750.300 144.450 755.250 ;
        RECT 155.700 752.400 157.500 755.250 ;
        RECT 159.000 751.050 160.800 755.250 ;
        RECT 136.650 748.950 144.450 750.300 ;
        RECT 155.100 749.400 160.800 751.050 ;
        RECT 163.200 749.400 165.000 755.250 ;
        RECT 175.650 749.400 177.450 755.250 ;
        RECT 113.250 746.250 117.000 747.300 ;
        RECT 134.250 746.250 138.000 747.300 ;
        RECT 115.950 742.950 117.150 746.250 ;
        RECT 119.100 744.150 120.900 745.950 ;
        RECT 101.100 741.150 102.900 742.950 ;
        RECT 97.950 737.850 100.050 739.950 ;
        RECT 100.950 739.050 103.050 741.150 ;
        RECT 115.950 740.850 118.050 742.950 ;
        RECT 118.950 742.050 121.050 744.150 ;
        RECT 136.950 742.950 138.150 746.250 ;
        RECT 140.100 744.150 141.900 745.950 ;
        RECT 121.950 740.850 124.050 742.950 ;
        RECT 136.950 740.850 139.050 742.950 ;
        RECT 139.950 742.050 142.050 744.150 ;
        RECT 155.100 742.950 156.300 749.400 ;
        RECT 176.250 747.300 177.450 749.400 ;
        RECT 178.650 750.300 180.450 755.250 ;
        RECT 181.650 751.200 183.450 755.250 ;
        RECT 184.650 750.300 186.450 755.250 ;
        RECT 196.650 752.400 198.450 755.250 ;
        RECT 199.650 752.400 201.450 755.250 ;
        RECT 178.650 748.950 186.450 750.300 ;
        RECT 176.250 746.250 180.000 747.300 ;
        RECT 158.100 744.150 159.900 745.950 ;
        RECT 142.950 740.850 145.050 742.950 ;
        RECT 154.950 740.850 157.050 742.950 ;
        RECT 157.950 742.050 160.050 744.150 ;
        RECT 160.950 743.850 163.050 745.950 ;
        RECT 164.100 744.150 165.900 745.950 ;
        RECT 161.100 742.050 162.900 743.850 ;
        RECT 163.950 742.050 166.050 744.150 ;
        RECT 178.950 742.950 180.150 746.250 ;
        RECT 182.100 744.150 183.900 745.950 ;
        RECT 197.400 744.150 198.600 752.400 ;
        RECT 212.850 748.200 214.650 755.250 ;
        RECT 217.350 749.400 219.150 755.250 ;
        RECT 212.850 747.300 216.450 748.200 ;
        RECT 178.950 740.850 181.050 742.950 ;
        RECT 181.950 742.050 184.050 744.150 ;
        RECT 184.950 740.850 187.050 742.950 ;
        RECT 196.950 742.050 199.050 744.150 ;
        RECT 199.950 743.850 202.050 745.950 ;
        RECT 200.100 742.050 201.900 743.850 ;
        RECT 112.950 737.850 115.050 739.950 ;
        RECT 79.950 736.050 81.750 737.850 ;
        RECT 32.250 729.900 39.300 730.800 ;
        RECT 32.250 729.600 33.450 729.900 ;
        RECT 31.650 723.750 33.450 729.600 ;
        RECT 37.650 729.600 39.300 729.900 ;
        RECT 53.700 729.900 60.750 730.800 ;
        RECT 53.700 729.600 55.350 729.900 ;
        RECT 34.650 723.750 36.450 729.000 ;
        RECT 37.650 723.750 39.450 729.600 ;
        RECT 40.650 723.750 42.450 729.600 ;
        RECT 50.550 723.750 52.350 729.600 ;
        RECT 53.550 723.750 55.350 729.600 ;
        RECT 59.550 729.600 60.750 729.900 ;
        RECT 56.550 723.750 58.350 729.000 ;
        RECT 59.550 723.750 61.350 729.600 ;
        RECT 72.300 723.750 74.100 735.600 ;
        RECT 76.500 723.750 78.300 735.600 ;
        RECT 98.250 729.600 99.450 737.850 ;
        RECT 113.250 736.050 115.050 737.850 ;
        RECT 116.850 735.600 118.050 740.850 ;
        RECT 122.100 739.050 123.900 740.850 ;
        RECT 133.950 737.850 136.050 739.950 ;
        RECT 134.250 736.050 136.050 737.850 ;
        RECT 137.850 735.600 139.050 740.850 ;
        RECT 143.100 739.050 144.900 740.850 ;
        RECT 155.100 735.600 156.300 740.850 ;
        RECT 175.950 737.850 178.050 739.950 ;
        RECT 176.250 736.050 178.050 737.850 ;
        RECT 179.850 735.600 181.050 740.850 ;
        RECT 185.100 739.050 186.900 740.850 ;
        RECT 79.800 723.750 81.600 729.600 ;
        RECT 94.650 723.750 96.450 729.600 ;
        RECT 97.650 723.750 99.450 729.600 ;
        RECT 100.650 723.750 102.450 729.600 ;
        RECT 113.400 723.750 115.200 729.600 ;
        RECT 116.700 723.750 118.500 735.600 ;
        RECT 120.900 723.750 122.700 735.600 ;
        RECT 134.400 723.750 136.200 729.600 ;
        RECT 137.700 723.750 139.500 735.600 ;
        RECT 141.900 723.750 143.700 735.600 ;
        RECT 154.650 723.750 156.450 735.600 ;
        RECT 157.650 734.700 165.450 735.600 ;
        RECT 157.650 723.750 159.450 734.700 ;
        RECT 160.650 723.750 162.450 733.800 ;
        RECT 163.650 723.750 165.450 734.700 ;
        RECT 176.400 723.750 178.200 729.600 ;
        RECT 179.700 723.750 181.500 735.600 ;
        RECT 183.900 723.750 185.700 735.600 ;
        RECT 197.400 729.600 198.600 742.050 ;
        RECT 212.100 741.150 213.900 742.950 ;
        RECT 211.950 739.050 214.050 741.150 ;
        RECT 215.250 739.950 216.450 747.300 ;
        RECT 236.100 747.000 237.900 755.250 ;
        RECT 233.400 745.350 237.900 747.000 ;
        RECT 241.500 746.400 243.300 755.250 ;
        RECT 253.650 749.400 255.450 755.250 ;
        RECT 254.250 747.300 255.450 749.400 ;
        RECT 256.650 750.300 258.450 755.250 ;
        RECT 259.650 751.200 261.450 755.250 ;
        RECT 262.650 750.300 264.450 755.250 ;
        RECT 256.650 748.950 264.450 750.300 ;
        RECT 273.000 749.400 274.800 755.250 ;
        RECT 277.200 751.050 279.000 755.250 ;
        RECT 280.500 752.400 282.300 755.250 ;
        RECT 277.200 749.400 282.900 751.050 ;
        RECT 293.850 749.400 295.650 755.250 ;
        RECT 254.250 746.250 258.000 747.300 ;
        RECT 218.100 741.150 219.900 742.950 ;
        RECT 233.400 741.150 234.600 745.350 ;
        RECT 256.950 742.950 258.150 746.250 ;
        RECT 260.100 744.150 261.900 745.950 ;
        RECT 272.100 744.150 273.900 745.950 ;
        RECT 214.950 737.850 217.050 739.950 ;
        RECT 217.950 739.050 220.050 741.150 ;
        RECT 232.950 739.050 235.050 741.150 ;
        RECT 256.950 740.850 259.050 742.950 ;
        RECT 259.950 742.050 262.050 744.150 ;
        RECT 262.950 740.850 265.050 742.950 ;
        RECT 271.950 742.050 274.050 744.150 ;
        RECT 274.950 743.850 277.050 745.950 ;
        RECT 278.100 744.150 279.900 745.950 ;
        RECT 275.100 742.050 276.900 743.850 ;
        RECT 277.950 742.050 280.050 744.150 ;
        RECT 281.700 742.950 282.900 749.400 ;
        RECT 298.350 748.200 300.150 755.250 ;
        RECT 314.700 752.400 316.500 755.250 ;
        RECT 318.000 751.050 319.800 755.250 ;
        RECT 296.550 747.300 300.150 748.200 ;
        RECT 314.100 749.400 319.800 751.050 ;
        RECT 322.200 749.400 324.000 755.250 ;
        RECT 337.650 752.400 339.450 755.250 ;
        RECT 340.650 752.400 342.450 755.250 ;
        RECT 280.950 740.850 283.050 742.950 ;
        RECT 293.100 741.150 294.900 742.950 ;
        RECT 215.250 729.600 216.450 737.850 ;
        RECT 233.250 730.800 234.300 739.050 ;
        RECT 235.950 737.850 238.050 739.950 ;
        RECT 241.950 737.850 244.050 739.950 ;
        RECT 253.950 737.850 256.050 739.950 ;
        RECT 235.950 736.050 237.750 737.850 ;
        RECT 238.950 734.850 241.050 736.950 ;
        RECT 242.100 736.050 243.900 737.850 ;
        RECT 254.250 736.050 256.050 737.850 ;
        RECT 257.850 735.600 259.050 740.850 ;
        RECT 263.100 739.050 264.900 740.850 ;
        RECT 281.700 735.600 282.900 740.850 ;
        RECT 292.950 739.050 295.050 741.150 ;
        RECT 296.550 739.950 297.750 747.300 ;
        RECT 314.100 742.950 315.300 749.400 ;
        RECT 317.100 744.150 318.900 745.950 ;
        RECT 299.100 741.150 300.900 742.950 ;
        RECT 295.950 737.850 298.050 739.950 ;
        RECT 298.950 739.050 301.050 741.150 ;
        RECT 313.950 740.850 316.050 742.950 ;
        RECT 316.950 742.050 319.050 744.150 ;
        RECT 319.950 743.850 322.050 745.950 ;
        RECT 323.100 744.150 324.900 745.950 ;
        RECT 338.400 744.150 339.600 752.400 ;
        RECT 352.650 749.400 354.450 755.250 ;
        RECT 353.250 747.300 354.450 749.400 ;
        RECT 355.650 750.300 357.450 755.250 ;
        RECT 358.650 751.200 360.450 755.250 ;
        RECT 361.650 750.300 363.450 755.250 ;
        RECT 355.650 748.950 363.450 750.300 ;
        RECT 353.250 746.250 357.000 747.300 ;
        RECT 377.100 747.000 378.900 755.250 ;
        RECT 320.100 742.050 321.900 743.850 ;
        RECT 322.950 742.050 325.050 744.150 ;
        RECT 337.950 742.050 340.050 744.150 ;
        RECT 340.950 743.850 343.050 745.950 ;
        RECT 341.100 742.050 342.900 743.850 ;
        RECT 355.950 742.950 357.150 746.250 ;
        RECT 359.100 744.150 360.900 745.950 ;
        RECT 374.400 745.350 378.900 747.000 ;
        RECT 382.500 746.400 384.300 755.250 ;
        RECT 394.650 752.400 396.450 755.250 ;
        RECT 397.650 752.400 399.450 755.250 ;
        RECT 239.100 733.050 240.900 734.850 ;
        RECT 233.250 729.900 240.300 730.800 ;
        RECT 233.250 729.600 234.450 729.900 ;
        RECT 196.650 723.750 198.450 729.600 ;
        RECT 199.650 723.750 201.450 729.600 ;
        RECT 211.650 723.750 213.450 729.600 ;
        RECT 214.650 723.750 216.450 729.600 ;
        RECT 217.650 723.750 219.450 729.600 ;
        RECT 232.650 723.750 234.450 729.600 ;
        RECT 238.650 729.600 240.300 729.900 ;
        RECT 235.650 723.750 237.450 729.000 ;
        RECT 238.650 723.750 240.450 729.600 ;
        RECT 241.650 723.750 243.450 729.600 ;
        RECT 254.400 723.750 256.200 729.600 ;
        RECT 257.700 723.750 259.500 735.600 ;
        RECT 261.900 723.750 263.700 735.600 ;
        RECT 272.550 734.700 280.350 735.600 ;
        RECT 272.550 723.750 274.350 734.700 ;
        RECT 275.550 723.750 277.350 733.800 ;
        RECT 278.550 723.750 280.350 734.700 ;
        RECT 281.550 723.750 283.350 735.600 ;
        RECT 296.550 729.600 297.750 737.850 ;
        RECT 314.100 735.600 315.300 740.850 ;
        RECT 293.550 723.750 295.350 729.600 ;
        RECT 296.550 723.750 298.350 729.600 ;
        RECT 299.550 723.750 301.350 729.600 ;
        RECT 313.650 723.750 315.450 735.600 ;
        RECT 316.650 734.700 324.450 735.600 ;
        RECT 316.650 723.750 318.450 734.700 ;
        RECT 319.650 723.750 321.450 733.800 ;
        RECT 322.650 723.750 324.450 734.700 ;
        RECT 338.400 729.600 339.600 742.050 ;
        RECT 355.950 740.850 358.050 742.950 ;
        RECT 358.950 742.050 361.050 744.150 ;
        RECT 361.950 740.850 364.050 742.950 ;
        RECT 374.400 741.150 375.600 745.350 ;
        RECT 395.400 744.150 396.600 752.400 ;
        RECT 413.850 748.200 415.650 755.250 ;
        RECT 418.350 749.400 420.150 755.250 ;
        RECT 428.550 752.400 430.350 755.250 ;
        RECT 431.550 752.400 433.350 755.250 ;
        RECT 413.850 747.300 417.450 748.200 ;
        RECT 394.950 742.050 397.050 744.150 ;
        RECT 397.950 743.850 400.050 745.950 ;
        RECT 398.100 742.050 399.900 743.850 ;
        RECT 352.950 737.850 355.050 739.950 ;
        RECT 353.250 736.050 355.050 737.850 ;
        RECT 356.850 735.600 358.050 740.850 ;
        RECT 362.100 739.050 363.900 740.850 ;
        RECT 373.950 739.050 376.050 741.150 ;
        RECT 337.650 723.750 339.450 729.600 ;
        RECT 340.650 723.750 342.450 729.600 ;
        RECT 353.400 723.750 355.200 729.600 ;
        RECT 356.700 723.750 358.500 735.600 ;
        RECT 360.900 723.750 362.700 735.600 ;
        RECT 374.250 730.800 375.300 739.050 ;
        RECT 376.950 737.850 379.050 739.950 ;
        RECT 382.950 737.850 385.050 739.950 ;
        RECT 376.950 736.050 378.750 737.850 ;
        RECT 379.950 734.850 382.050 736.950 ;
        RECT 383.100 736.050 384.900 737.850 ;
        RECT 380.100 733.050 381.900 734.850 ;
        RECT 374.250 729.900 381.300 730.800 ;
        RECT 374.250 729.600 375.450 729.900 ;
        RECT 373.650 723.750 375.450 729.600 ;
        RECT 379.650 729.600 381.300 729.900 ;
        RECT 395.400 729.600 396.600 742.050 ;
        RECT 413.100 741.150 414.900 742.950 ;
        RECT 412.950 739.050 415.050 741.150 ;
        RECT 416.250 739.950 417.450 747.300 ;
        RECT 427.950 743.850 430.050 745.950 ;
        RECT 431.400 744.150 432.600 752.400 ;
        RECT 443.700 746.400 445.500 755.250 ;
        RECT 449.100 747.000 450.900 755.250 ;
        RECT 466.650 749.400 468.450 755.250 ;
        RECT 467.250 747.300 468.450 749.400 ;
        RECT 469.650 750.300 471.450 755.250 ;
        RECT 472.650 751.200 474.450 755.250 ;
        RECT 475.650 750.300 477.450 755.250 ;
        RECT 469.650 748.950 477.450 750.300 ;
        RECT 487.650 749.400 489.450 755.250 ;
        RECT 488.250 747.300 489.450 749.400 ;
        RECT 490.650 750.300 492.450 755.250 ;
        RECT 493.650 751.200 495.450 755.250 ;
        RECT 496.650 750.300 498.450 755.250 ;
        RECT 509.700 752.400 511.500 755.250 ;
        RECT 513.000 751.050 514.800 755.250 ;
        RECT 490.650 748.950 498.450 750.300 ;
        RECT 509.100 749.400 514.800 751.050 ;
        RECT 517.200 749.400 519.000 755.250 ;
        RECT 527.550 752.400 529.350 755.250 ;
        RECT 530.550 752.400 532.350 755.250 ;
        RECT 533.550 752.400 535.350 755.250 ;
        RECT 449.100 745.350 453.600 747.000 ;
        RECT 467.250 746.250 471.000 747.300 ;
        RECT 488.250 746.250 492.000 747.300 ;
        RECT 419.100 741.150 420.900 742.950 ;
        RECT 428.100 742.050 429.900 743.850 ;
        RECT 430.950 742.050 433.050 744.150 ;
        RECT 415.950 737.850 418.050 739.950 ;
        RECT 418.950 739.050 421.050 741.150 ;
        RECT 416.250 729.600 417.450 737.850 ;
        RECT 418.950 735.450 421.050 736.050 ;
        RECT 424.950 735.450 427.050 736.050 ;
        RECT 418.950 734.550 427.050 735.450 ;
        RECT 418.950 733.950 421.050 734.550 ;
        RECT 424.950 733.950 427.050 734.550 ;
        RECT 431.400 729.600 432.600 742.050 ;
        RECT 452.400 741.150 453.600 745.350 ;
        RECT 469.950 742.950 471.150 746.250 ;
        RECT 473.100 744.150 474.900 745.950 ;
        RECT 442.950 737.850 445.050 739.950 ;
        RECT 448.950 737.850 451.050 739.950 ;
        RECT 451.950 739.050 454.050 741.150 ;
        RECT 469.950 740.850 472.050 742.950 ;
        RECT 472.950 742.050 475.050 744.150 ;
        RECT 490.950 742.950 492.150 746.250 ;
        RECT 494.100 744.150 495.900 745.950 ;
        RECT 475.950 740.850 478.050 742.950 ;
        RECT 490.950 740.850 493.050 742.950 ;
        RECT 493.950 742.050 496.050 744.150 ;
        RECT 509.100 742.950 510.300 749.400 ;
        RECT 531.450 748.200 532.350 752.400 ;
        RECT 536.550 749.400 538.350 755.250 ;
        RECT 550.650 752.400 552.450 755.250 ;
        RECT 553.650 752.400 555.450 755.250 ;
        RECT 556.650 752.400 558.450 755.250 ;
        RECT 531.450 747.300 534.750 748.200 ;
        RECT 532.950 746.400 534.750 747.300 ;
        RECT 512.100 744.150 513.900 745.950 ;
        RECT 496.950 740.850 499.050 742.950 ;
        RECT 508.950 740.850 511.050 742.950 ;
        RECT 511.950 742.050 514.050 744.150 ;
        RECT 514.950 743.850 517.050 745.950 ;
        RECT 518.100 744.150 519.900 745.950 ;
        RECT 515.100 742.050 516.900 743.850 ;
        RECT 517.950 742.050 520.050 744.150 ;
        RECT 526.950 743.850 529.050 745.950 ;
        RECT 527.100 742.050 528.900 743.850 ;
        RECT 529.950 740.850 532.050 742.950 ;
        RECT 443.100 736.050 444.900 737.850 ;
        RECT 445.950 734.850 448.050 736.950 ;
        RECT 449.250 736.050 451.050 737.850 ;
        RECT 446.100 733.050 447.900 734.850 ;
        RECT 452.700 730.800 453.750 739.050 ;
        RECT 466.950 737.850 469.050 739.950 ;
        RECT 467.250 736.050 469.050 737.850 ;
        RECT 470.850 735.600 472.050 740.850 ;
        RECT 476.100 739.050 477.900 740.850 ;
        RECT 487.950 737.850 490.050 739.950 ;
        RECT 488.250 736.050 490.050 737.850 ;
        RECT 491.850 735.600 493.050 740.850 ;
        RECT 497.100 739.050 498.900 740.850 ;
        RECT 509.100 735.600 510.300 740.850 ;
        RECT 530.100 739.050 531.900 740.850 ;
        RECT 533.700 738.150 534.600 746.400 ;
        RECT 537.000 744.150 538.050 749.400 ;
        RECT 535.950 742.050 538.050 744.150 ;
        RECT 553.950 745.950 555.000 752.400 ;
        RECT 572.100 747.000 573.900 755.250 ;
        RECT 553.950 743.850 556.050 745.950 ;
        RECT 569.400 745.350 573.900 747.000 ;
        RECT 577.500 746.400 579.300 755.250 ;
        RECT 589.650 752.400 591.450 755.250 ;
        RECT 592.650 752.400 594.450 755.250 ;
        RECT 532.950 738.000 534.750 738.150 ;
        RECT 527.550 736.800 534.750 738.000 ;
        RECT 527.550 735.600 528.750 736.800 ;
        RECT 532.950 736.350 534.750 736.800 ;
        RECT 446.700 729.900 453.750 730.800 ;
        RECT 446.700 729.600 448.350 729.900 ;
        RECT 376.650 723.750 378.450 729.000 ;
        RECT 379.650 723.750 381.450 729.600 ;
        RECT 382.650 723.750 384.450 729.600 ;
        RECT 394.650 723.750 396.450 729.600 ;
        RECT 397.650 723.750 399.450 729.600 ;
        RECT 412.650 723.750 414.450 729.600 ;
        RECT 415.650 723.750 417.450 729.600 ;
        RECT 418.650 723.750 420.450 729.600 ;
        RECT 428.550 723.750 430.350 729.600 ;
        RECT 431.550 723.750 433.350 729.600 ;
        RECT 443.550 723.750 445.350 729.600 ;
        RECT 446.550 723.750 448.350 729.600 ;
        RECT 452.550 729.600 453.750 729.900 ;
        RECT 449.550 723.750 451.350 729.000 ;
        RECT 452.550 723.750 454.350 729.600 ;
        RECT 467.400 723.750 469.200 729.600 ;
        RECT 470.700 723.750 472.500 735.600 ;
        RECT 474.900 723.750 476.700 735.600 ;
        RECT 488.400 723.750 490.200 729.600 ;
        RECT 491.700 723.750 493.500 735.600 ;
        RECT 495.900 723.750 497.700 735.600 ;
        RECT 508.650 723.750 510.450 735.600 ;
        RECT 511.650 734.700 519.450 735.600 ;
        RECT 511.650 723.750 513.450 734.700 ;
        RECT 514.650 723.750 516.450 733.800 ;
        RECT 517.650 723.750 519.450 734.700 ;
        RECT 527.550 723.750 529.350 735.600 ;
        RECT 536.100 735.450 537.450 742.050 ;
        RECT 550.950 740.850 553.050 742.950 ;
        RECT 551.100 739.050 552.900 740.850 ;
        RECT 553.950 736.650 555.000 743.850 ;
        RECT 556.950 740.850 559.050 742.950 ;
        RECT 569.400 741.150 570.600 745.350 ;
        RECT 590.400 744.150 591.600 752.400 ;
        RECT 602.700 746.400 604.500 755.250 ;
        RECT 608.100 747.000 609.900 755.250 ;
        RECT 589.950 742.050 592.050 744.150 ;
        RECT 592.950 743.850 595.050 745.950 ;
        RECT 608.100 745.350 612.600 747.000 ;
        RECT 623.700 746.400 625.500 755.250 ;
        RECT 629.100 747.000 630.900 755.250 ;
        RECT 648.150 750.900 649.950 755.250 ;
        RECT 646.650 749.400 649.950 750.900 ;
        RECT 651.150 749.400 652.950 755.250 ;
        RECT 629.100 745.350 633.600 747.000 ;
        RECT 593.100 742.050 594.900 743.850 ;
        RECT 557.100 739.050 558.900 740.850 ;
        RECT 568.950 739.050 571.050 741.150 ;
        RECT 532.050 723.750 533.850 735.450 ;
        RECT 535.050 734.100 537.450 735.450 ;
        RECT 552.450 735.600 555.000 736.650 ;
        RECT 535.050 723.750 536.850 734.100 ;
        RECT 552.450 723.750 554.250 735.600 ;
        RECT 556.650 723.750 558.450 735.600 ;
        RECT 569.250 730.800 570.300 739.050 ;
        RECT 571.950 737.850 574.050 739.950 ;
        RECT 577.950 737.850 580.050 739.950 ;
        RECT 571.950 736.050 573.750 737.850 ;
        RECT 574.950 734.850 577.050 736.950 ;
        RECT 578.100 736.050 579.900 737.850 ;
        RECT 575.100 733.050 576.900 734.850 ;
        RECT 569.250 729.900 576.300 730.800 ;
        RECT 569.250 729.600 570.450 729.900 ;
        RECT 568.650 723.750 570.450 729.600 ;
        RECT 574.650 729.600 576.300 729.900 ;
        RECT 590.400 729.600 591.600 742.050 ;
        RECT 611.400 741.150 612.600 745.350 ;
        RECT 616.950 744.450 619.050 745.050 ;
        RECT 625.950 744.450 628.050 745.050 ;
        RECT 616.950 743.550 628.050 744.450 ;
        RECT 616.950 742.950 619.050 743.550 ;
        RECT 625.950 742.950 628.050 743.550 ;
        RECT 632.400 741.150 633.600 745.350 ;
        RECT 646.650 742.950 647.850 749.400 ;
        RECT 649.950 747.900 651.750 748.500 ;
        RECT 655.650 747.900 657.450 755.250 ;
        RECT 668.550 752.400 670.350 755.250 ;
        RECT 671.550 752.400 673.350 755.250 ;
        RECT 674.550 752.400 676.350 755.250 ;
        RECT 649.950 746.700 657.450 747.900 ;
        RECT 672.450 748.200 673.350 752.400 ;
        RECT 677.550 749.400 679.350 755.250 ;
        RECT 689.550 752.400 691.350 755.250 ;
        RECT 692.550 752.400 694.350 755.250 ;
        RECT 695.550 752.400 697.350 755.250 ;
        RECT 672.450 747.300 675.750 748.200 ;
        RECT 601.950 737.850 604.050 739.950 ;
        RECT 607.950 737.850 610.050 739.950 ;
        RECT 610.950 739.050 613.050 741.150 ;
        RECT 602.100 736.050 603.900 737.850 ;
        RECT 604.950 734.850 607.050 736.950 ;
        RECT 608.250 736.050 610.050 737.850 ;
        RECT 605.100 733.050 606.900 734.850 ;
        RECT 611.700 730.800 612.750 739.050 ;
        RECT 622.950 737.850 625.050 739.950 ;
        RECT 628.950 737.850 631.050 739.950 ;
        RECT 631.950 739.050 634.050 741.150 ;
        RECT 646.650 740.850 649.050 742.950 ;
        RECT 650.100 741.150 651.900 742.950 ;
        RECT 623.100 736.050 624.900 737.850 ;
        RECT 625.950 734.850 628.050 736.950 ;
        RECT 629.250 736.050 631.050 737.850 ;
        RECT 626.100 733.050 627.900 734.850 ;
        RECT 632.700 730.800 633.750 739.050 ;
        RECT 646.650 735.600 647.850 740.850 ;
        RECT 649.950 739.050 652.050 741.150 ;
        RECT 605.700 729.900 612.750 730.800 ;
        RECT 605.700 729.600 607.350 729.900 ;
        RECT 571.650 723.750 573.450 729.000 ;
        RECT 574.650 723.750 576.450 729.600 ;
        RECT 577.650 723.750 579.450 729.600 ;
        RECT 589.650 723.750 591.450 729.600 ;
        RECT 592.650 723.750 594.450 729.600 ;
        RECT 602.550 723.750 604.350 729.600 ;
        RECT 605.550 723.750 607.350 729.600 ;
        RECT 611.550 729.600 612.750 729.900 ;
        RECT 626.700 729.900 633.750 730.800 ;
        RECT 626.700 729.600 628.350 729.900 ;
        RECT 608.550 723.750 610.350 729.000 ;
        RECT 611.550 723.750 613.350 729.600 ;
        RECT 623.550 723.750 625.350 729.600 ;
        RECT 626.550 723.750 628.350 729.600 ;
        RECT 632.550 729.600 633.750 729.900 ;
        RECT 629.550 723.750 631.350 729.000 ;
        RECT 632.550 723.750 634.350 729.600 ;
        RECT 646.050 723.750 647.850 735.600 ;
        RECT 649.050 723.750 650.850 735.600 ;
        RECT 653.100 729.600 654.300 746.700 ;
        RECT 673.950 746.400 675.750 747.300 ;
        RECT 667.950 743.850 670.050 745.950 ;
        RECT 655.950 740.850 658.050 742.950 ;
        RECT 668.100 742.050 669.900 743.850 ;
        RECT 670.950 740.850 673.050 742.950 ;
        RECT 656.100 739.050 657.900 740.850 ;
        RECT 671.100 739.050 672.900 740.850 ;
        RECT 674.700 738.150 675.600 746.400 ;
        RECT 678.000 744.150 679.050 749.400 ;
        RECT 693.000 745.950 694.050 752.400 ;
        RECT 709.650 749.400 711.450 755.250 ;
        RECT 710.250 747.300 711.450 749.400 ;
        RECT 712.650 750.300 714.450 755.250 ;
        RECT 715.650 751.200 717.450 755.250 ;
        RECT 718.650 750.300 720.450 755.250 ;
        RECT 712.650 748.950 720.450 750.300 ;
        RECT 722.550 749.400 724.350 755.250 ;
        RECT 725.850 752.400 727.650 755.250 ;
        RECT 730.350 752.400 732.150 755.250 ;
        RECT 734.550 752.400 736.350 755.250 ;
        RECT 738.450 752.400 740.250 755.250 ;
        RECT 741.750 752.400 743.550 755.250 ;
        RECT 746.250 753.300 748.050 755.250 ;
        RECT 746.250 752.400 750.000 753.300 ;
        RECT 751.050 752.400 752.850 755.250 ;
        RECT 730.650 751.500 731.700 752.400 ;
        RECT 727.950 750.300 731.700 751.500 ;
        RECT 739.200 750.600 740.250 752.400 ;
        RECT 748.950 751.500 750.000 752.400 ;
        RECT 727.950 749.400 730.050 750.300 ;
        RECT 710.250 746.250 714.000 747.300 ;
        RECT 722.550 747.150 723.750 749.400 ;
        RECT 735.150 748.200 736.950 750.000 ;
        RECT 739.200 749.550 744.150 750.600 ;
        RECT 742.350 748.800 744.150 749.550 ;
        RECT 745.650 748.800 747.450 750.600 ;
        RECT 748.950 749.400 751.050 751.500 ;
        RECT 754.050 749.400 755.850 755.250 ;
        RECT 736.050 747.900 736.950 748.200 ;
        RECT 746.100 747.900 747.150 748.800 ;
        RECT 676.950 742.050 679.050 744.150 ;
        RECT 691.950 743.850 694.050 745.950 ;
        RECT 673.950 738.000 675.750 738.150 ;
        RECT 668.550 736.800 675.750 738.000 ;
        RECT 668.550 735.600 669.750 736.800 ;
        RECT 673.950 736.350 675.750 736.800 ;
        RECT 652.650 723.750 654.450 729.600 ;
        RECT 655.650 723.750 657.450 729.600 ;
        RECT 668.550 723.750 670.350 735.600 ;
        RECT 677.100 735.450 678.450 742.050 ;
        RECT 688.950 740.850 691.050 742.950 ;
        RECT 689.100 739.050 690.900 740.850 ;
        RECT 693.000 736.650 694.050 743.850 ;
        RECT 712.950 742.950 714.150 746.250 ;
        RECT 716.100 744.150 717.900 745.950 ;
        RECT 722.550 745.050 727.050 747.150 ;
        RECT 736.050 747.000 747.150 747.900 ;
        RECT 694.950 740.850 697.050 742.950 ;
        RECT 712.950 740.850 715.050 742.950 ;
        RECT 715.950 742.050 718.050 744.150 ;
        RECT 718.950 740.850 721.050 742.950 ;
        RECT 695.100 739.050 696.900 740.850 ;
        RECT 709.950 737.850 712.050 739.950 ;
        RECT 693.000 735.600 695.550 736.650 ;
        RECT 710.250 736.050 712.050 737.850 ;
        RECT 713.850 735.600 715.050 740.850 ;
        RECT 719.100 739.050 720.900 740.850 ;
        RECT 722.550 735.600 723.750 745.050 ;
        RECT 724.950 743.250 728.850 745.050 ;
        RECT 724.950 742.950 727.050 743.250 ;
        RECT 736.050 742.950 736.950 747.000 ;
        RECT 746.100 745.800 747.150 747.000 ;
        RECT 746.100 744.600 753.000 745.800 ;
        RECT 746.100 744.000 747.900 744.600 ;
        RECT 752.100 743.850 753.000 744.600 ;
        RECT 749.100 742.950 750.900 743.700 ;
        RECT 736.050 740.850 739.050 742.950 ;
        RECT 742.950 741.900 750.900 742.950 ;
        RECT 752.100 742.050 753.900 743.850 ;
        RECT 742.950 740.850 745.050 741.900 ;
        RECT 724.950 737.400 726.750 739.200 ;
        RECT 725.850 736.200 730.050 737.400 ;
        RECT 736.050 736.200 736.950 740.850 ;
        RECT 744.750 737.100 746.550 737.400 ;
        RECT 673.050 723.750 674.850 735.450 ;
        RECT 676.050 734.100 678.450 735.450 ;
        RECT 676.050 723.750 677.850 734.100 ;
        RECT 689.550 723.750 691.350 735.600 ;
        RECT 693.750 723.750 695.550 735.600 ;
        RECT 710.400 723.750 712.200 729.600 ;
        RECT 713.700 723.750 715.500 735.600 ;
        RECT 717.900 723.750 719.700 735.600 ;
        RECT 722.550 723.750 724.350 735.600 ;
        RECT 727.950 735.300 730.050 736.200 ;
        RECT 730.950 735.300 736.950 736.200 ;
        RECT 738.150 736.800 746.550 737.100 ;
        RECT 754.950 736.800 755.850 749.400 ;
        RECT 764.550 750.300 766.350 755.250 ;
        RECT 767.550 751.200 769.350 755.250 ;
        RECT 770.550 750.300 772.350 755.250 ;
        RECT 764.550 748.950 772.350 750.300 ;
        RECT 773.550 749.400 775.350 755.250 ;
        RECT 779.550 749.400 781.350 755.250 ;
        RECT 782.850 752.400 784.650 755.250 ;
        RECT 787.350 752.400 789.150 755.250 ;
        RECT 791.550 752.400 793.350 755.250 ;
        RECT 795.450 752.400 797.250 755.250 ;
        RECT 798.750 752.400 800.550 755.250 ;
        RECT 803.250 753.300 805.050 755.250 ;
        RECT 803.250 752.400 807.000 753.300 ;
        RECT 808.050 752.400 809.850 755.250 ;
        RECT 787.650 751.500 788.700 752.400 ;
        RECT 784.950 750.300 788.700 751.500 ;
        RECT 796.200 750.600 797.250 752.400 ;
        RECT 805.950 751.500 807.000 752.400 ;
        RECT 784.950 749.400 787.050 750.300 ;
        RECT 773.550 747.300 774.750 749.400 ;
        RECT 771.000 746.250 774.750 747.300 ;
        RECT 779.550 747.150 780.750 749.400 ;
        RECT 792.150 748.200 793.950 750.000 ;
        RECT 796.200 749.550 801.150 750.600 ;
        RECT 799.350 748.800 801.150 749.550 ;
        RECT 802.650 748.800 804.450 750.600 ;
        RECT 805.950 749.400 808.050 751.500 ;
        RECT 811.050 749.400 812.850 755.250 ;
        RECT 793.050 747.900 793.950 748.200 ;
        RECT 803.100 747.900 804.150 748.800 ;
        RECT 767.100 744.150 768.900 745.950 ;
        RECT 763.950 740.850 766.050 742.950 ;
        RECT 766.950 742.050 769.050 744.150 ;
        RECT 770.850 742.950 772.050 746.250 ;
        RECT 769.950 740.850 772.050 742.950 ;
        RECT 779.550 745.050 784.050 747.150 ;
        RECT 793.050 747.000 804.150 747.900 ;
        RECT 764.100 739.050 765.900 740.850 ;
        RECT 738.150 736.200 755.850 736.800 ;
        RECT 730.950 734.400 731.850 735.300 ;
        RECT 729.150 732.600 731.850 734.400 ;
        RECT 732.750 734.100 734.550 734.400 ;
        RECT 738.150 734.100 739.050 736.200 ;
        RECT 744.750 735.600 755.850 736.200 ;
        RECT 769.950 735.600 771.150 740.850 ;
        RECT 772.950 737.850 775.050 739.950 ;
        RECT 772.950 736.050 774.750 737.850 ;
        RECT 779.550 735.600 780.750 745.050 ;
        RECT 781.950 743.250 785.850 745.050 ;
        RECT 781.950 742.950 784.050 743.250 ;
        RECT 793.050 742.950 793.950 747.000 ;
        RECT 803.100 745.800 804.150 747.000 ;
        RECT 803.100 744.600 810.000 745.800 ;
        RECT 803.100 744.000 804.900 744.600 ;
        RECT 809.100 743.850 810.000 744.600 ;
        RECT 806.100 742.950 807.900 743.700 ;
        RECT 793.050 740.850 796.050 742.950 ;
        RECT 799.950 741.900 807.900 742.950 ;
        RECT 809.100 742.050 810.900 743.850 ;
        RECT 799.950 740.850 802.050 741.900 ;
        RECT 781.950 737.400 783.750 739.200 ;
        RECT 782.850 736.200 787.050 737.400 ;
        RECT 793.050 736.200 793.950 740.850 ;
        RECT 801.750 737.100 803.550 737.400 ;
        RECT 732.750 733.200 739.050 734.100 ;
        RECT 739.950 734.700 741.750 735.300 ;
        RECT 739.950 733.500 747.450 734.700 ;
        RECT 732.750 732.600 734.550 733.200 ;
        RECT 746.250 732.600 747.450 733.500 ;
        RECT 727.950 729.600 731.850 731.700 ;
        RECT 736.950 730.500 743.850 732.300 ;
        RECT 746.250 730.500 751.050 732.600 ;
        RECT 725.550 723.750 727.350 726.600 ;
        RECT 730.050 723.750 731.850 729.600 ;
        RECT 734.250 723.750 736.050 729.600 ;
        RECT 738.150 723.750 739.950 730.500 ;
        RECT 746.250 729.600 747.450 730.500 ;
        RECT 741.150 723.750 742.950 729.600 ;
        RECT 745.950 723.750 747.750 729.600 ;
        RECT 751.050 723.750 752.850 729.600 ;
        RECT 754.050 723.750 755.850 735.600 ;
        RECT 765.300 723.750 767.100 735.600 ;
        RECT 769.500 723.750 771.300 735.600 ;
        RECT 772.800 723.750 774.600 729.600 ;
        RECT 779.550 723.750 781.350 735.600 ;
        RECT 784.950 735.300 787.050 736.200 ;
        RECT 787.950 735.300 793.950 736.200 ;
        RECT 795.150 736.800 803.550 737.100 ;
        RECT 811.950 736.800 812.850 749.400 ;
        RECT 824.850 748.200 826.650 755.250 ;
        RECT 829.350 749.400 831.150 755.250 ;
        RECT 839.850 749.400 841.650 755.250 ;
        RECT 844.350 748.200 846.150 755.250 ;
        RECT 860.850 749.400 862.650 755.250 ;
        RECT 865.350 748.200 867.150 755.250 ;
        RECT 824.850 747.300 828.450 748.200 ;
        RECT 824.100 741.150 825.900 742.950 ;
        RECT 823.950 739.050 826.050 741.150 ;
        RECT 827.250 739.950 828.450 747.300 ;
        RECT 832.950 745.950 835.050 748.050 ;
        RECT 838.950 747.450 841.050 748.050 ;
        RECT 836.550 746.550 841.050 747.450 ;
        RECT 830.100 741.150 831.900 742.950 ;
        RECT 826.950 737.850 829.050 739.950 ;
        RECT 829.950 739.050 832.050 741.150 ;
        RECT 795.150 736.200 812.850 736.800 ;
        RECT 787.950 734.400 788.850 735.300 ;
        RECT 786.150 732.600 788.850 734.400 ;
        RECT 789.750 734.100 791.550 734.400 ;
        RECT 795.150 734.100 796.050 736.200 ;
        RECT 801.750 735.600 812.850 736.200 ;
        RECT 789.750 733.200 796.050 734.100 ;
        RECT 796.950 734.700 798.750 735.300 ;
        RECT 796.950 733.500 804.450 734.700 ;
        RECT 789.750 732.600 791.550 733.200 ;
        RECT 803.250 732.600 804.450 733.500 ;
        RECT 784.950 729.600 788.850 731.700 ;
        RECT 793.950 730.500 800.850 732.300 ;
        RECT 803.250 730.500 808.050 732.600 ;
        RECT 782.550 723.750 784.350 726.600 ;
        RECT 787.050 723.750 788.850 729.600 ;
        RECT 791.250 723.750 793.050 729.600 ;
        RECT 795.150 723.750 796.950 730.500 ;
        RECT 803.250 729.600 804.450 730.500 ;
        RECT 798.150 723.750 799.950 729.600 ;
        RECT 802.950 723.750 804.750 729.600 ;
        RECT 808.050 723.750 809.850 729.600 ;
        RECT 811.050 723.750 812.850 735.600 ;
        RECT 827.250 729.600 828.450 737.850 ;
        RECT 829.950 735.450 832.050 736.050 ;
        RECT 833.550 735.450 834.450 745.950 ;
        RECT 829.950 734.550 834.450 735.450 ;
        RECT 836.550 735.450 837.450 746.550 ;
        RECT 838.950 745.950 841.050 746.550 ;
        RECT 842.550 747.300 846.150 748.200 ;
        RECT 863.550 747.300 867.150 748.200 ;
        RECT 839.100 741.150 840.900 742.950 ;
        RECT 838.950 739.050 841.050 741.150 ;
        RECT 842.550 739.950 843.750 747.300 ;
        RECT 845.100 741.150 846.900 742.950 ;
        RECT 860.100 741.150 861.900 742.950 ;
        RECT 841.950 737.850 844.050 739.950 ;
        RECT 844.950 739.050 847.050 741.150 ;
        RECT 859.950 739.050 862.050 741.150 ;
        RECT 863.550 739.950 864.750 747.300 ;
        RECT 866.100 741.150 867.900 742.950 ;
        RECT 862.950 737.850 865.050 739.950 ;
        RECT 865.950 739.050 868.050 741.150 ;
        RECT 836.550 734.550 840.450 735.450 ;
        RECT 829.950 733.950 832.050 734.550 ;
        RECT 839.550 733.050 840.450 734.550 ;
        RECT 838.950 730.950 841.050 733.050 ;
        RECT 842.550 729.600 843.750 737.850 ;
        RECT 863.550 729.600 864.750 737.850 ;
        RECT 823.650 723.750 825.450 729.600 ;
        RECT 826.650 723.750 828.450 729.600 ;
        RECT 829.650 723.750 831.450 729.600 ;
        RECT 839.550 723.750 841.350 729.600 ;
        RECT 842.550 723.750 844.350 729.600 ;
        RECT 845.550 723.750 847.350 729.600 ;
        RECT 860.550 723.750 862.350 729.600 ;
        RECT 863.550 723.750 865.350 729.600 ;
        RECT 866.550 723.750 868.350 729.600 ;
        RECT 10.650 707.400 12.450 719.250 ;
        RECT 13.650 708.300 15.450 719.250 ;
        RECT 16.650 709.200 18.450 719.250 ;
        RECT 19.650 708.300 21.450 719.250 ;
        RECT 31.650 713.400 33.450 719.250 ;
        RECT 34.650 714.000 36.450 719.250 ;
        RECT 13.650 707.400 21.450 708.300 ;
        RECT 32.250 713.100 33.450 713.400 ;
        RECT 37.650 713.400 39.450 719.250 ;
        RECT 40.650 713.400 42.450 719.250 ;
        RECT 37.650 713.100 39.300 713.400 ;
        RECT 32.250 712.200 39.300 713.100 ;
        RECT 11.100 702.150 12.300 707.400 ;
        RECT 32.250 703.950 33.300 712.200 ;
        RECT 38.100 708.150 39.900 709.950 ;
        RECT 50.550 708.300 52.350 719.250 ;
        RECT 53.550 709.200 55.350 719.250 ;
        RECT 56.550 708.300 58.350 719.250 ;
        RECT 34.950 705.150 36.750 706.950 ;
        RECT 37.950 706.050 40.050 708.150 ;
        RECT 50.550 707.400 58.350 708.300 ;
        RECT 59.550 707.400 61.350 719.250 ;
        RECT 71.550 713.400 73.350 719.250 ;
        RECT 74.550 713.400 76.350 719.250 ;
        RECT 77.550 713.400 79.350 719.250 ;
        RECT 91.650 713.400 93.450 719.250 ;
        RECT 94.650 714.000 96.450 719.250 ;
        RECT 41.100 705.150 42.900 706.950 ;
        RECT 10.950 700.050 13.050 702.150 ;
        RECT 31.950 701.850 34.050 703.950 ;
        RECT 34.950 703.050 37.050 705.150 ;
        RECT 40.950 703.050 43.050 705.150 ;
        RECT 59.700 702.150 60.900 707.400 ;
        RECT 74.550 705.150 75.750 713.400 ;
        RECT 92.250 713.100 93.450 713.400 ;
        RECT 97.650 713.400 99.450 719.250 ;
        RECT 100.650 713.400 102.450 719.250 ;
        RECT 115.650 713.400 117.450 719.250 ;
        RECT 118.650 714.000 120.450 719.250 ;
        RECT 97.650 713.100 99.300 713.400 ;
        RECT 92.250 712.200 99.300 713.100 ;
        RECT 116.250 713.100 117.450 713.400 ;
        RECT 121.650 713.400 123.450 719.250 ;
        RECT 124.650 713.400 126.450 719.250 ;
        RECT 134.550 713.400 136.350 719.250 ;
        RECT 137.550 713.400 139.350 719.250 ;
        RECT 149.550 713.400 151.350 719.250 ;
        RECT 152.550 713.400 154.350 719.250 ;
        RECT 166.650 713.400 168.450 719.250 ;
        RECT 169.650 713.400 171.450 719.250 ;
        RECT 182.400 713.400 184.200 719.250 ;
        RECT 121.650 713.100 123.300 713.400 ;
        RECT 116.250 712.200 123.300 713.100 ;
        RECT 11.100 693.600 12.300 700.050 ;
        RECT 13.950 698.850 16.050 700.950 ;
        RECT 17.100 699.150 18.900 700.950 ;
        RECT 14.100 697.050 15.900 698.850 ;
        RECT 16.950 697.050 19.050 699.150 ;
        RECT 19.950 698.850 22.050 700.950 ;
        RECT 20.100 697.050 21.900 698.850 ;
        RECT 32.400 697.650 33.600 701.850 ;
        RECT 49.950 698.850 52.050 700.950 ;
        RECT 53.100 699.150 54.900 700.950 ;
        RECT 32.400 696.000 36.900 697.650 ;
        RECT 50.100 697.050 51.900 698.850 ;
        RECT 52.950 697.050 55.050 699.150 ;
        RECT 55.950 698.850 58.050 700.950 ;
        RECT 58.950 700.050 61.050 702.150 ;
        RECT 70.950 701.850 73.050 703.950 ;
        RECT 73.950 703.050 76.050 705.150 ;
        RECT 92.250 703.950 93.300 712.200 ;
        RECT 98.100 708.150 99.900 709.950 ;
        RECT 94.950 705.150 96.750 706.950 ;
        RECT 97.950 706.050 100.050 708.150 ;
        RECT 101.100 705.150 102.900 706.950 ;
        RECT 71.100 700.050 72.900 701.850 ;
        RECT 56.100 697.050 57.900 698.850 ;
        RECT 11.100 691.950 16.800 693.600 ;
        RECT 11.700 687.750 13.500 690.600 ;
        RECT 15.000 687.750 16.800 691.950 ;
        RECT 19.200 687.750 21.000 693.600 ;
        RECT 35.100 687.750 36.900 696.000 ;
        RECT 40.500 687.750 42.300 696.600 ;
        RECT 59.700 693.600 60.900 700.050 ;
        RECT 74.550 695.700 75.750 703.050 ;
        RECT 76.950 701.850 79.050 703.950 ;
        RECT 91.950 701.850 94.050 703.950 ;
        RECT 94.950 703.050 97.050 705.150 ;
        RECT 100.950 703.050 103.050 705.150 ;
        RECT 116.250 703.950 117.300 712.200 ;
        RECT 122.100 708.150 123.900 709.950 ;
        RECT 118.950 705.150 120.750 706.950 ;
        RECT 121.950 706.050 124.050 708.150 ;
        RECT 125.100 705.150 126.900 706.950 ;
        RECT 115.950 701.850 118.050 703.950 ;
        RECT 118.950 703.050 121.050 705.150 ;
        RECT 124.950 703.050 127.050 705.150 ;
        RECT 77.100 700.050 78.900 701.850 ;
        RECT 92.400 697.650 93.600 701.850 ;
        RECT 116.400 697.650 117.600 701.850 ;
        RECT 137.400 700.950 138.600 713.400 ;
        RECT 152.400 700.950 153.600 713.400 ;
        RECT 167.400 700.950 168.600 713.400 ;
        RECT 185.700 707.400 187.500 719.250 ;
        RECT 189.900 707.400 191.700 719.250 ;
        RECT 201.300 707.400 203.100 719.250 ;
        RECT 205.500 707.400 207.300 719.250 ;
        RECT 208.800 713.400 210.600 719.250 ;
        RECT 221.550 713.400 223.350 719.250 ;
        RECT 224.550 713.400 226.350 719.250 ;
        RECT 236.550 713.400 238.350 719.250 ;
        RECT 239.550 713.400 241.350 719.250 ;
        RECT 242.550 714.000 244.350 719.250 ;
        RECT 182.250 705.150 184.050 706.950 ;
        RECT 181.950 703.050 184.050 705.150 ;
        RECT 185.850 702.150 187.050 707.400 ;
        RECT 191.100 702.150 192.900 703.950 ;
        RECT 200.100 702.150 201.900 703.950 ;
        RECT 205.950 702.150 207.150 707.400 ;
        RECT 208.950 705.150 210.750 706.950 ;
        RECT 208.950 703.050 211.050 705.150 ;
        RECT 134.100 699.150 135.900 700.950 ;
        RECT 92.400 696.000 96.900 697.650 ;
        RECT 74.550 694.800 78.150 695.700 ;
        RECT 51.000 687.750 52.800 693.600 ;
        RECT 55.200 691.950 60.900 693.600 ;
        RECT 55.200 687.750 57.000 691.950 ;
        RECT 58.500 687.750 60.300 690.600 ;
        RECT 71.850 687.750 73.650 693.600 ;
        RECT 76.350 687.750 78.150 694.800 ;
        RECT 95.100 687.750 96.900 696.000 ;
        RECT 100.500 687.750 102.300 696.600 ;
        RECT 116.400 696.000 120.900 697.650 ;
        RECT 133.950 697.050 136.050 699.150 ;
        RECT 136.950 698.850 139.050 700.950 ;
        RECT 149.100 699.150 150.900 700.950 ;
        RECT 119.100 687.750 120.900 696.000 ;
        RECT 124.500 687.750 126.300 696.600 ;
        RECT 137.400 690.600 138.600 698.850 ;
        RECT 148.950 697.050 151.050 699.150 ;
        RECT 151.950 698.850 154.050 700.950 ;
        RECT 166.950 698.850 169.050 700.950 ;
        RECT 170.100 699.150 171.900 700.950 ;
        RECT 184.950 700.050 187.050 702.150 ;
        RECT 152.400 690.600 153.600 698.850 ;
        RECT 167.400 690.600 168.600 698.850 ;
        RECT 169.950 697.050 172.050 699.150 ;
        RECT 184.950 696.750 186.150 700.050 ;
        RECT 187.950 698.850 190.050 700.950 ;
        RECT 190.950 700.050 193.050 702.150 ;
        RECT 199.950 700.050 202.050 702.150 ;
        RECT 202.950 698.850 205.050 700.950 ;
        RECT 205.950 700.050 208.050 702.150 ;
        RECT 224.400 700.950 225.600 713.400 ;
        RECT 239.700 713.100 241.350 713.400 ;
        RECT 245.550 713.400 247.350 719.250 ;
        RECT 260.400 713.400 262.200 719.250 ;
        RECT 245.550 713.100 246.750 713.400 ;
        RECT 239.700 712.200 246.750 713.100 ;
        RECT 239.100 708.150 240.900 709.950 ;
        RECT 236.100 705.150 237.900 706.950 ;
        RECT 238.950 706.050 241.050 708.150 ;
        RECT 242.250 705.150 244.050 706.950 ;
        RECT 235.950 703.050 238.050 705.150 ;
        RECT 241.950 703.050 244.050 705.150 ;
        RECT 245.700 703.950 246.750 712.200 ;
        RECT 263.700 707.400 265.500 719.250 ;
        RECT 267.900 707.400 269.700 719.250 ;
        RECT 280.650 713.400 282.450 719.250 ;
        RECT 283.650 713.400 285.450 719.250 ;
        RECT 286.650 713.400 288.450 719.250 ;
        RECT 260.250 705.150 262.050 706.950 ;
        RECT 244.950 701.850 247.050 703.950 ;
        RECT 259.950 703.050 262.050 705.150 ;
        RECT 263.850 702.150 265.050 707.400 ;
        RECT 284.250 705.150 285.450 713.400 ;
        RECT 297.300 707.400 299.100 719.250 ;
        RECT 301.500 707.400 303.300 719.250 ;
        RECT 304.800 713.400 306.600 719.250 ;
        RECT 319.650 713.400 321.450 719.250 ;
        RECT 322.650 714.000 324.450 719.250 ;
        RECT 320.250 713.100 321.450 713.400 ;
        RECT 325.650 713.400 327.450 719.250 ;
        RECT 328.650 713.400 330.450 719.250 ;
        RECT 325.650 713.100 327.300 713.400 ;
        RECT 320.250 712.200 327.300 713.100 ;
        RECT 269.100 702.150 270.900 703.950 ;
        RECT 188.100 697.050 189.900 698.850 ;
        RECT 203.100 697.050 204.900 698.850 ;
        RECT 206.850 696.750 208.050 700.050 ;
        RECT 221.100 699.150 222.900 700.950 ;
        RECT 220.950 697.050 223.050 699.150 ;
        RECT 223.950 698.850 226.050 700.950 ;
        RECT 182.250 695.700 186.000 696.750 ;
        RECT 207.000 695.700 210.750 696.750 ;
        RECT 182.250 693.600 183.450 695.700 ;
        RECT 134.550 687.750 136.350 690.600 ;
        RECT 137.550 687.750 139.350 690.600 ;
        RECT 149.550 687.750 151.350 690.600 ;
        RECT 152.550 687.750 154.350 690.600 ;
        RECT 166.650 687.750 168.450 690.600 ;
        RECT 169.650 687.750 171.450 690.600 ;
        RECT 181.650 687.750 183.450 693.600 ;
        RECT 184.650 692.700 192.450 694.050 ;
        RECT 184.650 687.750 186.450 692.700 ;
        RECT 187.650 687.750 189.450 691.800 ;
        RECT 190.650 687.750 192.450 692.700 ;
        RECT 200.550 692.700 208.350 694.050 ;
        RECT 200.550 687.750 202.350 692.700 ;
        RECT 203.550 687.750 205.350 691.800 ;
        RECT 206.550 687.750 208.350 692.700 ;
        RECT 209.550 693.600 210.750 695.700 ;
        RECT 209.550 687.750 211.350 693.600 ;
        RECT 224.400 690.600 225.600 698.850 ;
        RECT 245.400 697.650 246.600 701.850 ;
        RECT 221.550 687.750 223.350 690.600 ;
        RECT 224.550 687.750 226.350 690.600 ;
        RECT 236.700 687.750 238.500 696.600 ;
        RECT 242.100 696.000 246.600 697.650 ;
        RECT 262.950 700.050 265.050 702.150 ;
        RECT 262.950 696.750 264.150 700.050 ;
        RECT 265.950 698.850 268.050 700.950 ;
        RECT 268.950 700.050 271.050 702.150 ;
        RECT 280.950 701.850 283.050 703.950 ;
        RECT 283.950 703.050 286.050 705.150 ;
        RECT 281.100 700.050 282.900 701.850 ;
        RECT 266.100 697.050 267.900 698.850 ;
        RECT 242.100 687.750 243.900 696.000 ;
        RECT 260.250 695.700 264.000 696.750 ;
        RECT 284.250 695.700 285.450 703.050 ;
        RECT 286.950 701.850 289.050 703.950 ;
        RECT 296.100 702.150 297.900 703.950 ;
        RECT 301.950 702.150 303.150 707.400 ;
        RECT 304.950 705.150 306.750 706.950 ;
        RECT 304.950 703.050 307.050 705.150 ;
        RECT 320.250 703.950 321.300 712.200 ;
        RECT 326.100 708.150 327.900 709.950 ;
        RECT 322.950 705.150 324.750 706.950 ;
        RECT 325.950 706.050 328.050 708.150 ;
        RECT 340.350 707.400 342.150 719.250 ;
        RECT 343.350 707.400 345.150 719.250 ;
        RECT 346.650 713.400 348.450 719.250 ;
        RECT 356.550 713.400 358.350 719.250 ;
        RECT 359.550 713.400 361.350 719.250 ;
        RECT 362.550 713.400 364.350 719.250 ;
        RECT 374.550 713.400 376.350 719.250 ;
        RECT 377.550 713.400 379.350 719.250 ;
        RECT 380.550 713.400 382.350 719.250 ;
        RECT 329.100 705.150 330.900 706.950 ;
        RECT 287.100 700.050 288.900 701.850 ;
        RECT 295.950 700.050 298.050 702.150 ;
        RECT 298.950 698.850 301.050 700.950 ;
        RECT 301.950 700.050 304.050 702.150 ;
        RECT 319.950 701.850 322.050 703.950 ;
        RECT 322.950 703.050 325.050 705.150 ;
        RECT 328.950 703.050 331.050 705.150 ;
        RECT 340.650 702.150 341.850 707.400 ;
        RECT 347.250 706.500 348.450 713.400 ;
        RECT 342.750 705.600 348.450 706.500 ;
        RECT 342.750 704.700 345.000 705.600 ;
        RECT 359.550 705.150 360.750 713.400 ;
        RECT 377.550 705.150 378.750 713.400 ;
        RECT 394.350 707.400 396.150 719.250 ;
        RECT 397.350 707.400 399.150 719.250 ;
        RECT 400.650 713.400 402.450 719.250 ;
        RECT 410.550 713.400 412.350 719.250 ;
        RECT 413.550 713.400 415.350 719.250 ;
        RECT 416.550 714.000 418.350 719.250 ;
        RECT 299.100 697.050 300.900 698.850 ;
        RECT 302.850 696.750 304.050 700.050 ;
        RECT 320.400 697.650 321.600 701.850 ;
        RECT 340.650 700.050 343.050 702.150 ;
        RECT 303.000 695.700 306.750 696.750 ;
        RECT 320.400 696.000 324.900 697.650 ;
        RECT 260.250 693.600 261.450 695.700 ;
        RECT 281.850 694.800 285.450 695.700 ;
        RECT 259.650 687.750 261.450 693.600 ;
        RECT 262.650 692.700 270.450 694.050 ;
        RECT 262.650 687.750 264.450 692.700 ;
        RECT 265.650 687.750 267.450 691.800 ;
        RECT 268.650 687.750 270.450 692.700 ;
        RECT 281.850 687.750 283.650 694.800 ;
        RECT 286.350 687.750 288.150 693.600 ;
        RECT 296.550 692.700 304.350 694.050 ;
        RECT 296.550 687.750 298.350 692.700 ;
        RECT 299.550 687.750 301.350 691.800 ;
        RECT 302.550 687.750 304.350 692.700 ;
        RECT 305.550 693.600 306.750 695.700 ;
        RECT 305.550 687.750 307.350 693.600 ;
        RECT 323.100 687.750 324.900 696.000 ;
        RECT 328.500 687.750 330.300 696.600 ;
        RECT 340.650 693.600 341.850 700.050 ;
        RECT 343.950 696.300 345.000 704.700 ;
        RECT 347.100 702.150 348.900 703.950 ;
        RECT 346.950 700.050 349.050 702.150 ;
        RECT 355.950 701.850 358.050 703.950 ;
        RECT 358.950 703.050 361.050 705.150 ;
        RECT 356.100 700.050 357.900 701.850 ;
        RECT 342.750 695.400 345.000 696.300 ;
        RECT 359.550 695.700 360.750 703.050 ;
        RECT 361.950 701.850 364.050 703.950 ;
        RECT 373.950 701.850 376.050 703.950 ;
        RECT 376.950 703.050 379.050 705.150 ;
        RECT 362.100 700.050 363.900 701.850 ;
        RECT 374.100 700.050 375.900 701.850 ;
        RECT 377.550 695.700 378.750 703.050 ;
        RECT 379.950 701.850 382.050 703.950 ;
        RECT 394.650 702.150 395.850 707.400 ;
        RECT 401.250 706.500 402.450 713.400 ;
        RECT 413.700 713.100 415.350 713.400 ;
        RECT 419.550 713.400 421.350 719.250 ;
        RECT 419.550 713.100 420.750 713.400 ;
        RECT 413.700 712.200 420.750 713.100 ;
        RECT 413.100 708.150 414.900 709.950 ;
        RECT 396.750 705.600 402.450 706.500 ;
        RECT 396.750 704.700 399.000 705.600 ;
        RECT 410.100 705.150 411.900 706.950 ;
        RECT 412.950 706.050 415.050 708.150 ;
        RECT 416.250 705.150 418.050 706.950 ;
        RECT 380.100 700.050 381.900 701.850 ;
        RECT 394.650 700.050 397.050 702.150 ;
        RECT 342.750 694.500 347.850 695.400 ;
        RECT 359.550 694.800 363.150 695.700 ;
        RECT 377.550 694.800 381.150 695.700 ;
        RECT 340.350 687.750 342.150 693.600 ;
        RECT 343.350 687.750 345.150 693.600 ;
        RECT 346.650 690.600 347.850 694.500 ;
        RECT 346.650 687.750 348.450 690.600 ;
        RECT 356.850 687.750 358.650 693.600 ;
        RECT 361.350 687.750 363.150 694.800 ;
        RECT 374.850 687.750 376.650 693.600 ;
        RECT 379.350 687.750 381.150 694.800 ;
        RECT 394.650 693.600 395.850 700.050 ;
        RECT 397.950 696.300 399.000 704.700 ;
        RECT 401.100 702.150 402.900 703.950 ;
        RECT 409.950 703.050 412.050 705.150 ;
        RECT 415.950 703.050 418.050 705.150 ;
        RECT 419.700 703.950 420.750 712.200 ;
        RECT 435.450 707.400 437.250 719.250 ;
        RECT 439.650 707.400 441.450 719.250 ;
        RECT 452.550 707.400 454.350 719.250 ;
        RECT 457.050 707.400 460.350 719.250 ;
        RECT 463.050 707.400 464.850 719.250 ;
        RECT 478.650 713.400 480.450 719.250 ;
        RECT 481.650 713.400 483.450 719.250 ;
        RECT 484.650 713.400 486.450 719.250 ;
        RECT 496.650 713.400 498.450 719.250 ;
        RECT 499.650 714.000 501.450 719.250 ;
        RECT 435.450 706.350 438.000 707.400 ;
        RECT 400.950 700.050 403.050 702.150 ;
        RECT 418.950 701.850 421.050 703.950 ;
        RECT 434.100 702.150 435.900 703.950 ;
        RECT 419.400 697.650 420.600 701.850 ;
        RECT 433.950 700.050 436.050 702.150 ;
        RECT 396.750 695.400 399.000 696.300 ;
        RECT 396.750 694.500 401.850 695.400 ;
        RECT 394.350 687.750 396.150 693.600 ;
        RECT 397.350 687.750 399.150 693.600 ;
        RECT 400.650 690.600 401.850 694.500 ;
        RECT 400.650 687.750 402.450 690.600 ;
        RECT 410.700 687.750 412.500 696.600 ;
        RECT 416.100 696.000 420.600 697.650 ;
        RECT 436.950 699.150 438.000 706.350 ;
        RECT 440.100 702.150 441.900 703.950 ;
        RECT 452.100 702.150 453.900 703.950 ;
        RECT 458.550 702.150 459.750 707.400 ;
        RECT 482.250 705.150 483.450 713.400 ;
        RECT 497.250 713.100 498.450 713.400 ;
        RECT 502.650 713.400 504.450 719.250 ;
        RECT 505.650 713.400 507.450 719.250 ;
        RECT 502.650 713.100 504.300 713.400 ;
        RECT 497.250 712.200 504.300 713.100 ;
        RECT 463.950 702.150 465.750 703.950 ;
        RECT 439.950 700.050 442.050 702.150 ;
        RECT 451.950 700.050 454.050 702.150 ;
        RECT 436.950 697.050 439.050 699.150 ;
        RECT 454.950 698.850 457.050 700.950 ;
        RECT 457.950 700.050 460.050 702.150 ;
        RECT 455.100 697.050 456.900 698.850 ;
        RECT 416.100 687.750 417.900 696.000 ;
        RECT 436.950 690.600 438.000 697.050 ;
        RECT 458.400 696.150 459.600 700.050 ;
        RECT 460.950 698.850 463.050 700.950 ;
        RECT 463.950 700.050 466.050 702.150 ;
        RECT 478.950 701.850 481.050 703.950 ;
        RECT 481.950 703.050 484.050 705.150 ;
        RECT 497.250 703.950 498.300 712.200 ;
        RECT 503.100 708.150 504.900 709.950 ;
        RECT 499.950 705.150 501.750 706.950 ;
        RECT 502.950 706.050 505.050 708.150 ;
        RECT 517.650 707.400 519.450 719.250 ;
        RECT 520.650 708.300 522.450 719.250 ;
        RECT 523.650 709.200 525.450 719.250 ;
        RECT 526.650 708.300 528.450 719.250 ;
        RECT 538.650 713.400 540.450 719.250 ;
        RECT 541.650 714.000 543.450 719.250 ;
        RECT 520.650 707.400 528.450 708.300 ;
        RECT 539.250 713.100 540.450 713.400 ;
        RECT 544.650 713.400 546.450 719.250 ;
        RECT 547.650 713.400 549.450 719.250 ;
        RECT 544.650 713.100 546.300 713.400 ;
        RECT 539.250 712.200 546.300 713.100 ;
        RECT 506.100 705.150 507.900 706.950 ;
        RECT 479.100 700.050 480.900 701.850 ;
        RECT 460.500 697.050 462.300 698.850 ;
        RECT 458.400 695.100 462.750 696.150 ;
        RECT 482.250 695.700 483.450 703.050 ;
        RECT 484.950 701.850 487.050 703.950 ;
        RECT 496.950 701.850 499.050 703.950 ;
        RECT 499.950 703.050 502.050 705.150 ;
        RECT 505.950 703.050 508.050 705.150 ;
        RECT 518.100 702.150 519.300 707.400 ;
        RECT 539.250 703.950 540.300 712.200 ;
        RECT 545.100 708.150 546.900 709.950 ;
        RECT 541.950 705.150 543.750 706.950 ;
        RECT 544.950 706.050 547.050 708.150 ;
        RECT 559.650 707.400 561.450 719.250 ;
        RECT 562.650 708.300 564.450 719.250 ;
        RECT 565.650 709.200 567.450 719.250 ;
        RECT 568.650 708.300 570.450 719.250 ;
        RECT 578.550 713.400 580.350 719.250 ;
        RECT 581.550 713.400 583.350 719.250 ;
        RECT 584.550 714.000 586.350 719.250 ;
        RECT 581.700 713.100 583.350 713.400 ;
        RECT 587.550 713.400 589.350 719.250 ;
        RECT 599.550 713.400 601.350 719.250 ;
        RECT 602.550 713.400 604.350 719.250 ;
        RECT 605.550 714.000 607.350 719.250 ;
        RECT 587.550 713.100 588.750 713.400 ;
        RECT 581.700 712.200 588.750 713.100 ;
        RECT 602.700 713.100 604.350 713.400 ;
        RECT 608.550 713.400 610.350 719.250 ;
        RECT 620.550 713.400 622.350 719.250 ;
        RECT 623.550 713.400 625.350 719.250 ;
        RECT 608.550 713.100 609.750 713.400 ;
        RECT 602.700 712.200 609.750 713.100 ;
        RECT 562.650 707.400 570.450 708.300 ;
        RECT 581.100 708.150 582.900 709.950 ;
        RECT 548.100 705.150 549.900 706.950 ;
        RECT 485.100 700.050 486.900 701.850 ;
        RECT 497.400 697.650 498.600 701.850 ;
        RECT 517.950 700.050 520.050 702.150 ;
        RECT 538.950 701.850 541.050 703.950 ;
        RECT 541.950 703.050 544.050 705.150 ;
        RECT 547.950 703.050 550.050 705.150 ;
        RECT 560.100 702.150 561.300 707.400 ;
        RECT 568.950 705.450 571.050 706.050 ;
        RECT 568.950 704.550 573.450 705.450 ;
        RECT 578.100 705.150 579.900 706.950 ;
        RECT 580.950 706.050 583.050 708.150 ;
        RECT 584.250 705.150 586.050 706.950 ;
        RECT 568.950 703.950 571.050 704.550 ;
        RECT 497.400 696.000 501.900 697.650 ;
        RECT 452.550 693.000 460.350 693.900 ;
        RECT 461.850 693.600 462.750 695.100 ;
        RECT 479.850 694.800 483.450 695.700 ;
        RECT 433.650 687.750 435.450 690.600 ;
        RECT 436.650 687.750 438.450 690.600 ;
        RECT 439.650 687.750 441.450 690.600 ;
        RECT 452.550 687.750 454.350 693.000 ;
        RECT 455.550 687.750 457.350 692.100 ;
        RECT 458.550 688.500 460.350 693.000 ;
        RECT 461.550 689.400 463.350 693.600 ;
        RECT 464.550 688.500 466.350 693.600 ;
        RECT 458.550 687.750 466.350 688.500 ;
        RECT 479.850 687.750 481.650 694.800 ;
        RECT 484.350 687.750 486.150 693.600 ;
        RECT 500.100 687.750 501.900 696.000 ;
        RECT 505.500 687.750 507.300 696.600 ;
        RECT 518.100 693.600 519.300 700.050 ;
        RECT 520.950 698.850 523.050 700.950 ;
        RECT 524.100 699.150 525.900 700.950 ;
        RECT 521.100 697.050 522.900 698.850 ;
        RECT 523.950 697.050 526.050 699.150 ;
        RECT 526.950 698.850 529.050 700.950 ;
        RECT 527.100 697.050 528.900 698.850 ;
        RECT 539.400 697.650 540.600 701.850 ;
        RECT 559.950 700.050 562.050 702.150 ;
        RECT 539.400 696.000 543.900 697.650 ;
        RECT 518.100 691.950 523.800 693.600 ;
        RECT 518.700 687.750 520.500 690.600 ;
        RECT 522.000 687.750 523.800 691.950 ;
        RECT 526.200 687.750 528.000 693.600 ;
        RECT 542.100 687.750 543.900 696.000 ;
        RECT 547.500 687.750 549.300 696.600 ;
        RECT 560.100 693.600 561.300 700.050 ;
        RECT 562.950 698.850 565.050 700.950 ;
        RECT 566.100 699.150 567.900 700.950 ;
        RECT 563.100 697.050 564.900 698.850 ;
        RECT 565.950 697.050 568.050 699.150 ;
        RECT 568.950 698.850 571.050 700.950 ;
        RECT 572.550 699.450 573.450 704.550 ;
        RECT 577.950 703.050 580.050 705.150 ;
        RECT 583.950 703.050 586.050 705.150 ;
        RECT 587.700 703.950 588.750 712.200 ;
        RECT 602.100 708.150 603.900 709.950 ;
        RECT 599.100 705.150 600.900 706.950 ;
        RECT 601.950 706.050 604.050 708.150 ;
        RECT 605.250 705.150 607.050 706.950 ;
        RECT 586.950 701.850 589.050 703.950 ;
        RECT 598.950 703.050 601.050 705.150 ;
        RECT 604.950 703.050 607.050 705.150 ;
        RECT 608.700 703.950 609.750 712.200 ;
        RECT 607.950 701.850 610.050 703.950 ;
        RECT 577.950 699.450 580.050 700.050 ;
        RECT 569.100 697.050 570.900 698.850 ;
        RECT 572.550 698.550 580.050 699.450 ;
        RECT 577.950 697.950 580.050 698.550 ;
        RECT 587.400 697.650 588.600 701.850 ;
        RECT 608.400 697.650 609.600 701.850 ;
        RECT 623.400 700.950 624.600 713.400 ;
        RECT 637.050 707.400 638.850 719.250 ;
        RECT 640.050 707.400 641.850 719.250 ;
        RECT 643.650 713.400 645.450 719.250 ;
        RECT 646.650 713.400 648.450 719.250 ;
        RECT 661.650 713.400 663.450 719.250 ;
        RECT 664.650 714.000 666.450 719.250 ;
        RECT 637.650 702.150 638.850 707.400 ;
        RECT 620.100 699.150 621.900 700.950 ;
        RECT 560.100 691.950 565.800 693.600 ;
        RECT 560.700 687.750 562.500 690.600 ;
        RECT 564.000 687.750 565.800 691.950 ;
        RECT 568.200 687.750 570.000 693.600 ;
        RECT 578.700 687.750 580.500 696.600 ;
        RECT 584.100 696.000 588.600 697.650 ;
        RECT 584.100 687.750 585.900 696.000 ;
        RECT 599.700 687.750 601.500 696.600 ;
        RECT 605.100 696.000 609.600 697.650 ;
        RECT 619.950 697.050 622.050 699.150 ;
        RECT 622.950 698.850 625.050 700.950 ;
        RECT 637.650 700.050 640.050 702.150 ;
        RECT 640.950 701.850 643.050 703.950 ;
        RECT 641.100 700.050 642.900 701.850 ;
        RECT 605.100 687.750 606.900 696.000 ;
        RECT 623.400 690.600 624.600 698.850 ;
        RECT 637.650 693.600 638.850 700.050 ;
        RECT 644.100 696.300 645.300 713.400 ;
        RECT 662.250 713.100 663.450 713.400 ;
        RECT 667.650 713.400 669.450 719.250 ;
        RECT 670.650 713.400 672.450 719.250 ;
        RECT 680.550 713.400 682.350 719.250 ;
        RECT 683.550 713.400 685.350 719.250 ;
        RECT 686.550 714.000 688.350 719.250 ;
        RECT 667.650 713.100 669.300 713.400 ;
        RECT 662.250 712.200 669.300 713.100 ;
        RECT 683.700 713.100 685.350 713.400 ;
        RECT 689.550 713.400 691.350 719.250 ;
        RECT 701.550 713.400 703.350 719.250 ;
        RECT 704.550 713.400 706.350 719.250 ;
        RECT 689.550 713.100 690.750 713.400 ;
        RECT 683.700 712.200 690.750 713.100 ;
        RECT 662.250 703.950 663.300 712.200 ;
        RECT 668.100 708.150 669.900 709.950 ;
        RECT 683.100 708.150 684.900 709.950 ;
        RECT 664.950 705.150 666.750 706.950 ;
        RECT 667.950 706.050 670.050 708.150 ;
        RECT 671.100 705.150 672.900 706.950 ;
        RECT 680.100 705.150 681.900 706.950 ;
        RECT 682.950 706.050 685.050 708.150 ;
        RECT 686.250 705.150 688.050 706.950 ;
        RECT 647.100 702.150 648.900 703.950 ;
        RECT 646.950 700.050 649.050 702.150 ;
        RECT 661.950 701.850 664.050 703.950 ;
        RECT 664.950 703.050 667.050 705.150 ;
        RECT 670.950 703.050 673.050 705.150 ;
        RECT 679.950 703.050 682.050 705.150 ;
        RECT 685.950 703.050 688.050 705.150 ;
        RECT 689.700 703.950 690.750 712.200 ;
        RECT 688.950 701.850 691.050 703.950 ;
        RECT 662.400 697.650 663.600 701.850 ;
        RECT 689.400 697.650 690.600 701.850 ;
        RECT 704.400 700.950 705.600 713.400 ;
        RECT 710.550 707.400 712.350 719.250 ;
        RECT 713.550 716.400 715.350 719.250 ;
        RECT 718.050 713.400 719.850 719.250 ;
        RECT 722.250 713.400 724.050 719.250 ;
        RECT 715.950 711.300 719.850 713.400 ;
        RECT 726.150 712.500 727.950 719.250 ;
        RECT 729.150 713.400 730.950 719.250 ;
        RECT 733.950 713.400 735.750 719.250 ;
        RECT 739.050 713.400 740.850 719.250 ;
        RECT 734.250 712.500 735.450 713.400 ;
        RECT 724.950 710.700 731.850 712.500 ;
        RECT 734.250 710.400 739.050 712.500 ;
        RECT 717.150 708.600 719.850 710.400 ;
        RECT 720.750 709.800 722.550 710.400 ;
        RECT 720.750 708.900 727.050 709.800 ;
        RECT 734.250 709.500 735.450 710.400 ;
        RECT 720.750 708.600 722.550 708.900 ;
        RECT 718.950 707.700 719.850 708.600 ;
        RECT 701.100 699.150 702.900 700.950 ;
        RECT 640.950 695.100 648.450 696.300 ;
        RECT 662.400 696.000 666.900 697.650 ;
        RECT 640.950 694.500 642.750 695.100 ;
        RECT 637.650 692.100 640.950 693.600 ;
        RECT 620.550 687.750 622.350 690.600 ;
        RECT 623.550 687.750 625.350 690.600 ;
        RECT 639.150 687.750 640.950 692.100 ;
        RECT 642.150 687.750 643.950 693.600 ;
        RECT 646.650 687.750 648.450 695.100 ;
        RECT 665.100 687.750 666.900 696.000 ;
        RECT 670.500 687.750 672.300 696.600 ;
        RECT 680.700 687.750 682.500 696.600 ;
        RECT 686.100 696.000 690.600 697.650 ;
        RECT 700.950 697.050 703.050 699.150 ;
        RECT 703.950 698.850 706.050 700.950 ;
        RECT 686.100 687.750 687.900 696.000 ;
        RECT 704.400 690.600 705.600 698.850 ;
        RECT 710.550 697.950 711.750 707.400 ;
        RECT 715.950 706.800 718.050 707.700 ;
        RECT 718.950 706.800 724.950 707.700 ;
        RECT 713.850 705.600 718.050 706.800 ;
        RECT 712.950 703.800 714.750 705.600 ;
        RECT 724.050 702.150 724.950 706.800 ;
        RECT 726.150 706.800 727.050 708.900 ;
        RECT 727.950 708.300 735.450 709.500 ;
        RECT 727.950 707.700 729.750 708.300 ;
        RECT 742.050 707.400 743.850 719.250 ;
        RECT 753.300 707.400 755.100 719.250 ;
        RECT 757.500 707.400 759.300 719.250 ;
        RECT 760.800 713.400 762.600 719.250 ;
        RECT 773.550 713.400 775.350 719.250 ;
        RECT 776.550 713.400 778.350 719.250 ;
        RECT 779.550 713.400 781.350 719.250 ;
        RECT 791.550 713.400 793.350 719.250 ;
        RECT 794.550 713.400 796.350 719.250 ;
        RECT 797.550 713.400 799.350 719.250 ;
        RECT 812.550 713.400 814.350 719.250 ;
        RECT 815.550 713.400 817.350 719.250 ;
        RECT 818.550 713.400 820.350 719.250 ;
        RECT 830.550 713.400 832.350 719.250 ;
        RECT 833.550 713.400 835.350 719.250 ;
        RECT 836.550 713.400 838.350 719.250 ;
        RECT 850.650 713.400 852.450 719.250 ;
        RECT 853.650 714.000 855.450 719.250 ;
        RECT 732.750 706.800 743.850 707.400 ;
        RECT 726.150 706.200 743.850 706.800 ;
        RECT 726.150 705.900 734.550 706.200 ;
        RECT 732.750 705.600 734.550 705.900 ;
        RECT 724.050 700.050 727.050 702.150 ;
        RECT 730.950 701.100 733.050 702.150 ;
        RECT 730.950 700.050 738.900 701.100 ;
        RECT 712.950 699.750 715.050 700.050 ;
        RECT 712.950 697.950 716.850 699.750 ;
        RECT 710.550 695.850 715.050 697.950 ;
        RECT 724.050 696.000 724.950 700.050 ;
        RECT 737.100 699.300 738.900 700.050 ;
        RECT 740.100 699.150 741.900 700.950 ;
        RECT 734.100 698.400 735.900 699.000 ;
        RECT 740.100 698.400 741.000 699.150 ;
        RECT 734.100 697.200 741.000 698.400 ;
        RECT 734.100 696.000 735.150 697.200 ;
        RECT 710.550 693.600 711.750 695.850 ;
        RECT 724.050 695.100 735.150 696.000 ;
        RECT 724.050 694.800 724.950 695.100 ;
        RECT 701.550 687.750 703.350 690.600 ;
        RECT 704.550 687.750 706.350 690.600 ;
        RECT 710.550 687.750 712.350 693.600 ;
        RECT 715.950 692.700 718.050 693.600 ;
        RECT 723.150 693.000 724.950 694.800 ;
        RECT 734.100 694.200 735.150 695.100 ;
        RECT 730.350 693.450 732.150 694.200 ;
        RECT 715.950 691.500 719.700 692.700 ;
        RECT 718.650 690.600 719.700 691.500 ;
        RECT 727.200 692.400 732.150 693.450 ;
        RECT 733.650 692.400 735.450 694.200 ;
        RECT 742.950 693.600 743.850 706.200 ;
        RECT 752.100 702.150 753.900 703.950 ;
        RECT 757.950 702.150 759.150 707.400 ;
        RECT 760.950 705.150 762.750 706.950 ;
        RECT 776.550 705.150 777.750 713.400 ;
        RECT 794.550 705.150 795.750 713.400 ;
        RECT 796.950 708.450 799.050 709.050 ;
        RECT 805.950 708.450 808.050 709.050 ;
        RECT 796.950 707.550 801.450 708.450 ;
        RECT 796.950 706.950 799.050 707.550 ;
        RECT 800.550 705.450 801.450 707.550 ;
        RECT 805.950 707.550 810.450 708.450 ;
        RECT 805.950 706.950 808.050 707.550 ;
        RECT 805.950 705.450 808.050 706.050 ;
        RECT 760.950 703.050 763.050 705.150 ;
        RECT 751.950 700.050 754.050 702.150 ;
        RECT 754.950 698.850 757.050 700.950 ;
        RECT 757.950 700.050 760.050 702.150 ;
        RECT 772.950 701.850 775.050 703.950 ;
        RECT 775.950 703.050 778.050 705.150 ;
        RECT 773.100 700.050 774.900 701.850 ;
        RECT 755.100 697.050 756.900 698.850 ;
        RECT 758.850 696.750 760.050 700.050 ;
        RECT 759.000 695.700 762.750 696.750 ;
        RECT 727.200 690.600 728.250 692.400 ;
        RECT 736.950 691.500 739.050 693.600 ;
        RECT 736.950 690.600 738.000 691.500 ;
        RECT 713.850 687.750 715.650 690.600 ;
        RECT 718.350 687.750 720.150 690.600 ;
        RECT 722.550 687.750 724.350 690.600 ;
        RECT 726.450 687.750 728.250 690.600 ;
        RECT 729.750 687.750 731.550 690.600 ;
        RECT 734.250 689.700 738.000 690.600 ;
        RECT 734.250 687.750 736.050 689.700 ;
        RECT 739.050 687.750 740.850 690.600 ;
        RECT 742.050 687.750 743.850 693.600 ;
        RECT 752.550 692.700 760.350 694.050 ;
        RECT 752.550 687.750 754.350 692.700 ;
        RECT 755.550 687.750 757.350 691.800 ;
        RECT 758.550 687.750 760.350 692.700 ;
        RECT 761.550 693.600 762.750 695.700 ;
        RECT 776.550 695.700 777.750 703.050 ;
        RECT 778.950 701.850 781.050 703.950 ;
        RECT 790.950 701.850 793.050 703.950 ;
        RECT 793.950 703.050 796.050 705.150 ;
        RECT 800.550 704.550 808.050 705.450 ;
        RECT 805.950 703.950 808.050 704.550 ;
        RECT 779.100 700.050 780.900 701.850 ;
        RECT 791.100 700.050 792.900 701.850 ;
        RECT 794.550 695.700 795.750 703.050 ;
        RECT 796.950 701.850 799.050 703.950 ;
        RECT 797.100 700.050 798.900 701.850 ;
        RECT 809.550 696.450 810.450 707.550 ;
        RECT 815.550 705.150 816.750 713.400 ;
        RECT 823.950 708.450 826.050 709.050 ;
        RECT 829.950 708.450 832.050 709.050 ;
        RECT 823.950 707.550 832.050 708.450 ;
        RECT 823.950 706.950 826.050 707.550 ;
        RECT 829.950 706.950 832.050 707.550 ;
        RECT 833.550 705.150 834.750 713.400 ;
        RECT 851.250 713.100 852.450 713.400 ;
        RECT 856.650 713.400 858.450 719.250 ;
        RECT 859.650 713.400 861.450 719.250 ;
        RECT 856.650 713.100 858.300 713.400 ;
        RECT 851.250 712.200 858.300 713.100 ;
        RECT 838.950 708.450 841.050 709.050 ;
        RECT 847.950 708.450 850.050 709.050 ;
        RECT 838.950 707.550 850.050 708.450 ;
        RECT 838.950 706.950 841.050 707.550 ;
        RECT 847.950 706.950 850.050 707.550 ;
        RECT 811.950 701.850 814.050 703.950 ;
        RECT 814.950 703.050 817.050 705.150 ;
        RECT 812.100 700.050 813.900 701.850 ;
        RECT 811.950 696.450 814.050 697.050 ;
        RECT 776.550 694.800 780.150 695.700 ;
        RECT 794.550 694.800 798.150 695.700 ;
        RECT 809.550 695.550 814.050 696.450 ;
        RECT 811.950 694.950 814.050 695.550 ;
        RECT 815.550 695.700 816.750 703.050 ;
        RECT 817.950 701.850 820.050 703.950 ;
        RECT 829.950 701.850 832.050 703.950 ;
        RECT 832.950 703.050 835.050 705.150 ;
        RECT 851.250 703.950 852.300 712.200 ;
        RECT 857.100 708.150 858.900 709.950 ;
        RECT 853.950 705.150 855.750 706.950 ;
        RECT 856.950 706.050 859.050 708.150 ;
        RECT 860.100 705.150 861.900 706.950 ;
        RECT 818.100 700.050 819.900 701.850 ;
        RECT 830.100 700.050 831.900 701.850 ;
        RECT 833.550 695.700 834.750 703.050 ;
        RECT 835.950 701.850 838.050 703.950 ;
        RECT 850.950 701.850 853.050 703.950 ;
        RECT 853.950 703.050 856.050 705.150 ;
        RECT 859.950 703.050 862.050 705.150 ;
        RECT 836.100 700.050 837.900 701.850 ;
        RECT 851.400 697.650 852.600 701.850 ;
        RECT 851.400 696.000 855.900 697.650 ;
        RECT 815.550 694.800 819.150 695.700 ;
        RECT 833.550 694.800 837.150 695.700 ;
        RECT 761.550 687.750 763.350 693.600 ;
        RECT 773.850 687.750 775.650 693.600 ;
        RECT 778.350 687.750 780.150 694.800 ;
        RECT 791.850 687.750 793.650 693.600 ;
        RECT 796.350 687.750 798.150 694.800 ;
        RECT 812.850 687.750 814.650 693.600 ;
        RECT 817.350 687.750 819.150 694.800 ;
        RECT 830.850 687.750 832.650 693.600 ;
        RECT 835.350 687.750 837.150 694.800 ;
        RECT 854.100 687.750 855.900 696.000 ;
        RECT 859.500 687.750 861.300 696.600 ;
        RECT 10.650 677.400 12.450 683.250 ;
        RECT 11.250 675.300 12.450 677.400 ;
        RECT 13.650 678.300 15.450 683.250 ;
        RECT 16.650 679.200 18.450 683.250 ;
        RECT 19.650 678.300 21.450 683.250 ;
        RECT 13.650 676.950 21.450 678.300 ;
        RECT 22.950 678.450 25.050 679.050 ;
        RECT 28.950 678.450 31.050 679.050 ;
        RECT 22.950 677.550 31.050 678.450 ;
        RECT 22.950 676.950 25.050 677.550 ;
        RECT 28.950 676.950 31.050 677.550 ;
        RECT 11.250 674.250 15.000 675.300 ;
        RECT 35.100 675.000 36.900 683.250 ;
        RECT 13.950 670.950 15.150 674.250 ;
        RECT 17.100 672.150 18.900 673.950 ;
        RECT 32.400 673.350 36.900 675.000 ;
        RECT 40.500 674.400 42.300 683.250 ;
        RECT 51.000 677.400 52.800 683.250 ;
        RECT 55.200 679.050 57.000 683.250 ;
        RECT 58.500 680.400 60.300 683.250 ;
        RECT 55.200 677.400 60.900 679.050 ;
        RECT 76.650 677.400 78.450 683.250 ;
        RECT 13.950 668.850 16.050 670.950 ;
        RECT 16.950 670.050 19.050 672.150 ;
        RECT 19.950 668.850 22.050 670.950 ;
        RECT 32.400 669.150 33.600 673.350 ;
        RECT 40.950 672.450 43.050 673.050 ;
        RECT 46.950 672.450 49.050 673.050 ;
        RECT 40.950 671.550 49.050 672.450 ;
        RECT 50.100 672.150 51.900 673.950 ;
        RECT 40.950 670.950 43.050 671.550 ;
        RECT 46.950 670.950 49.050 671.550 ;
        RECT 49.950 670.050 52.050 672.150 ;
        RECT 52.950 671.850 55.050 673.950 ;
        RECT 56.100 672.150 57.900 673.950 ;
        RECT 53.100 670.050 54.900 671.850 ;
        RECT 55.950 670.050 58.050 672.150 ;
        RECT 59.700 670.950 60.900 677.400 ;
        RECT 77.250 675.300 78.450 677.400 ;
        RECT 79.650 678.300 81.450 683.250 ;
        RECT 82.650 679.200 84.450 683.250 ;
        RECT 85.650 678.300 87.450 683.250 ;
        RECT 79.650 676.950 87.450 678.300 ;
        RECT 97.650 677.400 99.450 683.250 ;
        RECT 98.250 675.300 99.450 677.400 ;
        RECT 100.650 678.300 102.450 683.250 ;
        RECT 103.650 679.200 105.450 683.250 ;
        RECT 106.650 678.300 108.450 683.250 ;
        RECT 116.550 680.400 118.350 683.250 ;
        RECT 119.550 680.400 121.350 683.250 ;
        RECT 100.650 676.950 108.450 678.300 ;
        RECT 77.250 674.250 81.000 675.300 ;
        RECT 98.250 674.250 102.000 675.300 ;
        RECT 79.950 670.950 81.150 674.250 ;
        RECT 83.100 672.150 84.900 673.950 ;
        RECT 10.950 665.850 13.050 667.950 ;
        RECT 11.250 664.050 13.050 665.850 ;
        RECT 14.850 663.600 16.050 668.850 ;
        RECT 20.100 667.050 21.900 668.850 ;
        RECT 31.950 667.050 34.050 669.150 ;
        RECT 58.950 668.850 61.050 670.950 ;
        RECT 79.950 668.850 82.050 670.950 ;
        RECT 82.950 670.050 85.050 672.150 ;
        RECT 100.950 670.950 102.150 674.250 ;
        RECT 104.100 672.150 105.900 673.950 ;
        RECT 85.950 668.850 88.050 670.950 ;
        RECT 100.950 668.850 103.050 670.950 ;
        RECT 103.950 670.050 106.050 672.150 ;
        RECT 115.950 671.850 118.050 673.950 ;
        RECT 119.400 672.150 120.600 680.400 ;
        RECT 132.000 677.400 133.800 683.250 ;
        RECT 136.200 679.050 138.000 683.250 ;
        RECT 139.500 680.400 141.300 683.250 ;
        RECT 154.650 680.400 156.450 683.250 ;
        RECT 157.650 680.400 159.450 683.250 ;
        RECT 136.200 677.400 141.900 679.050 ;
        RECT 131.100 672.150 132.900 673.950 ;
        RECT 106.950 668.850 109.050 670.950 ;
        RECT 116.100 670.050 117.900 671.850 ;
        RECT 118.950 670.050 121.050 672.150 ;
        RECT 130.950 670.050 133.050 672.150 ;
        RECT 133.950 671.850 136.050 673.950 ;
        RECT 137.100 672.150 138.900 673.950 ;
        RECT 134.100 670.050 135.900 671.850 ;
        RECT 136.950 670.050 139.050 672.150 ;
        RECT 140.700 670.950 141.900 677.400 ;
        RECT 155.400 672.150 156.600 680.400 ;
        RECT 173.100 675.000 174.900 683.250 ;
        RECT 11.400 651.750 13.200 657.600 ;
        RECT 14.700 651.750 16.500 663.600 ;
        RECT 18.900 651.750 20.700 663.600 ;
        RECT 32.250 658.800 33.300 667.050 ;
        RECT 34.950 665.850 37.050 667.950 ;
        RECT 40.950 665.850 43.050 667.950 ;
        RECT 34.950 664.050 36.750 665.850 ;
        RECT 37.950 662.850 40.050 664.950 ;
        RECT 41.100 664.050 42.900 665.850 ;
        RECT 59.700 663.600 60.900 668.850 ;
        RECT 76.950 665.850 79.050 667.950 ;
        RECT 77.250 664.050 79.050 665.850 ;
        RECT 80.850 663.600 82.050 668.850 ;
        RECT 86.100 667.050 87.900 668.850 ;
        RECT 97.950 665.850 100.050 667.950 ;
        RECT 98.250 664.050 100.050 665.850 ;
        RECT 101.850 663.600 103.050 668.850 ;
        RECT 107.100 667.050 108.900 668.850 ;
        RECT 38.100 661.050 39.900 662.850 ;
        RECT 50.550 662.700 58.350 663.600 ;
        RECT 32.250 657.900 39.300 658.800 ;
        RECT 32.250 657.600 33.450 657.900 ;
        RECT 31.650 651.750 33.450 657.600 ;
        RECT 37.650 657.600 39.300 657.900 ;
        RECT 34.650 651.750 36.450 657.000 ;
        RECT 37.650 651.750 39.450 657.600 ;
        RECT 40.650 651.750 42.450 657.600 ;
        RECT 50.550 651.750 52.350 662.700 ;
        RECT 53.550 651.750 55.350 661.800 ;
        RECT 56.550 651.750 58.350 662.700 ;
        RECT 59.550 651.750 61.350 663.600 ;
        RECT 77.400 651.750 79.200 657.600 ;
        RECT 80.700 651.750 82.500 663.600 ;
        RECT 84.900 651.750 86.700 663.600 ;
        RECT 98.400 651.750 100.200 657.600 ;
        RECT 101.700 651.750 103.500 663.600 ;
        RECT 105.900 651.750 107.700 663.600 ;
        RECT 119.400 657.600 120.600 670.050 ;
        RECT 139.950 668.850 142.050 670.950 ;
        RECT 154.950 670.050 157.050 672.150 ;
        RECT 157.950 671.850 160.050 673.950 ;
        RECT 170.400 673.350 174.900 675.000 ;
        RECT 178.500 674.400 180.300 683.250 ;
        RECT 191.700 680.400 193.500 683.250 ;
        RECT 195.000 679.050 196.800 683.250 ;
        RECT 191.100 677.400 196.800 679.050 ;
        RECT 199.200 677.400 201.000 683.250 ;
        RECT 211.650 680.400 213.450 683.250 ;
        RECT 214.650 680.400 216.450 683.250 ;
        RECT 158.100 670.050 159.900 671.850 ;
        RECT 140.700 663.600 141.900 668.850 ;
        RECT 131.550 662.700 139.350 663.600 ;
        RECT 116.550 651.750 118.350 657.600 ;
        RECT 119.550 651.750 121.350 657.600 ;
        RECT 131.550 651.750 133.350 662.700 ;
        RECT 134.550 651.750 136.350 661.800 ;
        RECT 137.550 651.750 139.350 662.700 ;
        RECT 140.550 651.750 142.350 663.600 ;
        RECT 155.400 657.600 156.600 670.050 ;
        RECT 170.400 669.150 171.600 673.350 ;
        RECT 191.100 670.950 192.300 677.400 ;
        RECT 194.100 672.150 195.900 673.950 ;
        RECT 169.950 667.050 172.050 669.150 ;
        RECT 190.950 668.850 193.050 670.950 ;
        RECT 193.950 670.050 196.050 672.150 ;
        RECT 196.950 671.850 199.050 673.950 ;
        RECT 200.100 672.150 201.900 673.950 ;
        RECT 212.400 672.150 213.600 680.400 ;
        RECT 224.550 678.300 226.350 683.250 ;
        RECT 227.550 679.200 229.350 683.250 ;
        RECT 230.550 678.300 232.350 683.250 ;
        RECT 224.550 676.950 232.350 678.300 ;
        RECT 233.550 677.400 235.350 683.250 ;
        RECT 233.550 675.300 234.750 677.400 ;
        RECT 248.850 676.200 250.650 683.250 ;
        RECT 253.350 677.400 255.150 683.250 ;
        RECT 248.850 675.300 252.450 676.200 ;
        RECT 231.000 674.250 234.750 675.300 ;
        RECT 197.100 670.050 198.900 671.850 ;
        RECT 199.950 670.050 202.050 672.150 ;
        RECT 211.950 670.050 214.050 672.150 ;
        RECT 214.950 671.850 217.050 673.950 ;
        RECT 227.100 672.150 228.900 673.950 ;
        RECT 215.100 670.050 216.900 671.850 ;
        RECT 170.250 658.800 171.300 667.050 ;
        RECT 172.950 665.850 175.050 667.950 ;
        RECT 178.950 665.850 181.050 667.950 ;
        RECT 172.950 664.050 174.750 665.850 ;
        RECT 175.950 662.850 178.050 664.950 ;
        RECT 179.100 664.050 180.900 665.850 ;
        RECT 191.100 663.600 192.300 668.850 ;
        RECT 176.100 661.050 177.900 662.850 ;
        RECT 170.250 657.900 177.300 658.800 ;
        RECT 170.250 657.600 171.450 657.900 ;
        RECT 154.650 651.750 156.450 657.600 ;
        RECT 157.650 651.750 159.450 657.600 ;
        RECT 169.650 651.750 171.450 657.600 ;
        RECT 175.650 657.600 177.300 657.900 ;
        RECT 172.650 651.750 174.450 657.000 ;
        RECT 175.650 651.750 177.450 657.600 ;
        RECT 178.650 651.750 180.450 657.600 ;
        RECT 190.650 651.750 192.450 663.600 ;
        RECT 193.650 662.700 201.450 663.600 ;
        RECT 193.650 651.750 195.450 662.700 ;
        RECT 196.650 651.750 198.450 661.800 ;
        RECT 199.650 651.750 201.450 662.700 ;
        RECT 212.400 657.600 213.600 670.050 ;
        RECT 223.950 668.850 226.050 670.950 ;
        RECT 226.950 670.050 229.050 672.150 ;
        RECT 230.850 670.950 232.050 674.250 ;
        RECT 229.950 668.850 232.050 670.950 ;
        RECT 248.100 669.150 249.900 670.950 ;
        RECT 224.100 667.050 225.900 668.850 ;
        RECT 229.950 663.600 231.150 668.850 ;
        RECT 232.950 665.850 235.050 667.950 ;
        RECT 247.950 667.050 250.050 669.150 ;
        RECT 251.250 667.950 252.450 675.300 ;
        RECT 269.100 675.000 270.900 683.250 ;
        RECT 266.400 673.350 270.900 675.000 ;
        RECT 274.500 674.400 276.300 683.250 ;
        RECT 286.650 680.400 288.450 683.250 ;
        RECT 289.650 680.400 291.450 683.250 ;
        RECT 292.650 680.400 294.450 683.250 ;
        RECT 289.950 673.950 291.000 680.400 ;
        RECT 292.950 675.450 295.050 676.050 ;
        RECT 301.950 675.450 304.050 676.050 ;
        RECT 292.950 674.550 304.050 675.450 ;
        RECT 308.100 675.000 309.900 683.250 ;
        RECT 292.950 673.950 295.050 674.550 ;
        RECT 301.950 673.950 304.050 674.550 ;
        RECT 254.100 669.150 255.900 670.950 ;
        RECT 266.400 669.150 267.600 673.350 ;
        RECT 289.950 671.850 292.050 673.950 ;
        RECT 305.400 673.350 309.900 675.000 ;
        RECT 313.500 674.400 315.300 683.250 ;
        RECT 332.100 675.000 333.900 683.250 ;
        RECT 329.400 673.350 333.900 675.000 ;
        RECT 337.500 674.400 339.300 683.250 ;
        RECT 350.850 676.200 352.650 683.250 ;
        RECT 355.350 677.400 357.150 683.250 ;
        RECT 350.850 675.300 354.450 676.200 ;
        RECT 250.950 665.850 253.050 667.950 ;
        RECT 253.950 667.050 256.050 669.150 ;
        RECT 265.950 667.050 268.050 669.150 ;
        RECT 286.950 668.850 289.050 670.950 ;
        RECT 232.950 664.050 234.750 665.850 ;
        RECT 211.650 651.750 213.450 657.600 ;
        RECT 214.650 651.750 216.450 657.600 ;
        RECT 225.300 651.750 227.100 663.600 ;
        RECT 229.500 651.750 231.300 663.600 ;
        RECT 251.250 657.600 252.450 665.850 ;
        RECT 266.250 658.800 267.300 667.050 ;
        RECT 268.950 665.850 271.050 667.950 ;
        RECT 274.950 665.850 277.050 667.950 ;
        RECT 287.100 667.050 288.900 668.850 ;
        RECT 268.950 664.050 270.750 665.850 ;
        RECT 271.950 662.850 274.050 664.950 ;
        RECT 275.100 664.050 276.900 665.850 ;
        RECT 289.950 664.650 291.000 671.850 ;
        RECT 292.950 668.850 295.050 670.950 ;
        RECT 305.400 669.150 306.600 673.350 ;
        RECT 329.400 669.150 330.600 673.350 ;
        RECT 350.100 669.150 351.900 670.950 ;
        RECT 293.100 667.050 294.900 668.850 ;
        RECT 304.950 667.050 307.050 669.150 ;
        RECT 288.450 663.600 291.000 664.650 ;
        RECT 272.100 661.050 273.900 662.850 ;
        RECT 266.250 657.900 273.300 658.800 ;
        RECT 266.250 657.600 267.450 657.900 ;
        RECT 232.800 651.750 234.600 657.600 ;
        RECT 247.650 651.750 249.450 657.600 ;
        RECT 250.650 651.750 252.450 657.600 ;
        RECT 253.650 651.750 255.450 657.600 ;
        RECT 265.650 651.750 267.450 657.600 ;
        RECT 271.650 657.600 273.300 657.900 ;
        RECT 268.650 651.750 270.450 657.000 ;
        RECT 271.650 651.750 273.450 657.600 ;
        RECT 274.650 651.750 276.450 657.600 ;
        RECT 288.450 651.750 290.250 663.600 ;
        RECT 292.650 651.750 294.450 663.600 ;
        RECT 305.250 658.800 306.300 667.050 ;
        RECT 307.950 665.850 310.050 667.950 ;
        RECT 313.950 665.850 316.050 667.950 ;
        RECT 328.950 667.050 331.050 669.150 ;
        RECT 307.950 664.050 309.750 665.850 ;
        RECT 310.950 662.850 313.050 664.950 ;
        RECT 314.100 664.050 315.900 665.850 ;
        RECT 311.100 661.050 312.900 662.850 ;
        RECT 329.250 658.800 330.300 667.050 ;
        RECT 331.950 665.850 334.050 667.950 ;
        RECT 337.950 665.850 340.050 667.950 ;
        RECT 349.950 667.050 352.050 669.150 ;
        RECT 353.250 667.950 354.450 675.300 ;
        RECT 371.100 675.000 372.900 683.250 ;
        RECT 368.400 673.350 372.900 675.000 ;
        RECT 376.500 674.400 378.300 683.250 ;
        RECT 386.700 674.400 388.500 683.250 ;
        RECT 392.100 675.000 393.900 683.250 ;
        RECT 409.650 680.400 411.450 683.250 ;
        RECT 412.650 680.400 414.450 683.250 ;
        RECT 424.650 680.400 426.450 683.250 ;
        RECT 427.650 680.400 429.450 683.250 ;
        RECT 430.650 680.400 432.450 683.250 ;
        RECT 392.100 673.350 396.600 675.000 ;
        RECT 356.100 669.150 357.900 670.950 ;
        RECT 368.400 669.150 369.600 673.350 ;
        RECT 395.400 669.150 396.600 673.350 ;
        RECT 410.400 672.150 411.600 680.400 ;
        RECT 427.950 673.950 429.000 680.400 ;
        RECT 446.100 675.000 447.900 683.250 ;
        RECT 409.950 670.050 412.050 672.150 ;
        RECT 412.950 671.850 415.050 673.950 ;
        RECT 427.950 671.850 430.050 673.950 ;
        RECT 443.400 673.350 447.900 675.000 ;
        RECT 451.500 674.400 453.300 683.250 ;
        RECT 467.100 675.000 468.900 683.250 ;
        RECT 464.400 673.350 468.900 675.000 ;
        RECT 472.500 674.400 474.300 683.250 ;
        RECT 482.550 680.400 484.350 683.250 ;
        RECT 485.550 680.400 487.350 683.250 ;
        RECT 413.100 670.050 414.900 671.850 ;
        RECT 352.950 665.850 355.050 667.950 ;
        RECT 355.950 667.050 358.050 669.150 ;
        RECT 367.950 667.050 370.050 669.150 ;
        RECT 331.950 664.050 333.750 665.850 ;
        RECT 334.950 662.850 337.050 664.950 ;
        RECT 338.100 664.050 339.900 665.850 ;
        RECT 335.100 661.050 336.900 662.850 ;
        RECT 305.250 657.900 312.300 658.800 ;
        RECT 305.250 657.600 306.450 657.900 ;
        RECT 304.650 651.750 306.450 657.600 ;
        RECT 310.650 657.600 312.300 657.900 ;
        RECT 329.250 657.900 336.300 658.800 ;
        RECT 329.250 657.600 330.450 657.900 ;
        RECT 307.650 651.750 309.450 657.000 ;
        RECT 310.650 651.750 312.450 657.600 ;
        RECT 313.650 651.750 315.450 657.600 ;
        RECT 328.650 651.750 330.450 657.600 ;
        RECT 334.650 657.600 336.300 657.900 ;
        RECT 353.250 657.600 354.450 665.850 ;
        RECT 368.250 658.800 369.300 667.050 ;
        RECT 370.950 665.850 373.050 667.950 ;
        RECT 376.950 665.850 379.050 667.950 ;
        RECT 385.950 665.850 388.050 667.950 ;
        RECT 391.950 665.850 394.050 667.950 ;
        RECT 394.950 667.050 397.050 669.150 ;
        RECT 370.950 664.050 372.750 665.850 ;
        RECT 373.950 662.850 376.050 664.950 ;
        RECT 377.100 664.050 378.900 665.850 ;
        RECT 386.100 664.050 387.900 665.850 ;
        RECT 388.950 662.850 391.050 664.950 ;
        RECT 392.250 664.050 394.050 665.850 ;
        RECT 374.100 661.050 375.900 662.850 ;
        RECT 389.100 661.050 390.900 662.850 ;
        RECT 395.700 658.800 396.750 667.050 ;
        RECT 368.250 657.900 375.300 658.800 ;
        RECT 368.250 657.600 369.450 657.900 ;
        RECT 331.650 651.750 333.450 657.000 ;
        RECT 334.650 651.750 336.450 657.600 ;
        RECT 337.650 651.750 339.450 657.600 ;
        RECT 349.650 651.750 351.450 657.600 ;
        RECT 352.650 651.750 354.450 657.600 ;
        RECT 355.650 651.750 357.450 657.600 ;
        RECT 367.650 651.750 369.450 657.600 ;
        RECT 373.650 657.600 375.300 657.900 ;
        RECT 389.700 657.900 396.750 658.800 ;
        RECT 389.700 657.600 391.350 657.900 ;
        RECT 370.650 651.750 372.450 657.000 ;
        RECT 373.650 651.750 375.450 657.600 ;
        RECT 376.650 651.750 378.450 657.600 ;
        RECT 386.550 651.750 388.350 657.600 ;
        RECT 389.550 651.750 391.350 657.600 ;
        RECT 395.550 657.600 396.750 657.900 ;
        RECT 410.400 657.600 411.600 670.050 ;
        RECT 424.950 668.850 427.050 670.950 ;
        RECT 425.100 667.050 426.900 668.850 ;
        RECT 427.950 664.650 429.000 671.850 ;
        RECT 430.950 668.850 433.050 670.950 ;
        RECT 443.400 669.150 444.600 673.350 ;
        RECT 464.400 669.150 465.600 673.350 ;
        RECT 481.950 671.850 484.050 673.950 ;
        RECT 485.400 672.150 486.600 680.400 ;
        RECT 497.550 678.300 499.350 683.250 ;
        RECT 500.550 679.200 502.350 683.250 ;
        RECT 503.550 678.300 505.350 683.250 ;
        RECT 497.550 676.950 505.350 678.300 ;
        RECT 506.550 677.400 508.350 683.250 ;
        RECT 522.150 678.900 523.950 683.250 ;
        RECT 520.650 677.400 523.950 678.900 ;
        RECT 525.150 677.400 526.950 683.250 ;
        RECT 506.550 675.300 507.750 677.400 ;
        RECT 504.000 674.250 507.750 675.300 ;
        RECT 500.100 672.150 501.900 673.950 ;
        RECT 482.100 670.050 483.900 671.850 ;
        RECT 484.950 670.050 487.050 672.150 ;
        RECT 431.100 667.050 432.900 668.850 ;
        RECT 442.950 667.050 445.050 669.150 ;
        RECT 426.450 663.600 429.000 664.650 ;
        RECT 392.550 651.750 394.350 657.000 ;
        RECT 395.550 651.750 397.350 657.600 ;
        RECT 409.650 651.750 411.450 657.600 ;
        RECT 412.650 651.750 414.450 657.600 ;
        RECT 426.450 651.750 428.250 663.600 ;
        RECT 430.650 651.750 432.450 663.600 ;
        RECT 443.250 658.800 444.300 667.050 ;
        RECT 445.950 665.850 448.050 667.950 ;
        RECT 451.950 665.850 454.050 667.950 ;
        RECT 463.950 667.050 466.050 669.150 ;
        RECT 445.950 664.050 447.750 665.850 ;
        RECT 448.950 662.850 451.050 664.950 ;
        RECT 452.100 664.050 453.900 665.850 ;
        RECT 449.100 661.050 450.900 662.850 ;
        RECT 464.250 658.800 465.300 667.050 ;
        RECT 466.950 665.850 469.050 667.950 ;
        RECT 472.950 665.850 475.050 667.950 ;
        RECT 466.950 664.050 468.750 665.850 ;
        RECT 469.950 662.850 472.050 664.950 ;
        RECT 473.100 664.050 474.900 665.850 ;
        RECT 470.100 661.050 471.900 662.850 ;
        RECT 443.250 657.900 450.300 658.800 ;
        RECT 443.250 657.600 444.450 657.900 ;
        RECT 442.650 651.750 444.450 657.600 ;
        RECT 448.650 657.600 450.300 657.900 ;
        RECT 464.250 657.900 471.300 658.800 ;
        RECT 464.250 657.600 465.450 657.900 ;
        RECT 445.650 651.750 447.450 657.000 ;
        RECT 448.650 651.750 450.450 657.600 ;
        RECT 451.650 651.750 453.450 657.600 ;
        RECT 463.650 651.750 465.450 657.600 ;
        RECT 469.650 657.600 471.300 657.900 ;
        RECT 485.400 657.600 486.600 670.050 ;
        RECT 496.950 668.850 499.050 670.950 ;
        RECT 499.950 670.050 502.050 672.150 ;
        RECT 503.850 670.950 505.050 674.250 ;
        RECT 502.950 668.850 505.050 670.950 ;
        RECT 520.650 670.950 521.850 677.400 ;
        RECT 523.950 675.900 525.750 676.500 ;
        RECT 529.650 675.900 531.450 683.250 ;
        RECT 542.850 677.400 544.650 683.250 ;
        RECT 547.350 676.200 549.150 683.250 ;
        RECT 562.650 677.400 564.450 683.250 ;
        RECT 565.650 680.400 567.450 683.250 ;
        RECT 568.650 680.400 570.450 683.250 ;
        RECT 571.650 680.400 573.450 683.250 ;
        RECT 523.950 674.700 531.450 675.900 ;
        RECT 545.550 675.300 549.150 676.200 ;
        RECT 520.650 668.850 523.050 670.950 ;
        RECT 524.100 669.150 525.900 670.950 ;
        RECT 497.100 667.050 498.900 668.850 ;
        RECT 502.950 663.600 504.150 668.850 ;
        RECT 505.950 665.850 508.050 667.950 ;
        RECT 505.950 664.050 507.750 665.850 ;
        RECT 520.650 663.600 521.850 668.850 ;
        RECT 523.950 667.050 526.050 669.150 ;
        RECT 466.650 651.750 468.450 657.000 ;
        RECT 469.650 651.750 471.450 657.600 ;
        RECT 472.650 651.750 474.450 657.600 ;
        RECT 482.550 651.750 484.350 657.600 ;
        RECT 485.550 651.750 487.350 657.600 ;
        RECT 498.300 651.750 500.100 663.600 ;
        RECT 502.500 651.750 504.300 663.600 ;
        RECT 505.800 651.750 507.600 657.600 ;
        RECT 520.050 651.750 521.850 663.600 ;
        RECT 523.050 651.750 524.850 663.600 ;
        RECT 527.100 657.600 528.300 674.700 ;
        RECT 529.950 668.850 532.050 670.950 ;
        RECT 542.100 669.150 543.900 670.950 ;
        RECT 530.100 667.050 531.900 668.850 ;
        RECT 541.950 667.050 544.050 669.150 ;
        RECT 545.550 667.950 546.750 675.300 ;
        RECT 562.950 672.150 564.000 677.400 ;
        RECT 568.650 676.200 569.550 680.400 ;
        RECT 581.850 677.400 583.650 683.250 ;
        RECT 586.350 676.200 588.150 683.250 ;
        RECT 601.350 677.400 603.150 683.250 ;
        RECT 604.350 677.400 606.150 683.250 ;
        RECT 607.650 680.400 609.450 683.250 ;
        RECT 566.250 675.300 569.550 676.200 ;
        RECT 584.550 675.300 588.150 676.200 ;
        RECT 566.250 674.400 568.050 675.300 ;
        RECT 548.100 669.150 549.900 670.950 ;
        RECT 562.950 670.050 565.050 672.150 ;
        RECT 544.950 665.850 547.050 667.950 ;
        RECT 547.950 667.050 550.050 669.150 ;
        RECT 545.550 657.600 546.750 665.850 ;
        RECT 563.550 663.450 564.900 670.050 ;
        RECT 566.400 666.150 567.300 674.400 ;
        RECT 571.950 671.850 574.050 673.950 ;
        RECT 568.950 668.850 571.050 670.950 ;
        RECT 572.100 670.050 573.900 671.850 ;
        RECT 581.100 669.150 582.900 670.950 ;
        RECT 569.100 667.050 570.900 668.850 ;
        RECT 580.950 667.050 583.050 669.150 ;
        RECT 584.550 667.950 585.750 675.300 ;
        RECT 601.650 670.950 602.850 677.400 ;
        RECT 607.650 676.500 608.850 680.400 ;
        RECT 603.750 675.600 608.850 676.500 ;
        RECT 617.550 675.900 619.350 683.250 ;
        RECT 622.050 677.400 623.850 683.250 ;
        RECT 625.050 678.900 626.850 683.250 ;
        RECT 625.050 677.400 628.350 678.900 ;
        RECT 623.250 675.900 625.050 676.500 ;
        RECT 603.750 674.700 606.000 675.600 ;
        RECT 617.550 674.700 625.050 675.900 ;
        RECT 587.100 669.150 588.900 670.950 ;
        RECT 566.250 666.000 568.050 666.150 ;
        RECT 566.250 664.800 573.450 666.000 ;
        RECT 583.950 665.850 586.050 667.950 ;
        RECT 586.950 667.050 589.050 669.150 ;
        RECT 601.650 668.850 604.050 670.950 ;
        RECT 566.250 664.350 568.050 664.800 ;
        RECT 572.250 663.600 573.450 664.800 ;
        RECT 563.550 662.100 565.950 663.450 ;
        RECT 526.650 651.750 528.450 657.600 ;
        RECT 529.650 651.750 531.450 657.600 ;
        RECT 542.550 651.750 544.350 657.600 ;
        RECT 545.550 651.750 547.350 657.600 ;
        RECT 548.550 651.750 550.350 657.600 ;
        RECT 564.150 651.750 565.950 662.100 ;
        RECT 567.150 651.750 568.950 663.450 ;
        RECT 571.650 651.750 573.450 663.600 ;
        RECT 584.550 657.600 585.750 665.850 ;
        RECT 601.650 663.600 602.850 668.850 ;
        RECT 604.950 666.300 606.000 674.700 ;
        RECT 607.950 668.850 610.050 670.950 ;
        RECT 616.950 668.850 619.050 670.950 ;
        RECT 608.100 667.050 609.900 668.850 ;
        RECT 617.100 667.050 618.900 668.850 ;
        RECT 603.750 665.400 606.000 666.300 ;
        RECT 603.750 664.500 609.450 665.400 ;
        RECT 581.550 651.750 583.350 657.600 ;
        RECT 584.550 651.750 586.350 657.600 ;
        RECT 587.550 651.750 589.350 657.600 ;
        RECT 601.350 651.750 603.150 663.600 ;
        RECT 604.350 651.750 606.150 663.600 ;
        RECT 608.250 657.600 609.450 664.500 ;
        RECT 620.700 657.600 621.900 674.700 ;
        RECT 627.150 670.950 628.350 677.400 ;
        RECT 641.850 676.200 643.650 683.250 ;
        RECT 646.350 677.400 648.150 683.250 ;
        RECT 658.650 677.400 660.450 683.250 ;
        RECT 641.850 675.300 645.450 676.200 ;
        RECT 623.100 669.150 624.900 670.950 ;
        RECT 622.950 667.050 625.050 669.150 ;
        RECT 625.950 668.850 628.350 670.950 ;
        RECT 641.100 669.150 642.900 670.950 ;
        RECT 627.150 663.600 628.350 668.850 ;
        RECT 640.950 667.050 643.050 669.150 ;
        RECT 644.250 667.950 645.450 675.300 ;
        RECT 659.250 675.300 660.450 677.400 ;
        RECT 661.650 678.300 663.450 683.250 ;
        RECT 664.650 679.200 666.450 683.250 ;
        RECT 667.650 678.300 669.450 683.250 ;
        RECT 661.650 676.950 669.450 678.300 ;
        RECT 677.850 677.400 679.650 683.250 ;
        RECT 682.350 676.200 684.150 683.250 ;
        RECT 680.550 675.300 684.150 676.200 ;
        RECT 698.850 676.200 700.650 683.250 ;
        RECT 703.350 677.400 705.150 683.250 ;
        RECT 713.550 680.400 715.350 683.250 ;
        RECT 716.550 680.400 718.350 683.250 ;
        RECT 698.850 675.300 702.450 676.200 ;
        RECT 659.250 674.250 663.000 675.300 ;
        RECT 661.950 670.950 663.150 674.250 ;
        RECT 665.100 672.150 666.900 673.950 ;
        RECT 647.100 669.150 648.900 670.950 ;
        RECT 643.950 665.850 646.050 667.950 ;
        RECT 646.950 667.050 649.050 669.150 ;
        RECT 661.950 668.850 664.050 670.950 ;
        RECT 664.950 670.050 667.050 672.150 ;
        RECT 667.950 668.850 670.050 670.950 ;
        RECT 677.100 669.150 678.900 670.950 ;
        RECT 658.950 665.850 661.050 667.950 ;
        RECT 607.650 651.750 609.450 657.600 ;
        RECT 617.550 651.750 619.350 657.600 ;
        RECT 620.550 651.750 622.350 657.600 ;
        RECT 624.150 651.750 625.950 663.600 ;
        RECT 627.150 651.750 628.950 663.600 ;
        RECT 644.250 657.600 645.450 665.850 ;
        RECT 659.250 664.050 661.050 665.850 ;
        RECT 662.850 663.600 664.050 668.850 ;
        RECT 668.100 667.050 669.900 668.850 ;
        RECT 676.950 667.050 679.050 669.150 ;
        RECT 680.550 667.950 681.750 675.300 ;
        RECT 683.100 669.150 684.900 670.950 ;
        RECT 698.100 669.150 699.900 670.950 ;
        RECT 679.950 665.850 682.050 667.950 ;
        RECT 682.950 667.050 685.050 669.150 ;
        RECT 697.950 667.050 700.050 669.150 ;
        RECT 701.250 667.950 702.450 675.300 ;
        RECT 712.950 671.850 715.050 673.950 ;
        RECT 716.400 672.150 717.600 680.400 ;
        RECT 728.850 677.400 730.650 683.250 ;
        RECT 733.350 676.200 735.150 683.250 ;
        RECT 746.550 678.300 748.350 683.250 ;
        RECT 749.550 679.200 751.350 683.250 ;
        RECT 752.550 678.300 754.350 683.250 ;
        RECT 746.550 676.950 754.350 678.300 ;
        RECT 755.550 677.400 757.350 683.250 ;
        RECT 761.550 677.400 763.350 683.250 ;
        RECT 764.850 680.400 766.650 683.250 ;
        RECT 769.350 680.400 771.150 683.250 ;
        RECT 773.550 680.400 775.350 683.250 ;
        RECT 777.450 680.400 779.250 683.250 ;
        RECT 780.750 680.400 782.550 683.250 ;
        RECT 785.250 681.300 787.050 683.250 ;
        RECT 785.250 680.400 789.000 681.300 ;
        RECT 790.050 680.400 791.850 683.250 ;
        RECT 769.650 679.500 770.700 680.400 ;
        RECT 766.950 678.300 770.700 679.500 ;
        RECT 778.200 678.600 779.250 680.400 ;
        RECT 787.950 679.500 789.000 680.400 ;
        RECT 766.950 677.400 769.050 678.300 ;
        RECT 731.550 675.300 735.150 676.200 ;
        RECT 755.550 675.300 756.750 677.400 ;
        RECT 704.100 669.150 705.900 670.950 ;
        RECT 713.100 670.050 714.900 671.850 ;
        RECT 715.950 670.050 718.050 672.150 ;
        RECT 700.950 665.850 703.050 667.950 ;
        RECT 703.950 667.050 706.050 669.150 ;
        RECT 640.650 651.750 642.450 657.600 ;
        RECT 643.650 651.750 645.450 657.600 ;
        RECT 646.650 651.750 648.450 657.600 ;
        RECT 659.400 651.750 661.200 657.600 ;
        RECT 662.700 651.750 664.500 663.600 ;
        RECT 666.900 651.750 668.700 663.600 ;
        RECT 680.550 657.600 681.750 665.850 ;
        RECT 701.250 657.600 702.450 665.850 ;
        RECT 716.400 657.600 717.600 670.050 ;
        RECT 728.100 669.150 729.900 670.950 ;
        RECT 727.950 667.050 730.050 669.150 ;
        RECT 731.550 667.950 732.750 675.300 ;
        RECT 753.000 674.250 756.750 675.300 ;
        RECT 761.550 675.150 762.750 677.400 ;
        RECT 774.150 676.200 775.950 678.000 ;
        RECT 778.200 677.550 783.150 678.600 ;
        RECT 781.350 676.800 783.150 677.550 ;
        RECT 784.650 676.800 786.450 678.600 ;
        RECT 787.950 677.400 790.050 679.500 ;
        RECT 793.050 677.400 794.850 683.250 ;
        RECT 775.050 675.900 775.950 676.200 ;
        RECT 785.100 675.900 786.150 676.800 ;
        RECT 749.100 672.150 750.900 673.950 ;
        RECT 734.100 669.150 735.900 670.950 ;
        RECT 730.950 665.850 733.050 667.950 ;
        RECT 733.950 667.050 736.050 669.150 ;
        RECT 745.950 668.850 748.050 670.950 ;
        RECT 748.950 670.050 751.050 672.150 ;
        RECT 752.850 670.950 754.050 674.250 ;
        RECT 751.950 668.850 754.050 670.950 ;
        RECT 761.550 673.050 766.050 675.150 ;
        RECT 775.050 675.000 786.150 675.900 ;
        RECT 746.100 667.050 747.900 668.850 ;
        RECT 731.550 657.600 732.750 665.850 ;
        RECT 751.950 663.600 753.150 668.850 ;
        RECT 754.950 665.850 757.050 667.950 ;
        RECT 754.950 664.050 756.750 665.850 ;
        RECT 761.550 663.600 762.750 673.050 ;
        RECT 763.950 671.250 767.850 673.050 ;
        RECT 763.950 670.950 766.050 671.250 ;
        RECT 775.050 670.950 775.950 675.000 ;
        RECT 785.100 673.800 786.150 675.000 ;
        RECT 785.100 672.600 792.000 673.800 ;
        RECT 785.100 672.000 786.900 672.600 ;
        RECT 791.100 671.850 792.000 672.600 ;
        RECT 788.100 670.950 789.900 671.700 ;
        RECT 775.050 668.850 778.050 670.950 ;
        RECT 781.950 669.900 789.900 670.950 ;
        RECT 791.100 670.050 792.900 671.850 ;
        RECT 781.950 668.850 784.050 669.900 ;
        RECT 763.950 665.400 765.750 667.200 ;
        RECT 764.850 664.200 769.050 665.400 ;
        RECT 775.050 664.200 775.950 668.850 ;
        RECT 783.750 665.100 785.550 665.400 ;
        RECT 677.550 651.750 679.350 657.600 ;
        RECT 680.550 651.750 682.350 657.600 ;
        RECT 683.550 651.750 685.350 657.600 ;
        RECT 697.650 651.750 699.450 657.600 ;
        RECT 700.650 651.750 702.450 657.600 ;
        RECT 703.650 651.750 705.450 657.600 ;
        RECT 713.550 651.750 715.350 657.600 ;
        RECT 716.550 651.750 718.350 657.600 ;
        RECT 728.550 651.750 730.350 657.600 ;
        RECT 731.550 651.750 733.350 657.600 ;
        RECT 734.550 651.750 736.350 657.600 ;
        RECT 747.300 651.750 749.100 663.600 ;
        RECT 751.500 651.750 753.300 663.600 ;
        RECT 754.800 651.750 756.600 657.600 ;
        RECT 761.550 651.750 763.350 663.600 ;
        RECT 766.950 663.300 769.050 664.200 ;
        RECT 769.950 663.300 775.950 664.200 ;
        RECT 777.150 664.800 785.550 665.100 ;
        RECT 793.950 664.800 794.850 677.400 ;
        RECT 803.550 678.300 805.350 683.250 ;
        RECT 806.550 679.200 808.350 683.250 ;
        RECT 809.550 678.300 811.350 683.250 ;
        RECT 803.550 676.950 811.350 678.300 ;
        RECT 812.550 677.400 814.350 683.250 ;
        RECT 824.550 680.400 826.350 683.250 ;
        RECT 827.550 680.400 829.350 683.250 ;
        RECT 830.550 680.400 832.350 683.250 ;
        RECT 812.550 675.300 813.750 677.400 ;
        RECT 828.450 676.200 829.350 680.400 ;
        RECT 833.550 677.400 835.350 683.250 ;
        RECT 847.650 677.400 849.450 683.250 ;
        RECT 828.450 675.300 831.750 676.200 ;
        RECT 810.000 674.250 813.750 675.300 ;
        RECT 829.950 674.400 831.750 675.300 ;
        RECT 806.100 672.150 807.900 673.950 ;
        RECT 802.950 668.850 805.050 670.950 ;
        RECT 805.950 670.050 808.050 672.150 ;
        RECT 809.850 670.950 811.050 674.250 ;
        RECT 823.950 671.850 826.050 673.950 ;
        RECT 808.950 668.850 811.050 670.950 ;
        RECT 824.100 670.050 825.900 671.850 ;
        RECT 826.950 668.850 829.050 670.950 ;
        RECT 803.100 667.050 804.900 668.850 ;
        RECT 777.150 664.200 794.850 664.800 ;
        RECT 769.950 662.400 770.850 663.300 ;
        RECT 768.150 660.600 770.850 662.400 ;
        RECT 771.750 662.100 773.550 662.400 ;
        RECT 777.150 662.100 778.050 664.200 ;
        RECT 783.750 663.600 794.850 664.200 ;
        RECT 808.950 663.600 810.150 668.850 ;
        RECT 811.950 665.850 814.050 667.950 ;
        RECT 827.100 667.050 828.900 668.850 ;
        RECT 830.700 666.150 831.600 674.400 ;
        RECT 834.000 672.150 835.050 677.400 ;
        RECT 848.250 675.300 849.450 677.400 ;
        RECT 850.650 678.300 852.450 683.250 ;
        RECT 853.650 679.200 855.450 683.250 ;
        RECT 856.650 678.300 858.450 683.250 ;
        RECT 850.650 676.950 858.450 678.300 ;
        RECT 848.250 674.250 852.000 675.300 ;
        RECT 832.950 670.050 835.050 672.150 ;
        RECT 850.950 670.950 852.150 674.250 ;
        RECT 854.100 672.150 855.900 673.950 ;
        RECT 829.950 666.000 831.750 666.150 ;
        RECT 811.950 664.050 813.750 665.850 ;
        RECT 824.550 664.800 831.750 666.000 ;
        RECT 824.550 663.600 825.750 664.800 ;
        RECT 829.950 664.350 831.750 664.800 ;
        RECT 771.750 661.200 778.050 662.100 ;
        RECT 778.950 662.700 780.750 663.300 ;
        RECT 778.950 661.500 786.450 662.700 ;
        RECT 771.750 660.600 773.550 661.200 ;
        RECT 785.250 660.600 786.450 661.500 ;
        RECT 766.950 657.600 770.850 659.700 ;
        RECT 775.950 658.500 782.850 660.300 ;
        RECT 785.250 658.500 790.050 660.600 ;
        RECT 764.550 651.750 766.350 654.600 ;
        RECT 769.050 651.750 770.850 657.600 ;
        RECT 773.250 651.750 775.050 657.600 ;
        RECT 777.150 651.750 778.950 658.500 ;
        RECT 785.250 657.600 786.450 658.500 ;
        RECT 780.150 651.750 781.950 657.600 ;
        RECT 784.950 651.750 786.750 657.600 ;
        RECT 790.050 651.750 791.850 657.600 ;
        RECT 793.050 651.750 794.850 663.600 ;
        RECT 804.300 651.750 806.100 663.600 ;
        RECT 808.500 651.750 810.300 663.600 ;
        RECT 811.800 651.750 813.600 657.600 ;
        RECT 824.550 651.750 826.350 663.600 ;
        RECT 833.100 663.450 834.450 670.050 ;
        RECT 850.950 668.850 853.050 670.950 ;
        RECT 853.950 670.050 856.050 672.150 ;
        RECT 856.950 668.850 859.050 670.950 ;
        RECT 847.950 665.850 850.050 667.950 ;
        RECT 848.250 664.050 850.050 665.850 ;
        RECT 851.850 663.600 853.050 668.850 ;
        RECT 857.100 667.050 858.900 668.850 ;
        RECT 829.050 651.750 830.850 663.450 ;
        RECT 832.050 662.100 834.450 663.450 ;
        RECT 832.050 651.750 833.850 662.100 ;
        RECT 848.400 651.750 850.200 657.600 ;
        RECT 851.700 651.750 853.500 663.600 ;
        RECT 855.900 651.750 857.700 663.600 ;
        RECT 14.400 641.400 16.200 647.250 ;
        RECT 17.700 635.400 19.500 647.250 ;
        RECT 21.900 635.400 23.700 647.250 ;
        RECT 35.400 641.400 37.200 647.250 ;
        RECT 38.700 635.400 40.500 647.250 ;
        RECT 42.900 635.400 44.700 647.250 ;
        RECT 58.650 641.400 60.450 647.250 ;
        RECT 61.650 642.000 63.450 647.250 ;
        RECT 59.250 641.100 60.450 641.400 ;
        RECT 64.650 641.400 66.450 647.250 ;
        RECT 67.650 641.400 69.450 647.250 ;
        RECT 79.650 641.400 81.450 647.250 ;
        RECT 82.650 642.000 84.450 647.250 ;
        RECT 64.650 641.100 66.300 641.400 ;
        RECT 59.250 640.200 66.300 641.100 ;
        RECT 80.250 641.100 81.450 641.400 ;
        RECT 85.650 641.400 87.450 647.250 ;
        RECT 88.650 641.400 90.450 647.250 ;
        RECT 85.650 641.100 87.300 641.400 ;
        RECT 80.250 640.200 87.300 641.100 ;
        RECT 14.250 633.150 16.050 634.950 ;
        RECT 13.950 631.050 16.050 633.150 ;
        RECT 17.850 630.150 19.050 635.400 ;
        RECT 35.250 633.150 37.050 634.950 ;
        RECT 23.100 630.150 24.900 631.950 ;
        RECT 34.950 631.050 37.050 633.150 ;
        RECT 38.850 630.150 40.050 635.400 ;
        RECT 59.250 631.950 60.300 640.200 ;
        RECT 65.100 636.150 66.900 637.950 ;
        RECT 61.950 633.150 63.750 634.950 ;
        RECT 64.950 634.050 67.050 636.150 ;
        RECT 68.100 633.150 69.900 634.950 ;
        RECT 44.100 630.150 45.900 631.950 ;
        RECT 16.950 628.050 19.050 630.150 ;
        RECT 16.950 624.750 18.150 628.050 ;
        RECT 19.950 626.850 22.050 628.950 ;
        RECT 22.950 628.050 25.050 630.150 ;
        RECT 37.950 628.050 40.050 630.150 ;
        RECT 20.100 625.050 21.900 626.850 ;
        RECT 37.950 624.750 39.150 628.050 ;
        RECT 40.950 626.850 43.050 628.950 ;
        RECT 43.950 628.050 46.050 630.150 ;
        RECT 58.950 629.850 61.050 631.950 ;
        RECT 61.950 631.050 64.050 633.150 ;
        RECT 67.950 631.050 70.050 633.150 ;
        RECT 80.250 631.950 81.300 640.200 ;
        RECT 86.100 636.150 87.900 637.950 ;
        RECT 102.150 636.900 103.950 647.250 ;
        RECT 82.950 633.150 84.750 634.950 ;
        RECT 85.950 634.050 88.050 636.150 ;
        RECT 101.550 635.550 103.950 636.900 ;
        RECT 105.150 635.550 106.950 647.250 ;
        RECT 89.100 633.150 90.900 634.950 ;
        RECT 79.950 629.850 82.050 631.950 ;
        RECT 82.950 631.050 85.050 633.150 ;
        RECT 88.950 631.050 91.050 633.150 ;
        RECT 41.100 625.050 42.900 626.850 ;
        RECT 59.400 625.650 60.600 629.850 ;
        RECT 80.400 625.650 81.600 629.850 ;
        RECT 101.550 628.950 102.900 635.550 ;
        RECT 109.650 635.400 111.450 647.250 ;
        RECT 122.400 641.400 124.200 647.250 ;
        RECT 125.700 635.400 127.500 647.250 ;
        RECT 129.900 635.400 131.700 647.250 ;
        RECT 140.550 641.400 142.350 647.250 ;
        RECT 143.550 641.400 145.350 647.250 ;
        RECT 104.250 634.200 106.050 634.650 ;
        RECT 110.250 634.200 111.450 635.400 ;
        RECT 104.250 633.000 111.450 634.200 ;
        RECT 122.250 633.150 124.050 634.950 ;
        RECT 104.250 632.850 106.050 633.000 ;
        RECT 100.950 626.850 103.050 628.950 ;
        RECT 14.250 623.700 18.000 624.750 ;
        RECT 35.250 623.700 39.000 624.750 ;
        RECT 59.400 624.000 63.900 625.650 ;
        RECT 14.250 621.600 15.450 623.700 ;
        RECT 13.650 615.750 15.450 621.600 ;
        RECT 16.650 620.700 24.450 622.050 ;
        RECT 35.250 621.600 36.450 623.700 ;
        RECT 16.650 615.750 18.450 620.700 ;
        RECT 19.650 615.750 21.450 619.800 ;
        RECT 22.650 615.750 24.450 620.700 ;
        RECT 34.650 615.750 36.450 621.600 ;
        RECT 37.650 620.700 45.450 622.050 ;
        RECT 37.650 615.750 39.450 620.700 ;
        RECT 40.650 615.750 42.450 619.800 ;
        RECT 43.650 615.750 45.450 620.700 ;
        RECT 62.100 615.750 63.900 624.000 ;
        RECT 67.500 615.750 69.300 624.600 ;
        RECT 80.400 624.000 84.900 625.650 ;
        RECT 73.950 621.450 76.050 622.050 ;
        RECT 79.950 621.450 82.050 622.050 ;
        RECT 73.950 620.550 82.050 621.450 ;
        RECT 73.950 619.950 76.050 620.550 ;
        RECT 79.950 619.950 82.050 620.550 ;
        RECT 83.100 615.750 84.900 624.000 ;
        RECT 88.500 615.750 90.300 624.600 ;
        RECT 100.950 621.600 102.000 626.850 ;
        RECT 104.400 624.600 105.300 632.850 ;
        RECT 107.100 630.150 108.900 631.950 ;
        RECT 121.950 631.050 124.050 633.150 ;
        RECT 125.850 630.150 127.050 635.400 ;
        RECT 131.100 630.150 132.900 631.950 ;
        RECT 106.950 628.050 109.050 630.150 ;
        RECT 110.100 627.150 111.900 628.950 ;
        RECT 124.950 628.050 127.050 630.150 ;
        RECT 109.950 625.050 112.050 627.150 ;
        RECT 124.950 624.750 126.150 628.050 ;
        RECT 127.950 626.850 130.050 628.950 ;
        RECT 130.950 628.050 133.050 630.150 ;
        RECT 143.400 628.950 144.600 641.400 ;
        RECT 157.650 635.400 159.450 647.250 ;
        RECT 160.650 636.300 162.450 647.250 ;
        RECT 163.650 637.200 165.450 647.250 ;
        RECT 166.650 636.300 168.450 647.250 ;
        RECT 181.650 641.400 183.450 647.250 ;
        RECT 184.650 642.000 186.450 647.250 ;
        RECT 160.650 635.400 168.450 636.300 ;
        RECT 182.250 641.100 183.450 641.400 ;
        RECT 187.650 641.400 189.450 647.250 ;
        RECT 190.650 641.400 192.450 647.250 ;
        RECT 202.650 641.400 204.450 647.250 ;
        RECT 205.650 641.400 207.450 647.250 ;
        RECT 208.650 641.400 210.450 647.250 ;
        RECT 220.650 641.400 222.450 647.250 ;
        RECT 223.650 641.400 225.450 647.250 ;
        RECT 226.650 641.400 228.450 647.250 ;
        RECT 187.650 641.100 189.300 641.400 ;
        RECT 182.250 640.200 189.300 641.100 ;
        RECT 158.100 630.150 159.300 635.400 ;
        RECT 182.250 631.950 183.300 640.200 ;
        RECT 188.100 636.150 189.900 637.950 ;
        RECT 184.950 633.150 186.750 634.950 ;
        RECT 187.950 634.050 190.050 636.150 ;
        RECT 191.100 633.150 192.900 634.950 ;
        RECT 206.250 633.150 207.450 641.400 ;
        RECT 224.250 633.150 225.450 641.400 ;
        RECT 240.450 635.400 242.250 647.250 ;
        RECT 244.650 635.400 246.450 647.250 ;
        RECT 256.650 641.400 258.450 647.250 ;
        RECT 259.650 642.000 261.450 647.250 ;
        RECT 257.250 641.100 258.450 641.400 ;
        RECT 262.650 641.400 264.450 647.250 ;
        RECT 265.650 641.400 267.450 647.250 ;
        RECT 277.650 641.400 279.450 647.250 ;
        RECT 280.650 642.000 282.450 647.250 ;
        RECT 262.650 641.100 264.300 641.400 ;
        RECT 257.250 640.200 264.300 641.100 ;
        RECT 278.250 641.100 279.450 641.400 ;
        RECT 283.650 641.400 285.450 647.250 ;
        RECT 286.650 641.400 288.450 647.250 ;
        RECT 296.550 641.400 298.350 647.250 ;
        RECT 299.550 641.400 301.350 647.250 ;
        RECT 302.550 642.000 304.350 647.250 ;
        RECT 283.650 641.100 285.300 641.400 ;
        RECT 278.250 640.200 285.300 641.100 ;
        RECT 299.700 641.100 301.350 641.400 ;
        RECT 305.550 641.400 307.350 647.250 ;
        RECT 317.550 641.400 319.350 647.250 ;
        RECT 320.550 641.400 322.350 647.250 ;
        RECT 323.550 642.000 325.350 647.250 ;
        RECT 305.550 641.100 306.750 641.400 ;
        RECT 299.700 640.200 306.750 641.100 ;
        RECT 320.700 641.100 322.350 641.400 ;
        RECT 326.550 641.400 328.350 647.250 ;
        RECT 326.550 641.100 327.750 641.400 ;
        RECT 320.700 640.200 327.750 641.100 ;
        RECT 240.450 634.350 243.000 635.400 ;
        RECT 140.100 627.150 141.900 628.950 ;
        RECT 128.100 625.050 129.900 626.850 ;
        RECT 139.950 625.050 142.050 627.150 ;
        RECT 142.950 626.850 145.050 628.950 ;
        RECT 157.950 628.050 160.050 630.150 ;
        RECT 181.950 629.850 184.050 631.950 ;
        RECT 184.950 631.050 187.050 633.150 ;
        RECT 190.950 631.050 193.050 633.150 ;
        RECT 202.950 629.850 205.050 631.950 ;
        RECT 205.950 631.050 208.050 633.150 ;
        RECT 104.250 623.700 106.050 624.600 ;
        RECT 122.250 623.700 126.000 624.750 ;
        RECT 104.250 622.800 107.550 623.700 ;
        RECT 100.650 615.750 102.450 621.600 ;
        RECT 106.650 618.600 107.550 622.800 ;
        RECT 122.250 621.600 123.450 623.700 ;
        RECT 103.650 615.750 105.450 618.600 ;
        RECT 106.650 615.750 108.450 618.600 ;
        RECT 109.650 615.750 111.450 618.600 ;
        RECT 121.650 615.750 123.450 621.600 ;
        RECT 124.650 620.700 132.450 622.050 ;
        RECT 124.650 615.750 126.450 620.700 ;
        RECT 127.650 615.750 129.450 619.800 ;
        RECT 130.650 615.750 132.450 620.700 ;
        RECT 143.400 618.600 144.600 626.850 ;
        RECT 158.100 621.600 159.300 628.050 ;
        RECT 160.950 626.850 163.050 628.950 ;
        RECT 164.100 627.150 165.900 628.950 ;
        RECT 161.100 625.050 162.900 626.850 ;
        RECT 163.950 625.050 166.050 627.150 ;
        RECT 166.950 626.850 169.050 628.950 ;
        RECT 167.100 625.050 168.900 626.850 ;
        RECT 182.400 625.650 183.600 629.850 ;
        RECT 203.100 628.050 204.900 629.850 ;
        RECT 182.400 624.000 186.900 625.650 ;
        RECT 158.100 619.950 163.800 621.600 ;
        RECT 140.550 615.750 142.350 618.600 ;
        RECT 143.550 615.750 145.350 618.600 ;
        RECT 158.700 615.750 160.500 618.600 ;
        RECT 162.000 615.750 163.800 619.950 ;
        RECT 166.200 615.750 168.000 621.600 ;
        RECT 185.100 615.750 186.900 624.000 ;
        RECT 190.500 615.750 192.300 624.600 ;
        RECT 206.250 623.700 207.450 631.050 ;
        RECT 208.950 629.850 211.050 631.950 ;
        RECT 220.950 629.850 223.050 631.950 ;
        RECT 223.950 631.050 226.050 633.150 ;
        RECT 209.100 628.050 210.900 629.850 ;
        RECT 221.100 628.050 222.900 629.850 ;
        RECT 224.250 623.700 225.450 631.050 ;
        RECT 226.950 629.850 229.050 631.950 ;
        RECT 239.100 630.150 240.900 631.950 ;
        RECT 227.100 628.050 228.900 629.850 ;
        RECT 238.950 628.050 241.050 630.150 ;
        RECT 203.850 622.800 207.450 623.700 ;
        RECT 221.850 622.800 225.450 623.700 ;
        RECT 241.950 627.150 243.000 634.350 ;
        RECT 257.250 631.950 258.300 640.200 ;
        RECT 263.100 636.150 264.900 637.950 ;
        RECT 259.950 633.150 261.750 634.950 ;
        RECT 262.950 634.050 265.050 636.150 ;
        RECT 266.100 633.150 267.900 634.950 ;
        RECT 245.100 630.150 246.900 631.950 ;
        RECT 244.950 628.050 247.050 630.150 ;
        RECT 256.950 629.850 259.050 631.950 ;
        RECT 259.950 631.050 262.050 633.150 ;
        RECT 265.950 631.050 268.050 633.150 ;
        RECT 278.250 631.950 279.300 640.200 ;
        RECT 284.100 636.150 285.900 637.950 ;
        RECT 299.100 636.150 300.900 637.950 ;
        RECT 280.950 633.150 282.750 634.950 ;
        RECT 283.950 634.050 286.050 636.150 ;
        RECT 287.100 633.150 288.900 634.950 ;
        RECT 296.100 633.150 297.900 634.950 ;
        RECT 298.950 634.050 301.050 636.150 ;
        RECT 302.250 633.150 304.050 634.950 ;
        RECT 277.950 629.850 280.050 631.950 ;
        RECT 280.950 631.050 283.050 633.150 ;
        RECT 286.950 631.050 289.050 633.150 ;
        RECT 295.950 631.050 298.050 633.150 ;
        RECT 301.950 631.050 304.050 633.150 ;
        RECT 305.700 631.950 306.750 640.200 ;
        RECT 320.100 636.150 321.900 637.950 ;
        RECT 317.100 633.150 318.900 634.950 ;
        RECT 319.950 634.050 322.050 636.150 ;
        RECT 323.250 633.150 325.050 634.950 ;
        RECT 304.950 629.850 307.050 631.950 ;
        RECT 316.950 631.050 319.050 633.150 ;
        RECT 322.950 631.050 325.050 633.150 ;
        RECT 326.700 631.950 327.750 640.200 ;
        RECT 342.450 635.400 344.250 647.250 ;
        RECT 346.650 635.400 348.450 647.250 ;
        RECT 362.400 641.400 364.200 647.250 ;
        RECT 365.700 635.400 367.500 647.250 ;
        RECT 369.900 635.400 371.700 647.250 ;
        RECT 385.650 641.400 387.450 647.250 ;
        RECT 388.650 642.000 390.450 647.250 ;
        RECT 386.250 641.100 387.450 641.400 ;
        RECT 391.650 641.400 393.450 647.250 ;
        RECT 394.650 641.400 396.450 647.250 ;
        RECT 404.550 641.400 406.350 647.250 ;
        RECT 407.550 641.400 409.350 647.250 ;
        RECT 422.550 641.400 424.350 647.250 ;
        RECT 425.550 641.400 427.350 647.250 ;
        RECT 428.550 642.000 430.350 647.250 ;
        RECT 391.650 641.100 393.300 641.400 ;
        RECT 386.250 640.200 393.300 641.100 ;
        RECT 342.450 634.350 345.000 635.400 ;
        RECT 325.950 629.850 328.050 631.950 ;
        RECT 341.100 630.150 342.900 631.950 ;
        RECT 241.950 625.050 244.050 627.150 ;
        RECT 257.400 625.650 258.600 629.850 ;
        RECT 278.400 625.650 279.600 629.850 ;
        RECT 305.400 625.650 306.600 629.850 ;
        RECT 326.400 625.650 327.600 629.850 ;
        RECT 340.950 628.050 343.050 630.150 ;
        RECT 203.850 615.750 205.650 622.800 ;
        RECT 208.350 615.750 210.150 621.600 ;
        RECT 221.850 615.750 223.650 622.800 ;
        RECT 226.350 615.750 228.150 621.600 ;
        RECT 241.950 618.600 243.000 625.050 ;
        RECT 257.400 624.000 261.900 625.650 ;
        RECT 238.650 615.750 240.450 618.600 ;
        RECT 241.650 615.750 243.450 618.600 ;
        RECT 244.650 615.750 246.450 618.600 ;
        RECT 260.100 615.750 261.900 624.000 ;
        RECT 265.500 615.750 267.300 624.600 ;
        RECT 278.400 624.000 282.900 625.650 ;
        RECT 281.100 615.750 282.900 624.000 ;
        RECT 286.500 615.750 288.300 624.600 ;
        RECT 296.700 615.750 298.500 624.600 ;
        RECT 302.100 624.000 306.600 625.650 ;
        RECT 302.100 615.750 303.900 624.000 ;
        RECT 317.700 615.750 319.500 624.600 ;
        RECT 323.100 624.000 327.600 625.650 ;
        RECT 343.950 627.150 345.000 634.350 ;
        RECT 362.250 633.150 364.050 634.950 ;
        RECT 347.100 630.150 348.900 631.950 ;
        RECT 361.950 631.050 364.050 633.150 ;
        RECT 365.850 630.150 367.050 635.400 ;
        RECT 386.250 631.950 387.300 640.200 ;
        RECT 392.100 636.150 393.900 637.950 ;
        RECT 388.950 633.150 390.750 634.950 ;
        RECT 391.950 634.050 394.050 636.150 ;
        RECT 395.100 633.150 396.900 634.950 ;
        RECT 371.100 630.150 372.900 631.950 ;
        RECT 346.950 628.050 349.050 630.150 ;
        RECT 364.950 628.050 367.050 630.150 ;
        RECT 343.950 625.050 346.050 627.150 ;
        RECT 323.100 615.750 324.900 624.000 ;
        RECT 343.950 618.600 345.000 625.050 ;
        RECT 364.950 624.750 366.150 628.050 ;
        RECT 367.950 626.850 370.050 628.950 ;
        RECT 370.950 628.050 373.050 630.150 ;
        RECT 385.950 629.850 388.050 631.950 ;
        RECT 388.950 631.050 391.050 633.150 ;
        RECT 394.950 631.050 397.050 633.150 ;
        RECT 368.100 625.050 369.900 626.850 ;
        RECT 386.400 625.650 387.600 629.850 ;
        RECT 407.400 628.950 408.600 641.400 ;
        RECT 425.700 641.100 427.350 641.400 ;
        RECT 431.550 641.400 433.350 647.250 ;
        RECT 443.550 641.400 445.350 647.250 ;
        RECT 446.550 641.400 448.350 647.250 ;
        RECT 449.550 641.400 451.350 647.250 ;
        RECT 431.550 641.100 432.750 641.400 ;
        RECT 425.700 640.200 432.750 641.100 ;
        RECT 425.100 636.150 426.900 637.950 ;
        RECT 422.100 633.150 423.900 634.950 ;
        RECT 424.950 634.050 427.050 636.150 ;
        RECT 428.250 633.150 430.050 634.950 ;
        RECT 421.950 631.050 424.050 633.150 ;
        RECT 427.950 631.050 430.050 633.150 ;
        RECT 431.700 631.950 432.750 640.200 ;
        RECT 446.550 633.150 447.750 641.400 ;
        RECT 461.550 636.300 463.350 647.250 ;
        RECT 464.550 637.200 466.350 647.250 ;
        RECT 467.550 636.300 469.350 647.250 ;
        RECT 461.550 635.400 469.350 636.300 ;
        RECT 470.550 635.400 472.350 647.250 ;
        RECT 482.550 636.300 484.350 647.250 ;
        RECT 485.550 637.200 487.350 647.250 ;
        RECT 488.550 636.300 490.350 647.250 ;
        RECT 482.550 635.400 490.350 636.300 ;
        RECT 491.550 635.400 493.350 647.250 ;
        RECT 504.300 635.400 506.100 647.250 ;
        RECT 508.500 635.400 510.300 647.250 ;
        RECT 511.800 641.400 513.600 647.250 ;
        RECT 527.550 641.400 529.350 647.250 ;
        RECT 530.550 641.400 532.350 647.250 ;
        RECT 542.550 641.400 544.350 647.250 ;
        RECT 545.550 641.400 547.350 647.250 ;
        RECT 548.550 642.000 550.350 647.250 ;
        RECT 430.950 629.850 433.050 631.950 ;
        RECT 442.950 629.850 445.050 631.950 ;
        RECT 445.950 631.050 448.050 633.150 ;
        RECT 404.100 627.150 405.900 628.950 ;
        RECT 362.250 623.700 366.000 624.750 ;
        RECT 386.400 624.000 390.900 625.650 ;
        RECT 403.950 625.050 406.050 627.150 ;
        RECT 406.950 626.850 409.050 628.950 ;
        RECT 362.250 621.600 363.450 623.700 ;
        RECT 340.650 615.750 342.450 618.600 ;
        RECT 343.650 615.750 345.450 618.600 ;
        RECT 346.650 615.750 348.450 618.600 ;
        RECT 361.650 615.750 363.450 621.600 ;
        RECT 364.650 620.700 372.450 622.050 ;
        RECT 364.650 615.750 366.450 620.700 ;
        RECT 367.650 615.750 369.450 619.800 ;
        RECT 370.650 615.750 372.450 620.700 ;
        RECT 389.100 615.750 390.900 624.000 ;
        RECT 394.500 615.750 396.300 624.600 ;
        RECT 407.400 618.600 408.600 626.850 ;
        RECT 431.400 625.650 432.600 629.850 ;
        RECT 443.100 628.050 444.900 629.850 ;
        RECT 404.550 615.750 406.350 618.600 ;
        RECT 407.550 615.750 409.350 618.600 ;
        RECT 422.700 615.750 424.500 624.600 ;
        RECT 428.100 624.000 432.600 625.650 ;
        RECT 428.100 615.750 429.900 624.000 ;
        RECT 446.550 623.700 447.750 631.050 ;
        RECT 448.950 629.850 451.050 631.950 ;
        RECT 470.700 630.150 471.900 635.400 ;
        RECT 491.700 630.150 492.900 635.400 ;
        RECT 503.100 630.150 504.900 631.950 ;
        RECT 508.950 630.150 510.150 635.400 ;
        RECT 511.950 633.150 513.750 634.950 ;
        RECT 511.950 631.050 514.050 633.150 ;
        RECT 449.100 628.050 450.900 629.850 ;
        RECT 460.950 626.850 463.050 628.950 ;
        RECT 464.100 627.150 465.900 628.950 ;
        RECT 461.100 625.050 462.900 626.850 ;
        RECT 463.950 625.050 466.050 627.150 ;
        RECT 466.950 626.850 469.050 628.950 ;
        RECT 469.950 628.050 472.050 630.150 ;
        RECT 467.100 625.050 468.900 626.850 ;
        RECT 446.550 622.800 450.150 623.700 ;
        RECT 443.850 615.750 445.650 621.600 ;
        RECT 448.350 615.750 450.150 622.800 ;
        RECT 470.700 621.600 471.900 628.050 ;
        RECT 481.950 626.850 484.050 628.950 ;
        RECT 485.100 627.150 486.900 628.950 ;
        RECT 482.100 625.050 483.900 626.850 ;
        RECT 484.950 625.050 487.050 627.150 ;
        RECT 487.950 626.850 490.050 628.950 ;
        RECT 490.950 628.050 493.050 630.150 ;
        RECT 502.950 628.050 505.050 630.150 ;
        RECT 488.100 625.050 489.900 626.850 ;
        RECT 491.700 621.600 492.900 628.050 ;
        RECT 505.950 626.850 508.050 628.950 ;
        RECT 508.950 628.050 511.050 630.150 ;
        RECT 530.400 628.950 531.600 641.400 ;
        RECT 545.700 641.100 547.350 641.400 ;
        RECT 551.550 641.400 553.350 647.250 ;
        RECT 563.550 641.400 565.350 647.250 ;
        RECT 566.550 641.400 568.350 647.250 ;
        RECT 569.550 642.000 571.350 647.250 ;
        RECT 551.550 641.100 552.750 641.400 ;
        RECT 545.700 640.200 552.750 641.100 ;
        RECT 566.700 641.100 568.350 641.400 ;
        RECT 572.550 641.400 574.350 647.250 ;
        RECT 586.650 641.400 588.450 647.250 ;
        RECT 589.650 641.400 591.450 647.250 ;
        RECT 592.650 641.400 594.450 647.250 ;
        RECT 607.650 641.400 609.450 647.250 ;
        RECT 610.650 641.400 612.450 647.250 ;
        RECT 613.650 641.400 615.450 647.250 ;
        RECT 625.650 641.400 627.450 647.250 ;
        RECT 628.650 641.400 630.450 647.250 ;
        RECT 631.650 641.400 633.450 647.250 ;
        RECT 644.400 641.400 646.200 647.250 ;
        RECT 572.550 641.100 573.750 641.400 ;
        RECT 566.700 640.200 573.750 641.100 ;
        RECT 545.100 636.150 546.900 637.950 ;
        RECT 542.100 633.150 543.900 634.950 ;
        RECT 544.950 634.050 547.050 636.150 ;
        RECT 548.250 633.150 550.050 634.950 ;
        RECT 541.950 631.050 544.050 633.150 ;
        RECT 547.950 631.050 550.050 633.150 ;
        RECT 551.700 631.950 552.750 640.200 ;
        RECT 566.100 636.150 567.900 637.950 ;
        RECT 563.100 633.150 564.900 634.950 ;
        RECT 565.950 634.050 568.050 636.150 ;
        RECT 569.250 633.150 571.050 634.950 ;
        RECT 550.950 629.850 553.050 631.950 ;
        RECT 562.950 631.050 565.050 633.150 ;
        RECT 568.950 631.050 571.050 633.150 ;
        RECT 572.700 631.950 573.750 640.200 ;
        RECT 590.250 633.150 591.450 641.400 ;
        RECT 611.250 633.150 612.450 641.400 ;
        RECT 629.250 633.150 630.450 641.400 ;
        RECT 647.700 635.400 649.500 647.250 ;
        RECT 651.900 635.400 653.700 647.250 ;
        RECT 662.550 635.400 664.350 647.250 ;
        RECT 667.050 635.550 668.850 647.250 ;
        RECT 670.050 636.900 671.850 647.250 ;
        RECT 686.400 641.400 688.200 647.250 ;
        RECT 670.050 635.550 672.450 636.900 ;
        RECT 644.250 633.150 646.050 634.950 ;
        RECT 571.950 629.850 574.050 631.950 ;
        RECT 586.950 629.850 589.050 631.950 ;
        RECT 589.950 631.050 592.050 633.150 ;
        RECT 506.100 625.050 507.900 626.850 ;
        RECT 509.850 624.750 511.050 628.050 ;
        RECT 527.100 627.150 528.900 628.950 ;
        RECT 526.950 625.050 529.050 627.150 ;
        RECT 529.950 626.850 532.050 628.950 ;
        RECT 510.000 623.700 513.750 624.750 ;
        RECT 462.000 615.750 463.800 621.600 ;
        RECT 466.200 619.950 471.900 621.600 ;
        RECT 466.200 615.750 468.000 619.950 ;
        RECT 469.500 615.750 471.300 618.600 ;
        RECT 483.000 615.750 484.800 621.600 ;
        RECT 487.200 619.950 492.900 621.600 ;
        RECT 503.550 620.700 511.350 622.050 ;
        RECT 487.200 615.750 489.000 619.950 ;
        RECT 490.500 615.750 492.300 618.600 ;
        RECT 503.550 615.750 505.350 620.700 ;
        RECT 506.550 615.750 508.350 619.800 ;
        RECT 509.550 615.750 511.350 620.700 ;
        RECT 512.550 621.600 513.750 623.700 ;
        RECT 512.550 615.750 514.350 621.600 ;
        RECT 530.400 618.600 531.600 626.850 ;
        RECT 551.400 625.650 552.600 629.850 ;
        RECT 572.400 625.650 573.600 629.850 ;
        RECT 587.100 628.050 588.900 629.850 ;
        RECT 527.550 615.750 529.350 618.600 ;
        RECT 530.550 615.750 532.350 618.600 ;
        RECT 542.700 615.750 544.500 624.600 ;
        RECT 548.100 624.000 552.600 625.650 ;
        RECT 548.100 615.750 549.900 624.000 ;
        RECT 563.700 615.750 565.500 624.600 ;
        RECT 569.100 624.000 573.600 625.650 ;
        RECT 569.100 615.750 570.900 624.000 ;
        RECT 590.250 623.700 591.450 631.050 ;
        RECT 592.950 629.850 595.050 631.950 ;
        RECT 607.950 629.850 610.050 631.950 ;
        RECT 610.950 631.050 613.050 633.150 ;
        RECT 593.100 628.050 594.900 629.850 ;
        RECT 608.100 628.050 609.900 629.850 ;
        RECT 611.250 623.700 612.450 631.050 ;
        RECT 613.950 629.850 616.050 631.950 ;
        RECT 625.950 629.850 628.050 631.950 ;
        RECT 628.950 631.050 631.050 633.150 ;
        RECT 614.100 628.050 615.900 629.850 ;
        RECT 626.100 628.050 627.900 629.850 ;
        RECT 629.250 623.700 630.450 631.050 ;
        RECT 631.950 629.850 634.050 631.950 ;
        RECT 643.950 631.050 646.050 633.150 ;
        RECT 647.850 630.150 649.050 635.400 ;
        RECT 662.550 634.200 663.750 635.400 ;
        RECT 667.950 634.200 669.750 634.650 ;
        RECT 662.550 633.000 669.750 634.200 ;
        RECT 667.950 632.850 669.750 633.000 ;
        RECT 653.100 630.150 654.900 631.950 ;
        RECT 665.100 630.150 666.900 631.950 ;
        RECT 632.100 628.050 633.900 629.850 ;
        RECT 646.950 628.050 649.050 630.150 ;
        RECT 646.950 624.750 648.150 628.050 ;
        RECT 649.950 626.850 652.050 628.950 ;
        RECT 652.950 628.050 655.050 630.150 ;
        RECT 662.100 627.150 663.900 628.950 ;
        RECT 664.950 628.050 667.050 630.150 ;
        RECT 650.100 625.050 651.900 626.850 ;
        RECT 661.950 625.050 664.050 627.150 ;
        RECT 587.850 622.800 591.450 623.700 ;
        RECT 608.850 622.800 612.450 623.700 ;
        RECT 626.850 622.800 630.450 623.700 ;
        RECT 644.250 623.700 648.000 624.750 ;
        RECT 668.700 624.600 669.600 632.850 ;
        RECT 671.100 628.950 672.450 635.550 ;
        RECT 689.700 635.400 691.500 647.250 ;
        RECT 693.900 635.400 695.700 647.250 ;
        RECT 708.300 635.400 710.100 647.250 ;
        RECT 712.500 635.400 714.300 647.250 ;
        RECT 715.800 641.400 717.600 647.250 ;
        RECT 728.550 635.400 730.350 647.250 ;
        RECT 732.750 635.400 734.550 647.250 ;
        RECT 746.550 641.400 748.350 647.250 ;
        RECT 749.550 641.400 751.350 647.250 ;
        RECT 686.250 633.150 688.050 634.950 ;
        RECT 685.950 631.050 688.050 633.150 ;
        RECT 689.850 630.150 691.050 635.400 ;
        RECT 695.100 630.150 696.900 631.950 ;
        RECT 707.100 630.150 708.900 631.950 ;
        RECT 712.950 630.150 714.150 635.400 ;
        RECT 715.950 633.150 717.750 634.950 ;
        RECT 732.000 634.350 734.550 635.400 ;
        RECT 715.950 631.050 718.050 633.150 ;
        RECT 728.100 630.150 729.900 631.950 ;
        RECT 670.950 626.850 673.050 628.950 ;
        RECT 667.950 623.700 669.750 624.600 ;
        RECT 587.850 615.750 589.650 622.800 ;
        RECT 592.350 615.750 594.150 621.600 ;
        RECT 608.850 615.750 610.650 622.800 ;
        RECT 613.350 615.750 615.150 621.600 ;
        RECT 626.850 615.750 628.650 622.800 ;
        RECT 644.250 621.600 645.450 623.700 ;
        RECT 666.450 622.800 669.750 623.700 ;
        RECT 631.350 615.750 633.150 621.600 ;
        RECT 643.650 615.750 645.450 621.600 ;
        RECT 646.650 620.700 654.450 622.050 ;
        RECT 646.650 615.750 648.450 620.700 ;
        RECT 649.650 615.750 651.450 619.800 ;
        RECT 652.650 615.750 654.450 620.700 ;
        RECT 666.450 618.600 667.350 622.800 ;
        RECT 672.000 621.600 673.050 626.850 ;
        RECT 688.950 628.050 691.050 630.150 ;
        RECT 688.950 624.750 690.150 628.050 ;
        RECT 691.950 626.850 694.050 628.950 ;
        RECT 694.950 628.050 697.050 630.150 ;
        RECT 706.950 628.050 709.050 630.150 ;
        RECT 709.950 626.850 712.050 628.950 ;
        RECT 712.950 628.050 715.050 630.150 ;
        RECT 727.950 628.050 730.050 630.150 ;
        RECT 692.100 625.050 693.900 626.850 ;
        RECT 710.100 625.050 711.900 626.850 ;
        RECT 713.850 624.750 715.050 628.050 ;
        RECT 732.000 627.150 733.050 634.350 ;
        RECT 734.100 630.150 735.900 631.950 ;
        RECT 733.950 628.050 736.050 630.150 ;
        RECT 749.400 628.950 750.600 641.400 ;
        RECT 764.550 636.300 766.350 647.250 ;
        RECT 767.550 637.200 769.350 647.250 ;
        RECT 770.550 636.300 772.350 647.250 ;
        RECT 764.550 635.400 772.350 636.300 ;
        RECT 773.550 635.400 775.350 647.250 ;
        RECT 786.300 635.400 788.100 647.250 ;
        RECT 790.500 635.400 792.300 647.250 ;
        RECT 793.800 641.400 795.600 647.250 ;
        RECT 806.550 641.400 808.350 647.250 ;
        RECT 809.550 641.400 811.350 647.250 ;
        RECT 757.950 633.450 760.050 634.050 ;
        RECT 769.950 633.450 772.050 634.050 ;
        RECT 757.950 632.550 772.050 633.450 ;
        RECT 757.950 631.950 760.050 632.550 ;
        RECT 769.950 631.950 772.050 632.550 ;
        RECT 773.700 630.150 774.900 635.400 ;
        RECT 785.100 630.150 786.900 631.950 ;
        RECT 790.950 630.150 792.150 635.400 ;
        RECT 793.950 633.150 795.750 634.950 ;
        RECT 793.950 631.050 796.050 633.150 ;
        RECT 746.100 627.150 747.900 628.950 ;
        RECT 730.950 625.050 733.050 627.150 ;
        RECT 745.950 625.050 748.050 627.150 ;
        RECT 748.950 626.850 751.050 628.950 ;
        RECT 763.950 626.850 766.050 628.950 ;
        RECT 767.100 627.150 768.900 628.950 ;
        RECT 686.250 623.700 690.000 624.750 ;
        RECT 714.000 623.700 717.750 624.750 ;
        RECT 686.250 621.600 687.450 623.700 ;
        RECT 662.550 615.750 664.350 618.600 ;
        RECT 665.550 615.750 667.350 618.600 ;
        RECT 668.550 615.750 670.350 618.600 ;
        RECT 671.550 615.750 673.350 621.600 ;
        RECT 685.650 615.750 687.450 621.600 ;
        RECT 688.650 620.700 696.450 622.050 ;
        RECT 688.650 615.750 690.450 620.700 ;
        RECT 691.650 615.750 693.450 619.800 ;
        RECT 694.650 615.750 696.450 620.700 ;
        RECT 707.550 620.700 715.350 622.050 ;
        RECT 707.550 615.750 709.350 620.700 ;
        RECT 710.550 615.750 712.350 619.800 ;
        RECT 713.550 615.750 715.350 620.700 ;
        RECT 716.550 621.600 717.750 623.700 ;
        RECT 716.550 615.750 718.350 621.600 ;
        RECT 732.000 618.600 733.050 625.050 ;
        RECT 749.400 618.600 750.600 626.850 ;
        RECT 764.100 625.050 765.900 626.850 ;
        RECT 766.950 625.050 769.050 627.150 ;
        RECT 769.950 626.850 772.050 628.950 ;
        RECT 772.950 628.050 775.050 630.150 ;
        RECT 784.950 628.050 787.050 630.150 ;
        RECT 770.100 625.050 771.900 626.850 ;
        RECT 773.700 621.600 774.900 628.050 ;
        RECT 787.950 626.850 790.050 628.950 ;
        RECT 790.950 628.050 793.050 630.150 ;
        RECT 809.400 628.950 810.600 641.400 ;
        RECT 822.300 635.400 824.100 647.250 ;
        RECT 826.500 635.400 828.300 647.250 ;
        RECT 829.800 641.400 831.600 647.250 ;
        RECT 837.150 635.400 838.950 647.250 ;
        RECT 840.150 641.400 841.950 647.250 ;
        RECT 845.250 641.400 847.050 647.250 ;
        RECT 850.050 641.400 851.850 647.250 ;
        RECT 845.550 640.500 846.750 641.400 ;
        RECT 853.050 640.500 854.850 647.250 ;
        RECT 856.950 641.400 858.750 647.250 ;
        RECT 861.150 641.400 862.950 647.250 ;
        RECT 865.650 644.400 867.450 647.250 ;
        RECT 841.950 638.400 846.750 640.500 ;
        RECT 849.150 638.700 856.050 640.500 ;
        RECT 861.150 639.300 865.050 641.400 ;
        RECT 845.550 637.500 846.750 638.400 ;
        RECT 858.450 637.800 860.250 638.400 ;
        RECT 845.550 636.300 853.050 637.500 ;
        RECT 851.250 635.700 853.050 636.300 ;
        RECT 853.950 636.900 860.250 637.800 ;
        RECT 821.100 630.150 822.900 631.950 ;
        RECT 826.950 630.150 828.150 635.400 ;
        RECT 829.950 633.150 831.750 634.950 ;
        RECT 837.150 634.800 848.250 635.400 ;
        RECT 853.950 634.800 854.850 636.900 ;
        RECT 858.450 636.600 860.250 636.900 ;
        RECT 861.150 636.600 863.850 638.400 ;
        RECT 861.150 635.700 862.050 636.600 ;
        RECT 837.150 634.200 854.850 634.800 ;
        RECT 829.950 631.050 832.050 633.150 ;
        RECT 788.100 625.050 789.900 626.850 ;
        RECT 791.850 624.750 793.050 628.050 ;
        RECT 806.100 627.150 807.900 628.950 ;
        RECT 805.950 625.050 808.050 627.150 ;
        RECT 808.950 626.850 811.050 628.950 ;
        RECT 820.950 628.050 823.050 630.150 ;
        RECT 823.950 626.850 826.050 628.950 ;
        RECT 826.950 628.050 829.050 630.150 ;
        RECT 792.000 623.700 795.750 624.750 ;
        RECT 728.550 615.750 730.350 618.600 ;
        RECT 731.550 615.750 733.350 618.600 ;
        RECT 734.550 615.750 736.350 618.600 ;
        RECT 746.550 615.750 748.350 618.600 ;
        RECT 749.550 615.750 751.350 618.600 ;
        RECT 765.000 615.750 766.800 621.600 ;
        RECT 769.200 619.950 774.900 621.600 ;
        RECT 785.550 620.700 793.350 622.050 ;
        RECT 769.200 615.750 771.000 619.950 ;
        RECT 772.500 615.750 774.300 618.600 ;
        RECT 785.550 615.750 787.350 620.700 ;
        RECT 788.550 615.750 790.350 619.800 ;
        RECT 791.550 615.750 793.350 620.700 ;
        RECT 794.550 621.600 795.750 623.700 ;
        RECT 794.550 615.750 796.350 621.600 ;
        RECT 809.400 618.600 810.600 626.850 ;
        RECT 824.100 625.050 825.900 626.850 ;
        RECT 827.850 624.750 829.050 628.050 ;
        RECT 828.000 623.700 831.750 624.750 ;
        RECT 821.550 620.700 829.350 622.050 ;
        RECT 806.550 615.750 808.350 618.600 ;
        RECT 809.550 615.750 811.350 618.600 ;
        RECT 821.550 615.750 823.350 620.700 ;
        RECT 824.550 615.750 826.350 619.800 ;
        RECT 827.550 615.750 829.350 620.700 ;
        RECT 830.550 621.600 831.750 623.700 ;
        RECT 837.150 621.600 838.050 634.200 ;
        RECT 846.450 633.900 854.850 634.200 ;
        RECT 856.050 634.800 862.050 635.700 ;
        RECT 862.950 634.800 865.050 635.700 ;
        RECT 868.650 635.400 870.450 647.250 ;
        RECT 846.450 633.600 848.250 633.900 ;
        RECT 856.050 630.150 856.950 634.800 ;
        RECT 862.950 633.600 867.150 634.800 ;
        RECT 866.250 631.800 868.050 633.600 ;
        RECT 847.950 629.100 850.050 630.150 ;
        RECT 839.100 627.150 840.900 628.950 ;
        RECT 842.100 628.050 850.050 629.100 ;
        RECT 853.950 628.050 856.950 630.150 ;
        RECT 842.100 627.300 843.900 628.050 ;
        RECT 840.000 626.400 840.900 627.150 ;
        RECT 845.100 626.400 846.900 627.000 ;
        RECT 840.000 625.200 846.900 626.400 ;
        RECT 845.850 624.000 846.900 625.200 ;
        RECT 856.050 624.000 856.950 628.050 ;
        RECT 865.950 627.750 868.050 628.050 ;
        RECT 864.150 625.950 868.050 627.750 ;
        RECT 869.250 625.950 870.450 635.400 ;
        RECT 845.850 623.100 856.950 624.000 ;
        RECT 865.950 623.850 870.450 625.950 ;
        RECT 845.850 622.200 846.900 623.100 ;
        RECT 856.050 622.800 856.950 623.100 ;
        RECT 830.550 615.750 832.350 621.600 ;
        RECT 837.150 615.750 838.950 621.600 ;
        RECT 841.950 619.500 844.050 621.600 ;
        RECT 845.550 620.400 847.350 622.200 ;
        RECT 848.850 621.450 850.650 622.200 ;
        RECT 848.850 620.400 853.800 621.450 ;
        RECT 856.050 621.000 857.850 622.800 ;
        RECT 869.250 621.600 870.450 623.850 ;
        RECT 862.950 620.700 865.050 621.600 ;
        RECT 843.000 618.600 844.050 619.500 ;
        RECT 852.750 618.600 853.800 620.400 ;
        RECT 861.300 619.500 865.050 620.700 ;
        RECT 861.300 618.600 862.350 619.500 ;
        RECT 840.150 615.750 841.950 618.600 ;
        RECT 843.000 617.700 846.750 618.600 ;
        RECT 844.950 615.750 846.750 617.700 ;
        RECT 849.450 615.750 851.250 618.600 ;
        RECT 852.750 615.750 854.550 618.600 ;
        RECT 856.650 615.750 858.450 618.600 ;
        RECT 860.850 615.750 862.650 618.600 ;
        RECT 865.350 615.750 867.150 618.600 ;
        RECT 868.650 615.750 870.450 621.600 ;
        RECT 10.650 608.400 12.450 611.250 ;
        RECT 13.650 608.400 15.450 611.250 ;
        RECT 11.400 600.150 12.600 608.400 ;
        RECT 26.550 606.300 28.350 611.250 ;
        RECT 29.550 607.200 31.350 611.250 ;
        RECT 32.550 606.300 34.350 611.250 ;
        RECT 26.550 604.950 34.350 606.300 ;
        RECT 35.550 605.400 37.350 611.250 ;
        RECT 49.650 608.400 51.450 611.250 ;
        RECT 52.650 608.400 54.450 611.250 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 35.550 603.300 36.750 605.400 ;
        RECT 33.000 602.250 36.750 603.300 ;
        RECT 10.950 598.050 13.050 600.150 ;
        RECT 13.950 599.850 16.050 601.950 ;
        RECT 14.100 598.050 15.900 599.850 ;
        RECT 11.400 585.600 12.600 598.050 ;
        RECT 13.950 591.450 16.050 592.050 ;
        RECT 19.950 591.450 22.050 592.050 ;
        RECT 13.950 590.550 22.050 591.450 ;
        RECT 13.950 589.950 16.050 590.550 ;
        RECT 19.950 589.950 22.050 590.550 ;
        RECT 13.950 588.450 16.050 589.050 ;
        RECT 23.550 588.450 24.450 601.950 ;
        RECT 29.100 600.150 30.900 601.950 ;
        RECT 25.950 596.850 28.050 598.950 ;
        RECT 28.950 598.050 31.050 600.150 ;
        RECT 32.850 598.950 34.050 602.250 ;
        RECT 50.400 600.150 51.600 608.400 ;
        RECT 66.000 605.400 67.800 611.250 ;
        RECT 70.200 607.050 72.000 611.250 ;
        RECT 73.500 608.400 75.300 611.250 ;
        RECT 88.650 608.400 90.450 611.250 ;
        RECT 91.650 608.400 93.450 611.250 ;
        RECT 94.650 608.400 96.450 611.250 ;
        RECT 109.650 608.400 111.450 611.250 ;
        RECT 112.650 608.400 114.450 611.250 ;
        RECT 70.200 605.400 75.900 607.050 ;
        RECT 31.950 596.850 34.050 598.950 ;
        RECT 49.950 598.050 52.050 600.150 ;
        RECT 52.950 599.850 55.050 601.950 ;
        RECT 65.100 600.150 66.900 601.950 ;
        RECT 53.100 598.050 54.900 599.850 ;
        RECT 64.950 598.050 67.050 600.150 ;
        RECT 67.950 599.850 70.050 601.950 ;
        RECT 71.100 600.150 72.900 601.950 ;
        RECT 68.100 598.050 69.900 599.850 ;
        RECT 70.950 598.050 73.050 600.150 ;
        RECT 74.700 598.950 75.900 605.400 ;
        RECT 91.950 601.950 93.000 608.400 ;
        RECT 91.950 599.850 94.050 601.950 ;
        RECT 110.400 600.150 111.600 608.400 ;
        RECT 122.550 606.300 124.350 611.250 ;
        RECT 125.550 607.200 127.350 611.250 ;
        RECT 128.550 606.300 130.350 611.250 ;
        RECT 122.550 604.950 130.350 606.300 ;
        RECT 131.550 605.400 133.350 611.250 ;
        RECT 143.550 608.400 145.350 611.250 ;
        RECT 146.550 608.400 148.350 611.250 ;
        RECT 131.550 603.300 132.750 605.400 ;
        RECT 129.000 602.250 132.750 603.300 ;
        RECT 26.100 595.050 27.900 596.850 ;
        RECT 31.950 591.600 33.150 596.850 ;
        RECT 34.950 593.850 37.050 595.950 ;
        RECT 34.950 592.050 36.750 593.850 ;
        RECT 13.950 587.550 24.450 588.450 ;
        RECT 13.950 586.950 16.050 587.550 ;
        RECT 10.650 579.750 12.450 585.600 ;
        RECT 13.650 579.750 15.450 585.600 ;
        RECT 27.300 579.750 29.100 591.600 ;
        RECT 31.500 579.750 33.300 591.600 ;
        RECT 50.400 585.600 51.600 598.050 ;
        RECT 73.950 596.850 76.050 598.950 ;
        RECT 88.950 596.850 91.050 598.950 ;
        RECT 74.700 591.600 75.900 596.850 ;
        RECT 89.100 595.050 90.900 596.850 ;
        RECT 91.950 592.650 93.000 599.850 ;
        RECT 94.950 596.850 97.050 598.950 ;
        RECT 109.950 598.050 112.050 600.150 ;
        RECT 112.950 599.850 115.050 601.950 ;
        RECT 125.100 600.150 126.900 601.950 ;
        RECT 113.100 598.050 114.900 599.850 ;
        RECT 95.100 595.050 96.900 596.850 ;
        RECT 90.450 591.600 93.000 592.650 ;
        RECT 65.550 590.700 73.350 591.600 ;
        RECT 34.800 579.750 36.600 585.600 ;
        RECT 49.650 579.750 51.450 585.600 ;
        RECT 52.650 579.750 54.450 585.600 ;
        RECT 65.550 579.750 67.350 590.700 ;
        RECT 68.550 579.750 70.350 589.800 ;
        RECT 71.550 579.750 73.350 590.700 ;
        RECT 74.550 579.750 76.350 591.600 ;
        RECT 90.450 579.750 92.250 591.600 ;
        RECT 94.650 579.750 96.450 591.600 ;
        RECT 110.400 585.600 111.600 598.050 ;
        RECT 121.950 596.850 124.050 598.950 ;
        RECT 124.950 598.050 127.050 600.150 ;
        RECT 128.850 598.950 130.050 602.250 ;
        RECT 142.950 599.850 145.050 601.950 ;
        RECT 146.400 600.150 147.600 608.400 ;
        RECT 158.700 602.400 160.500 611.250 ;
        RECT 164.100 603.000 165.900 611.250 ;
        RECT 180.000 605.400 181.800 611.250 ;
        RECT 184.200 605.400 186.000 611.250 ;
        RECT 188.400 605.400 190.200 611.250 ;
        RECT 206.850 605.400 208.650 611.250 ;
        RECT 164.100 601.350 168.600 603.000 ;
        RECT 127.950 596.850 130.050 598.950 ;
        RECT 143.100 598.050 144.900 599.850 ;
        RECT 145.950 598.050 148.050 600.150 ;
        RECT 122.100 595.050 123.900 596.850 ;
        RECT 127.950 591.600 129.150 596.850 ;
        RECT 130.950 593.850 133.050 595.950 ;
        RECT 130.950 592.050 132.750 593.850 ;
        RECT 109.650 579.750 111.450 585.600 ;
        RECT 112.650 579.750 114.450 585.600 ;
        RECT 123.300 579.750 125.100 591.600 ;
        RECT 127.500 579.750 129.300 591.600 ;
        RECT 146.400 585.600 147.600 598.050 ;
        RECT 167.400 597.150 168.600 601.350 ;
        RECT 182.250 600.150 184.050 601.950 ;
        RECT 157.950 593.850 160.050 595.950 ;
        RECT 163.950 593.850 166.050 595.950 ;
        RECT 166.950 595.050 169.050 597.150 ;
        RECT 178.950 596.850 181.050 598.950 ;
        RECT 181.950 598.050 184.050 600.150 ;
        RECT 184.950 598.950 186.000 605.400 ;
        RECT 211.350 604.200 213.150 611.250 ;
        RECT 226.650 608.400 228.450 611.250 ;
        RECT 229.650 608.400 231.450 611.250 ;
        RECT 241.650 608.400 243.450 611.250 ;
        RECT 244.650 608.400 246.450 611.250 ;
        RECT 247.650 608.400 249.450 611.250 ;
        RECT 259.650 608.400 261.450 611.250 ;
        RECT 262.650 608.400 264.450 611.250 ;
        RECT 209.550 603.300 213.150 604.200 ;
        RECT 187.950 600.150 189.750 601.950 ;
        RECT 184.950 596.850 187.050 598.950 ;
        RECT 187.950 598.050 190.050 600.150 ;
        RECT 190.950 596.850 193.050 598.950 ;
        RECT 206.100 597.150 207.900 598.950 ;
        RECT 179.250 595.050 181.050 596.850 ;
        RECT 158.100 592.050 159.900 593.850 ;
        RECT 160.950 590.850 163.050 592.950 ;
        RECT 164.250 592.050 166.050 593.850 ;
        RECT 161.100 589.050 162.900 590.850 ;
        RECT 167.700 586.800 168.750 595.050 ;
        RECT 186.150 593.400 187.050 596.850 ;
        RECT 191.100 595.050 192.900 596.850 ;
        RECT 205.950 595.050 208.050 597.150 ;
        RECT 209.550 595.950 210.750 603.300 ;
        RECT 227.400 600.150 228.600 608.400 ;
        RECT 244.950 601.950 246.000 608.400 ;
        RECT 247.950 606.450 250.050 607.050 ;
        RECT 253.950 606.450 256.050 607.050 ;
        RECT 247.950 605.550 256.050 606.450 ;
        RECT 247.950 604.950 250.050 605.550 ;
        RECT 253.950 604.950 256.050 605.550 ;
        RECT 212.100 597.150 213.900 598.950 ;
        RECT 226.950 598.050 229.050 600.150 ;
        RECT 229.950 599.850 232.050 601.950 ;
        RECT 244.950 599.850 247.050 601.950 ;
        RECT 260.400 600.150 261.600 608.400 ;
        RECT 272.700 602.400 274.500 611.250 ;
        RECT 278.100 603.000 279.900 611.250 ;
        RECT 295.650 605.400 297.450 611.250 ;
        RECT 296.250 603.300 297.450 605.400 ;
        RECT 298.650 606.300 300.450 611.250 ;
        RECT 301.650 607.200 303.450 611.250 ;
        RECT 304.650 606.300 306.450 611.250 ;
        RECT 298.650 604.950 306.450 606.300 ;
        RECT 230.100 598.050 231.900 599.850 ;
        RECT 208.950 593.850 211.050 595.950 ;
        RECT 211.950 595.050 214.050 597.150 ;
        RECT 186.150 592.500 190.200 593.400 ;
        RECT 188.400 591.600 190.200 592.500 ;
        RECT 161.700 585.900 168.750 586.800 ;
        RECT 161.700 585.600 163.350 585.900 ;
        RECT 130.800 579.750 132.600 585.600 ;
        RECT 143.550 579.750 145.350 585.600 ;
        RECT 146.550 579.750 148.350 585.600 ;
        RECT 158.550 579.750 160.350 585.600 ;
        RECT 161.550 579.750 163.350 585.600 ;
        RECT 167.550 585.600 168.750 585.900 ;
        RECT 179.550 590.400 187.350 591.300 ;
        RECT 164.550 579.750 166.350 585.000 ;
        RECT 167.550 579.750 169.350 585.600 ;
        RECT 179.550 579.750 181.350 590.400 ;
        RECT 182.550 579.750 184.350 589.500 ;
        RECT 185.550 580.500 187.350 590.400 ;
        RECT 188.550 581.400 190.350 591.600 ;
        RECT 191.550 580.500 193.350 591.600 ;
        RECT 209.550 585.600 210.750 593.850 ;
        RECT 227.400 585.600 228.600 598.050 ;
        RECT 241.950 596.850 244.050 598.950 ;
        RECT 242.100 595.050 243.900 596.850 ;
        RECT 244.950 592.650 246.000 599.850 ;
        RECT 247.950 596.850 250.050 598.950 ;
        RECT 259.950 598.050 262.050 600.150 ;
        RECT 262.950 599.850 265.050 601.950 ;
        RECT 278.100 601.350 282.600 603.000 ;
        RECT 296.250 602.250 300.000 603.300 ;
        RECT 323.100 603.000 324.900 611.250 ;
        RECT 263.100 598.050 264.900 599.850 ;
        RECT 248.100 595.050 249.900 596.850 ;
        RECT 243.450 591.600 246.000 592.650 ;
        RECT 185.550 579.750 193.350 580.500 ;
        RECT 206.550 579.750 208.350 585.600 ;
        RECT 209.550 579.750 211.350 585.600 ;
        RECT 212.550 579.750 214.350 585.600 ;
        RECT 226.650 579.750 228.450 585.600 ;
        RECT 229.650 579.750 231.450 585.600 ;
        RECT 243.450 579.750 245.250 591.600 ;
        RECT 247.650 579.750 249.450 591.600 ;
        RECT 260.400 585.600 261.600 598.050 ;
        RECT 281.400 597.150 282.600 601.350 ;
        RECT 298.950 598.950 300.150 602.250 ;
        RECT 302.100 600.150 303.900 601.950 ;
        RECT 320.400 601.350 324.900 603.000 ;
        RECT 328.500 602.400 330.300 611.250 ;
        RECT 338.700 602.400 340.500 611.250 ;
        RECT 344.100 603.000 345.900 611.250 ;
        RECT 361.650 605.400 363.450 611.250 ;
        RECT 362.250 603.300 363.450 605.400 ;
        RECT 364.650 606.300 366.450 611.250 ;
        RECT 367.650 607.200 369.450 611.250 ;
        RECT 370.650 606.300 372.450 611.250 ;
        RECT 364.650 604.950 372.450 606.300 ;
        RECT 383.850 604.200 385.650 611.250 ;
        RECT 388.350 605.400 390.150 611.250 ;
        RECT 398.850 605.400 400.650 611.250 ;
        RECT 403.350 604.200 405.150 611.250 ;
        RECT 383.850 603.300 387.450 604.200 ;
        RECT 344.100 601.350 348.600 603.000 ;
        RECT 362.250 602.250 366.000 603.300 ;
        RECT 271.950 593.850 274.050 595.950 ;
        RECT 277.950 593.850 280.050 595.950 ;
        RECT 280.950 595.050 283.050 597.150 ;
        RECT 298.950 596.850 301.050 598.950 ;
        RECT 301.950 598.050 304.050 600.150 ;
        RECT 304.950 596.850 307.050 598.950 ;
        RECT 320.400 597.150 321.600 601.350 ;
        RECT 347.400 597.150 348.600 601.350 ;
        RECT 364.950 598.950 366.150 602.250 ;
        RECT 368.100 600.150 369.900 601.950 ;
        RECT 272.100 592.050 273.900 593.850 ;
        RECT 274.950 590.850 277.050 592.950 ;
        RECT 278.250 592.050 280.050 593.850 ;
        RECT 275.100 589.050 276.900 590.850 ;
        RECT 281.700 586.800 282.750 595.050 ;
        RECT 295.950 593.850 298.050 595.950 ;
        RECT 296.250 592.050 298.050 593.850 ;
        RECT 299.850 591.600 301.050 596.850 ;
        RECT 305.100 595.050 306.900 596.850 ;
        RECT 319.950 595.050 322.050 597.150 ;
        RECT 275.700 585.900 282.750 586.800 ;
        RECT 275.700 585.600 277.350 585.900 ;
        RECT 259.650 579.750 261.450 585.600 ;
        RECT 262.650 579.750 264.450 585.600 ;
        RECT 272.550 579.750 274.350 585.600 ;
        RECT 275.550 579.750 277.350 585.600 ;
        RECT 281.550 585.600 282.750 585.900 ;
        RECT 278.550 579.750 280.350 585.000 ;
        RECT 281.550 579.750 283.350 585.600 ;
        RECT 296.400 579.750 298.200 585.600 ;
        RECT 299.700 579.750 301.500 591.600 ;
        RECT 303.900 579.750 305.700 591.600 ;
        RECT 320.250 586.800 321.300 595.050 ;
        RECT 322.950 593.850 325.050 595.950 ;
        RECT 328.950 593.850 331.050 595.950 ;
        RECT 337.950 593.850 340.050 595.950 ;
        RECT 343.950 593.850 346.050 595.950 ;
        RECT 346.950 595.050 349.050 597.150 ;
        RECT 364.950 596.850 367.050 598.950 ;
        RECT 367.950 598.050 370.050 600.150 ;
        RECT 370.950 596.850 373.050 598.950 ;
        RECT 383.100 597.150 384.900 598.950 ;
        RECT 322.950 592.050 324.750 593.850 ;
        RECT 325.950 590.850 328.050 592.950 ;
        RECT 329.100 592.050 330.900 593.850 ;
        RECT 338.100 592.050 339.900 593.850 ;
        RECT 340.950 590.850 343.050 592.950 ;
        RECT 344.250 592.050 346.050 593.850 ;
        RECT 326.100 589.050 327.900 590.850 ;
        RECT 341.100 589.050 342.900 590.850 ;
        RECT 347.700 586.800 348.750 595.050 ;
        RECT 361.950 593.850 364.050 595.950 ;
        RECT 362.250 592.050 364.050 593.850 ;
        RECT 365.850 591.600 367.050 596.850 ;
        RECT 371.100 595.050 372.900 596.850 ;
        RECT 382.950 595.050 385.050 597.150 ;
        RECT 386.250 595.950 387.450 603.300 ;
        RECT 388.950 603.450 391.050 604.050 ;
        RECT 388.950 602.550 393.450 603.450 ;
        RECT 388.950 601.950 391.050 602.550 ;
        RECT 389.100 597.150 390.900 598.950 ;
        RECT 385.950 593.850 388.050 595.950 ;
        RECT 388.950 595.050 391.050 597.150 ;
        RECT 392.550 595.050 393.450 602.550 ;
        RECT 401.550 603.300 405.150 604.200 ;
        RECT 394.950 595.950 397.050 598.050 ;
        RECT 398.100 597.150 399.900 598.950 ;
        RECT 320.250 585.900 327.300 586.800 ;
        RECT 320.250 585.600 321.450 585.900 ;
        RECT 319.650 579.750 321.450 585.600 ;
        RECT 325.650 585.600 327.300 585.900 ;
        RECT 341.700 585.900 348.750 586.800 ;
        RECT 341.700 585.600 343.350 585.900 ;
        RECT 322.650 579.750 324.450 585.000 ;
        RECT 325.650 579.750 327.450 585.600 ;
        RECT 328.650 579.750 330.450 585.600 ;
        RECT 338.550 579.750 340.350 585.600 ;
        RECT 341.550 579.750 343.350 585.600 ;
        RECT 347.550 585.600 348.750 585.900 ;
        RECT 344.550 579.750 346.350 585.000 ;
        RECT 347.550 579.750 349.350 585.600 ;
        RECT 362.400 579.750 364.200 585.600 ;
        RECT 365.700 579.750 367.500 591.600 ;
        RECT 369.900 579.750 371.700 591.600 ;
        RECT 386.250 585.600 387.450 593.850 ;
        RECT 391.950 592.950 394.050 595.050 ;
        RECT 388.950 591.450 391.050 592.050 ;
        RECT 395.550 591.450 396.450 595.950 ;
        RECT 397.950 595.050 400.050 597.150 ;
        RECT 401.550 595.950 402.750 603.300 ;
        RECT 416.700 602.400 418.500 611.250 ;
        RECT 422.100 603.000 423.900 611.250 ;
        RECT 422.100 601.350 426.600 603.000 ;
        RECT 437.700 602.400 439.500 611.250 ;
        RECT 443.100 603.000 444.900 611.250 ;
        RECT 460.650 608.400 462.450 611.250 ;
        RECT 463.650 608.400 465.450 611.250 ;
        RECT 443.100 601.350 447.600 603.000 ;
        RECT 404.100 597.150 405.900 598.950 ;
        RECT 425.400 597.150 426.600 601.350 ;
        RECT 446.400 597.150 447.600 601.350 ;
        RECT 461.400 600.150 462.600 608.400 ;
        RECT 479.100 603.000 480.900 611.250 ;
        RECT 460.950 598.050 463.050 600.150 ;
        RECT 463.950 599.850 466.050 601.950 ;
        RECT 476.400 601.350 480.900 603.000 ;
        RECT 484.500 602.400 486.300 611.250 ;
        RECT 496.650 608.400 498.450 611.250 ;
        RECT 499.650 608.400 501.450 611.250 ;
        RECT 464.100 598.050 465.900 599.850 ;
        RECT 400.950 593.850 403.050 595.950 ;
        RECT 403.950 595.050 406.050 597.150 ;
        RECT 415.950 593.850 418.050 595.950 ;
        RECT 421.950 593.850 424.050 595.950 ;
        RECT 424.950 595.050 427.050 597.150 ;
        RECT 388.950 590.550 396.450 591.450 ;
        RECT 388.950 589.950 391.050 590.550 ;
        RECT 401.550 585.600 402.750 593.850 ;
        RECT 416.100 592.050 417.900 593.850 ;
        RECT 418.950 590.850 421.050 592.950 ;
        RECT 422.250 592.050 424.050 593.850 ;
        RECT 419.100 589.050 420.900 590.850 ;
        RECT 425.700 586.800 426.750 595.050 ;
        RECT 436.950 593.850 439.050 595.950 ;
        RECT 442.950 593.850 445.050 595.950 ;
        RECT 445.950 595.050 448.050 597.150 ;
        RECT 437.100 592.050 438.900 593.850 ;
        RECT 439.950 590.850 442.050 592.950 ;
        RECT 443.250 592.050 445.050 593.850 ;
        RECT 440.100 589.050 441.900 590.850 ;
        RECT 446.700 586.800 447.750 595.050 ;
        RECT 419.700 585.900 426.750 586.800 ;
        RECT 419.700 585.600 421.350 585.900 ;
        RECT 382.650 579.750 384.450 585.600 ;
        RECT 385.650 579.750 387.450 585.600 ;
        RECT 388.650 579.750 390.450 585.600 ;
        RECT 398.550 579.750 400.350 585.600 ;
        RECT 401.550 579.750 403.350 585.600 ;
        RECT 404.550 579.750 406.350 585.600 ;
        RECT 416.550 579.750 418.350 585.600 ;
        RECT 419.550 579.750 421.350 585.600 ;
        RECT 425.550 585.600 426.750 585.900 ;
        RECT 440.700 585.900 447.750 586.800 ;
        RECT 440.700 585.600 442.350 585.900 ;
        RECT 422.550 579.750 424.350 585.000 ;
        RECT 425.550 579.750 427.350 585.600 ;
        RECT 437.550 579.750 439.350 585.600 ;
        RECT 440.550 579.750 442.350 585.600 ;
        RECT 446.550 585.600 447.750 585.900 ;
        RECT 461.400 585.600 462.600 598.050 ;
        RECT 476.400 597.150 477.600 601.350 ;
        RECT 497.400 600.150 498.600 608.400 ;
        RECT 511.650 605.400 513.450 611.250 ;
        RECT 512.250 603.300 513.450 605.400 ;
        RECT 514.650 606.300 516.450 611.250 ;
        RECT 517.650 607.200 519.450 611.250 ;
        RECT 520.650 606.300 522.450 611.250 ;
        RECT 514.650 604.950 522.450 606.300 ;
        RECT 530.850 605.400 532.650 611.250 ;
        RECT 535.350 604.200 537.150 611.250 ;
        RECT 550.650 605.400 552.450 611.250 ;
        RECT 553.650 608.400 555.450 611.250 ;
        RECT 556.650 608.400 558.450 611.250 ;
        RECT 559.650 608.400 561.450 611.250 ;
        RECT 533.550 603.300 537.150 604.200 ;
        RECT 512.250 602.250 516.000 603.300 ;
        RECT 496.950 598.050 499.050 600.150 ;
        RECT 499.950 599.850 502.050 601.950 ;
        RECT 500.100 598.050 501.900 599.850 ;
        RECT 514.950 598.950 516.150 602.250 ;
        RECT 518.100 600.150 519.900 601.950 ;
        RECT 475.950 595.050 478.050 597.150 ;
        RECT 476.250 586.800 477.300 595.050 ;
        RECT 478.950 593.850 481.050 595.950 ;
        RECT 484.950 593.850 487.050 595.950 ;
        RECT 478.950 592.050 480.750 593.850 ;
        RECT 481.950 590.850 484.050 592.950 ;
        RECT 485.100 592.050 486.900 593.850 ;
        RECT 482.100 589.050 483.900 590.850 ;
        RECT 476.250 585.900 483.300 586.800 ;
        RECT 476.250 585.600 477.450 585.900 ;
        RECT 443.550 579.750 445.350 585.000 ;
        RECT 446.550 579.750 448.350 585.600 ;
        RECT 460.650 579.750 462.450 585.600 ;
        RECT 463.650 579.750 465.450 585.600 ;
        RECT 475.650 579.750 477.450 585.600 ;
        RECT 481.650 585.600 483.300 585.900 ;
        RECT 497.400 585.600 498.600 598.050 ;
        RECT 514.950 596.850 517.050 598.950 ;
        RECT 517.950 598.050 520.050 600.150 ;
        RECT 520.950 596.850 523.050 598.950 ;
        RECT 530.100 597.150 531.900 598.950 ;
        RECT 511.950 593.850 514.050 595.950 ;
        RECT 512.250 592.050 514.050 593.850 ;
        RECT 515.850 591.600 517.050 596.850 ;
        RECT 521.100 595.050 522.900 596.850 ;
        RECT 529.950 595.050 532.050 597.150 ;
        RECT 533.550 595.950 534.750 603.300 ;
        RECT 550.950 600.150 552.000 605.400 ;
        RECT 556.650 604.200 557.550 608.400 ;
        RECT 572.850 605.400 574.650 611.250 ;
        RECT 577.350 604.200 579.150 611.250 ;
        RECT 592.650 605.400 594.450 611.250 ;
        RECT 554.250 603.300 557.550 604.200 ;
        RECT 575.550 603.300 579.150 604.200 ;
        RECT 593.250 603.300 594.450 605.400 ;
        RECT 595.650 606.300 597.450 611.250 ;
        RECT 598.650 607.200 600.450 611.250 ;
        RECT 601.650 606.300 603.450 611.250 ;
        RECT 614.700 608.400 616.500 611.250 ;
        RECT 618.000 607.050 619.800 611.250 ;
        RECT 595.650 604.950 603.450 606.300 ;
        RECT 614.100 605.400 619.800 607.050 ;
        RECT 622.200 605.400 624.000 611.250 ;
        RECT 632.850 605.400 634.650 611.250 ;
        RECT 554.250 602.400 556.050 603.300 ;
        RECT 536.100 597.150 537.900 598.950 ;
        RECT 550.950 598.050 553.050 600.150 ;
        RECT 532.950 593.850 535.050 595.950 ;
        RECT 535.950 595.050 538.050 597.150 ;
        RECT 478.650 579.750 480.450 585.000 ;
        RECT 481.650 579.750 483.450 585.600 ;
        RECT 484.650 579.750 486.450 585.600 ;
        RECT 496.650 579.750 498.450 585.600 ;
        RECT 499.650 579.750 501.450 585.600 ;
        RECT 512.400 579.750 514.200 585.600 ;
        RECT 515.700 579.750 517.500 591.600 ;
        RECT 519.900 579.750 521.700 591.600 ;
        RECT 533.550 585.600 534.750 593.850 ;
        RECT 551.550 591.450 552.900 598.050 ;
        RECT 554.400 594.150 555.300 602.400 ;
        RECT 559.950 599.850 562.050 601.950 ;
        RECT 556.950 596.850 559.050 598.950 ;
        RECT 560.100 598.050 561.900 599.850 ;
        RECT 572.100 597.150 573.900 598.950 ;
        RECT 557.100 595.050 558.900 596.850 ;
        RECT 571.950 595.050 574.050 597.150 ;
        RECT 575.550 595.950 576.750 603.300 ;
        RECT 593.250 602.250 597.000 603.300 ;
        RECT 595.950 598.950 597.150 602.250 ;
        RECT 599.100 600.150 600.900 601.950 ;
        RECT 578.100 597.150 579.900 598.950 ;
        RECT 554.250 594.000 556.050 594.150 ;
        RECT 554.250 592.800 561.450 594.000 ;
        RECT 574.950 593.850 577.050 595.950 ;
        RECT 577.950 595.050 580.050 597.150 ;
        RECT 595.950 596.850 598.050 598.950 ;
        RECT 598.950 598.050 601.050 600.150 ;
        RECT 614.100 598.950 615.300 605.400 ;
        RECT 637.350 604.200 639.150 611.250 ;
        RECT 650.550 606.300 652.350 611.250 ;
        RECT 653.550 607.200 655.350 611.250 ;
        RECT 656.550 606.300 658.350 611.250 ;
        RECT 650.550 604.950 658.350 606.300 ;
        RECT 659.550 605.400 661.350 611.250 ;
        RECT 671.550 606.300 673.350 611.250 ;
        RECT 674.550 607.200 676.350 611.250 ;
        RECT 677.550 606.300 679.350 611.250 ;
        RECT 635.550 603.300 639.150 604.200 ;
        RECT 659.550 603.300 660.750 605.400 ;
        RECT 671.550 604.950 679.350 606.300 ;
        RECT 680.550 605.400 682.350 611.250 ;
        RECT 692.550 608.400 694.350 611.250 ;
        RECT 695.550 608.400 697.350 611.250 ;
        RECT 698.550 608.400 700.350 611.250 ;
        RECT 680.550 603.300 681.750 605.400 ;
        RECT 696.450 604.200 697.350 608.400 ;
        RECT 701.550 605.400 703.350 611.250 ;
        RECT 696.450 603.300 699.750 604.200 ;
        RECT 617.100 600.150 618.900 601.950 ;
        RECT 601.950 596.850 604.050 598.950 ;
        RECT 613.950 596.850 616.050 598.950 ;
        RECT 616.950 598.050 619.050 600.150 ;
        RECT 619.950 599.850 622.050 601.950 ;
        RECT 623.100 600.150 624.900 601.950 ;
        RECT 620.100 598.050 621.900 599.850 ;
        RECT 622.950 598.050 625.050 600.150 ;
        RECT 632.100 597.150 633.900 598.950 ;
        RECT 592.950 593.850 595.050 595.950 ;
        RECT 554.250 592.350 556.050 592.800 ;
        RECT 560.250 591.600 561.450 592.800 ;
        RECT 551.550 590.100 553.950 591.450 ;
        RECT 530.550 579.750 532.350 585.600 ;
        RECT 533.550 579.750 535.350 585.600 ;
        RECT 536.550 579.750 538.350 585.600 ;
        RECT 552.150 579.750 553.950 590.100 ;
        RECT 555.150 579.750 556.950 591.450 ;
        RECT 559.650 579.750 561.450 591.600 ;
        RECT 575.550 585.600 576.750 593.850 ;
        RECT 593.250 592.050 595.050 593.850 ;
        RECT 596.850 591.600 598.050 596.850 ;
        RECT 602.100 595.050 603.900 596.850 ;
        RECT 614.100 591.600 615.300 596.850 ;
        RECT 631.950 595.050 634.050 597.150 ;
        RECT 635.550 595.950 636.750 603.300 ;
        RECT 657.000 602.250 660.750 603.300 ;
        RECT 678.000 602.250 681.750 603.300 ;
        RECT 697.950 602.400 699.750 603.300 ;
        RECT 653.100 600.150 654.900 601.950 ;
        RECT 638.100 597.150 639.900 598.950 ;
        RECT 634.950 593.850 637.050 595.950 ;
        RECT 637.950 595.050 640.050 597.150 ;
        RECT 649.950 596.850 652.050 598.950 ;
        RECT 652.950 598.050 655.050 600.150 ;
        RECT 656.850 598.950 658.050 602.250 ;
        RECT 674.100 600.150 675.900 601.950 ;
        RECT 655.950 596.850 658.050 598.950 ;
        RECT 670.950 596.850 673.050 598.950 ;
        RECT 673.950 598.050 676.050 600.150 ;
        RECT 677.850 598.950 679.050 602.250 ;
        RECT 691.950 599.850 694.050 601.950 ;
        RECT 676.950 596.850 679.050 598.950 ;
        RECT 692.100 598.050 693.900 599.850 ;
        RECT 694.950 596.850 697.050 598.950 ;
        RECT 650.100 595.050 651.900 596.850 ;
        RECT 572.550 579.750 574.350 585.600 ;
        RECT 575.550 579.750 577.350 585.600 ;
        RECT 578.550 579.750 580.350 585.600 ;
        RECT 593.400 579.750 595.200 585.600 ;
        RECT 596.700 579.750 598.500 591.600 ;
        RECT 600.900 579.750 602.700 591.600 ;
        RECT 613.650 579.750 615.450 591.600 ;
        RECT 616.650 590.700 624.450 591.600 ;
        RECT 616.650 579.750 618.450 590.700 ;
        RECT 619.650 579.750 621.450 589.800 ;
        RECT 622.650 579.750 624.450 590.700 ;
        RECT 635.550 585.600 636.750 593.850 ;
        RECT 655.950 591.600 657.150 596.850 ;
        RECT 658.950 593.850 661.050 595.950 ;
        RECT 671.100 595.050 672.900 596.850 ;
        RECT 658.950 592.050 660.750 593.850 ;
        RECT 676.950 591.600 678.150 596.850 ;
        RECT 679.950 593.850 682.050 595.950 ;
        RECT 695.100 595.050 696.900 596.850 ;
        RECT 698.700 594.150 699.600 602.400 ;
        RECT 702.000 600.150 703.050 605.400 ;
        RECT 716.850 604.200 718.650 611.250 ;
        RECT 721.350 605.400 723.150 611.250 ;
        RECT 716.850 603.300 720.450 604.200 ;
        RECT 700.950 598.050 703.050 600.150 ;
        RECT 697.950 594.000 699.750 594.150 ;
        RECT 679.950 592.050 681.750 593.850 ;
        RECT 692.550 592.800 699.750 594.000 ;
        RECT 692.550 591.600 693.750 592.800 ;
        RECT 697.950 592.350 699.750 592.800 ;
        RECT 632.550 579.750 634.350 585.600 ;
        RECT 635.550 579.750 637.350 585.600 ;
        RECT 638.550 579.750 640.350 585.600 ;
        RECT 651.300 579.750 653.100 591.600 ;
        RECT 655.500 579.750 657.300 591.600 ;
        RECT 658.800 579.750 660.600 585.600 ;
        RECT 672.300 579.750 674.100 591.600 ;
        RECT 676.500 579.750 678.300 591.600 ;
        RECT 679.800 579.750 681.600 585.600 ;
        RECT 692.550 579.750 694.350 591.600 ;
        RECT 701.100 591.450 702.450 598.050 ;
        RECT 716.100 597.150 717.900 598.950 ;
        RECT 715.950 595.050 718.050 597.150 ;
        RECT 719.250 595.950 720.450 603.300 ;
        RECT 731.700 602.400 733.500 611.250 ;
        RECT 737.100 603.000 738.900 611.250 ;
        RECT 752.550 608.400 754.350 611.250 ;
        RECT 755.550 608.400 757.350 611.250 ;
        RECT 769.650 608.400 771.450 611.250 ;
        RECT 772.650 608.400 774.450 611.250 ;
        RECT 737.100 601.350 741.600 603.000 ;
        RECT 722.100 597.150 723.900 598.950 ;
        RECT 740.400 597.150 741.600 601.350 ;
        RECT 751.950 599.850 754.050 601.950 ;
        RECT 755.400 600.150 756.600 608.400 ;
        RECT 770.400 600.150 771.600 608.400 ;
        RECT 776.550 605.400 778.350 611.250 ;
        RECT 779.850 608.400 781.650 611.250 ;
        RECT 784.350 608.400 786.150 611.250 ;
        RECT 788.550 608.400 790.350 611.250 ;
        RECT 792.450 608.400 794.250 611.250 ;
        RECT 795.750 608.400 797.550 611.250 ;
        RECT 800.250 609.300 802.050 611.250 ;
        RECT 800.250 608.400 804.000 609.300 ;
        RECT 805.050 608.400 806.850 611.250 ;
        RECT 784.650 607.500 785.700 608.400 ;
        RECT 781.950 606.300 785.700 607.500 ;
        RECT 793.200 606.600 794.250 608.400 ;
        RECT 802.950 607.500 804.000 608.400 ;
        RECT 781.950 605.400 784.050 606.300 ;
        RECT 776.550 603.150 777.750 605.400 ;
        RECT 789.150 604.200 790.950 606.000 ;
        RECT 793.200 605.550 798.150 606.600 ;
        RECT 796.350 604.800 798.150 605.550 ;
        RECT 799.650 604.800 801.450 606.600 ;
        RECT 802.950 605.400 805.050 607.500 ;
        RECT 808.050 605.400 809.850 611.250 ;
        RECT 790.050 603.900 790.950 604.200 ;
        RECT 800.100 603.900 801.150 604.800 ;
        RECT 752.100 598.050 753.900 599.850 ;
        RECT 754.950 598.050 757.050 600.150 ;
        RECT 769.950 598.050 772.050 600.150 ;
        RECT 772.950 599.850 775.050 601.950 ;
        RECT 776.550 601.050 781.050 603.150 ;
        RECT 790.050 603.000 801.150 603.900 ;
        RECT 773.100 598.050 774.900 599.850 ;
        RECT 718.950 593.850 721.050 595.950 ;
        RECT 721.950 595.050 724.050 597.150 ;
        RECT 730.950 593.850 733.050 595.950 ;
        RECT 736.950 593.850 739.050 595.950 ;
        RECT 739.950 595.050 742.050 597.150 ;
        RECT 697.050 579.750 698.850 591.450 ;
        RECT 700.050 590.100 702.450 591.450 ;
        RECT 700.050 579.750 701.850 590.100 ;
        RECT 719.250 585.600 720.450 593.850 ;
        RECT 731.100 592.050 732.900 593.850 ;
        RECT 733.950 590.850 736.050 592.950 ;
        RECT 737.250 592.050 739.050 593.850 ;
        RECT 734.100 589.050 735.900 590.850 ;
        RECT 740.700 586.800 741.750 595.050 ;
        RECT 734.700 585.900 741.750 586.800 ;
        RECT 734.700 585.600 736.350 585.900 ;
        RECT 715.650 579.750 717.450 585.600 ;
        RECT 718.650 579.750 720.450 585.600 ;
        RECT 721.650 579.750 723.450 585.600 ;
        RECT 731.550 579.750 733.350 585.600 ;
        RECT 734.550 579.750 736.350 585.600 ;
        RECT 740.550 585.600 741.750 585.900 ;
        RECT 755.400 585.600 756.600 598.050 ;
        RECT 770.400 585.600 771.600 598.050 ;
        RECT 776.550 591.600 777.750 601.050 ;
        RECT 778.950 599.250 782.850 601.050 ;
        RECT 778.950 598.950 781.050 599.250 ;
        RECT 790.050 598.950 790.950 603.000 ;
        RECT 800.100 601.800 801.150 603.000 ;
        RECT 800.100 600.600 807.000 601.800 ;
        RECT 800.100 600.000 801.900 600.600 ;
        RECT 806.100 599.850 807.000 600.600 ;
        RECT 803.100 598.950 804.900 599.700 ;
        RECT 790.050 596.850 793.050 598.950 ;
        RECT 796.950 597.900 804.900 598.950 ;
        RECT 806.100 598.050 807.900 599.850 ;
        RECT 796.950 596.850 799.050 597.900 ;
        RECT 778.950 593.400 780.750 595.200 ;
        RECT 779.850 592.200 784.050 593.400 ;
        RECT 790.050 592.200 790.950 596.850 ;
        RECT 798.750 593.100 800.550 593.400 ;
        RECT 737.550 579.750 739.350 585.000 ;
        RECT 740.550 579.750 742.350 585.600 ;
        RECT 752.550 579.750 754.350 585.600 ;
        RECT 755.550 579.750 757.350 585.600 ;
        RECT 769.650 579.750 771.450 585.600 ;
        RECT 772.650 579.750 774.450 585.600 ;
        RECT 776.550 579.750 778.350 591.600 ;
        RECT 781.950 591.300 784.050 592.200 ;
        RECT 784.950 591.300 790.950 592.200 ;
        RECT 792.150 592.800 800.550 593.100 ;
        RECT 808.950 592.800 809.850 605.400 ;
        RECT 792.150 592.200 809.850 592.800 ;
        RECT 784.950 590.400 785.850 591.300 ;
        RECT 783.150 588.600 785.850 590.400 ;
        RECT 786.750 590.100 788.550 590.400 ;
        RECT 792.150 590.100 793.050 592.200 ;
        RECT 798.750 591.600 809.850 592.200 ;
        RECT 786.750 589.200 793.050 590.100 ;
        RECT 793.950 590.700 795.750 591.300 ;
        RECT 793.950 589.500 801.450 590.700 ;
        RECT 786.750 588.600 788.550 589.200 ;
        RECT 800.250 588.600 801.450 589.500 ;
        RECT 781.950 585.600 785.850 587.700 ;
        RECT 790.950 586.500 797.850 588.300 ;
        RECT 800.250 586.500 805.050 588.600 ;
        RECT 779.550 579.750 781.350 582.600 ;
        RECT 784.050 579.750 785.850 585.600 ;
        RECT 788.250 579.750 790.050 585.600 ;
        RECT 792.150 579.750 793.950 586.500 ;
        RECT 800.250 585.600 801.450 586.500 ;
        RECT 795.150 579.750 796.950 585.600 ;
        RECT 799.950 579.750 801.750 585.600 ;
        RECT 805.050 579.750 806.850 585.600 ;
        RECT 808.050 579.750 809.850 591.600 ;
        RECT 812.550 605.400 814.350 611.250 ;
        RECT 815.850 608.400 817.650 611.250 ;
        RECT 820.350 608.400 822.150 611.250 ;
        RECT 824.550 608.400 826.350 611.250 ;
        RECT 828.450 608.400 830.250 611.250 ;
        RECT 831.750 608.400 833.550 611.250 ;
        RECT 836.250 609.300 838.050 611.250 ;
        RECT 836.250 608.400 840.000 609.300 ;
        RECT 841.050 608.400 842.850 611.250 ;
        RECT 820.650 607.500 821.700 608.400 ;
        RECT 817.950 606.300 821.700 607.500 ;
        RECT 829.200 606.600 830.250 608.400 ;
        RECT 838.950 607.500 840.000 608.400 ;
        RECT 817.950 605.400 820.050 606.300 ;
        RECT 812.550 603.150 813.750 605.400 ;
        RECT 825.150 604.200 826.950 606.000 ;
        RECT 829.200 605.550 834.150 606.600 ;
        RECT 832.350 604.800 834.150 605.550 ;
        RECT 835.650 604.800 837.450 606.600 ;
        RECT 838.950 605.400 841.050 607.500 ;
        RECT 844.050 605.400 845.850 611.250 ;
        RECT 826.050 603.900 826.950 604.200 ;
        RECT 836.100 603.900 837.150 604.800 ;
        RECT 812.550 601.050 817.050 603.150 ;
        RECT 826.050 603.000 837.150 603.900 ;
        RECT 812.550 591.600 813.750 601.050 ;
        RECT 814.950 599.250 818.850 601.050 ;
        RECT 814.950 598.950 817.050 599.250 ;
        RECT 826.050 598.950 826.950 603.000 ;
        RECT 836.100 601.800 837.150 603.000 ;
        RECT 836.100 600.600 843.000 601.800 ;
        RECT 836.100 600.000 837.900 600.600 ;
        RECT 842.100 599.850 843.000 600.600 ;
        RECT 839.100 598.950 840.900 599.700 ;
        RECT 826.050 596.850 829.050 598.950 ;
        RECT 832.950 597.900 840.900 598.950 ;
        RECT 842.100 598.050 843.900 599.850 ;
        RECT 832.950 596.850 835.050 597.900 ;
        RECT 814.950 593.400 816.750 595.200 ;
        RECT 815.850 592.200 820.050 593.400 ;
        RECT 826.050 592.200 826.950 596.850 ;
        RECT 834.750 593.100 836.550 593.400 ;
        RECT 812.550 579.750 814.350 591.600 ;
        RECT 817.950 591.300 820.050 592.200 ;
        RECT 820.950 591.300 826.950 592.200 ;
        RECT 828.150 592.800 836.550 593.100 ;
        RECT 844.950 592.800 845.850 605.400 ;
        RECT 854.550 606.300 856.350 611.250 ;
        RECT 857.550 607.200 859.350 611.250 ;
        RECT 860.550 606.300 862.350 611.250 ;
        RECT 854.550 604.950 862.350 606.300 ;
        RECT 863.550 605.400 865.350 611.250 ;
        RECT 863.550 603.300 864.750 605.400 ;
        RECT 861.000 602.250 864.750 603.300 ;
        RECT 857.100 600.150 858.900 601.950 ;
        RECT 853.950 596.850 856.050 598.950 ;
        RECT 856.950 598.050 859.050 600.150 ;
        RECT 860.850 598.950 862.050 602.250 ;
        RECT 859.950 596.850 862.050 598.950 ;
        RECT 854.100 595.050 855.900 596.850 ;
        RECT 828.150 592.200 845.850 592.800 ;
        RECT 820.950 590.400 821.850 591.300 ;
        RECT 819.150 588.600 821.850 590.400 ;
        RECT 822.750 590.100 824.550 590.400 ;
        RECT 828.150 590.100 829.050 592.200 ;
        RECT 834.750 591.600 845.850 592.200 ;
        RECT 859.950 591.600 861.150 596.850 ;
        RECT 862.950 593.850 865.050 595.950 ;
        RECT 862.950 592.050 864.750 593.850 ;
        RECT 822.750 589.200 829.050 590.100 ;
        RECT 829.950 590.700 831.750 591.300 ;
        RECT 829.950 589.500 837.450 590.700 ;
        RECT 822.750 588.600 824.550 589.200 ;
        RECT 836.250 588.600 837.450 589.500 ;
        RECT 817.950 585.600 821.850 587.700 ;
        RECT 826.950 586.500 833.850 588.300 ;
        RECT 836.250 586.500 841.050 588.600 ;
        RECT 815.550 579.750 817.350 582.600 ;
        RECT 820.050 579.750 821.850 585.600 ;
        RECT 824.250 579.750 826.050 585.600 ;
        RECT 828.150 579.750 829.950 586.500 ;
        RECT 836.250 585.600 837.450 586.500 ;
        RECT 831.150 579.750 832.950 585.600 ;
        RECT 835.950 579.750 837.750 585.600 ;
        RECT 841.050 579.750 842.850 585.600 ;
        RECT 844.050 579.750 845.850 591.600 ;
        RECT 855.300 579.750 857.100 591.600 ;
        RECT 859.500 579.750 861.300 591.600 ;
        RECT 862.800 579.750 864.600 585.600 ;
        RECT 10.650 569.400 12.450 575.250 ;
        RECT 13.650 569.400 15.450 575.250 ;
        RECT 16.650 569.400 18.450 575.250 ;
        RECT 28.650 569.400 30.450 575.250 ;
        RECT 31.650 570.000 33.450 575.250 ;
        RECT 14.250 561.150 15.450 569.400 ;
        RECT 29.250 569.100 30.450 569.400 ;
        RECT 34.650 569.400 36.450 575.250 ;
        RECT 37.650 569.400 39.450 575.250 ;
        RECT 49.050 574.500 56.850 575.250 ;
        RECT 34.650 569.100 36.300 569.400 ;
        RECT 29.250 568.200 36.300 569.100 ;
        RECT 10.950 557.850 13.050 559.950 ;
        RECT 13.950 559.050 16.050 561.150 ;
        RECT 29.250 559.950 30.300 568.200 ;
        RECT 35.100 564.150 36.900 565.950 ;
        RECT 49.050 565.200 50.850 574.500 ;
        RECT 52.050 565.800 53.850 573.600 ;
        RECT 31.950 561.150 33.750 562.950 ;
        RECT 34.950 562.050 37.050 564.150 ;
        RECT 52.650 563.400 53.850 565.800 ;
        RECT 55.050 565.800 56.850 574.500 ;
        RECT 58.650 574.500 66.450 575.250 ;
        RECT 58.650 566.700 60.450 574.500 ;
        RECT 61.650 565.800 63.450 573.600 ;
        RECT 55.050 564.900 63.450 565.800 ;
        RECT 64.650 565.500 66.450 574.500 ;
        RECT 67.650 566.400 69.450 575.250 ;
        RECT 70.650 565.500 72.450 575.250 ;
        RECT 83.400 569.400 85.200 575.250 ;
        RECT 64.650 564.600 72.450 565.500 ;
        RECT 86.700 563.400 88.500 575.250 ;
        RECT 90.900 563.400 92.700 575.250 ;
        RECT 103.650 569.400 105.450 575.250 ;
        RECT 106.650 569.400 108.450 575.250 ;
        RECT 109.650 569.400 111.450 575.250 ;
        RECT 38.100 561.150 39.900 562.950 ;
        RECT 52.650 562.200 56.100 563.400 ;
        RECT 11.100 556.050 12.900 557.850 ;
        RECT 14.250 551.700 15.450 559.050 ;
        RECT 16.950 557.850 19.050 559.950 ;
        RECT 28.950 557.850 31.050 559.950 ;
        RECT 31.950 559.050 34.050 561.150 ;
        RECT 37.950 559.050 40.050 561.150 ;
        RECT 17.100 556.050 18.900 557.850 ;
        RECT 29.400 553.650 30.600 557.850 ;
        RECT 54.900 556.950 56.100 562.200 ;
        RECT 83.250 561.150 85.050 562.950 ;
        RECT 59.100 558.150 60.900 559.950 ;
        RECT 68.100 558.150 69.900 559.950 ;
        RECT 82.950 559.050 85.050 561.150 ;
        RECT 86.850 558.150 88.050 563.400 ;
        RECT 107.250 561.150 108.450 569.400 ;
        RECT 120.300 563.400 122.100 575.250 ;
        RECT 124.500 563.400 126.300 575.250 ;
        RECT 127.800 569.400 129.600 575.250 ;
        RECT 145.650 574.500 153.450 575.250 ;
        RECT 145.650 563.400 147.450 574.500 ;
        RECT 148.650 563.400 150.450 573.600 ;
        RECT 151.650 564.600 153.450 574.500 ;
        RECT 154.650 565.500 156.450 575.250 ;
        RECT 157.650 564.600 159.450 575.250 ;
        RECT 167.550 569.400 169.350 575.250 ;
        RECT 170.550 569.400 172.350 575.250 ;
        RECT 173.550 569.400 175.350 575.250 ;
        RECT 185.550 569.400 187.350 575.250 ;
        RECT 188.550 569.400 190.350 575.250 ;
        RECT 191.550 570.000 193.350 575.250 ;
        RECT 151.650 563.700 159.450 564.600 ;
        RECT 92.100 558.150 93.900 559.950 ;
        RECT 52.950 554.850 56.100 556.950 ;
        RECT 58.950 556.050 61.050 558.150 ;
        RECT 61.950 554.850 64.050 556.950 ;
        RECT 67.950 556.050 70.050 558.150 ;
        RECT 85.950 556.050 88.050 558.150 ;
        RECT 29.400 552.000 33.900 553.650 ;
        RECT 11.850 550.800 15.450 551.700 ;
        RECT 11.850 543.750 13.650 550.800 ;
        RECT 16.350 543.750 18.150 549.600 ;
        RECT 32.100 543.750 33.900 552.000 ;
        RECT 37.500 543.750 39.300 552.600 ;
        RECT 54.900 548.400 56.100 554.850 ;
        RECT 62.100 553.050 63.900 554.850 ;
        RECT 85.950 552.750 87.150 556.050 ;
        RECT 88.950 554.850 91.050 556.950 ;
        RECT 91.950 556.050 94.050 558.150 ;
        RECT 103.950 557.850 106.050 559.950 ;
        RECT 106.950 559.050 109.050 561.150 ;
        RECT 104.100 556.050 105.900 557.850 ;
        RECT 89.100 553.050 90.900 554.850 ;
        RECT 83.250 551.700 87.000 552.750 ;
        RECT 107.250 551.700 108.450 559.050 ;
        RECT 109.950 557.850 112.050 559.950 ;
        RECT 119.100 558.150 120.900 559.950 ;
        RECT 124.950 558.150 126.150 563.400 ;
        RECT 127.950 561.150 129.750 562.950 ;
        RECT 148.800 562.500 150.600 563.400 ;
        RECT 148.800 561.600 152.850 562.500 ;
        RECT 127.950 559.050 130.050 561.150 ;
        RECT 146.100 558.150 147.900 559.950 ;
        RECT 151.950 558.150 152.850 561.600 ;
        RECT 170.550 561.150 171.750 569.400 ;
        RECT 188.700 569.100 190.350 569.400 ;
        RECT 194.550 569.400 196.350 575.250 ;
        RECT 194.550 569.100 195.750 569.400 ;
        RECT 188.700 568.200 195.750 569.100 ;
        RECT 188.100 564.150 189.900 565.950 ;
        RECT 185.100 561.150 186.900 562.950 ;
        RECT 187.950 562.050 190.050 564.150 ;
        RECT 191.250 561.150 193.050 562.950 ;
        RECT 157.950 558.150 159.750 559.950 ;
        RECT 110.100 556.050 111.900 557.850 ;
        RECT 118.950 556.050 121.050 558.150 ;
        RECT 121.950 554.850 124.050 556.950 ;
        RECT 124.950 556.050 127.050 558.150 ;
        RECT 145.950 556.050 148.050 558.150 ;
        RECT 122.100 553.050 123.900 554.850 ;
        RECT 125.850 552.750 127.050 556.050 ;
        RECT 148.950 554.850 151.050 556.950 ;
        RECT 151.950 556.050 154.050 558.150 ;
        RECT 149.250 553.050 151.050 554.850 ;
        RECT 126.000 551.700 129.750 552.750 ;
        RECT 83.250 549.600 84.450 551.700 ;
        RECT 104.850 550.800 108.450 551.700 ;
        RECT 54.900 547.500 65.700 548.400 ;
        RECT 58.650 546.600 59.700 547.500 ;
        RECT 64.650 546.600 65.700 547.500 ;
        RECT 58.650 543.750 60.450 546.600 ;
        RECT 61.650 543.750 63.450 546.600 ;
        RECT 64.650 543.750 66.450 546.600 ;
        RECT 67.650 543.750 69.750 546.600 ;
        RECT 82.650 543.750 84.450 549.600 ;
        RECT 85.650 548.700 93.450 550.050 ;
        RECT 85.650 543.750 87.450 548.700 ;
        RECT 88.650 543.750 90.450 547.800 ;
        RECT 91.650 543.750 93.450 548.700 ;
        RECT 104.850 543.750 106.650 550.800 ;
        RECT 109.350 543.750 111.150 549.600 ;
        RECT 119.550 548.700 127.350 550.050 ;
        RECT 119.550 543.750 121.350 548.700 ;
        RECT 122.550 543.750 124.350 547.800 ;
        RECT 125.550 543.750 127.350 548.700 ;
        RECT 128.550 549.600 129.750 551.700 ;
        RECT 153.000 549.600 154.050 556.050 ;
        RECT 154.950 554.850 157.050 556.950 ;
        RECT 157.950 556.050 160.050 558.150 ;
        RECT 166.950 557.850 169.050 559.950 ;
        RECT 169.950 559.050 172.050 561.150 ;
        RECT 167.100 556.050 168.900 557.850 ;
        RECT 154.950 553.050 156.750 554.850 ;
        RECT 170.550 551.700 171.750 559.050 ;
        RECT 172.950 557.850 175.050 559.950 ;
        RECT 184.950 559.050 187.050 561.150 ;
        RECT 190.950 559.050 193.050 561.150 ;
        RECT 194.700 559.950 195.750 568.200 ;
        RECT 206.550 564.300 208.350 575.250 ;
        RECT 209.550 565.200 211.350 575.250 ;
        RECT 212.550 564.300 214.350 575.250 ;
        RECT 206.550 563.400 214.350 564.300 ;
        RECT 215.550 563.400 217.350 575.250 ;
        RECT 228.300 563.400 230.100 575.250 ;
        RECT 232.500 563.400 234.300 575.250 ;
        RECT 235.800 569.400 237.600 575.250 ;
        RECT 248.550 569.400 250.350 575.250 ;
        RECT 251.550 569.400 253.350 575.250 ;
        RECT 265.650 569.400 267.450 575.250 ;
        RECT 268.650 569.400 270.450 575.250 ;
        RECT 271.650 569.400 273.450 575.250 ;
        RECT 281.550 569.400 283.350 575.250 ;
        RECT 284.550 569.400 286.350 575.250 ;
        RECT 287.550 569.400 289.350 575.250 ;
        RECT 202.950 561.450 205.050 562.050 ;
        RECT 211.950 561.450 214.050 562.050 ;
        RECT 202.950 560.550 214.050 561.450 ;
        RECT 202.950 559.950 205.050 560.550 ;
        RECT 211.950 559.950 214.050 560.550 ;
        RECT 193.950 557.850 196.050 559.950 ;
        RECT 215.700 558.150 216.900 563.400 ;
        RECT 227.100 558.150 228.900 559.950 ;
        RECT 232.950 558.150 234.150 563.400 ;
        RECT 235.950 561.150 237.750 562.950 ;
        RECT 235.950 559.050 238.050 561.150 ;
        RECT 173.100 556.050 174.900 557.850 ;
        RECT 194.400 553.650 195.600 557.850 ;
        RECT 205.950 554.850 208.050 556.950 ;
        RECT 209.100 555.150 210.900 556.950 ;
        RECT 170.550 550.800 174.150 551.700 ;
        RECT 128.550 543.750 130.350 549.600 ;
        RECT 148.800 543.750 150.600 549.600 ;
        RECT 153.000 543.750 154.800 549.600 ;
        RECT 157.200 543.750 159.000 549.600 ;
        RECT 167.850 543.750 169.650 549.600 ;
        RECT 172.350 543.750 174.150 550.800 ;
        RECT 185.700 543.750 187.500 552.600 ;
        RECT 191.100 552.000 195.600 553.650 ;
        RECT 206.100 553.050 207.900 554.850 ;
        RECT 208.950 553.050 211.050 555.150 ;
        RECT 211.950 554.850 214.050 556.950 ;
        RECT 214.950 556.050 217.050 558.150 ;
        RECT 226.950 556.050 229.050 558.150 ;
        RECT 212.100 553.050 213.900 554.850 ;
        RECT 191.100 543.750 192.900 552.000 ;
        RECT 215.700 549.600 216.900 556.050 ;
        RECT 229.950 554.850 232.050 556.950 ;
        RECT 232.950 556.050 235.050 558.150 ;
        RECT 251.400 556.950 252.600 569.400 ;
        RECT 269.250 561.150 270.450 569.400 ;
        RECT 284.550 561.150 285.750 569.400 ;
        RECT 299.550 563.400 301.350 575.250 ;
        RECT 304.050 563.550 305.850 575.250 ;
        RECT 307.050 564.900 308.850 575.250 ;
        RECT 320.550 569.400 322.350 575.250 ;
        RECT 323.550 569.400 325.350 575.250 ;
        RECT 326.550 569.400 328.350 575.250 ;
        RECT 338.550 569.400 340.350 575.250 ;
        RECT 341.550 569.400 343.350 575.250 ;
        RECT 344.550 570.000 346.350 575.250 ;
        RECT 307.050 563.550 309.450 564.900 ;
        RECT 299.550 562.200 300.750 563.400 ;
        RECT 304.950 562.200 306.750 562.650 ;
        RECT 265.950 557.850 268.050 559.950 ;
        RECT 268.950 559.050 271.050 561.150 ;
        RECT 230.100 553.050 231.900 554.850 ;
        RECT 233.850 552.750 235.050 556.050 ;
        RECT 248.100 555.150 249.900 556.950 ;
        RECT 247.950 553.050 250.050 555.150 ;
        RECT 250.950 554.850 253.050 556.950 ;
        RECT 266.100 556.050 267.900 557.850 ;
        RECT 234.000 551.700 237.750 552.750 ;
        RECT 207.000 543.750 208.800 549.600 ;
        RECT 211.200 547.950 216.900 549.600 ;
        RECT 227.550 548.700 235.350 550.050 ;
        RECT 211.200 543.750 213.000 547.950 ;
        RECT 214.500 543.750 216.300 546.600 ;
        RECT 227.550 543.750 229.350 548.700 ;
        RECT 230.550 543.750 232.350 547.800 ;
        RECT 233.550 543.750 235.350 548.700 ;
        RECT 236.550 549.600 237.750 551.700 ;
        RECT 236.550 543.750 238.350 549.600 ;
        RECT 251.400 546.600 252.600 554.850 ;
        RECT 269.250 551.700 270.450 559.050 ;
        RECT 271.950 557.850 274.050 559.950 ;
        RECT 280.950 557.850 283.050 559.950 ;
        RECT 283.950 559.050 286.050 561.150 ;
        RECT 299.550 561.000 306.750 562.200 ;
        RECT 304.950 560.850 306.750 561.000 ;
        RECT 272.100 556.050 273.900 557.850 ;
        RECT 281.100 556.050 282.900 557.850 ;
        RECT 266.850 550.800 270.450 551.700 ;
        RECT 284.550 551.700 285.750 559.050 ;
        RECT 286.950 557.850 289.050 559.950 ;
        RECT 302.100 558.150 303.900 559.950 ;
        RECT 287.100 556.050 288.900 557.850 ;
        RECT 299.100 555.150 300.900 556.950 ;
        RECT 301.950 556.050 304.050 558.150 ;
        RECT 298.950 553.050 301.050 555.150 ;
        RECT 305.700 552.600 306.600 560.850 ;
        RECT 308.100 556.950 309.450 563.550 ;
        RECT 323.550 561.150 324.750 569.400 ;
        RECT 341.700 569.100 343.350 569.400 ;
        RECT 347.550 569.400 349.350 575.250 ;
        RECT 362.400 569.400 364.200 575.250 ;
        RECT 347.550 569.100 348.750 569.400 ;
        RECT 341.700 568.200 348.750 569.100 ;
        RECT 341.100 564.150 342.900 565.950 ;
        RECT 338.100 561.150 339.900 562.950 ;
        RECT 340.950 562.050 343.050 564.150 ;
        RECT 344.250 561.150 346.050 562.950 ;
        RECT 319.950 557.850 322.050 559.950 ;
        RECT 322.950 559.050 325.050 561.150 ;
        RECT 307.950 554.850 310.050 556.950 ;
        RECT 320.100 556.050 321.900 557.850 ;
        RECT 304.950 551.700 306.750 552.600 ;
        RECT 284.550 550.800 288.150 551.700 ;
        RECT 248.550 543.750 250.350 546.600 ;
        RECT 251.550 543.750 253.350 546.600 ;
        RECT 266.850 543.750 268.650 550.800 ;
        RECT 271.350 543.750 273.150 549.600 ;
        RECT 281.850 543.750 283.650 549.600 ;
        RECT 286.350 543.750 288.150 550.800 ;
        RECT 303.450 550.800 306.750 551.700 ;
        RECT 303.450 546.600 304.350 550.800 ;
        RECT 309.000 549.600 310.050 554.850 ;
        RECT 323.550 551.700 324.750 559.050 ;
        RECT 325.950 557.850 328.050 559.950 ;
        RECT 337.950 559.050 340.050 561.150 ;
        RECT 343.950 559.050 346.050 561.150 ;
        RECT 347.700 559.950 348.750 568.200 ;
        RECT 365.700 563.400 367.500 575.250 ;
        RECT 369.900 563.400 371.700 575.250 ;
        RECT 380.550 569.400 382.350 575.250 ;
        RECT 383.550 569.400 385.350 575.250 ;
        RECT 386.550 569.400 388.350 575.250 ;
        RECT 362.250 561.150 364.050 562.950 ;
        RECT 346.950 557.850 349.050 559.950 ;
        RECT 361.950 559.050 364.050 561.150 ;
        RECT 365.850 558.150 367.050 563.400 ;
        RECT 383.550 561.150 384.750 569.400 ;
        RECT 399.300 563.400 401.100 575.250 ;
        RECT 403.500 563.400 405.300 575.250 ;
        RECT 406.800 569.400 408.600 575.250 ;
        RECT 421.650 569.400 423.450 575.250 ;
        RECT 424.650 569.400 426.450 575.250 ;
        RECT 437.400 569.400 439.200 575.250 ;
        RECT 371.100 558.150 372.900 559.950 ;
        RECT 326.100 556.050 327.900 557.850 ;
        RECT 347.400 553.650 348.600 557.850 ;
        RECT 323.550 550.800 327.150 551.700 ;
        RECT 299.550 543.750 301.350 546.600 ;
        RECT 302.550 543.750 304.350 546.600 ;
        RECT 305.550 543.750 307.350 546.600 ;
        RECT 308.550 543.750 310.350 549.600 ;
        RECT 320.850 543.750 322.650 549.600 ;
        RECT 325.350 543.750 327.150 550.800 ;
        RECT 338.700 543.750 340.500 552.600 ;
        RECT 344.100 552.000 348.600 553.650 ;
        RECT 364.950 556.050 367.050 558.150 ;
        RECT 364.950 552.750 366.150 556.050 ;
        RECT 367.950 554.850 370.050 556.950 ;
        RECT 370.950 556.050 373.050 558.150 ;
        RECT 379.950 557.850 382.050 559.950 ;
        RECT 382.950 559.050 385.050 561.150 ;
        RECT 380.100 556.050 381.900 557.850 ;
        RECT 368.100 553.050 369.900 554.850 ;
        RECT 344.100 543.750 345.900 552.000 ;
        RECT 362.250 551.700 366.000 552.750 ;
        RECT 383.550 551.700 384.750 559.050 ;
        RECT 385.950 557.850 388.050 559.950 ;
        RECT 398.100 558.150 399.900 559.950 ;
        RECT 403.950 558.150 405.150 563.400 ;
        RECT 406.950 561.150 408.750 562.950 ;
        RECT 406.950 559.050 409.050 561.150 ;
        RECT 386.100 556.050 387.900 557.850 ;
        RECT 397.950 556.050 400.050 558.150 ;
        RECT 400.950 554.850 403.050 556.950 ;
        RECT 403.950 556.050 406.050 558.150 ;
        RECT 422.400 556.950 423.600 569.400 ;
        RECT 440.700 563.400 442.500 575.250 ;
        RECT 444.900 563.400 446.700 575.250 ;
        RECT 455.550 569.400 457.350 575.250 ;
        RECT 458.550 569.400 460.350 575.250 ;
        RECT 461.550 569.400 463.350 575.250 ;
        RECT 478.650 569.400 480.450 575.250 ;
        RECT 481.650 569.400 483.450 575.250 ;
        RECT 484.650 569.400 486.450 575.250 ;
        RECT 496.650 569.400 498.450 575.250 ;
        RECT 499.650 569.400 501.450 575.250 ;
        RECT 509.550 569.400 511.350 575.250 ;
        RECT 512.550 569.400 514.350 575.250 ;
        RECT 515.550 570.000 517.350 575.250 ;
        RECT 437.250 561.150 439.050 562.950 ;
        RECT 436.950 559.050 439.050 561.150 ;
        RECT 440.850 558.150 442.050 563.400 ;
        RECT 458.550 561.150 459.750 569.400 ;
        RECT 460.950 564.450 463.050 565.050 ;
        RECT 478.950 564.450 481.050 565.050 ;
        RECT 460.950 563.550 481.050 564.450 ;
        RECT 460.950 562.950 463.050 563.550 ;
        RECT 478.950 562.950 481.050 563.550 ;
        RECT 482.250 561.150 483.450 569.400 ;
        RECT 446.100 558.150 447.900 559.950 ;
        RECT 401.100 553.050 402.900 554.850 ;
        RECT 404.850 552.750 406.050 556.050 ;
        RECT 421.950 554.850 424.050 556.950 ;
        RECT 425.100 555.150 426.900 556.950 ;
        RECT 439.950 556.050 442.050 558.150 ;
        RECT 405.000 551.700 408.750 552.750 ;
        RECT 362.250 549.600 363.450 551.700 ;
        RECT 383.550 550.800 387.150 551.700 ;
        RECT 361.650 543.750 363.450 549.600 ;
        RECT 364.650 548.700 372.450 550.050 ;
        RECT 364.650 543.750 366.450 548.700 ;
        RECT 367.650 543.750 369.450 547.800 ;
        RECT 370.650 543.750 372.450 548.700 ;
        RECT 380.850 543.750 382.650 549.600 ;
        RECT 385.350 543.750 387.150 550.800 ;
        RECT 398.550 548.700 406.350 550.050 ;
        RECT 398.550 543.750 400.350 548.700 ;
        RECT 401.550 543.750 403.350 547.800 ;
        RECT 404.550 543.750 406.350 548.700 ;
        RECT 407.550 549.600 408.750 551.700 ;
        RECT 407.550 543.750 409.350 549.600 ;
        RECT 422.400 546.600 423.600 554.850 ;
        RECT 424.950 553.050 427.050 555.150 ;
        RECT 439.950 552.750 441.150 556.050 ;
        RECT 442.950 554.850 445.050 556.950 ;
        RECT 445.950 556.050 448.050 558.150 ;
        RECT 454.950 557.850 457.050 559.950 ;
        RECT 457.950 559.050 460.050 561.150 ;
        RECT 455.100 556.050 456.900 557.850 ;
        RECT 443.100 553.050 444.900 554.850 ;
        RECT 437.250 551.700 441.000 552.750 ;
        RECT 458.550 551.700 459.750 559.050 ;
        RECT 460.950 557.850 463.050 559.950 ;
        RECT 478.950 557.850 481.050 559.950 ;
        RECT 481.950 559.050 484.050 561.150 ;
        RECT 461.100 556.050 462.900 557.850 ;
        RECT 479.100 556.050 480.900 557.850 ;
        RECT 482.250 551.700 483.450 559.050 ;
        RECT 484.950 557.850 487.050 559.950 ;
        RECT 485.100 556.050 486.900 557.850 ;
        RECT 497.400 556.950 498.600 569.400 ;
        RECT 512.700 569.100 514.350 569.400 ;
        RECT 518.550 569.400 520.350 575.250 ;
        RECT 530.550 569.400 532.350 575.250 ;
        RECT 533.550 569.400 535.350 575.250 ;
        RECT 518.550 569.100 519.750 569.400 ;
        RECT 512.700 568.200 519.750 569.100 ;
        RECT 502.950 567.450 505.050 568.050 ;
        RECT 508.950 567.450 511.050 568.050 ;
        RECT 502.950 566.550 511.050 567.450 ;
        RECT 502.950 565.950 505.050 566.550 ;
        RECT 508.950 565.950 511.050 566.550 ;
        RECT 512.100 564.150 513.900 565.950 ;
        RECT 509.100 561.150 510.900 562.950 ;
        RECT 511.950 562.050 514.050 564.150 ;
        RECT 515.250 561.150 517.050 562.950 ;
        RECT 508.950 559.050 511.050 561.150 ;
        RECT 514.950 559.050 517.050 561.150 ;
        RECT 518.700 559.950 519.750 568.200 ;
        RECT 517.950 557.850 520.050 559.950 ;
        RECT 496.950 554.850 499.050 556.950 ;
        RECT 500.100 555.150 501.900 556.950 ;
        RECT 437.250 549.600 438.450 551.700 ;
        RECT 458.550 550.800 462.150 551.700 ;
        RECT 421.650 543.750 423.450 546.600 ;
        RECT 424.650 543.750 426.450 546.600 ;
        RECT 436.650 543.750 438.450 549.600 ;
        RECT 439.650 548.700 447.450 550.050 ;
        RECT 439.650 543.750 441.450 548.700 ;
        RECT 442.650 543.750 444.450 547.800 ;
        RECT 445.650 543.750 447.450 548.700 ;
        RECT 455.850 543.750 457.650 549.600 ;
        RECT 460.350 543.750 462.150 550.800 ;
        RECT 479.850 550.800 483.450 551.700 ;
        RECT 479.850 543.750 481.650 550.800 ;
        RECT 484.350 543.750 486.150 549.600 ;
        RECT 497.400 546.600 498.600 554.850 ;
        RECT 499.950 553.050 502.050 555.150 ;
        RECT 518.400 553.650 519.600 557.850 ;
        RECT 533.400 556.950 534.600 569.400 ;
        RECT 549.450 563.400 551.250 575.250 ;
        RECT 553.650 563.400 555.450 575.250 ;
        RECT 566.550 569.400 568.350 575.250 ;
        RECT 569.550 569.400 571.350 575.250 ;
        RECT 572.550 569.400 574.350 575.250 ;
        RECT 584.550 569.400 586.350 575.250 ;
        RECT 587.550 569.400 589.350 575.250 ;
        RECT 601.650 569.400 603.450 575.250 ;
        RECT 604.650 569.400 606.450 575.250 ;
        RECT 549.450 562.350 552.000 563.400 ;
        RECT 548.100 558.150 549.900 559.950 ;
        RECT 530.100 555.150 531.900 556.950 ;
        RECT 496.650 543.750 498.450 546.600 ;
        RECT 499.650 543.750 501.450 546.600 ;
        RECT 509.700 543.750 511.500 552.600 ;
        RECT 515.100 552.000 519.600 553.650 ;
        RECT 529.950 553.050 532.050 555.150 ;
        RECT 532.950 554.850 535.050 556.950 ;
        RECT 547.950 556.050 550.050 558.150 ;
        RECT 550.950 555.150 552.000 562.350 ;
        RECT 569.550 561.150 570.750 569.400 ;
        RECT 554.100 558.150 555.900 559.950 ;
        RECT 553.950 556.050 556.050 558.150 ;
        RECT 565.950 557.850 568.050 559.950 ;
        RECT 568.950 559.050 571.050 561.150 ;
        RECT 566.100 556.050 567.900 557.850 ;
        RECT 515.100 543.750 516.900 552.000 ;
        RECT 533.400 546.600 534.600 554.850 ;
        RECT 550.950 553.050 553.050 555.150 ;
        RECT 550.950 546.600 552.000 553.050 ;
        RECT 569.550 551.700 570.750 559.050 ;
        RECT 571.950 557.850 574.050 559.950 ;
        RECT 572.100 556.050 573.900 557.850 ;
        RECT 587.400 556.950 588.600 569.400 ;
        RECT 602.400 556.950 603.600 569.400 ;
        RECT 608.550 563.400 610.350 575.250 ;
        RECT 611.550 572.400 613.350 575.250 ;
        RECT 616.050 569.400 617.850 575.250 ;
        RECT 620.250 569.400 622.050 575.250 ;
        RECT 613.950 567.300 617.850 569.400 ;
        RECT 624.150 568.500 625.950 575.250 ;
        RECT 627.150 569.400 628.950 575.250 ;
        RECT 631.950 569.400 633.750 575.250 ;
        RECT 637.050 569.400 638.850 575.250 ;
        RECT 632.250 568.500 633.450 569.400 ;
        RECT 622.950 566.700 629.850 568.500 ;
        RECT 632.250 566.400 637.050 568.500 ;
        RECT 615.150 564.600 617.850 566.400 ;
        RECT 618.750 565.800 620.550 566.400 ;
        RECT 618.750 564.900 625.050 565.800 ;
        RECT 632.250 565.500 633.450 566.400 ;
        RECT 618.750 564.600 620.550 564.900 ;
        RECT 616.950 563.700 617.850 564.600 ;
        RECT 584.100 555.150 585.900 556.950 ;
        RECT 583.950 553.050 586.050 555.150 ;
        RECT 586.950 554.850 589.050 556.950 ;
        RECT 601.950 554.850 604.050 556.950 ;
        RECT 605.100 555.150 606.900 556.950 ;
        RECT 569.550 550.800 573.150 551.700 ;
        RECT 530.550 543.750 532.350 546.600 ;
        RECT 533.550 543.750 535.350 546.600 ;
        RECT 547.650 543.750 549.450 546.600 ;
        RECT 550.650 543.750 552.450 546.600 ;
        RECT 553.650 543.750 555.450 546.600 ;
        RECT 566.850 543.750 568.650 549.600 ;
        RECT 571.350 543.750 573.150 550.800 ;
        RECT 587.400 546.600 588.600 554.850 ;
        RECT 602.400 546.600 603.600 554.850 ;
        RECT 604.950 553.050 607.050 555.150 ;
        RECT 608.550 553.950 609.750 563.400 ;
        RECT 613.950 562.800 616.050 563.700 ;
        RECT 616.950 562.800 622.950 563.700 ;
        RECT 611.850 561.600 616.050 562.800 ;
        RECT 610.950 559.800 612.750 561.600 ;
        RECT 622.050 558.150 622.950 562.800 ;
        RECT 624.150 562.800 625.050 564.900 ;
        RECT 625.950 564.300 633.450 565.500 ;
        RECT 625.950 563.700 627.750 564.300 ;
        RECT 640.050 563.400 641.850 575.250 ;
        RECT 654.150 563.400 655.950 575.250 ;
        RECT 658.650 563.400 661.950 575.250 ;
        RECT 664.650 563.400 666.450 575.250 ;
        RECT 674.550 569.400 676.350 575.250 ;
        RECT 677.550 569.400 679.350 575.250 ;
        RECT 680.550 569.400 682.350 575.250 ;
        RECT 630.750 562.800 641.850 563.400 ;
        RECT 624.150 562.200 641.850 562.800 ;
        RECT 624.150 561.900 632.550 562.200 ;
        RECT 630.750 561.600 632.550 561.900 ;
        RECT 622.050 556.050 625.050 558.150 ;
        RECT 628.950 557.100 631.050 558.150 ;
        RECT 628.950 556.050 636.900 557.100 ;
        RECT 610.950 555.750 613.050 556.050 ;
        RECT 610.950 553.950 614.850 555.750 ;
        RECT 608.550 551.850 613.050 553.950 ;
        RECT 622.050 552.000 622.950 556.050 ;
        RECT 635.100 555.300 636.900 556.050 ;
        RECT 638.100 555.150 639.900 556.950 ;
        RECT 632.100 554.400 633.900 555.000 ;
        RECT 638.100 554.400 639.000 555.150 ;
        RECT 632.100 553.200 639.000 554.400 ;
        RECT 632.100 552.000 633.150 553.200 ;
        RECT 608.550 549.600 609.750 551.850 ;
        RECT 622.050 551.100 633.150 552.000 ;
        RECT 622.050 550.800 622.950 551.100 ;
        RECT 584.550 543.750 586.350 546.600 ;
        RECT 587.550 543.750 589.350 546.600 ;
        RECT 601.650 543.750 603.450 546.600 ;
        RECT 604.650 543.750 606.450 546.600 ;
        RECT 608.550 543.750 610.350 549.600 ;
        RECT 613.950 548.700 616.050 549.600 ;
        RECT 621.150 549.000 622.950 550.800 ;
        RECT 632.100 550.200 633.150 551.100 ;
        RECT 628.350 549.450 630.150 550.200 ;
        RECT 613.950 547.500 617.700 548.700 ;
        RECT 616.650 546.600 617.700 547.500 ;
        RECT 625.200 548.400 630.150 549.450 ;
        RECT 631.650 548.400 633.450 550.200 ;
        RECT 640.950 549.600 641.850 562.200 ;
        RECT 653.250 558.150 655.050 559.950 ;
        RECT 659.250 558.150 660.450 563.400 ;
        RECT 677.550 561.150 678.750 569.400 ;
        RECT 692.550 563.400 694.350 575.250 ;
        RECT 696.750 563.400 698.550 575.250 ;
        RECT 711.300 563.400 713.100 575.250 ;
        RECT 715.500 563.400 717.300 575.250 ;
        RECT 718.800 569.400 720.600 575.250 ;
        RECT 731.550 563.400 733.350 575.250 ;
        RECT 734.550 563.400 736.350 575.250 ;
        RECT 751.650 569.400 753.450 575.250 ;
        RECT 754.650 569.400 756.450 575.250 ;
        RECT 757.650 569.400 759.450 575.250 ;
        RECT 767.550 569.400 769.350 575.250 ;
        RECT 770.550 569.400 772.350 575.250 ;
        RECT 696.000 562.350 698.550 563.400 ;
        RECT 665.100 558.150 666.900 559.950 ;
        RECT 652.950 556.050 655.050 558.150 ;
        RECT 655.950 554.850 658.050 556.950 ;
        RECT 658.950 556.050 661.050 558.150 ;
        RECT 656.700 553.050 658.500 554.850 ;
        RECT 659.400 552.150 660.600 556.050 ;
        RECT 661.950 554.850 664.050 556.950 ;
        RECT 664.950 556.050 667.050 558.150 ;
        RECT 673.950 557.850 676.050 559.950 ;
        RECT 676.950 559.050 679.050 561.150 ;
        RECT 674.100 556.050 675.900 557.850 ;
        RECT 662.100 553.050 663.900 554.850 ;
        RECT 656.250 551.100 660.600 552.150 ;
        RECT 677.550 551.700 678.750 559.050 ;
        RECT 679.950 557.850 682.050 559.950 ;
        RECT 692.100 558.150 693.900 559.950 ;
        RECT 680.100 556.050 681.900 557.850 ;
        RECT 691.950 556.050 694.050 558.150 ;
        RECT 696.000 555.150 697.050 562.350 ;
        RECT 698.100 558.150 699.900 559.950 ;
        RECT 710.100 558.150 711.900 559.950 ;
        RECT 715.950 558.150 717.150 563.400 ;
        RECT 718.950 561.150 720.750 562.950 ;
        RECT 724.950 561.450 727.050 562.050 ;
        RECT 730.950 561.450 733.050 562.050 ;
        RECT 718.950 559.050 721.050 561.150 ;
        RECT 724.950 560.550 733.050 561.450 ;
        RECT 724.950 559.950 727.050 560.550 ;
        RECT 730.950 559.950 733.050 560.550 ;
        RECT 734.400 558.150 735.600 563.400 ;
        RECT 755.250 561.150 756.450 569.400 ;
        RECT 697.950 556.050 700.050 558.150 ;
        RECT 709.950 556.050 712.050 558.150 ;
        RECT 694.950 553.050 697.050 555.150 ;
        RECT 712.950 554.850 715.050 556.950 ;
        RECT 715.950 556.050 718.050 558.150 ;
        RECT 713.100 553.050 714.900 554.850 ;
        RECT 656.250 549.600 657.150 551.100 ;
        RECT 677.550 550.800 681.150 551.700 ;
        RECT 625.200 546.600 626.250 548.400 ;
        RECT 634.950 547.500 637.050 549.600 ;
        RECT 634.950 546.600 636.000 547.500 ;
        RECT 611.850 543.750 613.650 546.600 ;
        RECT 616.350 543.750 618.150 546.600 ;
        RECT 620.550 543.750 622.350 546.600 ;
        RECT 624.450 543.750 626.250 546.600 ;
        RECT 627.750 543.750 629.550 546.600 ;
        RECT 632.250 545.700 636.000 546.600 ;
        RECT 632.250 543.750 634.050 545.700 ;
        RECT 637.050 543.750 638.850 546.600 ;
        RECT 640.050 543.750 641.850 549.600 ;
        RECT 652.650 544.500 654.450 549.600 ;
        RECT 655.650 545.400 657.450 549.600 ;
        RECT 658.650 549.000 666.450 549.900 ;
        RECT 658.650 544.500 660.450 549.000 ;
        RECT 652.650 543.750 660.450 544.500 ;
        RECT 661.650 543.750 663.450 548.100 ;
        RECT 664.650 543.750 666.450 549.000 ;
        RECT 674.850 543.750 676.650 549.600 ;
        RECT 679.350 543.750 681.150 550.800 ;
        RECT 696.000 546.600 697.050 553.050 ;
        RECT 716.850 552.750 718.050 556.050 ;
        RECT 730.950 554.850 733.050 556.950 ;
        RECT 733.950 556.050 736.050 558.150 ;
        RECT 751.950 557.850 754.050 559.950 ;
        RECT 754.950 559.050 757.050 561.150 ;
        RECT 752.100 556.050 753.900 557.850 ;
        RECT 731.100 553.050 732.900 554.850 ;
        RECT 717.000 551.700 720.750 552.750 ;
        RECT 710.550 548.700 718.350 550.050 ;
        RECT 692.550 543.750 694.350 546.600 ;
        RECT 695.550 543.750 697.350 546.600 ;
        RECT 698.550 543.750 700.350 546.600 ;
        RECT 710.550 543.750 712.350 548.700 ;
        RECT 713.550 543.750 715.350 547.800 ;
        RECT 716.550 543.750 718.350 548.700 ;
        RECT 719.550 549.600 720.750 551.700 ;
        RECT 734.400 549.600 735.600 556.050 ;
        RECT 755.250 551.700 756.450 559.050 ;
        RECT 757.950 557.850 760.050 559.950 ;
        RECT 758.100 556.050 759.900 557.850 ;
        RECT 770.400 556.950 771.600 569.400 ;
        RECT 784.650 563.400 786.450 575.250 ;
        RECT 787.650 562.500 789.450 575.250 ;
        RECT 790.650 563.400 792.450 575.250 ;
        RECT 793.650 562.500 795.450 575.250 ;
        RECT 796.650 563.400 798.450 575.250 ;
        RECT 799.650 562.500 801.450 575.250 ;
        RECT 802.650 563.400 804.450 575.250 ;
        RECT 805.650 562.500 807.450 575.250 ;
        RECT 808.650 563.400 810.450 575.250 ;
        RECT 812.550 563.400 814.350 575.250 ;
        RECT 815.550 572.400 817.350 575.250 ;
        RECT 820.050 569.400 821.850 575.250 ;
        RECT 824.250 569.400 826.050 575.250 ;
        RECT 817.950 567.300 821.850 569.400 ;
        RECT 828.150 568.500 829.950 575.250 ;
        RECT 831.150 569.400 832.950 575.250 ;
        RECT 835.950 569.400 837.750 575.250 ;
        RECT 841.050 569.400 842.850 575.250 ;
        RECT 836.250 568.500 837.450 569.400 ;
        RECT 826.950 566.700 833.850 568.500 ;
        RECT 836.250 566.400 841.050 568.500 ;
        RECT 819.150 564.600 821.850 566.400 ;
        RECT 822.750 565.800 824.550 566.400 ;
        RECT 822.750 564.900 829.050 565.800 ;
        RECT 836.250 565.500 837.450 566.400 ;
        RECT 822.750 564.600 824.550 564.900 ;
        RECT 820.950 563.700 821.850 564.600 ;
        RECT 786.750 561.300 789.450 562.500 ;
        RECT 791.700 561.300 795.450 562.500 ;
        RECT 797.700 561.300 801.450 562.500 ;
        RECT 803.550 561.300 807.450 562.500 ;
        RECT 786.750 556.950 787.800 561.300 ;
        RECT 767.100 555.150 768.900 556.950 ;
        RECT 766.950 553.050 769.050 555.150 ;
        RECT 769.950 554.850 772.050 556.950 ;
        RECT 784.950 554.850 787.800 556.950 ;
        RECT 752.850 550.800 756.450 551.700 ;
        RECT 719.550 543.750 721.350 549.600 ;
        RECT 731.550 543.750 733.350 549.600 ;
        RECT 734.550 543.750 736.350 549.600 ;
        RECT 752.850 543.750 754.650 550.800 ;
        RECT 757.350 543.750 759.150 549.600 ;
        RECT 770.400 546.600 771.600 554.850 ;
        RECT 786.750 551.700 787.800 554.850 ;
        RECT 791.700 554.400 792.900 561.300 ;
        RECT 797.700 554.400 798.900 561.300 ;
        RECT 803.550 554.400 804.750 561.300 ;
        RECT 805.950 554.850 808.050 556.950 ;
        RECT 788.700 552.600 792.900 554.400 ;
        RECT 794.700 552.600 798.900 554.400 ;
        RECT 800.700 552.600 804.750 554.400 ;
        RECT 806.100 553.050 807.900 554.850 ;
        RECT 812.550 553.950 813.750 563.400 ;
        RECT 817.950 562.800 820.050 563.700 ;
        RECT 820.950 562.800 826.950 563.700 ;
        RECT 815.850 561.600 820.050 562.800 ;
        RECT 814.950 559.800 816.750 561.600 ;
        RECT 826.050 558.150 826.950 562.800 ;
        RECT 828.150 562.800 829.050 564.900 ;
        RECT 829.950 564.300 837.450 565.500 ;
        RECT 829.950 563.700 831.750 564.300 ;
        RECT 844.050 563.400 845.850 575.250 ;
        RECT 856.650 569.400 858.450 575.250 ;
        RECT 859.650 569.400 861.450 575.250 ;
        RECT 862.650 569.400 864.450 575.250 ;
        RECT 834.750 562.800 845.850 563.400 ;
        RECT 828.150 562.200 845.850 562.800 ;
        RECT 828.150 561.900 836.550 562.200 ;
        RECT 834.750 561.600 836.550 561.900 ;
        RECT 826.050 556.050 829.050 558.150 ;
        RECT 832.950 557.100 835.050 558.150 ;
        RECT 832.950 556.050 840.900 557.100 ;
        RECT 814.950 555.750 817.050 556.050 ;
        RECT 814.950 553.950 818.850 555.750 ;
        RECT 791.700 551.700 792.900 552.600 ;
        RECT 797.700 551.700 798.900 552.600 ;
        RECT 803.550 551.700 804.750 552.600 ;
        RECT 812.550 551.850 817.050 553.950 ;
        RECT 826.050 552.000 826.950 556.050 ;
        RECT 839.100 555.300 840.900 556.050 ;
        RECT 842.100 555.150 843.900 556.950 ;
        RECT 836.100 554.400 837.900 555.000 ;
        RECT 842.100 554.400 843.000 555.150 ;
        RECT 836.100 553.200 843.000 554.400 ;
        RECT 836.100 552.000 837.150 553.200 ;
        RECT 786.750 550.650 789.600 551.700 ;
        RECT 786.900 550.500 789.600 550.650 ;
        RECT 791.700 550.500 795.600 551.700 ;
        RECT 797.700 550.500 801.450 551.700 ;
        RECT 803.550 550.500 807.600 551.700 ;
        RECT 787.800 549.600 789.600 550.500 ;
        RECT 793.800 549.600 795.600 550.500 ;
        RECT 767.550 543.750 769.350 546.600 ;
        RECT 770.550 543.750 772.350 546.600 ;
        RECT 784.650 543.750 786.450 549.600 ;
        RECT 787.650 543.750 789.450 549.600 ;
        RECT 790.650 543.750 792.450 549.600 ;
        RECT 793.650 543.750 795.450 549.600 ;
        RECT 796.650 543.750 798.450 549.600 ;
        RECT 799.650 543.750 801.450 550.500 ;
        RECT 805.800 549.600 807.600 550.500 ;
        RECT 812.550 549.600 813.750 551.850 ;
        RECT 826.050 551.100 837.150 552.000 ;
        RECT 826.050 550.800 826.950 551.100 ;
        RECT 802.650 543.750 804.450 549.600 ;
        RECT 805.650 543.750 807.450 549.600 ;
        RECT 808.650 543.750 810.450 549.600 ;
        RECT 812.550 543.750 814.350 549.600 ;
        RECT 817.950 548.700 820.050 549.600 ;
        RECT 825.150 549.000 826.950 550.800 ;
        RECT 836.100 550.200 837.150 551.100 ;
        RECT 832.350 549.450 834.150 550.200 ;
        RECT 817.950 547.500 821.700 548.700 ;
        RECT 820.650 546.600 821.700 547.500 ;
        RECT 829.200 548.400 834.150 549.450 ;
        RECT 835.650 548.400 837.450 550.200 ;
        RECT 844.950 549.600 845.850 562.200 ;
        RECT 860.250 561.150 861.450 569.400 ;
        RECT 856.950 557.850 859.050 559.950 ;
        RECT 859.950 559.050 862.050 561.150 ;
        RECT 857.100 556.050 858.900 557.850 ;
        RECT 860.250 551.700 861.450 559.050 ;
        RECT 862.950 557.850 865.050 559.950 ;
        RECT 863.100 556.050 864.900 557.850 ;
        RECT 829.200 546.600 830.250 548.400 ;
        RECT 838.950 547.500 841.050 549.600 ;
        RECT 838.950 546.600 840.000 547.500 ;
        RECT 815.850 543.750 817.650 546.600 ;
        RECT 820.350 543.750 822.150 546.600 ;
        RECT 824.550 543.750 826.350 546.600 ;
        RECT 828.450 543.750 830.250 546.600 ;
        RECT 831.750 543.750 833.550 546.600 ;
        RECT 836.250 545.700 840.000 546.600 ;
        RECT 836.250 543.750 838.050 545.700 ;
        RECT 841.050 543.750 842.850 546.600 ;
        RECT 844.050 543.750 845.850 549.600 ;
        RECT 857.850 550.800 861.450 551.700 ;
        RECT 857.850 543.750 859.650 550.800 ;
        RECT 862.350 543.750 864.150 549.600 ;
        RECT 10.650 533.400 12.450 539.250 ;
        RECT 11.250 531.300 12.450 533.400 ;
        RECT 13.650 534.300 15.450 539.250 ;
        RECT 16.650 535.200 18.450 539.250 ;
        RECT 19.650 534.300 21.450 539.250 ;
        RECT 13.650 532.950 21.450 534.300 ;
        RECT 30.000 533.400 31.800 539.250 ;
        RECT 34.200 535.050 36.000 539.250 ;
        RECT 37.500 536.400 39.300 539.250 ;
        RECT 50.550 536.400 52.350 539.250 ;
        RECT 53.550 536.400 55.350 539.250 ;
        RECT 34.200 533.400 39.900 535.050 ;
        RECT 11.250 530.250 15.000 531.300 ;
        RECT 10.950 528.450 13.050 529.050 ;
        RECT 8.550 527.550 13.050 528.450 ;
        RECT 8.550 516.450 9.450 527.550 ;
        RECT 10.950 526.950 13.050 527.550 ;
        RECT 13.950 526.950 15.150 530.250 ;
        RECT 17.100 528.150 18.900 529.950 ;
        RECT 29.100 528.150 30.900 529.950 ;
        RECT 13.950 524.850 16.050 526.950 ;
        RECT 16.950 526.050 19.050 528.150 ;
        RECT 19.950 524.850 22.050 526.950 ;
        RECT 28.950 526.050 31.050 528.150 ;
        RECT 31.950 527.850 34.050 529.950 ;
        RECT 35.100 528.150 36.900 529.950 ;
        RECT 32.100 526.050 33.900 527.850 ;
        RECT 34.950 526.050 37.050 528.150 ;
        RECT 38.700 526.950 39.900 533.400 ;
        RECT 49.950 527.850 52.050 529.950 ;
        RECT 53.400 528.150 54.600 536.400 ;
        RECT 65.550 534.300 67.350 539.250 ;
        RECT 68.550 535.200 70.350 539.250 ;
        RECT 71.550 534.300 73.350 539.250 ;
        RECT 65.550 532.950 73.350 534.300 ;
        RECT 74.550 533.400 76.350 539.250 ;
        RECT 74.550 531.300 75.750 533.400 ;
        RECT 72.000 530.250 75.750 531.300 ;
        RECT 86.700 530.400 88.500 539.250 ;
        RECT 92.100 531.000 93.900 539.250 ;
        RECT 113.850 532.200 115.650 539.250 ;
        RECT 118.350 533.400 120.150 539.250 ;
        RECT 131.850 532.200 133.650 539.250 ;
        RECT 136.350 533.400 138.150 539.250 ;
        RECT 146.550 534.300 148.350 539.250 ;
        RECT 149.550 535.200 151.350 539.250 ;
        RECT 152.550 534.300 154.350 539.250 ;
        RECT 146.550 532.950 154.350 534.300 ;
        RECT 155.550 533.400 157.350 539.250 ;
        RECT 113.850 531.300 117.450 532.200 ;
        RECT 131.850 531.300 135.450 532.200 ;
        RECT 155.550 531.300 156.750 533.400 ;
        RECT 68.100 528.150 69.900 529.950 ;
        RECT 37.950 524.850 40.050 526.950 ;
        RECT 50.100 526.050 51.900 527.850 ;
        RECT 52.950 526.050 55.050 528.150 ;
        RECT 10.950 521.850 13.050 523.950 ;
        RECT 11.250 520.050 13.050 521.850 ;
        RECT 14.850 519.600 16.050 524.850 ;
        RECT 20.100 523.050 21.900 524.850 ;
        RECT 38.700 519.600 39.900 524.850 ;
        RECT 10.950 516.450 13.050 517.050 ;
        RECT 8.550 515.550 13.050 516.450 ;
        RECT 10.950 514.950 13.050 515.550 ;
        RECT 11.400 507.750 13.200 513.600 ;
        RECT 14.700 507.750 16.500 519.600 ;
        RECT 18.900 507.750 20.700 519.600 ;
        RECT 29.550 518.700 37.350 519.600 ;
        RECT 29.550 507.750 31.350 518.700 ;
        RECT 32.550 507.750 34.350 517.800 ;
        RECT 35.550 507.750 37.350 518.700 ;
        RECT 38.550 507.750 40.350 519.600 ;
        RECT 53.400 513.600 54.600 526.050 ;
        RECT 64.950 524.850 67.050 526.950 ;
        RECT 67.950 526.050 70.050 528.150 ;
        RECT 71.850 526.950 73.050 530.250 ;
        RECT 92.100 529.350 96.600 531.000 ;
        RECT 70.950 524.850 73.050 526.950 ;
        RECT 95.400 525.150 96.600 529.350 ;
        RECT 113.100 525.150 114.900 526.950 ;
        RECT 65.100 523.050 66.900 524.850 ;
        RECT 70.950 519.600 72.150 524.850 ;
        RECT 73.950 521.850 76.050 523.950 ;
        RECT 85.950 521.850 88.050 523.950 ;
        RECT 91.950 521.850 94.050 523.950 ;
        RECT 94.950 523.050 97.050 525.150 ;
        RECT 112.950 523.050 115.050 525.150 ;
        RECT 116.250 523.950 117.450 531.300 ;
        RECT 119.100 525.150 120.900 526.950 ;
        RECT 131.100 525.150 132.900 526.950 ;
        RECT 73.950 520.050 75.750 521.850 ;
        RECT 86.100 520.050 87.900 521.850 ;
        RECT 50.550 507.750 52.350 513.600 ;
        RECT 53.550 507.750 55.350 513.600 ;
        RECT 66.300 507.750 68.100 519.600 ;
        RECT 70.500 507.750 72.300 519.600 ;
        RECT 88.950 518.850 91.050 520.950 ;
        RECT 92.250 520.050 94.050 521.850 ;
        RECT 89.100 517.050 90.900 518.850 ;
        RECT 95.700 514.800 96.750 523.050 ;
        RECT 115.950 521.850 118.050 523.950 ;
        RECT 118.950 523.050 121.050 525.150 ;
        RECT 130.950 523.050 133.050 525.150 ;
        RECT 134.250 523.950 135.450 531.300 ;
        RECT 153.000 530.250 156.750 531.300 ;
        RECT 173.100 531.000 174.900 539.250 ;
        RECT 149.100 528.150 150.900 529.950 ;
        RECT 137.100 525.150 138.900 526.950 ;
        RECT 133.950 521.850 136.050 523.950 ;
        RECT 136.950 523.050 139.050 525.150 ;
        RECT 145.950 524.850 148.050 526.950 ;
        RECT 148.950 526.050 151.050 528.150 ;
        RECT 152.850 526.950 154.050 530.250 ;
        RECT 151.950 524.850 154.050 526.950 ;
        RECT 170.400 529.350 174.900 531.000 ;
        RECT 178.500 530.400 180.300 539.250 ;
        RECT 188.850 533.400 190.650 539.250 ;
        RECT 193.350 532.200 195.150 539.250 ;
        RECT 191.550 531.300 195.150 532.200 ;
        RECT 170.400 525.150 171.600 529.350 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 146.100 523.050 147.900 524.850 ;
        RECT 89.700 513.900 96.750 514.800 ;
        RECT 89.700 513.600 91.350 513.900 ;
        RECT 73.800 507.750 75.600 513.600 ;
        RECT 86.550 507.750 88.350 513.600 ;
        RECT 89.550 507.750 91.350 513.600 ;
        RECT 95.550 513.600 96.750 513.900 ;
        RECT 116.250 513.600 117.450 521.850 ;
        RECT 134.250 513.600 135.450 521.850 ;
        RECT 151.950 519.600 153.150 524.850 ;
        RECT 154.950 521.850 157.050 523.950 ;
        RECT 169.950 523.050 172.050 525.150 ;
        RECT 154.950 520.050 156.750 521.850 ;
        RECT 92.550 507.750 94.350 513.000 ;
        RECT 95.550 507.750 97.350 513.600 ;
        RECT 112.650 507.750 114.450 513.600 ;
        RECT 115.650 507.750 117.450 513.600 ;
        RECT 118.650 507.750 120.450 513.600 ;
        RECT 130.650 507.750 132.450 513.600 ;
        RECT 133.650 507.750 135.450 513.600 ;
        RECT 136.650 507.750 138.450 513.600 ;
        RECT 147.300 507.750 149.100 519.600 ;
        RECT 151.500 507.750 153.300 519.600 ;
        RECT 170.250 514.800 171.300 523.050 ;
        RECT 172.950 521.850 175.050 523.950 ;
        RECT 178.950 521.850 181.050 523.950 ;
        RECT 172.950 520.050 174.750 521.850 ;
        RECT 175.950 518.850 178.050 520.950 ;
        RECT 179.100 520.050 180.900 521.850 ;
        RECT 182.550 519.450 183.450 526.950 ;
        RECT 188.100 525.150 189.900 526.950 ;
        RECT 187.950 523.050 190.050 525.150 ;
        RECT 191.550 523.950 192.750 531.300 ;
        RECT 212.100 531.000 213.900 539.250 ;
        RECT 209.400 529.350 213.900 531.000 ;
        RECT 217.500 530.400 219.300 539.250 ;
        RECT 227.550 534.300 229.350 539.250 ;
        RECT 230.550 535.200 232.350 539.250 ;
        RECT 233.550 534.300 235.350 539.250 ;
        RECT 227.550 532.950 235.350 534.300 ;
        RECT 236.550 533.400 238.350 539.250 ;
        RECT 251.700 536.400 253.500 539.250 ;
        RECT 255.000 535.050 256.800 539.250 ;
        RECT 251.100 533.400 256.800 535.050 ;
        RECT 259.200 533.400 261.000 539.250 ;
        RECT 236.550 531.300 237.750 533.400 ;
        RECT 234.000 530.250 237.750 531.300 ;
        RECT 194.100 525.150 195.900 526.950 ;
        RECT 209.400 525.150 210.600 529.350 ;
        RECT 230.100 528.150 231.900 529.950 ;
        RECT 190.950 521.850 193.050 523.950 ;
        RECT 193.950 523.050 196.050 525.150 ;
        RECT 208.950 523.050 211.050 525.150 ;
        RECT 226.950 524.850 229.050 526.950 ;
        RECT 229.950 526.050 232.050 528.150 ;
        RECT 233.850 526.950 235.050 530.250 ;
        RECT 251.100 526.950 252.300 533.400 ;
        RECT 275.100 531.000 276.900 539.250 ;
        RECT 254.100 528.150 255.900 529.950 ;
        RECT 232.950 524.850 235.050 526.950 ;
        RECT 250.950 524.850 253.050 526.950 ;
        RECT 253.950 526.050 256.050 528.150 ;
        RECT 256.950 527.850 259.050 529.950 ;
        RECT 260.100 528.150 261.900 529.950 ;
        RECT 272.400 529.350 276.900 531.000 ;
        RECT 280.500 530.400 282.300 539.250 ;
        RECT 291.000 533.400 292.800 539.250 ;
        RECT 295.200 535.050 297.000 539.250 ;
        RECT 298.500 536.400 300.300 539.250 ;
        RECT 295.200 533.400 300.900 535.050 ;
        RECT 313.650 533.400 315.450 539.250 ;
        RECT 257.100 526.050 258.900 527.850 ;
        RECT 259.950 526.050 262.050 528.150 ;
        RECT 272.400 525.150 273.600 529.350 ;
        RECT 290.100 528.150 291.900 529.950 ;
        RECT 289.950 526.050 292.050 528.150 ;
        RECT 292.950 527.850 295.050 529.950 ;
        RECT 296.100 528.150 297.900 529.950 ;
        RECT 293.100 526.050 294.900 527.850 ;
        RECT 295.950 526.050 298.050 528.150 ;
        RECT 299.700 526.950 300.900 533.400 ;
        RECT 314.250 531.300 315.450 533.400 ;
        RECT 316.650 534.300 318.450 539.250 ;
        RECT 319.650 535.200 321.450 539.250 ;
        RECT 322.650 534.300 324.450 539.250 ;
        RECT 316.650 532.950 324.450 534.300 ;
        RECT 335.550 534.300 337.350 539.250 ;
        RECT 338.550 535.200 340.350 539.250 ;
        RECT 341.550 534.300 343.350 539.250 ;
        RECT 335.550 532.950 343.350 534.300 ;
        RECT 344.550 533.400 346.350 539.250 ;
        RECT 359.700 536.400 361.500 539.250 ;
        RECT 363.000 535.050 364.800 539.250 ;
        RECT 359.100 533.400 364.800 535.050 ;
        RECT 367.200 533.400 369.000 539.250 ;
        RECT 381.150 534.900 382.950 539.250 ;
        RECT 379.650 533.400 382.950 534.900 ;
        RECT 384.150 533.400 385.950 539.250 ;
        RECT 322.950 531.450 325.050 532.050 ;
        RECT 328.950 531.450 331.050 532.050 ;
        RECT 314.250 530.250 318.000 531.300 ;
        RECT 322.950 530.550 331.050 531.450 ;
        RECT 344.550 531.300 345.750 533.400 ;
        RECT 316.950 526.950 318.150 530.250 ;
        RECT 322.950 529.950 325.050 530.550 ;
        RECT 328.950 529.950 331.050 530.550 ;
        RECT 342.000 530.250 345.750 531.300 ;
        RECT 320.100 528.150 321.900 529.950 ;
        RECT 338.100 528.150 339.900 529.950 ;
        RECT 187.950 519.450 190.050 520.050 ;
        RECT 176.100 517.050 177.900 518.850 ;
        RECT 182.550 518.550 190.050 519.450 ;
        RECT 187.950 517.950 190.050 518.550 ;
        RECT 170.250 513.900 177.300 514.800 ;
        RECT 170.250 513.600 171.450 513.900 ;
        RECT 154.800 507.750 156.600 513.600 ;
        RECT 169.650 507.750 171.450 513.600 ;
        RECT 175.650 513.600 177.300 513.900 ;
        RECT 191.550 513.600 192.750 521.850 ;
        RECT 209.250 514.800 210.300 523.050 ;
        RECT 211.950 521.850 214.050 523.950 ;
        RECT 217.950 521.850 220.050 523.950 ;
        RECT 227.100 523.050 228.900 524.850 ;
        RECT 211.950 520.050 213.750 521.850 ;
        RECT 214.950 518.850 217.050 520.950 ;
        RECT 218.100 520.050 219.900 521.850 ;
        RECT 232.950 519.600 234.150 524.850 ;
        RECT 235.950 521.850 238.050 523.950 ;
        RECT 235.950 520.050 237.750 521.850 ;
        RECT 251.100 519.600 252.300 524.850 ;
        RECT 271.950 523.050 274.050 525.150 ;
        RECT 298.950 524.850 301.050 526.950 ;
        RECT 316.950 524.850 319.050 526.950 ;
        RECT 319.950 526.050 322.050 528.150 ;
        RECT 322.950 524.850 325.050 526.950 ;
        RECT 334.950 524.850 337.050 526.950 ;
        RECT 337.950 526.050 340.050 528.150 ;
        RECT 341.850 526.950 343.050 530.250 ;
        RECT 359.100 526.950 360.300 533.400 ;
        RECT 362.100 528.150 363.900 529.950 ;
        RECT 340.950 524.850 343.050 526.950 ;
        RECT 358.950 524.850 361.050 526.950 ;
        RECT 361.950 526.050 364.050 528.150 ;
        RECT 364.950 527.850 367.050 529.950 ;
        RECT 368.100 528.150 369.900 529.950 ;
        RECT 365.100 526.050 366.900 527.850 ;
        RECT 367.950 526.050 370.050 528.150 ;
        RECT 379.650 526.950 380.850 533.400 ;
        RECT 382.950 531.900 384.750 532.500 ;
        RECT 388.650 531.900 390.450 539.250 ;
        RECT 398.850 533.400 400.650 539.250 ;
        RECT 403.350 532.200 405.150 539.250 ;
        RECT 418.650 533.400 420.450 539.250 ;
        RECT 382.950 530.700 390.450 531.900 ;
        RECT 401.550 531.300 405.150 532.200 ;
        RECT 419.250 531.300 420.450 533.400 ;
        RECT 421.650 534.300 423.450 539.250 ;
        RECT 424.650 535.200 426.450 539.250 ;
        RECT 427.650 534.300 429.450 539.250 ;
        RECT 421.650 532.950 429.450 534.300 ;
        RECT 442.350 533.400 444.150 539.250 ;
        RECT 445.350 533.400 447.150 539.250 ;
        RECT 448.650 536.400 450.450 539.250 ;
        RECT 379.650 524.850 382.050 526.950 ;
        RECT 383.100 525.150 384.900 526.950 ;
        RECT 215.100 517.050 216.900 518.850 ;
        RECT 209.250 513.900 216.300 514.800 ;
        RECT 209.250 513.600 210.450 513.900 ;
        RECT 172.650 507.750 174.450 513.000 ;
        RECT 175.650 507.750 177.450 513.600 ;
        RECT 178.650 507.750 180.450 513.600 ;
        RECT 188.550 507.750 190.350 513.600 ;
        RECT 191.550 507.750 193.350 513.600 ;
        RECT 194.550 507.750 196.350 513.600 ;
        RECT 208.650 507.750 210.450 513.600 ;
        RECT 214.650 513.600 216.300 513.900 ;
        RECT 211.650 507.750 213.450 513.000 ;
        RECT 214.650 507.750 216.450 513.600 ;
        RECT 217.650 507.750 219.450 513.600 ;
        RECT 228.300 507.750 230.100 519.600 ;
        RECT 232.500 507.750 234.300 519.600 ;
        RECT 235.800 507.750 237.600 513.600 ;
        RECT 250.650 507.750 252.450 519.600 ;
        RECT 253.650 518.700 261.450 519.600 ;
        RECT 253.650 507.750 255.450 518.700 ;
        RECT 256.650 507.750 258.450 517.800 ;
        RECT 259.650 507.750 261.450 518.700 ;
        RECT 272.250 514.800 273.300 523.050 ;
        RECT 274.950 521.850 277.050 523.950 ;
        RECT 280.950 521.850 283.050 523.950 ;
        RECT 274.950 520.050 276.750 521.850 ;
        RECT 277.950 518.850 280.050 520.950 ;
        RECT 281.100 520.050 282.900 521.850 ;
        RECT 299.700 519.600 300.900 524.850 ;
        RECT 313.950 521.850 316.050 523.950 ;
        RECT 314.250 520.050 316.050 521.850 ;
        RECT 317.850 519.600 319.050 524.850 ;
        RECT 323.100 523.050 324.900 524.850 ;
        RECT 335.100 523.050 336.900 524.850 ;
        RECT 340.950 519.600 342.150 524.850 ;
        RECT 343.950 521.850 346.050 523.950 ;
        RECT 343.950 520.050 345.750 521.850 ;
        RECT 359.100 519.600 360.300 524.850 ;
        RECT 379.650 519.600 380.850 524.850 ;
        RECT 382.950 523.050 385.050 525.150 ;
        RECT 278.100 517.050 279.900 518.850 ;
        RECT 290.550 518.700 298.350 519.600 ;
        RECT 272.250 513.900 279.300 514.800 ;
        RECT 272.250 513.600 273.450 513.900 ;
        RECT 271.650 507.750 273.450 513.600 ;
        RECT 277.650 513.600 279.300 513.900 ;
        RECT 274.650 507.750 276.450 513.000 ;
        RECT 277.650 507.750 279.450 513.600 ;
        RECT 280.650 507.750 282.450 513.600 ;
        RECT 290.550 507.750 292.350 518.700 ;
        RECT 293.550 507.750 295.350 517.800 ;
        RECT 296.550 507.750 298.350 518.700 ;
        RECT 299.550 507.750 301.350 519.600 ;
        RECT 314.400 507.750 316.200 513.600 ;
        RECT 317.700 507.750 319.500 519.600 ;
        RECT 321.900 507.750 323.700 519.600 ;
        RECT 336.300 507.750 338.100 519.600 ;
        RECT 340.500 507.750 342.300 519.600 ;
        RECT 343.800 507.750 345.600 513.600 ;
        RECT 358.650 507.750 360.450 519.600 ;
        RECT 361.650 518.700 369.450 519.600 ;
        RECT 361.650 507.750 363.450 518.700 ;
        RECT 364.650 507.750 366.450 517.800 ;
        RECT 367.650 507.750 369.450 518.700 ;
        RECT 379.050 507.750 380.850 519.600 ;
        RECT 382.050 507.750 383.850 519.600 ;
        RECT 386.100 513.600 387.300 530.700 ;
        RECT 388.950 524.850 391.050 526.950 ;
        RECT 398.100 525.150 399.900 526.950 ;
        RECT 389.100 523.050 390.900 524.850 ;
        RECT 397.950 523.050 400.050 525.150 ;
        RECT 401.550 523.950 402.750 531.300 ;
        RECT 419.250 530.250 423.000 531.300 ;
        RECT 421.950 526.950 423.150 530.250 ;
        RECT 425.100 528.150 426.900 529.950 ;
        RECT 404.100 525.150 405.900 526.950 ;
        RECT 400.950 521.850 403.050 523.950 ;
        RECT 403.950 523.050 406.050 525.150 ;
        RECT 421.950 524.850 424.050 526.950 ;
        RECT 424.950 526.050 427.050 528.150 ;
        RECT 442.650 526.950 443.850 533.400 ;
        RECT 448.650 532.500 449.850 536.400 ;
        RECT 444.750 531.600 449.850 532.500 ;
        RECT 461.850 532.200 463.650 539.250 ;
        RECT 466.350 533.400 468.150 539.250 ;
        RECT 444.750 530.700 447.000 531.600 ;
        RECT 461.850 531.300 465.450 532.200 ;
        RECT 427.950 524.850 430.050 526.950 ;
        RECT 442.650 524.850 445.050 526.950 ;
        RECT 418.950 521.850 421.050 523.950 ;
        RECT 401.550 513.600 402.750 521.850 ;
        RECT 419.250 520.050 421.050 521.850 ;
        RECT 422.850 519.600 424.050 524.850 ;
        RECT 428.100 523.050 429.900 524.850 ;
        RECT 442.650 519.600 443.850 524.850 ;
        RECT 445.950 522.300 447.000 530.700 ;
        RECT 448.950 524.850 451.050 526.950 ;
        RECT 461.100 525.150 462.900 526.950 ;
        RECT 449.100 523.050 450.900 524.850 ;
        RECT 460.950 523.050 463.050 525.150 ;
        RECT 464.250 523.950 465.450 531.300 ;
        RECT 476.700 530.400 478.500 539.250 ;
        RECT 482.100 531.000 483.900 539.250 ;
        RECT 503.100 531.000 504.900 539.250 ;
        RECT 482.100 529.350 486.600 531.000 ;
        RECT 467.100 525.150 468.900 526.950 ;
        RECT 485.400 525.150 486.600 529.350 ;
        RECT 500.400 529.350 504.900 531.000 ;
        RECT 508.500 530.400 510.300 539.250 ;
        RECT 520.650 533.400 522.450 539.250 ;
        RECT 521.250 531.300 522.450 533.400 ;
        RECT 523.650 534.300 525.450 539.250 ;
        RECT 526.650 535.200 528.450 539.250 ;
        RECT 529.650 534.300 531.450 539.250 ;
        RECT 523.650 532.950 531.450 534.300 ;
        RECT 541.650 533.400 543.450 539.250 ;
        RECT 542.250 531.300 543.450 533.400 ;
        RECT 544.650 534.300 546.450 539.250 ;
        RECT 547.650 535.200 549.450 539.250 ;
        RECT 550.650 534.300 552.450 539.250 ;
        RECT 564.150 534.900 565.950 539.250 ;
        RECT 544.650 532.950 552.450 534.300 ;
        RECT 562.650 533.400 565.950 534.900 ;
        RECT 567.150 533.400 568.950 539.250 ;
        RECT 521.250 530.250 525.000 531.300 ;
        RECT 542.250 530.250 546.000 531.300 ;
        RECT 500.400 525.150 501.600 529.350 ;
        RECT 508.950 528.450 511.050 529.050 ;
        RECT 514.950 528.450 517.050 529.050 ;
        RECT 508.950 527.550 517.050 528.450 ;
        RECT 508.950 526.950 511.050 527.550 ;
        RECT 514.950 526.950 517.050 527.550 ;
        RECT 523.950 526.950 525.150 530.250 ;
        RECT 527.100 528.150 528.900 529.950 ;
        RECT 444.750 521.400 447.000 522.300 ;
        RECT 463.950 521.850 466.050 523.950 ;
        RECT 466.950 523.050 469.050 525.150 ;
        RECT 475.950 521.850 478.050 523.950 ;
        RECT 481.950 521.850 484.050 523.950 ;
        RECT 484.950 523.050 487.050 525.150 ;
        RECT 499.950 523.050 502.050 525.150 ;
        RECT 523.950 524.850 526.050 526.950 ;
        RECT 526.950 526.050 529.050 528.150 ;
        RECT 544.950 526.950 546.150 530.250 ;
        RECT 548.100 528.150 549.900 529.950 ;
        RECT 529.950 524.850 532.050 526.950 ;
        RECT 544.950 524.850 547.050 526.950 ;
        RECT 547.950 526.050 550.050 528.150 ;
        RECT 562.650 526.950 563.850 533.400 ;
        RECT 565.950 531.900 567.750 532.500 ;
        RECT 571.650 531.900 573.450 539.250 ;
        RECT 581.550 536.400 583.350 539.250 ;
        RECT 584.550 536.400 586.350 539.250 ;
        RECT 587.550 536.400 589.350 539.250 ;
        RECT 565.950 530.700 573.450 531.900 ;
        RECT 550.950 524.850 553.050 526.950 ;
        RECT 562.650 524.850 565.050 526.950 ;
        RECT 566.100 525.150 567.900 526.950 ;
        RECT 444.750 520.500 450.450 521.400 ;
        RECT 385.650 507.750 387.450 513.600 ;
        RECT 388.650 507.750 390.450 513.600 ;
        RECT 398.550 507.750 400.350 513.600 ;
        RECT 401.550 507.750 403.350 513.600 ;
        RECT 404.550 507.750 406.350 513.600 ;
        RECT 419.400 507.750 421.200 513.600 ;
        RECT 422.700 507.750 424.500 519.600 ;
        RECT 426.900 507.750 428.700 519.600 ;
        RECT 442.350 507.750 444.150 519.600 ;
        RECT 445.350 507.750 447.150 519.600 ;
        RECT 449.250 513.600 450.450 520.500 ;
        RECT 464.250 513.600 465.450 521.850 ;
        RECT 476.100 520.050 477.900 521.850 ;
        RECT 478.950 518.850 481.050 520.950 ;
        RECT 482.250 520.050 484.050 521.850 ;
        RECT 479.100 517.050 480.900 518.850 ;
        RECT 485.700 514.800 486.750 523.050 ;
        RECT 479.700 513.900 486.750 514.800 ;
        RECT 479.700 513.600 481.350 513.900 ;
        RECT 448.650 507.750 450.450 513.600 ;
        RECT 460.650 507.750 462.450 513.600 ;
        RECT 463.650 507.750 465.450 513.600 ;
        RECT 466.650 507.750 468.450 513.600 ;
        RECT 476.550 507.750 478.350 513.600 ;
        RECT 479.550 507.750 481.350 513.600 ;
        RECT 485.550 513.600 486.750 513.900 ;
        RECT 500.250 514.800 501.300 523.050 ;
        RECT 502.950 521.850 505.050 523.950 ;
        RECT 508.950 521.850 511.050 523.950 ;
        RECT 520.950 521.850 523.050 523.950 ;
        RECT 502.950 520.050 504.750 521.850 ;
        RECT 505.950 518.850 508.050 520.950 ;
        RECT 509.100 520.050 510.900 521.850 ;
        RECT 521.250 520.050 523.050 521.850 ;
        RECT 524.850 519.600 526.050 524.850 ;
        RECT 530.100 523.050 531.900 524.850 ;
        RECT 541.950 521.850 544.050 523.950 ;
        RECT 542.250 520.050 544.050 521.850 ;
        RECT 545.850 519.600 547.050 524.850 ;
        RECT 551.100 523.050 552.900 524.850 ;
        RECT 562.650 519.600 563.850 524.850 ;
        RECT 565.950 523.050 568.050 525.150 ;
        RECT 506.100 517.050 507.900 518.850 ;
        RECT 500.250 513.900 507.300 514.800 ;
        RECT 500.250 513.600 501.450 513.900 ;
        RECT 482.550 507.750 484.350 513.000 ;
        RECT 485.550 507.750 487.350 513.600 ;
        RECT 499.650 507.750 501.450 513.600 ;
        RECT 505.650 513.600 507.300 513.900 ;
        RECT 502.650 507.750 504.450 513.000 ;
        RECT 505.650 507.750 507.450 513.600 ;
        RECT 508.650 507.750 510.450 513.600 ;
        RECT 521.400 507.750 523.200 513.600 ;
        RECT 524.700 507.750 526.500 519.600 ;
        RECT 528.900 507.750 530.700 519.600 ;
        RECT 542.400 507.750 544.200 513.600 ;
        RECT 545.700 507.750 547.500 519.600 ;
        RECT 549.900 507.750 551.700 519.600 ;
        RECT 562.050 507.750 563.850 519.600 ;
        RECT 565.050 507.750 566.850 519.600 ;
        RECT 569.100 513.600 570.300 530.700 ;
        RECT 585.000 529.950 586.050 536.400 ;
        RECT 604.650 533.400 606.450 539.250 ;
        RECT 605.250 531.300 606.450 533.400 ;
        RECT 607.650 534.300 609.450 539.250 ;
        RECT 610.650 535.200 612.450 539.250 ;
        RECT 613.650 534.300 615.450 539.250 ;
        RECT 623.550 536.400 625.350 539.250 ;
        RECT 626.550 536.400 628.350 539.250 ;
        RECT 607.650 532.950 615.450 534.300 ;
        RECT 605.250 530.250 609.000 531.300 ;
        RECT 583.950 527.850 586.050 529.950 ;
        RECT 571.950 524.850 574.050 526.950 ;
        RECT 580.950 524.850 583.050 526.950 ;
        RECT 572.100 523.050 573.900 524.850 ;
        RECT 581.100 523.050 582.900 524.850 ;
        RECT 585.000 520.650 586.050 527.850 ;
        RECT 607.950 526.950 609.150 530.250 ;
        RECT 611.100 528.150 612.900 529.950 ;
        RECT 586.950 524.850 589.050 526.950 ;
        RECT 607.950 524.850 610.050 526.950 ;
        RECT 610.950 526.050 613.050 528.150 ;
        RECT 622.950 527.850 625.050 529.950 ;
        RECT 626.400 528.150 627.600 536.400 ;
        RECT 638.550 534.300 640.350 539.250 ;
        RECT 641.550 535.200 643.350 539.250 ;
        RECT 644.550 534.300 646.350 539.250 ;
        RECT 638.550 532.950 646.350 534.300 ;
        RECT 647.550 533.400 649.350 539.250 ;
        RECT 647.550 531.300 648.750 533.400 ;
        RECT 662.850 532.200 664.650 539.250 ;
        RECT 667.350 533.400 669.150 539.250 ;
        RECT 677.850 533.400 679.650 539.250 ;
        RECT 682.350 532.200 684.150 539.250 ;
        RECT 645.000 530.250 648.750 531.300 ;
        RECT 649.950 531.450 652.050 532.050 ;
        RECT 658.950 531.450 661.050 532.050 ;
        RECT 649.950 530.550 661.050 531.450 ;
        RECT 662.850 531.300 666.450 532.200 ;
        RECT 641.100 528.150 642.900 529.950 ;
        RECT 613.950 524.850 616.050 526.950 ;
        RECT 623.100 526.050 624.900 527.850 ;
        RECT 625.950 526.050 628.050 528.150 ;
        RECT 587.100 523.050 588.900 524.850 ;
        RECT 604.950 521.850 607.050 523.950 ;
        RECT 585.000 519.600 587.550 520.650 ;
        RECT 605.250 520.050 607.050 521.850 ;
        RECT 608.850 519.600 610.050 524.850 ;
        RECT 614.100 523.050 615.900 524.850 ;
        RECT 568.650 507.750 570.450 513.600 ;
        RECT 571.650 507.750 573.450 513.600 ;
        RECT 581.550 507.750 583.350 519.600 ;
        RECT 585.750 507.750 587.550 519.600 ;
        RECT 605.400 507.750 607.200 513.600 ;
        RECT 608.700 507.750 610.500 519.600 ;
        RECT 612.900 507.750 614.700 519.600 ;
        RECT 626.400 513.600 627.600 526.050 ;
        RECT 637.950 524.850 640.050 526.950 ;
        RECT 640.950 526.050 643.050 528.150 ;
        RECT 644.850 526.950 646.050 530.250 ;
        RECT 649.950 529.950 652.050 530.550 ;
        RECT 658.950 529.950 661.050 530.550 ;
        RECT 643.950 524.850 646.050 526.950 ;
        RECT 662.100 525.150 663.900 526.950 ;
        RECT 638.100 523.050 639.900 524.850 ;
        RECT 643.950 519.600 645.150 524.850 ;
        RECT 646.950 521.850 649.050 523.950 ;
        RECT 661.950 523.050 664.050 525.150 ;
        RECT 665.250 523.950 666.450 531.300 ;
        RECT 680.550 531.300 684.150 532.200 ;
        RECT 689.550 533.400 691.350 539.250 ;
        RECT 692.850 536.400 694.650 539.250 ;
        RECT 697.350 536.400 699.150 539.250 ;
        RECT 701.550 536.400 703.350 539.250 ;
        RECT 705.450 536.400 707.250 539.250 ;
        RECT 708.750 536.400 710.550 539.250 ;
        RECT 713.250 537.300 715.050 539.250 ;
        RECT 713.250 536.400 717.000 537.300 ;
        RECT 718.050 536.400 719.850 539.250 ;
        RECT 697.650 535.500 698.700 536.400 ;
        RECT 694.950 534.300 698.700 535.500 ;
        RECT 706.200 534.600 707.250 536.400 ;
        RECT 715.950 535.500 717.000 536.400 ;
        RECT 694.950 533.400 697.050 534.300 ;
        RECT 668.100 525.150 669.900 526.950 ;
        RECT 677.100 525.150 678.900 526.950 ;
        RECT 664.950 521.850 667.050 523.950 ;
        RECT 667.950 523.050 670.050 525.150 ;
        RECT 676.950 523.050 679.050 525.150 ;
        RECT 680.550 523.950 681.750 531.300 ;
        RECT 689.550 531.150 690.750 533.400 ;
        RECT 702.150 532.200 703.950 534.000 ;
        RECT 706.200 533.550 711.150 534.600 ;
        RECT 709.350 532.800 711.150 533.550 ;
        RECT 712.650 532.800 714.450 534.600 ;
        RECT 715.950 533.400 718.050 535.500 ;
        RECT 721.050 533.400 722.850 539.250 ;
        RECT 703.050 531.900 703.950 532.200 ;
        RECT 713.100 531.900 714.150 532.800 ;
        RECT 689.550 529.050 694.050 531.150 ;
        RECT 703.050 531.000 714.150 531.900 ;
        RECT 683.100 525.150 684.900 526.950 ;
        RECT 679.950 521.850 682.050 523.950 ;
        RECT 682.950 523.050 685.050 525.150 ;
        RECT 646.950 520.050 648.750 521.850 ;
        RECT 623.550 507.750 625.350 513.600 ;
        RECT 626.550 507.750 628.350 513.600 ;
        RECT 639.300 507.750 641.100 519.600 ;
        RECT 643.500 507.750 645.300 519.600 ;
        RECT 665.250 513.600 666.450 521.850 ;
        RECT 680.550 513.600 681.750 521.850 ;
        RECT 689.550 519.600 690.750 529.050 ;
        RECT 691.950 527.250 695.850 529.050 ;
        RECT 691.950 526.950 694.050 527.250 ;
        RECT 703.050 526.950 703.950 531.000 ;
        RECT 713.100 529.800 714.150 531.000 ;
        RECT 713.100 528.600 720.000 529.800 ;
        RECT 713.100 528.000 714.900 528.600 ;
        RECT 719.100 527.850 720.000 528.600 ;
        RECT 716.100 526.950 717.900 527.700 ;
        RECT 703.050 524.850 706.050 526.950 ;
        RECT 709.950 525.900 717.900 526.950 ;
        RECT 719.100 526.050 720.900 527.850 ;
        RECT 709.950 524.850 712.050 525.900 ;
        RECT 691.950 521.400 693.750 523.200 ;
        RECT 692.850 520.200 697.050 521.400 ;
        RECT 703.050 520.200 703.950 524.850 ;
        RECT 711.750 521.100 713.550 521.400 ;
        RECT 646.800 507.750 648.600 513.600 ;
        RECT 661.650 507.750 663.450 513.600 ;
        RECT 664.650 507.750 666.450 513.600 ;
        RECT 667.650 507.750 669.450 513.600 ;
        RECT 677.550 507.750 679.350 513.600 ;
        RECT 680.550 507.750 682.350 513.600 ;
        RECT 683.550 507.750 685.350 513.600 ;
        RECT 689.550 507.750 691.350 519.600 ;
        RECT 694.950 519.300 697.050 520.200 ;
        RECT 697.950 519.300 703.950 520.200 ;
        RECT 705.150 520.800 713.550 521.100 ;
        RECT 721.950 520.800 722.850 533.400 ;
        RECT 734.850 532.200 736.650 539.250 ;
        RECT 739.350 533.400 741.150 539.250 ;
        RECT 751.650 533.400 753.450 539.250 ;
        RECT 734.850 531.300 738.450 532.200 ;
        RECT 734.100 525.150 735.900 526.950 ;
        RECT 733.950 523.050 736.050 525.150 ;
        RECT 737.250 523.950 738.450 531.300 ;
        RECT 752.250 531.300 753.450 533.400 ;
        RECT 754.650 534.300 756.450 539.250 ;
        RECT 757.650 535.200 759.450 539.250 ;
        RECT 760.650 534.300 762.450 539.250 ;
        RECT 754.650 532.950 762.450 534.300 ;
        RECT 773.850 533.400 775.650 539.250 ;
        RECT 778.350 532.200 780.150 539.250 ;
        RECT 776.550 531.300 780.150 532.200 ;
        RECT 786.150 533.400 787.950 539.250 ;
        RECT 789.150 536.400 790.950 539.250 ;
        RECT 793.950 537.300 795.750 539.250 ;
        RECT 792.000 536.400 795.750 537.300 ;
        RECT 798.450 536.400 800.250 539.250 ;
        RECT 801.750 536.400 803.550 539.250 ;
        RECT 805.650 536.400 807.450 539.250 ;
        RECT 809.850 536.400 811.650 539.250 ;
        RECT 814.350 536.400 816.150 539.250 ;
        RECT 792.000 535.500 793.050 536.400 ;
        RECT 790.950 533.400 793.050 535.500 ;
        RECT 801.750 534.600 802.800 536.400 ;
        RECT 752.250 530.250 756.000 531.300 ;
        RECT 754.950 526.950 756.150 530.250 ;
        RECT 758.100 528.150 759.900 529.950 ;
        RECT 740.100 525.150 741.900 526.950 ;
        RECT 736.950 521.850 739.050 523.950 ;
        RECT 739.950 523.050 742.050 525.150 ;
        RECT 754.950 524.850 757.050 526.950 ;
        RECT 757.950 526.050 760.050 528.150 ;
        RECT 760.950 524.850 763.050 526.950 ;
        RECT 773.100 525.150 774.900 526.950 ;
        RECT 751.950 521.850 754.050 523.950 ;
        RECT 705.150 520.200 722.850 520.800 ;
        RECT 697.950 518.400 698.850 519.300 ;
        RECT 696.150 516.600 698.850 518.400 ;
        RECT 699.750 518.100 701.550 518.400 ;
        RECT 705.150 518.100 706.050 520.200 ;
        RECT 711.750 519.600 722.850 520.200 ;
        RECT 699.750 517.200 706.050 518.100 ;
        RECT 706.950 518.700 708.750 519.300 ;
        RECT 706.950 517.500 714.450 518.700 ;
        RECT 699.750 516.600 701.550 517.200 ;
        RECT 713.250 516.600 714.450 517.500 ;
        RECT 694.950 513.600 698.850 515.700 ;
        RECT 703.950 514.500 710.850 516.300 ;
        RECT 713.250 514.500 718.050 516.600 ;
        RECT 692.550 507.750 694.350 510.600 ;
        RECT 697.050 507.750 698.850 513.600 ;
        RECT 701.250 507.750 703.050 513.600 ;
        RECT 705.150 507.750 706.950 514.500 ;
        RECT 713.250 513.600 714.450 514.500 ;
        RECT 708.150 507.750 709.950 513.600 ;
        RECT 712.950 507.750 714.750 513.600 ;
        RECT 718.050 507.750 719.850 513.600 ;
        RECT 721.050 507.750 722.850 519.600 ;
        RECT 737.250 513.600 738.450 521.850 ;
        RECT 752.250 520.050 754.050 521.850 ;
        RECT 755.850 519.600 757.050 524.850 ;
        RECT 761.100 523.050 762.900 524.850 ;
        RECT 772.950 523.050 775.050 525.150 ;
        RECT 776.550 523.950 777.750 531.300 ;
        RECT 779.100 525.150 780.900 526.950 ;
        RECT 775.950 521.850 778.050 523.950 ;
        RECT 778.950 523.050 781.050 525.150 ;
        RECT 733.650 507.750 735.450 513.600 ;
        RECT 736.650 507.750 738.450 513.600 ;
        RECT 739.650 507.750 741.450 513.600 ;
        RECT 752.400 507.750 754.200 513.600 ;
        RECT 755.700 507.750 757.500 519.600 ;
        RECT 759.900 507.750 761.700 519.600 ;
        RECT 776.550 513.600 777.750 521.850 ;
        RECT 786.150 520.800 787.050 533.400 ;
        RECT 794.550 532.800 796.350 534.600 ;
        RECT 797.850 533.550 802.800 534.600 ;
        RECT 810.300 535.500 811.350 536.400 ;
        RECT 810.300 534.300 814.050 535.500 ;
        RECT 797.850 532.800 799.650 533.550 ;
        RECT 794.850 531.900 795.900 532.800 ;
        RECT 805.050 532.200 806.850 534.000 ;
        RECT 811.950 533.400 814.050 534.300 ;
        RECT 817.650 533.400 819.450 539.250 ;
        RECT 805.050 531.900 805.950 532.200 ;
        RECT 794.850 531.000 805.950 531.900 ;
        RECT 818.250 531.150 819.450 533.400 ;
        RECT 830.850 532.200 832.650 539.250 ;
        RECT 835.350 533.400 837.150 539.250 ;
        RECT 845.550 534.300 847.350 539.250 ;
        RECT 848.550 535.200 850.350 539.250 ;
        RECT 851.550 534.300 853.350 539.250 ;
        RECT 845.550 532.950 853.350 534.300 ;
        RECT 854.550 533.400 856.350 539.250 ;
        RECT 830.850 531.300 834.450 532.200 ;
        RECT 854.550 531.300 855.750 533.400 ;
        RECT 794.850 529.800 795.900 531.000 ;
        RECT 789.000 528.600 795.900 529.800 ;
        RECT 789.000 527.850 789.900 528.600 ;
        RECT 794.100 528.000 795.900 528.600 ;
        RECT 788.100 526.050 789.900 527.850 ;
        RECT 791.100 526.950 792.900 527.700 ;
        RECT 805.050 526.950 805.950 531.000 ;
        RECT 814.950 529.050 819.450 531.150 ;
        RECT 813.150 527.250 817.050 529.050 ;
        RECT 814.950 526.950 817.050 527.250 ;
        RECT 791.100 525.900 799.050 526.950 ;
        RECT 796.950 524.850 799.050 525.900 ;
        RECT 802.950 524.850 805.950 526.950 ;
        RECT 795.450 521.100 797.250 521.400 ;
        RECT 795.450 520.800 803.850 521.100 ;
        RECT 786.150 520.200 803.850 520.800 ;
        RECT 786.150 519.600 797.250 520.200 ;
        RECT 773.550 507.750 775.350 513.600 ;
        RECT 776.550 507.750 778.350 513.600 ;
        RECT 779.550 507.750 781.350 513.600 ;
        RECT 786.150 507.750 787.950 519.600 ;
        RECT 800.250 518.700 802.050 519.300 ;
        RECT 794.550 517.500 802.050 518.700 ;
        RECT 802.950 518.100 803.850 520.200 ;
        RECT 805.050 520.200 805.950 524.850 ;
        RECT 815.250 521.400 817.050 523.200 ;
        RECT 811.950 520.200 816.150 521.400 ;
        RECT 805.050 519.300 811.050 520.200 ;
        RECT 811.950 519.300 814.050 520.200 ;
        RECT 818.250 519.600 819.450 529.050 ;
        RECT 830.100 525.150 831.900 526.950 ;
        RECT 829.950 523.050 832.050 525.150 ;
        RECT 833.250 523.950 834.450 531.300 ;
        RECT 852.000 530.250 855.750 531.300 ;
        RECT 848.100 528.150 849.900 529.950 ;
        RECT 836.100 525.150 837.900 526.950 ;
        RECT 832.950 521.850 835.050 523.950 ;
        RECT 835.950 523.050 838.050 525.150 ;
        RECT 844.950 524.850 847.050 526.950 ;
        RECT 847.950 526.050 850.050 528.150 ;
        RECT 851.850 526.950 853.050 530.250 ;
        RECT 850.950 524.850 853.050 526.950 ;
        RECT 845.100 523.050 846.900 524.850 ;
        RECT 810.150 518.400 811.050 519.300 ;
        RECT 807.450 518.100 809.250 518.400 ;
        RECT 794.550 516.600 795.750 517.500 ;
        RECT 802.950 517.200 809.250 518.100 ;
        RECT 807.450 516.600 809.250 517.200 ;
        RECT 810.150 516.600 812.850 518.400 ;
        RECT 790.950 514.500 795.750 516.600 ;
        RECT 798.150 514.500 805.050 516.300 ;
        RECT 794.550 513.600 795.750 514.500 ;
        RECT 789.150 507.750 790.950 513.600 ;
        RECT 794.250 507.750 796.050 513.600 ;
        RECT 799.050 507.750 800.850 513.600 ;
        RECT 802.050 507.750 803.850 514.500 ;
        RECT 810.150 513.600 814.050 515.700 ;
        RECT 805.950 507.750 807.750 513.600 ;
        RECT 810.150 507.750 811.950 513.600 ;
        RECT 814.650 507.750 816.450 510.600 ;
        RECT 817.650 507.750 819.450 519.600 ;
        RECT 833.250 513.600 834.450 521.850 ;
        RECT 850.950 519.600 852.150 524.850 ;
        RECT 853.950 521.850 856.050 523.950 ;
        RECT 853.950 520.050 855.750 521.850 ;
        RECT 829.650 507.750 831.450 513.600 ;
        RECT 832.650 507.750 834.450 513.600 ;
        RECT 835.650 507.750 837.450 513.600 ;
        RECT 846.300 507.750 848.100 519.600 ;
        RECT 850.500 507.750 852.300 519.600 ;
        RECT 853.800 507.750 855.600 513.600 ;
        RECT 10.650 497.400 12.450 503.250 ;
        RECT 13.650 497.400 15.450 503.250 ;
        RECT 26.400 497.400 28.200 503.250 ;
        RECT 11.400 484.950 12.600 497.400 ;
        RECT 29.700 491.400 31.500 503.250 ;
        RECT 33.900 491.400 35.700 503.250 ;
        RECT 46.650 497.400 48.450 503.250 ;
        RECT 49.650 497.400 51.450 503.250 ;
        RECT 59.550 497.400 61.350 503.250 ;
        RECT 62.550 497.400 64.350 503.250 ;
        RECT 65.550 497.400 67.350 503.250 ;
        RECT 13.950 489.450 16.050 490.050 ;
        RECT 13.950 488.550 18.450 489.450 ;
        RECT 26.250 489.150 28.050 490.950 ;
        RECT 13.950 487.950 16.050 488.550 ;
        RECT 10.950 482.850 13.050 484.950 ;
        RECT 14.100 483.150 15.900 484.950 ;
        RECT 11.400 474.600 12.600 482.850 ;
        RECT 13.950 481.050 16.050 483.150 ;
        RECT 13.950 477.450 16.050 478.050 ;
        RECT 17.550 477.450 18.450 488.550 ;
        RECT 25.950 487.050 28.050 489.150 ;
        RECT 29.850 486.150 31.050 491.400 ;
        RECT 35.100 486.150 36.900 487.950 ;
        RECT 28.950 484.050 31.050 486.150 ;
        RECT 28.950 480.750 30.150 484.050 ;
        RECT 31.950 482.850 34.050 484.950 ;
        RECT 34.950 484.050 37.050 486.150 ;
        RECT 47.400 484.950 48.600 497.400 ;
        RECT 62.550 489.150 63.750 497.400 ;
        RECT 77.550 492.300 79.350 503.250 ;
        RECT 80.550 493.200 82.350 503.250 ;
        RECT 83.550 492.300 85.350 503.250 ;
        RECT 77.550 491.400 85.350 492.300 ;
        RECT 86.550 491.400 88.350 503.250 ;
        RECT 98.550 497.400 100.350 503.250 ;
        RECT 101.550 497.400 103.350 503.250 ;
        RECT 58.950 485.850 61.050 487.950 ;
        RECT 61.950 487.050 64.050 489.150 ;
        RECT 46.950 482.850 49.050 484.950 ;
        RECT 50.100 483.150 51.900 484.950 ;
        RECT 59.100 484.050 60.900 485.850 ;
        RECT 32.100 481.050 33.900 482.850 ;
        RECT 26.250 479.700 30.000 480.750 ;
        RECT 26.250 477.600 27.450 479.700 ;
        RECT 13.950 476.550 18.450 477.450 ;
        RECT 13.950 475.950 16.050 476.550 ;
        RECT 10.650 471.750 12.450 474.600 ;
        RECT 13.650 471.750 15.450 474.600 ;
        RECT 25.650 471.750 27.450 477.600 ;
        RECT 28.650 476.700 36.450 478.050 ;
        RECT 28.650 471.750 30.450 476.700 ;
        RECT 31.650 471.750 33.450 475.800 ;
        RECT 34.650 471.750 36.450 476.700 ;
        RECT 47.400 474.600 48.600 482.850 ;
        RECT 49.950 481.050 52.050 483.150 ;
        RECT 62.550 479.700 63.750 487.050 ;
        RECT 64.950 485.850 67.050 487.950 ;
        RECT 86.700 486.150 87.900 491.400 ;
        RECT 98.100 486.150 99.900 487.950 ;
        RECT 65.100 484.050 66.900 485.850 ;
        RECT 76.950 482.850 79.050 484.950 ;
        RECT 80.100 483.150 81.900 484.950 ;
        RECT 77.100 481.050 78.900 482.850 ;
        RECT 79.950 481.050 82.050 483.150 ;
        RECT 82.950 482.850 85.050 484.950 ;
        RECT 85.950 484.050 88.050 486.150 ;
        RECT 97.950 484.050 100.050 486.150 ;
        RECT 83.100 481.050 84.900 482.850 ;
        RECT 62.550 478.800 66.150 479.700 ;
        RECT 46.650 471.750 48.450 474.600 ;
        RECT 49.650 471.750 51.450 474.600 ;
        RECT 59.850 471.750 61.650 477.600 ;
        RECT 64.350 471.750 66.150 478.800 ;
        RECT 86.700 477.600 87.900 484.050 ;
        RECT 101.700 480.300 102.900 497.400 ;
        RECT 105.150 491.400 106.950 503.250 ;
        RECT 108.150 491.400 109.950 503.250 ;
        RECT 124.650 497.400 126.450 503.250 ;
        RECT 127.650 497.400 129.450 503.250 ;
        RECT 130.650 497.400 132.450 503.250 ;
        RECT 142.650 497.400 144.450 503.250 ;
        RECT 145.650 498.000 147.450 503.250 ;
        RECT 103.950 485.850 106.050 487.950 ;
        RECT 108.150 486.150 109.350 491.400 ;
        RECT 128.250 489.150 129.450 497.400 ;
        RECT 143.250 497.100 144.450 497.400 ;
        RECT 148.650 497.400 150.450 503.250 ;
        RECT 151.650 497.400 153.450 503.250 ;
        RECT 163.650 497.400 165.450 503.250 ;
        RECT 166.650 498.000 168.450 503.250 ;
        RECT 148.650 497.100 150.300 497.400 ;
        RECT 143.250 496.200 150.300 497.100 ;
        RECT 164.250 497.100 165.450 497.400 ;
        RECT 169.650 497.400 171.450 503.250 ;
        RECT 172.650 497.400 174.450 503.250 ;
        RECT 169.650 497.100 171.300 497.400 ;
        RECT 164.250 496.200 171.300 497.100 ;
        RECT 104.100 484.050 105.900 485.850 ;
        RECT 106.950 484.050 109.350 486.150 ;
        RECT 124.950 485.850 127.050 487.950 ;
        RECT 127.950 487.050 130.050 489.150 ;
        RECT 143.250 487.950 144.300 496.200 ;
        RECT 149.100 492.150 150.900 493.950 ;
        RECT 145.950 489.150 147.750 490.950 ;
        RECT 148.950 490.050 151.050 492.150 ;
        RECT 152.100 489.150 153.900 490.950 ;
        RECT 125.100 484.050 126.900 485.850 ;
        RECT 78.000 471.750 79.800 477.600 ;
        RECT 82.200 475.950 87.900 477.600 ;
        RECT 98.550 479.100 106.050 480.300 ;
        RECT 82.200 471.750 84.000 475.950 ;
        RECT 85.500 471.750 87.300 474.600 ;
        RECT 98.550 471.750 100.350 479.100 ;
        RECT 104.250 478.500 106.050 479.100 ;
        RECT 108.150 477.600 109.350 484.050 ;
        RECT 128.250 479.700 129.450 487.050 ;
        RECT 130.950 485.850 133.050 487.950 ;
        RECT 142.950 485.850 145.050 487.950 ;
        RECT 145.950 487.050 148.050 489.150 ;
        RECT 151.950 487.050 154.050 489.150 ;
        RECT 164.250 487.950 165.300 496.200 ;
        RECT 170.100 492.150 171.900 493.950 ;
        RECT 182.550 492.300 184.350 503.250 ;
        RECT 185.550 493.200 187.350 503.250 ;
        RECT 188.550 492.300 190.350 503.250 ;
        RECT 166.950 489.150 168.750 490.950 ;
        RECT 169.950 490.050 172.050 492.150 ;
        RECT 182.550 491.400 190.350 492.300 ;
        RECT 191.550 491.400 193.350 503.250 ;
        RECT 205.650 497.400 207.450 503.250 ;
        RECT 208.650 497.400 210.450 503.250 ;
        RECT 220.650 497.400 222.450 503.250 ;
        RECT 223.650 498.000 225.450 503.250 ;
        RECT 173.100 489.150 174.900 490.950 ;
        RECT 163.950 485.850 166.050 487.950 ;
        RECT 166.950 487.050 169.050 489.150 ;
        RECT 172.950 487.050 175.050 489.150 ;
        RECT 191.700 486.150 192.900 491.400 ;
        RECT 131.100 484.050 132.900 485.850 ;
        RECT 143.400 481.650 144.600 485.850 ;
        RECT 164.400 481.650 165.600 485.850 ;
        RECT 181.950 482.850 184.050 484.950 ;
        RECT 185.100 483.150 186.900 484.950 ;
        RECT 143.400 480.000 147.900 481.650 ;
        RECT 103.050 471.750 104.850 477.600 ;
        RECT 106.050 476.100 109.350 477.600 ;
        RECT 125.850 478.800 129.450 479.700 ;
        RECT 106.050 471.750 107.850 476.100 ;
        RECT 125.850 471.750 127.650 478.800 ;
        RECT 130.350 471.750 132.150 477.600 ;
        RECT 146.100 471.750 147.900 480.000 ;
        RECT 151.500 471.750 153.300 480.600 ;
        RECT 164.400 480.000 168.900 481.650 ;
        RECT 182.100 481.050 183.900 482.850 ;
        RECT 184.950 481.050 187.050 483.150 ;
        RECT 187.950 482.850 190.050 484.950 ;
        RECT 190.950 484.050 193.050 486.150 ;
        RECT 206.400 484.950 207.600 497.400 ;
        RECT 221.250 497.100 222.450 497.400 ;
        RECT 226.650 497.400 228.450 503.250 ;
        RECT 229.650 497.400 231.450 503.250 ;
        RECT 241.650 497.400 243.450 503.250 ;
        RECT 244.650 498.000 246.450 503.250 ;
        RECT 226.650 497.100 228.300 497.400 ;
        RECT 221.250 496.200 228.300 497.100 ;
        RECT 242.250 497.100 243.450 497.400 ;
        RECT 247.650 497.400 249.450 503.250 ;
        RECT 250.650 497.400 252.450 503.250 ;
        RECT 247.650 497.100 249.300 497.400 ;
        RECT 242.250 496.200 249.300 497.100 ;
        RECT 221.250 487.950 222.300 496.200 ;
        RECT 227.100 492.150 228.900 493.950 ;
        RECT 223.950 489.150 225.750 490.950 ;
        RECT 226.950 490.050 229.050 492.150 ;
        RECT 230.100 489.150 231.900 490.950 ;
        RECT 220.950 485.850 223.050 487.950 ;
        RECT 223.950 487.050 226.050 489.150 ;
        RECT 229.950 487.050 232.050 489.150 ;
        RECT 242.250 487.950 243.300 496.200 ;
        RECT 248.100 492.150 249.900 493.950 ;
        RECT 244.950 489.150 246.750 490.950 ;
        RECT 247.950 490.050 250.050 492.150 ;
        RECT 262.650 491.400 264.450 503.250 ;
        RECT 265.650 492.300 267.450 503.250 ;
        RECT 268.650 493.200 270.450 503.250 ;
        RECT 271.650 492.300 273.450 503.250 ;
        RECT 286.650 497.400 288.450 503.250 ;
        RECT 289.650 497.400 291.450 503.250 ;
        RECT 292.650 497.400 294.450 503.250 ;
        RECT 277.950 495.450 280.050 496.050 ;
        RECT 283.950 495.450 286.050 496.050 ;
        RECT 277.950 494.550 286.050 495.450 ;
        RECT 277.950 493.950 280.050 494.550 ;
        RECT 283.950 493.950 286.050 494.550 ;
        RECT 265.650 491.400 273.450 492.300 ;
        RECT 251.100 489.150 252.900 490.950 ;
        RECT 241.950 485.850 244.050 487.950 ;
        RECT 244.950 487.050 247.050 489.150 ;
        RECT 250.950 487.050 253.050 489.150 ;
        RECT 263.100 486.150 264.300 491.400 ;
        RECT 290.250 489.150 291.450 497.400 ;
        RECT 304.650 491.400 306.450 503.250 ;
        RECT 307.650 492.300 309.450 503.250 ;
        RECT 310.650 493.200 312.450 503.250 ;
        RECT 313.650 492.300 315.450 503.250 ;
        RECT 323.550 497.400 325.350 503.250 ;
        RECT 326.550 497.400 328.350 503.250 ;
        RECT 329.550 497.400 331.350 503.250 ;
        RECT 307.650 491.400 315.450 492.300 ;
        RECT 188.100 481.050 189.900 482.850 ;
        RECT 167.100 471.750 168.900 480.000 ;
        RECT 172.500 471.750 174.300 480.600 ;
        RECT 191.700 477.600 192.900 484.050 ;
        RECT 205.950 482.850 208.050 484.950 ;
        RECT 209.100 483.150 210.900 484.950 ;
        RECT 183.000 471.750 184.800 477.600 ;
        RECT 187.200 475.950 192.900 477.600 ;
        RECT 187.200 471.750 189.000 475.950 ;
        RECT 206.400 474.600 207.600 482.850 ;
        RECT 208.950 481.050 211.050 483.150 ;
        RECT 221.400 481.650 222.600 485.850 ;
        RECT 242.400 481.650 243.600 485.850 ;
        RECT 262.950 484.050 265.050 486.150 ;
        RECT 286.950 485.850 289.050 487.950 ;
        RECT 289.950 487.050 292.050 489.150 ;
        RECT 221.400 480.000 225.900 481.650 ;
        RECT 190.500 471.750 192.300 474.600 ;
        RECT 205.650 471.750 207.450 474.600 ;
        RECT 208.650 471.750 210.450 474.600 ;
        RECT 224.100 471.750 225.900 480.000 ;
        RECT 229.500 471.750 231.300 480.600 ;
        RECT 242.400 480.000 246.900 481.650 ;
        RECT 245.100 471.750 246.900 480.000 ;
        RECT 250.500 471.750 252.300 480.600 ;
        RECT 263.100 477.600 264.300 484.050 ;
        RECT 265.950 482.850 268.050 484.950 ;
        RECT 269.100 483.150 270.900 484.950 ;
        RECT 266.100 481.050 267.900 482.850 ;
        RECT 268.950 481.050 271.050 483.150 ;
        RECT 271.950 482.850 274.050 484.950 ;
        RECT 287.100 484.050 288.900 485.850 ;
        RECT 272.100 481.050 273.900 482.850 ;
        RECT 290.250 479.700 291.450 487.050 ;
        RECT 292.950 485.850 295.050 487.950 ;
        RECT 305.100 486.150 306.300 491.400 ;
        RECT 326.550 489.150 327.750 497.400 ;
        RECT 343.050 491.400 344.850 503.250 ;
        RECT 346.050 491.400 347.850 503.250 ;
        RECT 349.650 497.400 351.450 503.250 ;
        RECT 352.650 497.400 354.450 503.250 ;
        RECT 362.550 497.400 364.350 503.250 ;
        RECT 365.550 497.400 367.350 503.250 ;
        RECT 368.550 497.400 370.350 503.250 ;
        RECT 383.400 497.400 385.200 503.250 ;
        RECT 293.100 484.050 294.900 485.850 ;
        RECT 304.950 484.050 307.050 486.150 ;
        RECT 322.950 485.850 325.050 487.950 ;
        RECT 325.950 487.050 328.050 489.150 ;
        RECT 287.850 478.800 291.450 479.700 ;
        RECT 263.100 475.950 268.800 477.600 ;
        RECT 263.700 471.750 265.500 474.600 ;
        RECT 267.000 471.750 268.800 475.950 ;
        RECT 271.200 471.750 273.000 477.600 ;
        RECT 287.850 471.750 289.650 478.800 ;
        RECT 305.100 477.600 306.300 484.050 ;
        RECT 307.950 482.850 310.050 484.950 ;
        RECT 311.100 483.150 312.900 484.950 ;
        RECT 308.100 481.050 309.900 482.850 ;
        RECT 310.950 481.050 313.050 483.150 ;
        RECT 313.950 482.850 316.050 484.950 ;
        RECT 323.100 484.050 324.900 485.850 ;
        RECT 314.100 481.050 315.900 482.850 ;
        RECT 326.550 479.700 327.750 487.050 ;
        RECT 328.950 485.850 331.050 487.950 ;
        RECT 343.650 486.150 344.850 491.400 ;
        RECT 329.100 484.050 330.900 485.850 ;
        RECT 343.650 484.050 346.050 486.150 ;
        RECT 346.950 485.850 349.050 487.950 ;
        RECT 347.100 484.050 348.900 485.850 ;
        RECT 326.550 478.800 330.150 479.700 ;
        RECT 292.350 471.750 294.150 477.600 ;
        RECT 305.100 475.950 310.800 477.600 ;
        RECT 305.700 471.750 307.500 474.600 ;
        RECT 309.000 471.750 310.800 475.950 ;
        RECT 313.200 471.750 315.000 477.600 ;
        RECT 323.850 471.750 325.650 477.600 ;
        RECT 328.350 471.750 330.150 478.800 ;
        RECT 343.650 477.600 344.850 484.050 ;
        RECT 350.100 480.300 351.300 497.400 ;
        RECT 365.550 489.150 366.750 497.400 ;
        RECT 386.700 491.400 388.500 503.250 ;
        RECT 390.900 491.400 392.700 503.250 ;
        RECT 403.650 491.400 405.450 503.250 ;
        RECT 406.650 492.300 408.450 503.250 ;
        RECT 409.650 493.200 411.450 503.250 ;
        RECT 412.650 492.300 414.450 503.250 ;
        RECT 422.550 497.400 424.350 503.250 ;
        RECT 425.550 497.400 427.350 503.250 ;
        RECT 428.550 498.000 430.350 503.250 ;
        RECT 425.700 497.100 427.350 497.400 ;
        RECT 431.550 497.400 433.350 503.250 ;
        RECT 443.550 497.400 445.350 503.250 ;
        RECT 446.550 497.400 448.350 503.250 ;
        RECT 449.550 498.000 451.350 503.250 ;
        RECT 431.550 497.100 432.750 497.400 ;
        RECT 425.700 496.200 432.750 497.100 ;
        RECT 446.700 497.100 448.350 497.400 ;
        RECT 452.550 497.400 454.350 503.250 ;
        RECT 466.650 497.400 468.450 503.250 ;
        RECT 469.650 497.400 471.450 503.250 ;
        RECT 472.650 497.400 474.450 503.250 ;
        RECT 487.650 497.400 489.450 503.250 ;
        RECT 490.650 497.400 492.450 503.250 ;
        RECT 493.650 497.400 495.450 503.250 ;
        RECT 503.550 497.400 505.350 503.250 ;
        RECT 506.550 497.400 508.350 503.250 ;
        RECT 520.650 497.400 522.450 503.250 ;
        RECT 523.650 498.000 525.450 503.250 ;
        RECT 452.550 497.100 453.750 497.400 ;
        RECT 446.700 496.200 453.750 497.100 ;
        RECT 406.650 491.400 414.450 492.300 ;
        RECT 425.100 492.150 426.900 493.950 ;
        RECT 383.250 489.150 385.050 490.950 ;
        RECT 353.100 486.150 354.900 487.950 ;
        RECT 352.950 484.050 355.050 486.150 ;
        RECT 361.950 485.850 364.050 487.950 ;
        RECT 364.950 487.050 367.050 489.150 ;
        RECT 362.100 484.050 363.900 485.850 ;
        RECT 346.950 479.100 354.450 480.300 ;
        RECT 346.950 478.500 348.750 479.100 ;
        RECT 343.650 476.100 346.950 477.600 ;
        RECT 345.150 471.750 346.950 476.100 ;
        RECT 348.150 471.750 349.950 477.600 ;
        RECT 352.650 471.750 354.450 479.100 ;
        RECT 365.550 479.700 366.750 487.050 ;
        RECT 367.950 485.850 370.050 487.950 ;
        RECT 382.950 487.050 385.050 489.150 ;
        RECT 386.850 486.150 388.050 491.400 ;
        RECT 392.100 486.150 393.900 487.950 ;
        RECT 404.100 486.150 405.300 491.400 ;
        RECT 422.100 489.150 423.900 490.950 ;
        RECT 424.950 490.050 427.050 492.150 ;
        RECT 428.250 489.150 430.050 490.950 ;
        RECT 421.950 487.050 424.050 489.150 ;
        RECT 427.950 487.050 430.050 489.150 ;
        RECT 431.700 487.950 432.750 496.200 ;
        RECT 446.100 492.150 447.900 493.950 ;
        RECT 443.100 489.150 444.900 490.950 ;
        RECT 445.950 490.050 448.050 492.150 ;
        RECT 449.250 489.150 451.050 490.950 ;
        RECT 368.100 484.050 369.900 485.850 ;
        RECT 385.950 484.050 388.050 486.150 ;
        RECT 385.950 480.750 387.150 484.050 ;
        RECT 388.950 482.850 391.050 484.950 ;
        RECT 391.950 484.050 394.050 486.150 ;
        RECT 403.950 484.050 406.050 486.150 ;
        RECT 430.950 485.850 433.050 487.950 ;
        RECT 442.950 487.050 445.050 489.150 ;
        RECT 448.950 487.050 451.050 489.150 ;
        RECT 452.700 487.950 453.750 496.200 ;
        RECT 470.250 489.150 471.450 497.400 ;
        RECT 491.250 489.150 492.450 497.400 ;
        RECT 451.950 485.850 454.050 487.950 ;
        RECT 466.950 485.850 469.050 487.950 ;
        RECT 469.950 487.050 472.050 489.150 ;
        RECT 389.100 481.050 390.900 482.850 ;
        RECT 383.250 479.700 387.000 480.750 ;
        RECT 365.550 478.800 369.150 479.700 ;
        RECT 362.850 471.750 364.650 477.600 ;
        RECT 367.350 471.750 369.150 478.800 ;
        RECT 383.250 477.600 384.450 479.700 ;
        RECT 382.650 471.750 384.450 477.600 ;
        RECT 385.650 476.700 393.450 478.050 ;
        RECT 385.650 471.750 387.450 476.700 ;
        RECT 388.650 471.750 390.450 475.800 ;
        RECT 391.650 471.750 393.450 476.700 ;
        RECT 404.100 477.600 405.300 484.050 ;
        RECT 406.950 482.850 409.050 484.950 ;
        RECT 410.100 483.150 411.900 484.950 ;
        RECT 407.100 481.050 408.900 482.850 ;
        RECT 409.950 481.050 412.050 483.150 ;
        RECT 412.950 482.850 415.050 484.950 ;
        RECT 418.950 483.450 421.050 484.050 ;
        RECT 424.950 483.450 427.050 484.050 ;
        RECT 413.100 481.050 414.900 482.850 ;
        RECT 418.950 482.550 427.050 483.450 ;
        RECT 418.950 481.950 421.050 482.550 ;
        RECT 424.950 481.950 427.050 482.550 ;
        RECT 431.400 481.650 432.600 485.850 ;
        RECT 439.950 483.450 442.050 484.050 ;
        RECT 445.950 483.450 448.050 484.050 ;
        RECT 439.950 482.550 448.050 483.450 ;
        RECT 439.950 481.950 442.050 482.550 ;
        RECT 445.950 481.950 448.050 482.550 ;
        RECT 452.400 481.650 453.600 485.850 ;
        RECT 467.100 484.050 468.900 485.850 ;
        RECT 404.100 475.950 409.800 477.600 ;
        RECT 404.700 471.750 406.500 474.600 ;
        RECT 408.000 471.750 409.800 475.950 ;
        RECT 412.200 471.750 414.000 477.600 ;
        RECT 422.700 471.750 424.500 480.600 ;
        RECT 428.100 480.000 432.600 481.650 ;
        RECT 428.100 471.750 429.900 480.000 ;
        RECT 430.950 477.450 433.050 478.050 ;
        RECT 439.950 477.450 442.050 478.050 ;
        RECT 430.950 476.550 442.050 477.450 ;
        RECT 430.950 475.950 433.050 476.550 ;
        RECT 439.950 475.950 442.050 476.550 ;
        RECT 443.700 471.750 445.500 480.600 ;
        RECT 449.100 480.000 453.600 481.650 ;
        RECT 449.100 471.750 450.900 480.000 ;
        RECT 470.250 479.700 471.450 487.050 ;
        RECT 472.950 485.850 475.050 487.950 ;
        RECT 487.950 485.850 490.050 487.950 ;
        RECT 490.950 487.050 493.050 489.150 ;
        RECT 473.100 484.050 474.900 485.850 ;
        RECT 488.100 484.050 489.900 485.850 ;
        RECT 491.250 479.700 492.450 487.050 ;
        RECT 493.950 485.850 496.050 487.950 ;
        RECT 494.100 484.050 495.900 485.850 ;
        RECT 506.400 484.950 507.600 497.400 ;
        RECT 521.250 497.100 522.450 497.400 ;
        RECT 526.650 497.400 528.450 503.250 ;
        RECT 529.650 497.400 531.450 503.250 ;
        RECT 526.650 497.100 528.300 497.400 ;
        RECT 521.250 496.200 528.300 497.100 ;
        RECT 521.250 487.950 522.300 496.200 ;
        RECT 527.100 492.150 528.900 493.950 ;
        RECT 539.550 492.300 541.350 503.250 ;
        RECT 542.550 493.200 544.350 503.250 ;
        RECT 545.550 492.300 547.350 503.250 ;
        RECT 523.950 489.150 525.750 490.950 ;
        RECT 526.950 490.050 529.050 492.150 ;
        RECT 539.550 491.400 547.350 492.300 ;
        RECT 548.550 491.400 550.350 503.250 ;
        RECT 563.400 497.400 565.200 503.250 ;
        RECT 566.700 491.400 568.500 503.250 ;
        RECT 570.900 491.400 572.700 503.250 ;
        RECT 581.550 497.400 583.350 503.250 ;
        RECT 584.550 497.400 586.350 503.250 ;
        RECT 530.100 489.150 531.900 490.950 ;
        RECT 520.950 485.850 523.050 487.950 ;
        RECT 523.950 487.050 526.050 489.150 ;
        RECT 529.950 487.050 532.050 489.150 ;
        RECT 548.700 486.150 549.900 491.400 ;
        RECT 563.250 489.150 565.050 490.950 ;
        RECT 562.950 487.050 565.050 489.150 ;
        RECT 566.850 486.150 568.050 491.400 ;
        RECT 572.100 486.150 573.900 487.950 ;
        RECT 503.100 483.150 504.900 484.950 ;
        RECT 502.950 481.050 505.050 483.150 ;
        RECT 505.950 482.850 508.050 484.950 ;
        RECT 467.850 478.800 471.450 479.700 ;
        RECT 488.850 478.800 492.450 479.700 ;
        RECT 467.850 471.750 469.650 478.800 ;
        RECT 472.350 471.750 474.150 477.600 ;
        RECT 488.850 471.750 490.650 478.800 ;
        RECT 493.350 471.750 495.150 477.600 ;
        RECT 506.400 474.600 507.600 482.850 ;
        RECT 521.400 481.650 522.600 485.850 ;
        RECT 538.950 482.850 541.050 484.950 ;
        RECT 542.100 483.150 543.900 484.950 ;
        RECT 521.400 480.000 525.900 481.650 ;
        RECT 539.100 481.050 540.900 482.850 ;
        RECT 541.950 481.050 544.050 483.150 ;
        RECT 544.950 482.850 547.050 484.950 ;
        RECT 547.950 484.050 550.050 486.150 ;
        RECT 565.950 484.050 568.050 486.150 ;
        RECT 545.100 481.050 546.900 482.850 ;
        RECT 503.550 471.750 505.350 474.600 ;
        RECT 506.550 471.750 508.350 474.600 ;
        RECT 524.100 471.750 525.900 480.000 ;
        RECT 529.500 471.750 531.300 480.600 ;
        RECT 548.700 477.600 549.900 484.050 ;
        RECT 565.950 480.750 567.150 484.050 ;
        RECT 568.950 482.850 571.050 484.950 ;
        RECT 571.950 484.050 574.050 486.150 ;
        RECT 584.400 484.950 585.600 497.400 ;
        RECT 590.550 491.400 592.350 503.250 ;
        RECT 593.550 500.400 595.350 503.250 ;
        RECT 598.050 497.400 599.850 503.250 ;
        RECT 602.250 497.400 604.050 503.250 ;
        RECT 595.950 495.300 599.850 497.400 ;
        RECT 606.150 496.500 607.950 503.250 ;
        RECT 609.150 497.400 610.950 503.250 ;
        RECT 613.950 497.400 615.750 503.250 ;
        RECT 619.050 497.400 620.850 503.250 ;
        RECT 614.250 496.500 615.450 497.400 ;
        RECT 604.950 494.700 611.850 496.500 ;
        RECT 614.250 494.400 619.050 496.500 ;
        RECT 597.150 492.600 599.850 494.400 ;
        RECT 600.750 493.800 602.550 494.400 ;
        RECT 600.750 492.900 607.050 493.800 ;
        RECT 614.250 493.500 615.450 494.400 ;
        RECT 600.750 492.600 602.550 492.900 ;
        RECT 598.950 491.700 599.850 492.600 ;
        RECT 581.100 483.150 582.900 484.950 ;
        RECT 569.100 481.050 570.900 482.850 ;
        RECT 580.950 481.050 583.050 483.150 ;
        RECT 583.950 482.850 586.050 484.950 ;
        RECT 563.250 479.700 567.000 480.750 ;
        RECT 563.250 477.600 564.450 479.700 ;
        RECT 540.000 471.750 541.800 477.600 ;
        RECT 544.200 475.950 549.900 477.600 ;
        RECT 544.200 471.750 546.000 475.950 ;
        RECT 547.500 471.750 549.300 474.600 ;
        RECT 562.650 471.750 564.450 477.600 ;
        RECT 565.650 476.700 573.450 478.050 ;
        RECT 565.650 471.750 567.450 476.700 ;
        RECT 568.650 471.750 570.450 475.800 ;
        RECT 571.650 471.750 573.450 476.700 ;
        RECT 584.400 474.600 585.600 482.850 ;
        RECT 590.550 481.950 591.750 491.400 ;
        RECT 595.950 490.800 598.050 491.700 ;
        RECT 598.950 490.800 604.950 491.700 ;
        RECT 593.850 489.600 598.050 490.800 ;
        RECT 592.950 487.800 594.750 489.600 ;
        RECT 604.050 486.150 604.950 490.800 ;
        RECT 606.150 490.800 607.050 492.900 ;
        RECT 607.950 492.300 615.450 493.500 ;
        RECT 607.950 491.700 609.750 492.300 ;
        RECT 622.050 491.400 623.850 503.250 ;
        RECT 633.300 491.400 635.100 503.250 ;
        RECT 637.500 491.400 639.300 503.250 ;
        RECT 640.800 497.400 642.600 503.250 ;
        RECT 654.300 491.400 656.100 503.250 ;
        RECT 658.500 491.400 660.300 503.250 ;
        RECT 661.800 497.400 663.600 503.250 ;
        RECT 668.550 491.400 670.350 503.250 ;
        RECT 671.550 500.400 673.350 503.250 ;
        RECT 676.050 497.400 677.850 503.250 ;
        RECT 680.250 497.400 682.050 503.250 ;
        RECT 673.950 495.300 677.850 497.400 ;
        RECT 684.150 496.500 685.950 503.250 ;
        RECT 687.150 497.400 688.950 503.250 ;
        RECT 691.950 497.400 693.750 503.250 ;
        RECT 697.050 497.400 698.850 503.250 ;
        RECT 692.250 496.500 693.450 497.400 ;
        RECT 682.950 494.700 689.850 496.500 ;
        RECT 692.250 494.400 697.050 496.500 ;
        RECT 675.150 492.600 677.850 494.400 ;
        RECT 678.750 493.800 680.550 494.400 ;
        RECT 678.750 492.900 685.050 493.800 ;
        RECT 692.250 493.500 693.450 494.400 ;
        RECT 678.750 492.600 680.550 492.900 ;
        RECT 676.950 491.700 677.850 492.600 ;
        RECT 612.750 490.800 623.850 491.400 ;
        RECT 606.150 490.200 623.850 490.800 ;
        RECT 606.150 489.900 614.550 490.200 ;
        RECT 612.750 489.600 614.550 489.900 ;
        RECT 604.050 484.050 607.050 486.150 ;
        RECT 610.950 485.100 613.050 486.150 ;
        RECT 610.950 484.050 618.900 485.100 ;
        RECT 592.950 483.750 595.050 484.050 ;
        RECT 592.950 481.950 596.850 483.750 ;
        RECT 590.550 479.850 595.050 481.950 ;
        RECT 604.050 480.000 604.950 484.050 ;
        RECT 617.100 483.300 618.900 484.050 ;
        RECT 620.100 483.150 621.900 484.950 ;
        RECT 614.100 482.400 615.900 483.000 ;
        RECT 620.100 482.400 621.000 483.150 ;
        RECT 614.100 481.200 621.000 482.400 ;
        RECT 614.100 480.000 615.150 481.200 ;
        RECT 590.550 477.600 591.750 479.850 ;
        RECT 604.050 479.100 615.150 480.000 ;
        RECT 604.050 478.800 604.950 479.100 ;
        RECT 581.550 471.750 583.350 474.600 ;
        RECT 584.550 471.750 586.350 474.600 ;
        RECT 590.550 471.750 592.350 477.600 ;
        RECT 595.950 476.700 598.050 477.600 ;
        RECT 603.150 477.000 604.950 478.800 ;
        RECT 614.100 478.200 615.150 479.100 ;
        RECT 610.350 477.450 612.150 478.200 ;
        RECT 595.950 475.500 599.700 476.700 ;
        RECT 598.650 474.600 599.700 475.500 ;
        RECT 607.200 476.400 612.150 477.450 ;
        RECT 613.650 476.400 615.450 478.200 ;
        RECT 622.950 477.600 623.850 490.200 ;
        RECT 632.100 486.150 633.900 487.950 ;
        RECT 637.950 486.150 639.150 491.400 ;
        RECT 640.950 489.150 642.750 490.950 ;
        RECT 640.950 487.050 643.050 489.150 ;
        RECT 653.100 486.150 654.900 487.950 ;
        RECT 658.950 486.150 660.150 491.400 ;
        RECT 661.950 489.150 663.750 490.950 ;
        RECT 661.950 487.050 664.050 489.150 ;
        RECT 631.950 484.050 634.050 486.150 ;
        RECT 634.950 482.850 637.050 484.950 ;
        RECT 637.950 484.050 640.050 486.150 ;
        RECT 652.950 484.050 655.050 486.150 ;
        RECT 635.100 481.050 636.900 482.850 ;
        RECT 638.850 480.750 640.050 484.050 ;
        RECT 655.950 482.850 658.050 484.950 ;
        RECT 658.950 484.050 661.050 486.150 ;
        RECT 656.100 481.050 657.900 482.850 ;
        RECT 659.850 480.750 661.050 484.050 ;
        RECT 668.550 481.950 669.750 491.400 ;
        RECT 673.950 490.800 676.050 491.700 ;
        RECT 676.950 490.800 682.950 491.700 ;
        RECT 671.850 489.600 676.050 490.800 ;
        RECT 670.950 487.800 672.750 489.600 ;
        RECT 682.050 486.150 682.950 490.800 ;
        RECT 684.150 490.800 685.050 492.900 ;
        RECT 685.950 492.300 693.450 493.500 ;
        RECT 685.950 491.700 687.750 492.300 ;
        RECT 700.050 491.400 701.850 503.250 ;
        RECT 711.300 491.400 713.100 503.250 ;
        RECT 715.500 491.400 717.300 503.250 ;
        RECT 718.800 497.400 720.600 503.250 ;
        RECT 733.650 497.400 735.450 503.250 ;
        RECT 736.650 497.400 738.450 503.250 ;
        RECT 739.650 497.400 741.450 503.250 ;
        RECT 752.400 497.400 754.200 503.250 ;
        RECT 690.750 490.800 701.850 491.400 ;
        RECT 684.150 490.200 701.850 490.800 ;
        RECT 684.150 489.900 692.550 490.200 ;
        RECT 690.750 489.600 692.550 489.900 ;
        RECT 682.050 484.050 685.050 486.150 ;
        RECT 688.950 485.100 691.050 486.150 ;
        RECT 688.950 484.050 696.900 485.100 ;
        RECT 670.950 483.750 673.050 484.050 ;
        RECT 670.950 481.950 674.850 483.750 ;
        RECT 639.000 479.700 642.750 480.750 ;
        RECT 660.000 479.700 663.750 480.750 ;
        RECT 607.200 474.600 608.250 476.400 ;
        RECT 616.950 475.500 619.050 477.600 ;
        RECT 616.950 474.600 618.000 475.500 ;
        RECT 593.850 471.750 595.650 474.600 ;
        RECT 598.350 471.750 600.150 474.600 ;
        RECT 602.550 471.750 604.350 474.600 ;
        RECT 606.450 471.750 608.250 474.600 ;
        RECT 609.750 471.750 611.550 474.600 ;
        RECT 614.250 473.700 618.000 474.600 ;
        RECT 614.250 471.750 616.050 473.700 ;
        RECT 619.050 471.750 620.850 474.600 ;
        RECT 622.050 471.750 623.850 477.600 ;
        RECT 632.550 476.700 640.350 478.050 ;
        RECT 632.550 471.750 634.350 476.700 ;
        RECT 635.550 471.750 637.350 475.800 ;
        RECT 638.550 471.750 640.350 476.700 ;
        RECT 641.550 477.600 642.750 479.700 ;
        RECT 641.550 471.750 643.350 477.600 ;
        RECT 653.550 476.700 661.350 478.050 ;
        RECT 653.550 471.750 655.350 476.700 ;
        RECT 656.550 471.750 658.350 475.800 ;
        RECT 659.550 471.750 661.350 476.700 ;
        RECT 662.550 477.600 663.750 479.700 ;
        RECT 668.550 479.850 673.050 481.950 ;
        RECT 682.050 480.000 682.950 484.050 ;
        RECT 695.100 483.300 696.900 484.050 ;
        RECT 698.100 483.150 699.900 484.950 ;
        RECT 692.100 482.400 693.900 483.000 ;
        RECT 698.100 482.400 699.000 483.150 ;
        RECT 692.100 481.200 699.000 482.400 ;
        RECT 692.100 480.000 693.150 481.200 ;
        RECT 668.550 477.600 669.750 479.850 ;
        RECT 682.050 479.100 693.150 480.000 ;
        RECT 682.050 478.800 682.950 479.100 ;
        RECT 662.550 471.750 664.350 477.600 ;
        RECT 668.550 471.750 670.350 477.600 ;
        RECT 673.950 476.700 676.050 477.600 ;
        RECT 681.150 477.000 682.950 478.800 ;
        RECT 692.100 478.200 693.150 479.100 ;
        RECT 688.350 477.450 690.150 478.200 ;
        RECT 673.950 475.500 677.700 476.700 ;
        RECT 676.650 474.600 677.700 475.500 ;
        RECT 685.200 476.400 690.150 477.450 ;
        RECT 691.650 476.400 693.450 478.200 ;
        RECT 700.950 477.600 701.850 490.200 ;
        RECT 710.100 486.150 711.900 487.950 ;
        RECT 715.950 486.150 717.150 491.400 ;
        RECT 718.950 489.150 720.750 490.950 ;
        RECT 737.250 489.150 738.450 497.400 ;
        RECT 755.700 491.400 757.500 503.250 ;
        RECT 759.900 491.400 761.700 503.250 ;
        RECT 772.650 497.400 774.450 503.250 ;
        RECT 775.650 497.400 777.450 503.250 ;
        RECT 787.650 497.400 789.450 503.250 ;
        RECT 790.650 497.400 792.450 503.250 ;
        RECT 793.650 497.400 795.450 503.250 ;
        RECT 803.550 497.400 805.350 503.250 ;
        RECT 806.550 497.400 808.350 503.250 ;
        RECT 752.250 489.150 754.050 490.950 ;
        RECT 718.950 487.050 721.050 489.150 ;
        RECT 709.950 484.050 712.050 486.150 ;
        RECT 712.950 482.850 715.050 484.950 ;
        RECT 715.950 484.050 718.050 486.150 ;
        RECT 733.950 485.850 736.050 487.950 ;
        RECT 736.950 487.050 739.050 489.150 ;
        RECT 734.100 484.050 735.900 485.850 ;
        RECT 713.100 481.050 714.900 482.850 ;
        RECT 716.850 480.750 718.050 484.050 ;
        RECT 717.000 479.700 720.750 480.750 ;
        RECT 737.250 479.700 738.450 487.050 ;
        RECT 739.950 485.850 742.050 487.950 ;
        RECT 751.950 487.050 754.050 489.150 ;
        RECT 755.850 486.150 757.050 491.400 ;
        RECT 761.100 486.150 762.900 487.950 ;
        RECT 740.100 484.050 741.900 485.850 ;
        RECT 754.950 484.050 757.050 486.150 ;
        RECT 754.950 480.750 756.150 484.050 ;
        RECT 757.950 482.850 760.050 484.950 ;
        RECT 760.950 484.050 763.050 486.150 ;
        RECT 773.400 484.950 774.600 497.400 ;
        RECT 791.250 489.150 792.450 497.400 ;
        RECT 787.950 485.850 790.050 487.950 ;
        RECT 790.950 487.050 793.050 489.150 ;
        RECT 772.950 482.850 775.050 484.950 ;
        RECT 776.100 483.150 777.900 484.950 ;
        RECT 788.100 484.050 789.900 485.850 ;
        RECT 758.100 481.050 759.900 482.850 ;
        RECT 685.200 474.600 686.250 476.400 ;
        RECT 694.950 475.500 697.050 477.600 ;
        RECT 694.950 474.600 696.000 475.500 ;
        RECT 671.850 471.750 673.650 474.600 ;
        RECT 676.350 471.750 678.150 474.600 ;
        RECT 680.550 471.750 682.350 474.600 ;
        RECT 684.450 471.750 686.250 474.600 ;
        RECT 687.750 471.750 689.550 474.600 ;
        RECT 692.250 473.700 696.000 474.600 ;
        RECT 692.250 471.750 694.050 473.700 ;
        RECT 697.050 471.750 698.850 474.600 ;
        RECT 700.050 471.750 701.850 477.600 ;
        RECT 710.550 476.700 718.350 478.050 ;
        RECT 710.550 471.750 712.350 476.700 ;
        RECT 713.550 471.750 715.350 475.800 ;
        RECT 716.550 471.750 718.350 476.700 ;
        RECT 719.550 477.600 720.750 479.700 ;
        RECT 734.850 478.800 738.450 479.700 ;
        RECT 752.250 479.700 756.000 480.750 ;
        RECT 719.550 471.750 721.350 477.600 ;
        RECT 734.850 471.750 736.650 478.800 ;
        RECT 752.250 477.600 753.450 479.700 ;
        RECT 739.350 471.750 741.150 477.600 ;
        RECT 751.650 471.750 753.450 477.600 ;
        RECT 754.650 476.700 762.450 478.050 ;
        RECT 754.650 471.750 756.450 476.700 ;
        RECT 757.650 471.750 759.450 475.800 ;
        RECT 760.650 471.750 762.450 476.700 ;
        RECT 773.400 474.600 774.600 482.850 ;
        RECT 775.950 481.050 778.050 483.150 ;
        RECT 791.250 479.700 792.450 487.050 ;
        RECT 793.950 485.850 796.050 487.950 ;
        RECT 794.100 484.050 795.900 485.850 ;
        RECT 806.400 484.950 807.600 497.400 ;
        RECT 822.300 491.400 824.100 503.250 ;
        RECT 826.500 491.400 828.300 503.250 ;
        RECT 829.800 497.400 831.600 503.250 ;
        RECT 847.650 497.400 849.450 503.250 ;
        RECT 850.650 497.400 852.450 503.250 ;
        RECT 853.650 497.400 855.450 503.250 ;
        RECT 821.100 486.150 822.900 487.950 ;
        RECT 826.950 486.150 828.150 491.400 ;
        RECT 829.950 489.150 831.750 490.950 ;
        RECT 851.250 489.150 852.450 497.400 ;
        RECT 829.950 487.050 832.050 489.150 ;
        RECT 803.100 483.150 804.900 484.950 ;
        RECT 802.950 481.050 805.050 483.150 ;
        RECT 805.950 482.850 808.050 484.950 ;
        RECT 820.950 484.050 823.050 486.150 ;
        RECT 823.950 482.850 826.050 484.950 ;
        RECT 826.950 484.050 829.050 486.150 ;
        RECT 847.950 485.850 850.050 487.950 ;
        RECT 850.950 487.050 853.050 489.150 ;
        RECT 848.100 484.050 849.900 485.850 ;
        RECT 788.850 478.800 792.450 479.700 ;
        RECT 772.650 471.750 774.450 474.600 ;
        RECT 775.650 471.750 777.450 474.600 ;
        RECT 788.850 471.750 790.650 478.800 ;
        RECT 793.350 471.750 795.150 477.600 ;
        RECT 806.400 474.600 807.600 482.850 ;
        RECT 824.100 481.050 825.900 482.850 ;
        RECT 827.850 480.750 829.050 484.050 ;
        RECT 828.000 479.700 831.750 480.750 ;
        RECT 851.250 479.700 852.450 487.050 ;
        RECT 853.950 485.850 856.050 487.950 ;
        RECT 854.100 484.050 855.900 485.850 ;
        RECT 821.550 476.700 829.350 478.050 ;
        RECT 803.550 471.750 805.350 474.600 ;
        RECT 806.550 471.750 808.350 474.600 ;
        RECT 821.550 471.750 823.350 476.700 ;
        RECT 824.550 471.750 826.350 475.800 ;
        RECT 827.550 471.750 829.350 476.700 ;
        RECT 830.550 477.600 831.750 479.700 ;
        RECT 848.850 478.800 852.450 479.700 ;
        RECT 830.550 471.750 832.350 477.600 ;
        RECT 848.850 471.750 850.650 478.800 ;
        RECT 853.350 471.750 855.150 477.600 ;
        RECT 15.150 462.900 16.950 467.250 ;
        RECT 13.650 461.400 16.950 462.900 ;
        RECT 18.150 461.400 19.950 467.250 ;
        RECT 13.650 454.950 14.850 461.400 ;
        RECT 16.950 459.900 18.750 460.500 ;
        RECT 22.650 459.900 24.450 467.250 ;
        RECT 16.950 458.700 24.450 459.900 ;
        RECT 13.650 452.850 16.050 454.950 ;
        RECT 17.100 453.150 18.900 454.950 ;
        RECT 13.650 447.600 14.850 452.850 ;
        RECT 16.950 451.050 19.050 453.150 ;
        RECT 13.050 435.750 14.850 447.600 ;
        RECT 16.050 435.750 17.850 447.600 ;
        RECT 20.100 441.600 21.300 458.700 ;
        RECT 35.700 458.400 37.500 467.250 ;
        RECT 41.100 459.000 42.900 467.250 ;
        RECT 56.850 461.400 58.650 467.250 ;
        RECT 61.350 460.200 63.150 467.250 ;
        RECT 76.650 461.400 78.450 467.250 ;
        RECT 59.550 459.300 63.150 460.200 ;
        RECT 77.250 459.300 78.450 461.400 ;
        RECT 79.650 462.300 81.450 467.250 ;
        RECT 82.650 463.200 84.450 467.250 ;
        RECT 85.650 462.300 87.450 467.250 ;
        RECT 79.650 460.950 87.450 462.300 ;
        RECT 95.550 462.300 97.350 467.250 ;
        RECT 98.550 463.200 100.350 467.250 ;
        RECT 101.550 462.300 103.350 467.250 ;
        RECT 95.550 460.950 103.350 462.300 ;
        RECT 104.550 461.400 106.350 467.250 ;
        RECT 116.550 462.300 118.350 467.250 ;
        RECT 119.550 463.200 121.350 467.250 ;
        RECT 122.550 462.300 124.350 467.250 ;
        RECT 104.550 459.300 105.750 461.400 ;
        RECT 116.550 460.950 124.350 462.300 ;
        RECT 125.550 461.400 127.350 467.250 ;
        RECT 137.550 462.300 139.350 467.250 ;
        RECT 140.550 463.200 142.350 467.250 ;
        RECT 143.550 462.300 145.350 467.250 ;
        RECT 125.550 459.300 126.750 461.400 ;
        RECT 137.550 460.950 145.350 462.300 ;
        RECT 146.550 461.400 148.350 467.250 ;
        RECT 146.550 459.300 147.750 461.400 ;
        RECT 161.850 460.200 163.650 467.250 ;
        RECT 166.350 461.400 168.150 467.250 ;
        RECT 181.650 464.400 183.450 467.250 ;
        RECT 184.650 464.400 186.450 467.250 ;
        RECT 187.650 464.400 189.450 467.250 ;
        RECT 161.850 459.300 165.450 460.200 ;
        RECT 41.100 457.350 45.600 459.000 ;
        RECT 22.950 452.850 25.050 454.950 ;
        RECT 44.400 453.150 45.600 457.350 ;
        RECT 56.100 453.150 57.900 454.950 ;
        RECT 23.100 451.050 24.900 452.850 ;
        RECT 34.950 449.850 37.050 451.950 ;
        RECT 40.950 449.850 43.050 451.950 ;
        RECT 43.950 451.050 46.050 453.150 ;
        RECT 55.950 451.050 58.050 453.150 ;
        RECT 59.550 451.950 60.750 459.300 ;
        RECT 77.250 458.250 81.000 459.300 ;
        RECT 102.000 458.250 105.750 459.300 ;
        RECT 123.000 458.250 126.750 459.300 ;
        RECT 144.000 458.250 147.750 459.300 ;
        RECT 79.950 454.950 81.150 458.250 ;
        RECT 83.100 456.150 84.900 457.950 ;
        RECT 98.100 456.150 99.900 457.950 ;
        RECT 62.100 453.150 63.900 454.950 ;
        RECT 35.100 448.050 36.900 449.850 ;
        RECT 37.950 446.850 40.050 448.950 ;
        RECT 41.250 448.050 43.050 449.850 ;
        RECT 38.100 445.050 39.900 446.850 ;
        RECT 44.700 442.800 45.750 451.050 ;
        RECT 58.950 449.850 61.050 451.950 ;
        RECT 61.950 451.050 64.050 453.150 ;
        RECT 79.950 452.850 82.050 454.950 ;
        RECT 82.950 454.050 85.050 456.150 ;
        RECT 85.950 452.850 88.050 454.950 ;
        RECT 94.950 452.850 97.050 454.950 ;
        RECT 97.950 454.050 100.050 456.150 ;
        RECT 101.850 454.950 103.050 458.250 ;
        RECT 119.100 456.150 120.900 457.950 ;
        RECT 100.950 452.850 103.050 454.950 ;
        RECT 115.950 452.850 118.050 454.950 ;
        RECT 118.950 454.050 121.050 456.150 ;
        RECT 122.850 454.950 124.050 458.250 ;
        RECT 140.100 456.150 141.900 457.950 ;
        RECT 121.950 452.850 124.050 454.950 ;
        RECT 136.950 452.850 139.050 454.950 ;
        RECT 139.950 454.050 142.050 456.150 ;
        RECT 143.850 454.950 145.050 458.250 ;
        RECT 145.950 456.450 148.050 457.050 ;
        RECT 151.950 456.450 154.050 457.050 ;
        RECT 145.950 455.550 154.050 456.450 ;
        RECT 145.950 454.950 148.050 455.550 ;
        RECT 151.950 454.950 154.050 455.550 ;
        RECT 142.950 452.850 145.050 454.950 ;
        RECT 161.100 453.150 162.900 454.950 ;
        RECT 76.950 449.850 79.050 451.950 ;
        RECT 38.700 441.900 45.750 442.800 ;
        RECT 38.700 441.600 40.350 441.900 ;
        RECT 19.650 435.750 21.450 441.600 ;
        RECT 22.650 435.750 24.450 441.600 ;
        RECT 35.550 435.750 37.350 441.600 ;
        RECT 38.550 435.750 40.350 441.600 ;
        RECT 44.550 441.600 45.750 441.900 ;
        RECT 59.550 441.600 60.750 449.850 ;
        RECT 77.250 448.050 79.050 449.850 ;
        RECT 80.850 447.600 82.050 452.850 ;
        RECT 86.100 451.050 87.900 452.850 ;
        RECT 95.100 451.050 96.900 452.850 ;
        RECT 100.950 447.600 102.150 452.850 ;
        RECT 103.950 449.850 106.050 451.950 ;
        RECT 116.100 451.050 117.900 452.850 ;
        RECT 103.950 448.050 105.750 449.850 ;
        RECT 121.950 447.600 123.150 452.850 ;
        RECT 124.950 449.850 127.050 451.950 ;
        RECT 137.100 451.050 138.900 452.850 ;
        RECT 124.950 448.050 126.750 449.850 ;
        RECT 142.950 447.600 144.150 452.850 ;
        RECT 145.950 449.850 148.050 451.950 ;
        RECT 160.950 451.050 163.050 453.150 ;
        RECT 164.250 451.950 165.450 459.300 ;
        RECT 184.950 457.950 186.000 464.400 ;
        RECT 197.550 462.300 199.350 467.250 ;
        RECT 200.550 463.200 202.350 467.250 ;
        RECT 203.550 462.300 205.350 467.250 ;
        RECT 197.550 460.950 205.350 462.300 ;
        RECT 206.550 461.400 208.350 467.250 ;
        RECT 206.550 459.300 207.750 461.400 ;
        RECT 204.000 458.250 207.750 459.300 ;
        RECT 224.100 459.000 225.900 467.250 ;
        RECT 184.950 455.850 187.050 457.950 ;
        RECT 200.100 456.150 201.900 457.950 ;
        RECT 167.100 453.150 168.900 454.950 ;
        RECT 163.950 449.850 166.050 451.950 ;
        RECT 166.950 451.050 169.050 453.150 ;
        RECT 181.950 452.850 184.050 454.950 ;
        RECT 182.100 451.050 183.900 452.850 ;
        RECT 145.950 448.050 147.750 449.850 ;
        RECT 41.550 435.750 43.350 441.000 ;
        RECT 44.550 435.750 46.350 441.600 ;
        RECT 56.550 435.750 58.350 441.600 ;
        RECT 59.550 435.750 61.350 441.600 ;
        RECT 62.550 435.750 64.350 441.600 ;
        RECT 77.400 435.750 79.200 441.600 ;
        RECT 80.700 435.750 82.500 447.600 ;
        RECT 84.900 435.750 86.700 447.600 ;
        RECT 96.300 435.750 98.100 447.600 ;
        RECT 100.500 435.750 102.300 447.600 ;
        RECT 103.800 435.750 105.600 441.600 ;
        RECT 117.300 435.750 119.100 447.600 ;
        RECT 121.500 435.750 123.300 447.600 ;
        RECT 124.800 435.750 126.600 441.600 ;
        RECT 138.300 435.750 140.100 447.600 ;
        RECT 142.500 435.750 144.300 447.600 ;
        RECT 164.250 441.600 165.450 449.850 ;
        RECT 184.950 448.650 186.000 455.850 ;
        RECT 187.950 452.850 190.050 454.950 ;
        RECT 196.950 452.850 199.050 454.950 ;
        RECT 199.950 454.050 202.050 456.150 ;
        RECT 203.850 454.950 205.050 458.250 ;
        RECT 202.950 452.850 205.050 454.950 ;
        RECT 221.400 457.350 225.900 459.000 ;
        RECT 229.500 458.400 231.300 467.250 ;
        RECT 245.700 464.400 247.500 467.250 ;
        RECT 249.000 463.050 250.800 467.250 ;
        RECT 245.100 461.400 250.800 463.050 ;
        RECT 253.200 461.400 255.000 467.250 ;
        RECT 265.650 461.400 267.450 467.250 ;
        RECT 221.400 453.150 222.600 457.350 ;
        RECT 245.100 454.950 246.300 461.400 ;
        RECT 266.250 459.300 267.450 461.400 ;
        RECT 268.650 462.300 270.450 467.250 ;
        RECT 271.650 463.200 273.450 467.250 ;
        RECT 274.650 462.300 276.450 467.250 ;
        RECT 268.650 460.950 276.450 462.300 ;
        RECT 284.550 462.300 286.350 467.250 ;
        RECT 287.550 463.200 289.350 467.250 ;
        RECT 290.550 462.300 292.350 467.250 ;
        RECT 284.550 460.950 292.350 462.300 ;
        RECT 293.550 461.400 295.350 467.250 ;
        RECT 310.650 461.400 312.450 467.250 ;
        RECT 293.550 459.300 294.750 461.400 ;
        RECT 266.250 458.250 270.000 459.300 ;
        RECT 291.000 458.250 294.750 459.300 ;
        RECT 311.250 459.300 312.450 461.400 ;
        RECT 313.650 462.300 315.450 467.250 ;
        RECT 316.650 463.200 318.450 467.250 ;
        RECT 319.650 462.300 321.450 467.250 ;
        RECT 313.650 460.950 321.450 462.300 ;
        RECT 331.650 461.400 333.450 467.250 ;
        RECT 332.250 459.300 333.450 461.400 ;
        RECT 334.650 462.300 336.450 467.250 ;
        RECT 337.650 463.200 339.450 467.250 ;
        RECT 340.650 462.300 342.450 467.250 ;
        RECT 356.700 464.400 358.500 467.250 ;
        RECT 360.000 463.050 361.800 467.250 ;
        RECT 334.650 460.950 342.450 462.300 ;
        RECT 356.100 461.400 361.800 463.050 ;
        RECT 364.200 461.400 366.000 467.250 ;
        RECT 377.700 464.400 379.500 467.250 ;
        RECT 381.000 463.050 382.800 467.250 ;
        RECT 377.100 461.400 382.800 463.050 ;
        RECT 385.200 461.400 387.000 467.250 ;
        RECT 400.800 461.400 402.600 467.250 ;
        RECT 405.000 461.400 406.800 467.250 ;
        RECT 409.200 461.400 411.000 467.250 ;
        RECT 421.650 461.400 423.450 467.250 ;
        RECT 424.650 464.400 426.450 467.250 ;
        RECT 427.650 464.400 429.450 467.250 ;
        RECT 430.650 464.400 432.450 467.250 ;
        RECT 440.550 464.400 442.350 467.250 ;
        RECT 443.550 464.400 445.350 467.250 ;
        RECT 446.550 464.400 448.350 467.250 ;
        RECT 311.250 458.250 315.000 459.300 ;
        RECT 332.250 458.250 336.000 459.300 ;
        RECT 248.100 456.150 249.900 457.950 ;
        RECT 188.100 451.050 189.900 452.850 ;
        RECT 197.100 451.050 198.900 452.850 ;
        RECT 183.450 447.600 186.000 448.650 ;
        RECT 202.950 447.600 204.150 452.850 ;
        RECT 205.950 449.850 208.050 451.950 ;
        RECT 220.950 451.050 223.050 453.150 ;
        RECT 244.950 452.850 247.050 454.950 ;
        RECT 247.950 454.050 250.050 456.150 ;
        RECT 250.950 455.850 253.050 457.950 ;
        RECT 254.100 456.150 255.900 457.950 ;
        RECT 251.100 454.050 252.900 455.850 ;
        RECT 253.950 454.050 256.050 456.150 ;
        RECT 268.950 454.950 270.150 458.250 ;
        RECT 272.100 456.150 273.900 457.950 ;
        RECT 287.100 456.150 288.900 457.950 ;
        RECT 268.950 452.850 271.050 454.950 ;
        RECT 271.950 454.050 274.050 456.150 ;
        RECT 274.950 452.850 277.050 454.950 ;
        RECT 283.950 452.850 286.050 454.950 ;
        RECT 286.950 454.050 289.050 456.150 ;
        RECT 290.850 454.950 292.050 458.250 ;
        RECT 289.950 452.850 292.050 454.950 ;
        RECT 313.950 454.950 315.150 458.250 ;
        RECT 317.100 456.150 318.900 457.950 ;
        RECT 313.950 452.850 316.050 454.950 ;
        RECT 316.950 454.050 319.050 456.150 ;
        RECT 334.950 454.950 336.150 458.250 ;
        RECT 338.100 456.150 339.900 457.950 ;
        RECT 319.950 452.850 322.050 454.950 ;
        RECT 334.950 452.850 337.050 454.950 ;
        RECT 337.950 454.050 340.050 456.150 ;
        RECT 356.100 454.950 357.300 461.400 ;
        RECT 359.100 456.150 360.900 457.950 ;
        RECT 340.950 452.850 343.050 454.950 ;
        RECT 355.950 452.850 358.050 454.950 ;
        RECT 358.950 454.050 361.050 456.150 ;
        RECT 361.950 455.850 364.050 457.950 ;
        RECT 365.100 456.150 366.900 457.950 ;
        RECT 362.100 454.050 363.900 455.850 ;
        RECT 364.950 454.050 367.050 456.150 ;
        RECT 377.100 454.950 378.300 461.400 ;
        RECT 380.100 456.150 381.900 457.950 ;
        RECT 376.950 452.850 379.050 454.950 ;
        RECT 379.950 454.050 382.050 456.150 ;
        RECT 382.950 455.850 385.050 457.950 ;
        RECT 386.100 456.150 387.900 457.950 ;
        RECT 401.250 456.150 403.050 457.950 ;
        RECT 383.100 454.050 384.900 455.850 ;
        RECT 385.950 454.050 388.050 456.150 ;
        RECT 397.950 452.850 400.050 454.950 ;
        RECT 400.950 454.050 403.050 456.150 ;
        RECT 405.000 454.950 406.050 461.400 ;
        RECT 403.950 452.850 406.050 454.950 ;
        RECT 406.950 456.150 408.750 457.950 ;
        RECT 421.950 456.150 423.000 461.400 ;
        RECT 427.650 460.200 428.550 464.400 ;
        RECT 425.250 459.300 428.550 460.200 ;
        RECT 425.250 458.400 427.050 459.300 ;
        RECT 406.950 454.050 409.050 456.150 ;
        RECT 409.950 452.850 412.050 454.950 ;
        RECT 421.950 454.050 424.050 456.150 ;
        RECT 205.950 448.050 207.750 449.850 ;
        RECT 145.800 435.750 147.600 441.600 ;
        RECT 160.650 435.750 162.450 441.600 ;
        RECT 163.650 435.750 165.450 441.600 ;
        RECT 166.650 435.750 168.450 441.600 ;
        RECT 183.450 435.750 185.250 447.600 ;
        RECT 187.650 435.750 189.450 447.600 ;
        RECT 198.300 435.750 200.100 447.600 ;
        RECT 202.500 435.750 204.300 447.600 ;
        RECT 221.250 442.800 222.300 451.050 ;
        RECT 223.950 449.850 226.050 451.950 ;
        RECT 229.950 449.850 232.050 451.950 ;
        RECT 223.950 448.050 225.750 449.850 ;
        RECT 226.950 446.850 229.050 448.950 ;
        RECT 230.100 448.050 231.900 449.850 ;
        RECT 245.100 447.600 246.300 452.850 ;
        RECT 265.950 449.850 268.050 451.950 ;
        RECT 266.250 448.050 268.050 449.850 ;
        RECT 269.850 447.600 271.050 452.850 ;
        RECT 275.100 451.050 276.900 452.850 ;
        RECT 284.100 451.050 285.900 452.850 ;
        RECT 289.950 447.600 291.150 452.850 ;
        RECT 292.950 449.850 295.050 451.950 ;
        RECT 310.950 449.850 313.050 451.950 ;
        RECT 292.950 448.050 294.750 449.850 ;
        RECT 311.250 448.050 313.050 449.850 ;
        RECT 314.850 447.600 316.050 452.850 ;
        RECT 320.100 451.050 321.900 452.850 ;
        RECT 331.950 449.850 334.050 451.950 ;
        RECT 332.250 448.050 334.050 449.850 ;
        RECT 335.850 447.600 337.050 452.850 ;
        RECT 341.100 451.050 342.900 452.850 ;
        RECT 356.100 447.600 357.300 452.850 ;
        RECT 377.100 447.600 378.300 452.850 ;
        RECT 398.100 451.050 399.900 452.850 ;
        RECT 379.950 450.450 382.050 451.050 ;
        RECT 388.950 450.450 391.050 451.050 ;
        RECT 379.950 449.550 391.050 450.450 ;
        RECT 379.950 448.950 382.050 449.550 ;
        RECT 388.950 448.950 391.050 449.550 ;
        RECT 403.950 449.400 404.850 452.850 ;
        RECT 409.950 451.050 411.750 452.850 ;
        RECT 400.800 448.500 404.850 449.400 ;
        RECT 400.800 447.600 402.600 448.500 ;
        RECT 227.100 445.050 228.900 446.850 ;
        RECT 221.250 441.900 228.300 442.800 ;
        RECT 221.250 441.600 222.450 441.900 ;
        RECT 205.800 435.750 207.600 441.600 ;
        RECT 220.650 435.750 222.450 441.600 ;
        RECT 226.650 441.600 228.300 441.900 ;
        RECT 223.650 435.750 225.450 441.000 ;
        RECT 226.650 435.750 228.450 441.600 ;
        RECT 229.650 435.750 231.450 441.600 ;
        RECT 244.650 435.750 246.450 447.600 ;
        RECT 247.650 446.700 255.450 447.600 ;
        RECT 247.650 435.750 249.450 446.700 ;
        RECT 250.650 435.750 252.450 445.800 ;
        RECT 253.650 435.750 255.450 446.700 ;
        RECT 266.400 435.750 268.200 441.600 ;
        RECT 269.700 435.750 271.500 447.600 ;
        RECT 273.900 435.750 275.700 447.600 ;
        RECT 285.300 435.750 287.100 447.600 ;
        RECT 289.500 435.750 291.300 447.600 ;
        RECT 292.800 435.750 294.600 441.600 ;
        RECT 311.400 435.750 313.200 441.600 ;
        RECT 314.700 435.750 316.500 447.600 ;
        RECT 318.900 435.750 320.700 447.600 ;
        RECT 332.400 435.750 334.200 441.600 ;
        RECT 335.700 435.750 337.500 447.600 ;
        RECT 339.900 435.750 341.700 447.600 ;
        RECT 355.650 435.750 357.450 447.600 ;
        RECT 358.650 446.700 366.450 447.600 ;
        RECT 358.650 435.750 360.450 446.700 ;
        RECT 361.650 435.750 363.450 445.800 ;
        RECT 364.650 435.750 366.450 446.700 ;
        RECT 376.650 435.750 378.450 447.600 ;
        RECT 379.650 446.700 387.450 447.600 ;
        RECT 379.650 435.750 381.450 446.700 ;
        RECT 382.650 435.750 384.450 445.800 ;
        RECT 385.650 435.750 387.450 446.700 ;
        RECT 397.650 436.500 399.450 447.600 ;
        RECT 400.650 437.400 402.450 447.600 ;
        RECT 422.550 447.450 423.900 454.050 ;
        RECT 425.400 450.150 426.300 458.400 ;
        RECT 444.000 457.950 445.050 464.400 ;
        RECT 461.850 461.400 463.650 467.250 ;
        RECT 466.350 460.200 468.150 467.250 ;
        RECT 483.150 462.900 484.950 467.250 ;
        RECT 430.950 455.850 433.050 457.950 ;
        RECT 442.950 455.850 445.050 457.950 ;
        RECT 427.950 452.850 430.050 454.950 ;
        RECT 431.100 454.050 432.900 455.850 ;
        RECT 439.950 452.850 442.050 454.950 ;
        RECT 428.100 451.050 429.900 452.850 ;
        RECT 440.100 451.050 441.900 452.850 ;
        RECT 425.250 450.000 427.050 450.150 ;
        RECT 425.250 448.800 432.450 450.000 ;
        RECT 425.250 448.350 427.050 448.800 ;
        RECT 431.250 447.600 432.450 448.800 ;
        RECT 444.000 448.650 445.050 455.850 ;
        RECT 464.550 459.300 468.150 460.200 ;
        RECT 481.650 461.400 484.950 462.900 ;
        RECT 486.150 461.400 487.950 467.250 ;
        RECT 445.950 452.850 448.050 454.950 ;
        RECT 461.100 453.150 462.900 454.950 ;
        RECT 446.100 451.050 447.900 452.850 ;
        RECT 460.950 451.050 463.050 453.150 ;
        RECT 464.550 451.950 465.750 459.300 ;
        RECT 481.650 454.950 482.850 461.400 ;
        RECT 484.950 459.900 486.750 460.500 ;
        RECT 490.650 459.900 492.450 467.250 ;
        RECT 500.550 464.400 502.350 467.250 ;
        RECT 503.550 464.400 505.350 467.250 ;
        RECT 506.550 464.400 508.350 467.250 ;
        RECT 484.950 458.700 492.450 459.900 ;
        RECT 504.450 460.200 505.350 464.400 ;
        RECT 509.550 461.400 511.350 467.250 ;
        RECT 523.650 461.400 525.450 467.250 ;
        RECT 504.450 459.300 507.750 460.200 ;
        RECT 467.100 453.150 468.900 454.950 ;
        RECT 463.950 449.850 466.050 451.950 ;
        RECT 466.950 451.050 469.050 453.150 ;
        RECT 481.650 452.850 484.050 454.950 ;
        RECT 485.100 453.150 486.900 454.950 ;
        RECT 444.000 447.600 446.550 448.650 ;
        RECT 403.650 446.400 411.450 447.300 ;
        RECT 403.650 436.500 405.450 446.400 ;
        RECT 397.650 435.750 405.450 436.500 ;
        RECT 406.650 435.750 408.450 445.500 ;
        RECT 409.650 435.750 411.450 446.400 ;
        RECT 422.550 446.100 424.950 447.450 ;
        RECT 423.150 435.750 424.950 446.100 ;
        RECT 426.150 435.750 427.950 447.450 ;
        RECT 430.650 435.750 432.450 447.600 ;
        RECT 440.550 435.750 442.350 447.600 ;
        RECT 444.750 435.750 446.550 447.600 ;
        RECT 464.550 441.600 465.750 449.850 ;
        RECT 466.950 447.450 469.050 448.050 ;
        RECT 472.950 447.450 475.050 448.050 ;
        RECT 481.650 447.600 482.850 452.850 ;
        RECT 484.950 451.050 487.050 453.150 ;
        RECT 466.950 446.550 475.050 447.450 ;
        RECT 466.950 445.950 469.050 446.550 ;
        RECT 472.950 445.950 475.050 446.550 ;
        RECT 461.550 435.750 463.350 441.600 ;
        RECT 464.550 435.750 466.350 441.600 ;
        RECT 467.550 435.750 469.350 441.600 ;
        RECT 481.050 435.750 482.850 447.600 ;
        RECT 484.050 435.750 485.850 447.600 ;
        RECT 488.100 441.600 489.300 458.700 ;
        RECT 505.950 458.400 507.750 459.300 ;
        RECT 499.950 455.850 502.050 457.950 ;
        RECT 490.950 452.850 493.050 454.950 ;
        RECT 500.100 454.050 501.900 455.850 ;
        RECT 502.950 452.850 505.050 454.950 ;
        RECT 491.100 451.050 492.900 452.850 ;
        RECT 503.100 451.050 504.900 452.850 ;
        RECT 506.700 450.150 507.600 458.400 ;
        RECT 510.000 456.150 511.050 461.400 ;
        RECT 524.250 459.300 525.450 461.400 ;
        RECT 526.650 462.300 528.450 467.250 ;
        RECT 529.650 463.200 531.450 467.250 ;
        RECT 532.650 462.300 534.450 467.250 ;
        RECT 526.650 460.950 534.450 462.300 ;
        RECT 544.650 461.400 546.450 467.250 ;
        RECT 545.250 459.300 546.450 461.400 ;
        RECT 547.650 462.300 549.450 467.250 ;
        RECT 550.650 463.200 552.450 467.250 ;
        RECT 553.650 462.300 555.450 467.250 ;
        RECT 547.650 460.950 555.450 462.300 ;
        RECT 565.650 461.400 567.450 467.250 ;
        RECT 568.650 464.400 570.450 467.250 ;
        RECT 571.650 464.400 573.450 467.250 ;
        RECT 574.650 464.400 576.450 467.250 ;
        RECT 524.250 458.250 528.000 459.300 ;
        RECT 545.250 458.250 549.000 459.300 ;
        RECT 508.950 454.050 511.050 456.150 ;
        RECT 526.950 454.950 528.150 458.250 ;
        RECT 530.100 456.150 531.900 457.950 ;
        RECT 505.950 450.000 507.750 450.150 ;
        RECT 500.550 448.800 507.750 450.000 ;
        RECT 500.550 447.600 501.750 448.800 ;
        RECT 505.950 448.350 507.750 448.800 ;
        RECT 487.650 435.750 489.450 441.600 ;
        RECT 490.650 435.750 492.450 441.600 ;
        RECT 500.550 435.750 502.350 447.600 ;
        RECT 509.100 447.450 510.450 454.050 ;
        RECT 526.950 452.850 529.050 454.950 ;
        RECT 529.950 454.050 532.050 456.150 ;
        RECT 547.950 454.950 549.150 458.250 ;
        RECT 551.100 456.150 552.900 457.950 ;
        RECT 565.950 456.150 567.000 461.400 ;
        RECT 571.650 460.200 572.550 464.400 ;
        RECT 591.150 462.900 592.950 467.250 ;
        RECT 569.250 459.300 572.550 460.200 ;
        RECT 589.650 461.400 592.950 462.900 ;
        RECT 594.150 461.400 595.950 467.250 ;
        RECT 569.250 458.400 571.050 459.300 ;
        RECT 532.950 452.850 535.050 454.950 ;
        RECT 547.950 452.850 550.050 454.950 ;
        RECT 550.950 454.050 553.050 456.150 ;
        RECT 553.950 452.850 556.050 454.950 ;
        RECT 565.950 454.050 568.050 456.150 ;
        RECT 523.950 449.850 526.050 451.950 ;
        RECT 524.250 448.050 526.050 449.850 ;
        RECT 527.850 447.600 529.050 452.850 ;
        RECT 533.100 451.050 534.900 452.850 ;
        RECT 544.950 449.850 547.050 451.950 ;
        RECT 545.250 448.050 547.050 449.850 ;
        RECT 548.850 447.600 550.050 452.850 ;
        RECT 554.100 451.050 555.900 452.850 ;
        RECT 505.050 435.750 506.850 447.450 ;
        RECT 508.050 446.100 510.450 447.450 ;
        RECT 508.050 435.750 509.850 446.100 ;
        RECT 524.400 435.750 526.200 441.600 ;
        RECT 527.700 435.750 529.500 447.600 ;
        RECT 531.900 435.750 533.700 447.600 ;
        RECT 545.400 435.750 547.200 441.600 ;
        RECT 548.700 435.750 550.500 447.600 ;
        RECT 552.900 435.750 554.700 447.600 ;
        RECT 566.550 447.450 567.900 454.050 ;
        RECT 569.400 450.150 570.300 458.400 ;
        RECT 574.950 455.850 577.050 457.950 ;
        RECT 571.950 452.850 574.050 454.950 ;
        RECT 575.100 454.050 576.900 455.850 ;
        RECT 589.650 454.950 590.850 461.400 ;
        RECT 592.950 459.900 594.750 460.500 ;
        RECT 598.650 459.900 600.450 467.250 ;
        RECT 608.550 464.400 610.350 467.250 ;
        RECT 611.550 464.400 613.350 467.250 ;
        RECT 614.550 464.400 616.350 467.250 ;
        RECT 592.950 458.700 600.450 459.900 ;
        RECT 589.650 452.850 592.050 454.950 ;
        RECT 593.100 453.150 594.900 454.950 ;
        RECT 572.100 451.050 573.900 452.850 ;
        RECT 569.250 450.000 571.050 450.150 ;
        RECT 569.250 448.800 576.450 450.000 ;
        RECT 569.250 448.350 571.050 448.800 ;
        RECT 575.250 447.600 576.450 448.800 ;
        RECT 589.650 447.600 590.850 452.850 ;
        RECT 592.950 451.050 595.050 453.150 ;
        RECT 566.550 446.100 568.950 447.450 ;
        RECT 567.150 435.750 568.950 446.100 ;
        RECT 570.150 435.750 571.950 447.450 ;
        RECT 574.650 435.750 576.450 447.600 ;
        RECT 589.050 435.750 590.850 447.600 ;
        RECT 592.050 435.750 593.850 447.600 ;
        RECT 596.100 441.600 597.300 458.700 ;
        RECT 612.000 457.950 613.050 464.400 ;
        RECT 626.700 458.400 628.500 467.250 ;
        RECT 632.100 459.000 633.900 467.250 ;
        RECT 642.150 461.400 643.950 467.250 ;
        RECT 645.150 464.400 646.950 467.250 ;
        RECT 649.950 465.300 651.750 467.250 ;
        RECT 648.000 464.400 651.750 465.300 ;
        RECT 654.450 464.400 656.250 467.250 ;
        RECT 657.750 464.400 659.550 467.250 ;
        RECT 661.650 464.400 663.450 467.250 ;
        RECT 665.850 464.400 667.650 467.250 ;
        RECT 670.350 464.400 672.150 467.250 ;
        RECT 648.000 463.500 649.050 464.400 ;
        RECT 646.950 461.400 649.050 463.500 ;
        RECT 657.750 462.600 658.800 464.400 ;
        RECT 610.950 455.850 613.050 457.950 ;
        RECT 632.100 457.350 636.600 459.000 ;
        RECT 598.950 452.850 601.050 454.950 ;
        RECT 607.950 452.850 610.050 454.950 ;
        RECT 599.100 451.050 600.900 452.850 ;
        RECT 608.100 451.050 609.900 452.850 ;
        RECT 612.000 448.650 613.050 455.850 ;
        RECT 613.950 452.850 616.050 454.950 ;
        RECT 635.400 453.150 636.600 457.350 ;
        RECT 614.100 451.050 615.900 452.850 ;
        RECT 625.950 449.850 628.050 451.950 ;
        RECT 631.950 449.850 634.050 451.950 ;
        RECT 634.950 451.050 637.050 453.150 ;
        RECT 612.000 447.600 614.550 448.650 ;
        RECT 626.100 448.050 627.900 449.850 ;
        RECT 595.650 435.750 597.450 441.600 ;
        RECT 598.650 435.750 600.450 441.600 ;
        RECT 608.550 435.750 610.350 447.600 ;
        RECT 612.750 435.750 614.550 447.600 ;
        RECT 628.950 446.850 631.050 448.950 ;
        RECT 632.250 448.050 634.050 449.850 ;
        RECT 629.100 445.050 630.900 446.850 ;
        RECT 635.700 442.800 636.750 451.050 ;
        RECT 629.700 441.900 636.750 442.800 ;
        RECT 629.700 441.600 631.350 441.900 ;
        RECT 626.550 435.750 628.350 441.600 ;
        RECT 629.550 435.750 631.350 441.600 ;
        RECT 635.550 441.600 636.750 441.900 ;
        RECT 642.150 448.800 643.050 461.400 ;
        RECT 650.550 460.800 652.350 462.600 ;
        RECT 653.850 461.550 658.800 462.600 ;
        RECT 666.300 463.500 667.350 464.400 ;
        RECT 666.300 462.300 670.050 463.500 ;
        RECT 653.850 460.800 655.650 461.550 ;
        RECT 650.850 459.900 651.900 460.800 ;
        RECT 661.050 460.200 662.850 462.000 ;
        RECT 667.950 461.400 670.050 462.300 ;
        RECT 673.650 461.400 675.450 467.250 ;
        RECT 661.050 459.900 661.950 460.200 ;
        RECT 650.850 459.000 661.950 459.900 ;
        RECT 674.250 459.150 675.450 461.400 ;
        RECT 686.550 462.300 688.350 467.250 ;
        RECT 689.550 463.200 691.350 467.250 ;
        RECT 692.550 462.300 694.350 467.250 ;
        RECT 686.550 460.950 694.350 462.300 ;
        RECT 695.550 461.400 697.350 467.250 ;
        RECT 707.550 462.300 709.350 467.250 ;
        RECT 710.550 463.200 712.350 467.250 ;
        RECT 713.550 462.300 715.350 467.250 ;
        RECT 695.550 459.300 696.750 461.400 ;
        RECT 707.550 460.950 715.350 462.300 ;
        RECT 716.550 461.400 718.350 467.250 ;
        RECT 716.550 459.300 717.750 461.400 ;
        RECT 731.850 460.200 733.650 467.250 ;
        RECT 736.350 461.400 738.150 467.250 ;
        RECT 746.850 461.400 748.650 467.250 ;
        RECT 751.350 460.200 753.150 467.250 ;
        RECT 731.850 459.300 735.450 460.200 ;
        RECT 650.850 457.800 651.900 459.000 ;
        RECT 645.000 456.600 651.900 457.800 ;
        RECT 645.000 455.850 645.900 456.600 ;
        RECT 650.100 456.000 651.900 456.600 ;
        RECT 644.100 454.050 645.900 455.850 ;
        RECT 647.100 454.950 648.900 455.700 ;
        RECT 661.050 454.950 661.950 459.000 ;
        RECT 670.950 457.050 675.450 459.150 ;
        RECT 693.000 458.250 696.750 459.300 ;
        RECT 714.000 458.250 717.750 459.300 ;
        RECT 669.150 455.250 673.050 457.050 ;
        RECT 670.950 454.950 673.050 455.250 ;
        RECT 647.100 453.900 655.050 454.950 ;
        RECT 652.950 452.850 655.050 453.900 ;
        RECT 658.950 452.850 661.950 454.950 ;
        RECT 651.450 449.100 653.250 449.400 ;
        RECT 651.450 448.800 659.850 449.100 ;
        RECT 642.150 448.200 659.850 448.800 ;
        RECT 642.150 447.600 653.250 448.200 ;
        RECT 632.550 435.750 634.350 441.000 ;
        RECT 635.550 435.750 637.350 441.600 ;
        RECT 642.150 435.750 643.950 447.600 ;
        RECT 656.250 446.700 658.050 447.300 ;
        RECT 650.550 445.500 658.050 446.700 ;
        RECT 658.950 446.100 659.850 448.200 ;
        RECT 661.050 448.200 661.950 452.850 ;
        RECT 671.250 449.400 673.050 451.200 ;
        RECT 667.950 448.200 672.150 449.400 ;
        RECT 661.050 447.300 667.050 448.200 ;
        RECT 667.950 447.300 670.050 448.200 ;
        RECT 674.250 447.600 675.450 457.050 ;
        RECT 689.100 456.150 690.900 457.950 ;
        RECT 685.950 452.850 688.050 454.950 ;
        RECT 688.950 454.050 691.050 456.150 ;
        RECT 692.850 454.950 694.050 458.250 ;
        RECT 710.100 456.150 711.900 457.950 ;
        RECT 691.950 452.850 694.050 454.950 ;
        RECT 706.950 452.850 709.050 454.950 ;
        RECT 709.950 454.050 712.050 456.150 ;
        RECT 713.850 454.950 715.050 458.250 ;
        RECT 712.950 452.850 715.050 454.950 ;
        RECT 731.100 453.150 732.900 454.950 ;
        RECT 686.100 451.050 687.900 452.850 ;
        RECT 691.950 447.600 693.150 452.850 ;
        RECT 694.950 449.850 697.050 451.950 ;
        RECT 707.100 451.050 708.900 452.850 ;
        RECT 694.950 448.050 696.750 449.850 ;
        RECT 712.950 447.600 714.150 452.850 ;
        RECT 715.950 449.850 718.050 451.950 ;
        RECT 730.950 451.050 733.050 453.150 ;
        RECT 734.250 451.950 735.450 459.300 ;
        RECT 749.550 459.300 753.150 460.200 ;
        RECT 759.150 461.400 760.950 467.250 ;
        RECT 762.150 464.400 763.950 467.250 ;
        RECT 766.950 465.300 768.750 467.250 ;
        RECT 765.000 464.400 768.750 465.300 ;
        RECT 771.450 464.400 773.250 467.250 ;
        RECT 774.750 464.400 776.550 467.250 ;
        RECT 778.650 464.400 780.450 467.250 ;
        RECT 782.850 464.400 784.650 467.250 ;
        RECT 787.350 464.400 789.150 467.250 ;
        RECT 765.000 463.500 766.050 464.400 ;
        RECT 763.950 461.400 766.050 463.500 ;
        RECT 774.750 462.600 775.800 464.400 ;
        RECT 737.100 453.150 738.900 454.950 ;
        RECT 746.100 453.150 747.900 454.950 ;
        RECT 733.950 449.850 736.050 451.950 ;
        RECT 736.950 451.050 739.050 453.150 ;
        RECT 745.950 451.050 748.050 453.150 ;
        RECT 749.550 451.950 750.750 459.300 ;
        RECT 752.100 453.150 753.900 454.950 ;
        RECT 748.950 449.850 751.050 451.950 ;
        RECT 751.950 451.050 754.050 453.150 ;
        RECT 715.950 448.050 717.750 449.850 ;
        RECT 666.150 446.400 667.050 447.300 ;
        RECT 663.450 446.100 665.250 446.400 ;
        RECT 650.550 444.600 651.750 445.500 ;
        RECT 658.950 445.200 665.250 446.100 ;
        RECT 663.450 444.600 665.250 445.200 ;
        RECT 666.150 444.600 668.850 446.400 ;
        RECT 646.950 442.500 651.750 444.600 ;
        RECT 654.150 442.500 661.050 444.300 ;
        RECT 650.550 441.600 651.750 442.500 ;
        RECT 645.150 435.750 646.950 441.600 ;
        RECT 650.250 435.750 652.050 441.600 ;
        RECT 655.050 435.750 656.850 441.600 ;
        RECT 658.050 435.750 659.850 442.500 ;
        RECT 666.150 441.600 670.050 443.700 ;
        RECT 661.950 435.750 663.750 441.600 ;
        RECT 666.150 435.750 667.950 441.600 ;
        RECT 670.650 435.750 672.450 438.600 ;
        RECT 673.650 435.750 675.450 447.600 ;
        RECT 687.300 435.750 689.100 447.600 ;
        RECT 691.500 435.750 693.300 447.600 ;
        RECT 694.800 435.750 696.600 441.600 ;
        RECT 708.300 435.750 710.100 447.600 ;
        RECT 712.500 435.750 714.300 447.600 ;
        RECT 734.250 441.600 735.450 449.850 ;
        RECT 749.550 441.600 750.750 449.850 ;
        RECT 759.150 448.800 760.050 461.400 ;
        RECT 767.550 460.800 769.350 462.600 ;
        RECT 770.850 461.550 775.800 462.600 ;
        RECT 783.300 463.500 784.350 464.400 ;
        RECT 783.300 462.300 787.050 463.500 ;
        RECT 770.850 460.800 772.650 461.550 ;
        RECT 767.850 459.900 768.900 460.800 ;
        RECT 778.050 460.200 779.850 462.000 ;
        RECT 784.950 461.400 787.050 462.300 ;
        RECT 790.650 461.400 792.450 467.250 ;
        RECT 802.650 461.400 804.450 467.250 ;
        RECT 805.650 461.400 807.450 467.250 ;
        RECT 808.650 461.400 810.450 467.250 ;
        RECT 811.650 461.400 813.450 467.250 ;
        RECT 814.650 461.400 816.450 467.250 ;
        RECT 778.050 459.900 778.950 460.200 ;
        RECT 767.850 459.000 778.950 459.900 ;
        RECT 791.250 459.150 792.450 461.400 ;
        RECT 805.800 460.500 807.600 461.400 ;
        RECT 811.800 460.500 813.600 461.400 ;
        RECT 817.650 460.500 819.450 467.250 ;
        RECT 820.650 461.400 822.450 467.250 ;
        RECT 823.650 461.400 825.450 467.250 ;
        RECT 826.650 461.400 828.450 467.250 ;
        RECT 830.550 461.400 832.350 467.250 ;
        RECT 833.850 464.400 835.650 467.250 ;
        RECT 838.350 464.400 840.150 467.250 ;
        RECT 842.550 464.400 844.350 467.250 ;
        RECT 846.450 464.400 848.250 467.250 ;
        RECT 849.750 464.400 851.550 467.250 ;
        RECT 854.250 465.300 856.050 467.250 ;
        RECT 854.250 464.400 858.000 465.300 ;
        RECT 859.050 464.400 860.850 467.250 ;
        RECT 838.650 463.500 839.700 464.400 ;
        RECT 835.950 462.300 839.700 463.500 ;
        RECT 847.200 462.600 848.250 464.400 ;
        RECT 856.950 463.500 858.000 464.400 ;
        RECT 835.950 461.400 838.050 462.300 ;
        RECT 823.800 460.500 825.600 461.400 ;
        RECT 804.900 460.350 807.600 460.500 ;
        RECT 767.850 457.800 768.900 459.000 ;
        RECT 762.000 456.600 768.900 457.800 ;
        RECT 762.000 455.850 762.900 456.600 ;
        RECT 767.100 456.000 768.900 456.600 ;
        RECT 761.100 454.050 762.900 455.850 ;
        RECT 764.100 454.950 765.900 455.700 ;
        RECT 778.050 454.950 778.950 459.000 ;
        RECT 787.950 457.050 792.450 459.150 ;
        RECT 786.150 455.250 790.050 457.050 ;
        RECT 787.950 454.950 790.050 455.250 ;
        RECT 764.100 453.900 772.050 454.950 ;
        RECT 769.950 452.850 772.050 453.900 ;
        RECT 775.950 452.850 778.950 454.950 ;
        RECT 768.450 449.100 770.250 449.400 ;
        RECT 768.450 448.800 776.850 449.100 ;
        RECT 759.150 448.200 776.850 448.800 ;
        RECT 759.150 447.600 770.250 448.200 ;
        RECT 715.800 435.750 717.600 441.600 ;
        RECT 730.650 435.750 732.450 441.600 ;
        RECT 733.650 435.750 735.450 441.600 ;
        RECT 736.650 435.750 738.450 441.600 ;
        RECT 746.550 435.750 748.350 441.600 ;
        RECT 749.550 435.750 751.350 441.600 ;
        RECT 752.550 435.750 754.350 441.600 ;
        RECT 759.150 435.750 760.950 447.600 ;
        RECT 773.250 446.700 775.050 447.300 ;
        RECT 767.550 445.500 775.050 446.700 ;
        RECT 775.950 446.100 776.850 448.200 ;
        RECT 778.050 448.200 778.950 452.850 ;
        RECT 788.250 449.400 790.050 451.200 ;
        RECT 784.950 448.200 789.150 449.400 ;
        RECT 778.050 447.300 784.050 448.200 ;
        RECT 784.950 447.300 787.050 448.200 ;
        RECT 791.250 447.600 792.450 457.050 ;
        RECT 804.750 459.300 807.600 460.350 ;
        RECT 809.700 459.300 813.600 460.500 ;
        RECT 815.700 459.300 819.450 460.500 ;
        RECT 821.550 459.300 825.600 460.500 ;
        RECT 804.750 456.150 805.800 459.300 ;
        RECT 809.700 458.400 810.900 459.300 ;
        RECT 815.700 458.400 816.900 459.300 ;
        RECT 821.550 458.400 822.750 459.300 ;
        RECT 806.700 456.600 810.900 458.400 ;
        RECT 812.700 456.600 816.900 458.400 ;
        RECT 818.700 456.600 822.750 458.400 ;
        RECT 830.550 459.150 831.750 461.400 ;
        RECT 843.150 460.200 844.950 462.000 ;
        RECT 847.200 461.550 852.150 462.600 ;
        RECT 850.350 460.800 852.150 461.550 ;
        RECT 853.650 460.800 855.450 462.600 ;
        RECT 856.950 461.400 859.050 463.500 ;
        RECT 862.050 461.400 863.850 467.250 ;
        RECT 844.050 459.900 844.950 460.200 ;
        RECT 854.100 459.900 855.150 460.800 ;
        RECT 802.950 454.050 805.800 456.150 ;
        RECT 804.750 449.700 805.800 454.050 ;
        RECT 809.700 449.700 810.900 456.600 ;
        RECT 815.700 449.700 816.900 456.600 ;
        RECT 821.550 449.700 822.750 456.600 ;
        RECT 824.100 456.150 825.900 457.950 ;
        RECT 830.550 457.050 835.050 459.150 ;
        RECT 844.050 459.000 855.150 459.900 ;
        RECT 823.950 454.050 826.050 456.150 ;
        RECT 804.750 448.500 807.450 449.700 ;
        RECT 809.700 448.500 813.450 449.700 ;
        RECT 815.700 448.500 819.450 449.700 ;
        RECT 821.550 448.500 825.450 449.700 ;
        RECT 783.150 446.400 784.050 447.300 ;
        RECT 780.450 446.100 782.250 446.400 ;
        RECT 767.550 444.600 768.750 445.500 ;
        RECT 775.950 445.200 782.250 446.100 ;
        RECT 780.450 444.600 782.250 445.200 ;
        RECT 783.150 444.600 785.850 446.400 ;
        RECT 763.950 442.500 768.750 444.600 ;
        RECT 771.150 442.500 778.050 444.300 ;
        RECT 767.550 441.600 768.750 442.500 ;
        RECT 762.150 435.750 763.950 441.600 ;
        RECT 767.250 435.750 769.050 441.600 ;
        RECT 772.050 435.750 773.850 441.600 ;
        RECT 775.050 435.750 776.850 442.500 ;
        RECT 783.150 441.600 787.050 443.700 ;
        RECT 778.950 435.750 780.750 441.600 ;
        RECT 783.150 435.750 784.950 441.600 ;
        RECT 787.650 435.750 789.450 438.600 ;
        RECT 790.650 435.750 792.450 447.600 ;
        RECT 802.650 435.750 804.450 447.600 ;
        RECT 805.650 435.750 807.450 448.500 ;
        RECT 808.650 435.750 810.450 447.600 ;
        RECT 811.650 435.750 813.450 448.500 ;
        RECT 814.650 435.750 816.450 447.600 ;
        RECT 817.650 435.750 819.450 448.500 ;
        RECT 820.650 435.750 822.450 447.600 ;
        RECT 823.650 435.750 825.450 448.500 ;
        RECT 830.550 447.600 831.750 457.050 ;
        RECT 832.950 455.250 836.850 457.050 ;
        RECT 832.950 454.950 835.050 455.250 ;
        RECT 844.050 454.950 844.950 459.000 ;
        RECT 854.100 457.800 855.150 459.000 ;
        RECT 854.100 456.600 861.000 457.800 ;
        RECT 854.100 456.000 855.900 456.600 ;
        RECT 860.100 455.850 861.000 456.600 ;
        RECT 857.100 454.950 858.900 455.700 ;
        RECT 844.050 452.850 847.050 454.950 ;
        RECT 850.950 453.900 858.900 454.950 ;
        RECT 860.100 454.050 861.900 455.850 ;
        RECT 850.950 452.850 853.050 453.900 ;
        RECT 832.950 449.400 834.750 451.200 ;
        RECT 833.850 448.200 838.050 449.400 ;
        RECT 844.050 448.200 844.950 452.850 ;
        RECT 852.750 449.100 854.550 449.400 ;
        RECT 826.650 435.750 828.450 447.600 ;
        RECT 830.550 435.750 832.350 447.600 ;
        RECT 835.950 447.300 838.050 448.200 ;
        RECT 838.950 447.300 844.950 448.200 ;
        RECT 846.150 448.800 854.550 449.100 ;
        RECT 862.950 448.800 863.850 461.400 ;
        RECT 846.150 448.200 863.850 448.800 ;
        RECT 838.950 446.400 839.850 447.300 ;
        RECT 837.150 444.600 839.850 446.400 ;
        RECT 840.750 446.100 842.550 446.400 ;
        RECT 846.150 446.100 847.050 448.200 ;
        RECT 852.750 447.600 863.850 448.200 ;
        RECT 840.750 445.200 847.050 446.100 ;
        RECT 847.950 446.700 849.750 447.300 ;
        RECT 847.950 445.500 855.450 446.700 ;
        RECT 840.750 444.600 842.550 445.200 ;
        RECT 854.250 444.600 855.450 445.500 ;
        RECT 835.950 441.600 839.850 443.700 ;
        RECT 844.950 442.500 851.850 444.300 ;
        RECT 854.250 442.500 859.050 444.600 ;
        RECT 833.550 435.750 835.350 438.600 ;
        RECT 838.050 435.750 839.850 441.600 ;
        RECT 842.250 435.750 844.050 441.600 ;
        RECT 846.150 435.750 847.950 442.500 ;
        RECT 854.250 441.600 855.450 442.500 ;
        RECT 849.150 435.750 850.950 441.600 ;
        RECT 853.950 435.750 855.750 441.600 ;
        RECT 859.050 435.750 860.850 441.600 ;
        RECT 862.050 435.750 863.850 447.600 ;
        RECT 10.650 425.400 12.450 431.250 ;
        RECT 13.650 425.400 15.450 431.250 ;
        RECT 16.650 425.400 18.450 431.250 ;
        RECT 14.250 417.150 15.450 425.400 ;
        RECT 27.300 419.400 29.100 431.250 ;
        RECT 31.500 419.400 33.300 431.250 ;
        RECT 34.800 425.400 36.600 431.250 ;
        RECT 49.650 425.400 51.450 431.250 ;
        RECT 52.650 425.400 54.450 431.250 ;
        RECT 10.950 413.850 13.050 415.950 ;
        RECT 13.950 415.050 16.050 417.150 ;
        RECT 11.100 412.050 12.900 413.850 ;
        RECT 14.250 407.700 15.450 415.050 ;
        RECT 16.950 413.850 19.050 415.950 ;
        RECT 26.100 414.150 27.900 415.950 ;
        RECT 31.950 414.150 33.150 419.400 ;
        RECT 34.950 417.150 36.750 418.950 ;
        RECT 34.950 415.050 37.050 417.150 ;
        RECT 17.100 412.050 18.900 413.850 ;
        RECT 25.950 412.050 28.050 414.150 ;
        RECT 28.950 410.850 31.050 412.950 ;
        RECT 31.950 412.050 34.050 414.150 ;
        RECT 50.400 412.950 51.600 425.400 ;
        RECT 62.550 420.300 64.350 431.250 ;
        RECT 65.550 421.200 67.350 431.250 ;
        RECT 68.550 420.300 70.350 431.250 ;
        RECT 62.550 419.400 70.350 420.300 ;
        RECT 71.550 419.400 73.350 431.250 ;
        RECT 85.650 425.400 87.450 431.250 ;
        RECT 88.650 425.400 90.450 431.250 ;
        RECT 91.650 425.400 93.450 431.250 ;
        RECT 101.550 425.400 103.350 431.250 ;
        RECT 104.550 425.400 106.350 431.250 ;
        RECT 71.700 414.150 72.900 419.400 ;
        RECT 89.250 417.150 90.450 425.400 ;
        RECT 29.100 409.050 30.900 410.850 ;
        RECT 32.850 408.750 34.050 412.050 ;
        RECT 49.950 410.850 52.050 412.950 ;
        RECT 53.100 411.150 54.900 412.950 ;
        RECT 33.000 407.700 36.750 408.750 ;
        RECT 11.850 406.800 15.450 407.700 ;
        RECT 11.850 399.750 13.650 406.800 ;
        RECT 16.350 399.750 18.150 405.600 ;
        RECT 26.550 404.700 34.350 406.050 ;
        RECT 26.550 399.750 28.350 404.700 ;
        RECT 29.550 399.750 31.350 403.800 ;
        RECT 32.550 399.750 34.350 404.700 ;
        RECT 35.550 405.600 36.750 407.700 ;
        RECT 35.550 399.750 37.350 405.600 ;
        RECT 50.400 402.600 51.600 410.850 ;
        RECT 52.950 409.050 55.050 411.150 ;
        RECT 61.950 410.850 64.050 412.950 ;
        RECT 65.100 411.150 66.900 412.950 ;
        RECT 62.100 409.050 63.900 410.850 ;
        RECT 64.950 409.050 67.050 411.150 ;
        RECT 67.950 410.850 70.050 412.950 ;
        RECT 70.950 412.050 73.050 414.150 ;
        RECT 85.950 413.850 88.050 415.950 ;
        RECT 88.950 415.050 91.050 417.150 ;
        RECT 86.100 412.050 87.900 413.850 ;
        RECT 68.100 409.050 69.900 410.850 ;
        RECT 71.700 405.600 72.900 412.050 ;
        RECT 89.250 407.700 90.450 415.050 ;
        RECT 91.950 413.850 94.050 415.950 ;
        RECT 101.100 414.150 102.900 415.950 ;
        RECT 92.100 412.050 93.900 413.850 ;
        RECT 100.950 412.050 103.050 414.150 ;
        RECT 104.700 408.300 105.900 425.400 ;
        RECT 108.150 419.400 109.950 431.250 ;
        RECT 111.150 419.400 112.950 431.250 ;
        RECT 122.550 425.400 124.350 431.250 ;
        RECT 125.550 425.400 127.350 431.250 ;
        RECT 128.550 425.400 130.350 431.250 ;
        RECT 106.950 413.850 109.050 415.950 ;
        RECT 111.150 414.150 112.350 419.400 ;
        RECT 125.550 417.150 126.750 425.400 ;
        RECT 140.550 420.300 142.350 431.250 ;
        RECT 143.550 421.200 145.350 431.250 ;
        RECT 146.550 420.300 148.350 431.250 ;
        RECT 140.550 419.400 148.350 420.300 ;
        RECT 149.550 419.400 151.350 431.250 ;
        RECT 161.550 425.400 163.350 431.250 ;
        RECT 164.550 425.400 166.350 431.250 ;
        RECT 167.550 425.400 169.350 431.250 ;
        RECT 185.400 425.400 187.200 431.250 ;
        RECT 107.100 412.050 108.900 413.850 ;
        RECT 109.950 412.050 112.350 414.150 ;
        RECT 121.950 413.850 124.050 415.950 ;
        RECT 124.950 415.050 127.050 417.150 ;
        RECT 122.100 412.050 123.900 413.850 ;
        RECT 49.650 399.750 51.450 402.600 ;
        RECT 52.650 399.750 54.450 402.600 ;
        RECT 63.000 399.750 64.800 405.600 ;
        RECT 67.200 403.950 72.900 405.600 ;
        RECT 86.850 406.800 90.450 407.700 ;
        RECT 101.550 407.100 109.050 408.300 ;
        RECT 67.200 399.750 69.000 403.950 ;
        RECT 70.500 399.750 72.300 402.600 ;
        RECT 86.850 399.750 88.650 406.800 ;
        RECT 91.350 399.750 93.150 405.600 ;
        RECT 101.550 399.750 103.350 407.100 ;
        RECT 107.250 406.500 109.050 407.100 ;
        RECT 111.150 405.600 112.350 412.050 ;
        RECT 125.550 407.700 126.750 415.050 ;
        RECT 127.950 413.850 130.050 415.950 ;
        RECT 149.700 414.150 150.900 419.400 ;
        RECT 164.550 417.150 165.750 425.400 ;
        RECT 188.700 419.400 190.500 431.250 ;
        RECT 192.900 419.400 194.700 431.250 ;
        RECT 204.300 419.400 206.100 431.250 ;
        RECT 208.500 419.400 210.300 431.250 ;
        RECT 211.800 425.400 213.600 431.250 ;
        RECT 228.150 420.900 229.950 431.250 ;
        RECT 227.550 419.550 229.950 420.900 ;
        RECT 231.150 419.550 232.950 431.250 ;
        RECT 185.250 417.150 187.050 418.950 ;
        RECT 128.100 412.050 129.900 413.850 ;
        RECT 139.950 410.850 142.050 412.950 ;
        RECT 143.100 411.150 144.900 412.950 ;
        RECT 140.100 409.050 141.900 410.850 ;
        RECT 142.950 409.050 145.050 411.150 ;
        RECT 145.950 410.850 148.050 412.950 ;
        RECT 148.950 412.050 151.050 414.150 ;
        RECT 160.950 413.850 163.050 415.950 ;
        RECT 163.950 415.050 166.050 417.150 ;
        RECT 161.100 412.050 162.900 413.850 ;
        RECT 146.100 409.050 147.900 410.850 ;
        RECT 125.550 406.800 129.150 407.700 ;
        RECT 106.050 399.750 107.850 405.600 ;
        RECT 109.050 404.100 112.350 405.600 ;
        RECT 109.050 399.750 110.850 404.100 ;
        RECT 122.850 399.750 124.650 405.600 ;
        RECT 127.350 399.750 129.150 406.800 ;
        RECT 149.700 405.600 150.900 412.050 ;
        RECT 164.550 407.700 165.750 415.050 ;
        RECT 166.950 413.850 169.050 415.950 ;
        RECT 184.950 415.050 187.050 417.150 ;
        RECT 188.850 414.150 190.050 419.400 ;
        RECT 194.100 414.150 195.900 415.950 ;
        RECT 203.100 414.150 204.900 415.950 ;
        RECT 208.950 414.150 210.150 419.400 ;
        RECT 211.950 417.150 213.750 418.950 ;
        RECT 211.950 415.050 214.050 417.150 ;
        RECT 167.100 412.050 168.900 413.850 ;
        RECT 187.950 412.050 190.050 414.150 ;
        RECT 187.950 408.750 189.150 412.050 ;
        RECT 190.950 410.850 193.050 412.950 ;
        RECT 193.950 412.050 196.050 414.150 ;
        RECT 202.950 412.050 205.050 414.150 ;
        RECT 205.950 410.850 208.050 412.950 ;
        RECT 208.950 412.050 211.050 414.150 ;
        RECT 227.550 412.950 228.900 419.550 ;
        RECT 235.650 419.400 237.450 431.250 ;
        RECT 245.550 419.400 247.350 431.250 ;
        RECT 249.750 419.400 251.550 431.250 ;
        RECT 265.050 419.400 266.850 431.250 ;
        RECT 268.050 419.400 269.850 431.250 ;
        RECT 271.650 425.400 273.450 431.250 ;
        RECT 274.650 425.400 276.450 431.250 ;
        RECT 289.650 425.400 291.450 431.250 ;
        RECT 292.650 425.400 294.450 431.250 ;
        RECT 295.650 425.400 297.450 431.250 ;
        RECT 230.250 418.200 232.050 418.650 ;
        RECT 236.250 418.200 237.450 419.400 ;
        RECT 230.250 417.000 237.450 418.200 ;
        RECT 249.000 418.350 251.550 419.400 ;
        RECT 230.250 416.850 232.050 417.000 ;
        RECT 191.100 409.050 192.900 410.850 ;
        RECT 206.100 409.050 207.900 410.850 ;
        RECT 209.850 408.750 211.050 412.050 ;
        RECT 226.950 410.850 229.050 412.950 ;
        RECT 185.250 407.700 189.000 408.750 ;
        RECT 210.000 407.700 213.750 408.750 ;
        RECT 164.550 406.800 168.150 407.700 ;
        RECT 141.000 399.750 142.800 405.600 ;
        RECT 145.200 403.950 150.900 405.600 ;
        RECT 145.200 399.750 147.000 403.950 ;
        RECT 148.500 399.750 150.300 402.600 ;
        RECT 161.850 399.750 163.650 405.600 ;
        RECT 166.350 399.750 168.150 406.800 ;
        RECT 185.250 405.600 186.450 407.700 ;
        RECT 184.650 399.750 186.450 405.600 ;
        RECT 187.650 404.700 195.450 406.050 ;
        RECT 187.650 399.750 189.450 404.700 ;
        RECT 190.650 399.750 192.450 403.800 ;
        RECT 193.650 399.750 195.450 404.700 ;
        RECT 203.550 404.700 211.350 406.050 ;
        RECT 203.550 399.750 205.350 404.700 ;
        RECT 206.550 399.750 208.350 403.800 ;
        RECT 209.550 399.750 211.350 404.700 ;
        RECT 212.550 405.600 213.750 407.700 ;
        RECT 226.950 405.600 228.000 410.850 ;
        RECT 230.400 408.600 231.300 416.850 ;
        RECT 233.100 414.150 234.900 415.950 ;
        RECT 245.100 414.150 246.900 415.950 ;
        RECT 232.950 412.050 235.050 414.150 ;
        RECT 236.100 411.150 237.900 412.950 ;
        RECT 244.950 412.050 247.050 414.150 ;
        RECT 249.000 411.150 250.050 418.350 ;
        RECT 251.100 414.150 252.900 415.950 ;
        RECT 265.650 414.150 266.850 419.400 ;
        RECT 250.950 412.050 253.050 414.150 ;
        RECT 265.650 412.050 268.050 414.150 ;
        RECT 268.950 413.850 271.050 415.950 ;
        RECT 269.100 412.050 270.900 413.850 ;
        RECT 235.950 409.050 238.050 411.150 ;
        RECT 247.950 409.050 250.050 411.150 ;
        RECT 230.250 407.700 232.050 408.600 ;
        RECT 230.250 406.800 233.550 407.700 ;
        RECT 212.550 399.750 214.350 405.600 ;
        RECT 226.650 399.750 228.450 405.600 ;
        RECT 232.650 402.600 233.550 406.800 ;
        RECT 238.950 405.450 241.050 406.050 ;
        RECT 244.950 405.450 247.050 406.050 ;
        RECT 238.950 404.550 247.050 405.450 ;
        RECT 238.950 403.950 241.050 404.550 ;
        RECT 244.950 403.950 247.050 404.550 ;
        RECT 249.000 402.600 250.050 409.050 ;
        RECT 265.650 405.600 266.850 412.050 ;
        RECT 272.100 408.300 273.300 425.400 ;
        RECT 293.250 417.150 294.450 425.400 ;
        RECT 306.300 419.400 308.100 431.250 ;
        RECT 310.500 419.400 312.300 431.250 ;
        RECT 313.800 425.400 315.600 431.250 ;
        RECT 328.050 419.400 329.850 431.250 ;
        RECT 331.050 419.400 332.850 431.250 ;
        RECT 334.650 425.400 336.450 431.250 ;
        RECT 337.650 425.400 339.450 431.250 ;
        RECT 349.650 425.400 351.450 431.250 ;
        RECT 352.650 425.400 354.450 431.250 ;
        RECT 355.650 425.400 357.450 431.250 ;
        RECT 275.100 414.150 276.900 415.950 ;
        RECT 274.950 412.050 277.050 414.150 ;
        RECT 289.950 413.850 292.050 415.950 ;
        RECT 292.950 415.050 295.050 417.150 ;
        RECT 290.100 412.050 291.900 413.850 ;
        RECT 268.950 407.100 276.450 408.300 ;
        RECT 293.250 407.700 294.450 415.050 ;
        RECT 295.950 413.850 298.050 415.950 ;
        RECT 305.100 414.150 306.900 415.950 ;
        RECT 310.950 414.150 312.150 419.400 ;
        RECT 313.950 417.150 315.750 418.950 ;
        RECT 313.950 415.050 316.050 417.150 ;
        RECT 328.650 414.150 329.850 419.400 ;
        RECT 296.100 412.050 297.900 413.850 ;
        RECT 304.950 412.050 307.050 414.150 ;
        RECT 307.950 410.850 310.050 412.950 ;
        RECT 310.950 412.050 313.050 414.150 ;
        RECT 308.100 409.050 309.900 410.850 ;
        RECT 311.850 408.750 313.050 412.050 ;
        RECT 328.650 412.050 331.050 414.150 ;
        RECT 331.950 413.850 334.050 415.950 ;
        RECT 332.100 412.050 333.900 413.850 ;
        RECT 312.000 407.700 315.750 408.750 ;
        RECT 268.950 406.500 270.750 407.100 ;
        RECT 265.650 404.100 268.950 405.600 ;
        RECT 229.650 399.750 231.450 402.600 ;
        RECT 232.650 399.750 234.450 402.600 ;
        RECT 235.650 399.750 237.450 402.600 ;
        RECT 245.550 399.750 247.350 402.600 ;
        RECT 248.550 399.750 250.350 402.600 ;
        RECT 251.550 399.750 253.350 402.600 ;
        RECT 267.150 399.750 268.950 404.100 ;
        RECT 270.150 399.750 271.950 405.600 ;
        RECT 274.650 399.750 276.450 407.100 ;
        RECT 290.850 406.800 294.450 407.700 ;
        RECT 290.850 399.750 292.650 406.800 ;
        RECT 295.350 399.750 297.150 405.600 ;
        RECT 305.550 404.700 313.350 406.050 ;
        RECT 305.550 399.750 307.350 404.700 ;
        RECT 308.550 399.750 310.350 403.800 ;
        RECT 311.550 399.750 313.350 404.700 ;
        RECT 314.550 405.600 315.750 407.700 ;
        RECT 328.650 405.600 329.850 412.050 ;
        RECT 335.100 408.300 336.300 425.400 ;
        RECT 353.250 417.150 354.450 425.400 ;
        RECT 368.550 419.400 370.350 431.250 ;
        RECT 372.750 419.400 374.550 431.250 ;
        RECT 388.650 425.400 390.450 431.250 ;
        RECT 391.650 426.000 393.450 431.250 ;
        RECT 372.000 418.350 374.550 419.400 ;
        RECT 389.250 425.100 390.450 425.400 ;
        RECT 394.650 425.400 396.450 431.250 ;
        RECT 397.650 425.400 399.450 431.250 ;
        RECT 394.650 425.100 396.300 425.400 ;
        RECT 389.250 424.200 396.300 425.100 ;
        RECT 338.100 414.150 339.900 415.950 ;
        RECT 337.950 412.050 340.050 414.150 ;
        RECT 349.950 413.850 352.050 415.950 ;
        RECT 352.950 415.050 355.050 417.150 ;
        RECT 350.100 412.050 351.900 413.850 ;
        RECT 331.950 407.100 339.450 408.300 ;
        RECT 353.250 407.700 354.450 415.050 ;
        RECT 355.950 413.850 358.050 415.950 ;
        RECT 368.100 414.150 369.900 415.950 ;
        RECT 356.100 412.050 357.900 413.850 ;
        RECT 367.950 412.050 370.050 414.150 ;
        RECT 372.000 411.150 373.050 418.350 ;
        RECT 389.250 415.950 390.300 424.200 ;
        RECT 395.100 420.150 396.900 421.950 ;
        RECT 391.950 417.150 393.750 418.950 ;
        RECT 394.950 418.050 397.050 420.150 ;
        RECT 409.050 419.400 410.850 431.250 ;
        RECT 412.050 419.400 413.850 431.250 ;
        RECT 415.650 425.400 417.450 431.250 ;
        RECT 418.650 425.400 420.450 431.250 ;
        RECT 398.100 417.150 399.900 418.950 ;
        RECT 374.100 414.150 375.900 415.950 ;
        RECT 373.950 412.050 376.050 414.150 ;
        RECT 388.950 413.850 391.050 415.950 ;
        RECT 391.950 415.050 394.050 417.150 ;
        RECT 397.950 415.050 400.050 417.150 ;
        RECT 409.650 414.150 410.850 419.400 ;
        RECT 370.950 409.050 373.050 411.150 ;
        RECT 331.950 406.500 333.750 407.100 ;
        RECT 314.550 399.750 316.350 405.600 ;
        RECT 328.650 404.100 331.950 405.600 ;
        RECT 330.150 399.750 331.950 404.100 ;
        RECT 333.150 399.750 334.950 405.600 ;
        RECT 337.650 399.750 339.450 407.100 ;
        RECT 350.850 406.800 354.450 407.700 ;
        RECT 358.950 408.450 361.050 409.050 ;
        RECT 367.950 408.450 370.050 409.050 ;
        RECT 358.950 407.550 370.050 408.450 ;
        RECT 358.950 406.950 361.050 407.550 ;
        RECT 367.950 406.950 370.050 407.550 ;
        RECT 350.850 399.750 352.650 406.800 ;
        RECT 355.350 399.750 357.150 405.600 ;
        RECT 372.000 402.600 373.050 409.050 ;
        RECT 389.400 409.650 390.600 413.850 ;
        RECT 409.650 412.050 412.050 414.150 ;
        RECT 412.950 413.850 415.050 415.950 ;
        RECT 413.100 412.050 414.900 413.850 ;
        RECT 389.400 408.000 393.900 409.650 ;
        RECT 368.550 399.750 370.350 402.600 ;
        RECT 371.550 399.750 373.350 402.600 ;
        RECT 374.550 399.750 376.350 402.600 ;
        RECT 392.100 399.750 393.900 408.000 ;
        RECT 397.500 399.750 399.300 408.600 ;
        RECT 409.650 405.600 410.850 412.050 ;
        RECT 416.100 408.300 417.300 425.400 ;
        RECT 432.300 419.400 434.100 431.250 ;
        RECT 436.500 419.400 438.300 431.250 ;
        RECT 439.800 425.400 441.600 431.250 ;
        RECT 454.650 425.400 456.450 431.250 ;
        RECT 457.650 426.000 459.450 431.250 ;
        RECT 455.250 425.100 456.450 425.400 ;
        RECT 460.650 425.400 462.450 431.250 ;
        RECT 463.650 425.400 465.450 431.250 ;
        RECT 473.550 425.400 475.350 431.250 ;
        RECT 476.550 425.400 478.350 431.250 ;
        RECT 479.550 425.400 481.350 431.250 ;
        RECT 494.400 425.400 496.200 431.250 ;
        RECT 460.650 425.100 462.300 425.400 ;
        RECT 455.250 424.200 462.300 425.100 ;
        RECT 419.100 414.150 420.900 415.950 ;
        RECT 431.100 414.150 432.900 415.950 ;
        RECT 436.950 414.150 438.150 419.400 ;
        RECT 439.950 417.150 441.750 418.950 ;
        RECT 439.950 415.050 442.050 417.150 ;
        RECT 455.250 415.950 456.300 424.200 ;
        RECT 461.100 420.150 462.900 421.950 ;
        RECT 457.950 417.150 459.750 418.950 ;
        RECT 460.950 418.050 463.050 420.150 ;
        RECT 464.100 417.150 465.900 418.950 ;
        RECT 476.550 417.150 477.750 425.400 ;
        RECT 478.950 420.450 481.050 421.050 ;
        RECT 484.950 420.450 487.050 421.050 ;
        RECT 478.950 419.550 487.050 420.450 ;
        RECT 478.950 418.950 481.050 419.550 ;
        RECT 484.950 418.950 487.050 419.550 ;
        RECT 497.700 419.400 499.500 431.250 ;
        RECT 501.900 419.400 503.700 431.250 ;
        RECT 514.050 419.400 515.850 431.250 ;
        RECT 517.050 419.400 518.850 431.250 ;
        RECT 520.650 425.400 522.450 431.250 ;
        RECT 523.650 425.400 525.450 431.250 ;
        RECT 494.250 417.150 496.050 418.950 ;
        RECT 418.950 412.050 421.050 414.150 ;
        RECT 430.950 412.050 433.050 414.150 ;
        RECT 433.950 410.850 436.050 412.950 ;
        RECT 436.950 412.050 439.050 414.150 ;
        RECT 454.950 413.850 457.050 415.950 ;
        RECT 457.950 415.050 460.050 417.150 ;
        RECT 463.950 415.050 466.050 417.150 ;
        RECT 472.950 413.850 475.050 415.950 ;
        RECT 475.950 415.050 478.050 417.150 ;
        RECT 434.100 409.050 435.900 410.850 ;
        RECT 437.850 408.750 439.050 412.050 ;
        RECT 455.400 409.650 456.600 413.850 ;
        RECT 473.100 412.050 474.900 413.850 ;
        RECT 412.950 407.100 420.450 408.300 ;
        RECT 438.000 407.700 441.750 408.750 ;
        RECT 455.400 408.000 459.900 409.650 ;
        RECT 412.950 406.500 414.750 407.100 ;
        RECT 409.650 404.100 412.950 405.600 ;
        RECT 411.150 399.750 412.950 404.100 ;
        RECT 414.150 399.750 415.950 405.600 ;
        RECT 418.650 399.750 420.450 407.100 ;
        RECT 431.550 404.700 439.350 406.050 ;
        RECT 431.550 399.750 433.350 404.700 ;
        RECT 434.550 399.750 436.350 403.800 ;
        RECT 437.550 399.750 439.350 404.700 ;
        RECT 440.550 405.600 441.750 407.700 ;
        RECT 440.550 399.750 442.350 405.600 ;
        RECT 458.100 399.750 459.900 408.000 ;
        RECT 463.500 399.750 465.300 408.600 ;
        RECT 476.550 407.700 477.750 415.050 ;
        RECT 478.950 413.850 481.050 415.950 ;
        RECT 493.950 415.050 496.050 417.150 ;
        RECT 497.850 414.150 499.050 419.400 ;
        RECT 503.100 414.150 504.900 415.950 ;
        RECT 514.650 414.150 515.850 419.400 ;
        RECT 479.100 412.050 480.900 413.850 ;
        RECT 496.950 412.050 499.050 414.150 ;
        RECT 496.950 408.750 498.150 412.050 ;
        RECT 499.950 410.850 502.050 412.950 ;
        RECT 502.950 412.050 505.050 414.150 ;
        RECT 514.650 412.050 517.050 414.150 ;
        RECT 517.950 413.850 520.050 415.950 ;
        RECT 518.100 412.050 519.900 413.850 ;
        RECT 500.100 409.050 501.900 410.850 ;
        RECT 494.250 407.700 498.000 408.750 ;
        RECT 476.550 406.800 480.150 407.700 ;
        RECT 473.850 399.750 475.650 405.600 ;
        RECT 478.350 399.750 480.150 406.800 ;
        RECT 494.250 405.600 495.450 407.700 ;
        RECT 493.650 399.750 495.450 405.600 ;
        RECT 496.650 404.700 504.450 406.050 ;
        RECT 496.650 399.750 498.450 404.700 ;
        RECT 499.650 399.750 501.450 403.800 ;
        RECT 502.650 399.750 504.450 404.700 ;
        RECT 514.650 405.600 515.850 412.050 ;
        RECT 521.100 408.300 522.300 425.400 ;
        RECT 533.550 419.400 535.350 431.250 ;
        RECT 537.750 419.400 539.550 431.250 ;
        RECT 551.550 425.400 553.350 431.250 ;
        RECT 554.550 425.400 556.350 431.250 ;
        RECT 557.550 426.000 559.350 431.250 ;
        RECT 554.700 425.100 556.350 425.400 ;
        RECT 560.550 425.400 562.350 431.250 ;
        RECT 572.550 425.400 574.350 431.250 ;
        RECT 575.550 425.400 577.350 431.250 ;
        RECT 578.550 425.400 580.350 431.250 ;
        RECT 560.550 425.100 561.750 425.400 ;
        RECT 554.700 424.200 561.750 425.100 ;
        RECT 554.100 420.150 555.900 421.950 ;
        RECT 537.000 418.350 539.550 419.400 ;
        RECT 524.100 414.150 525.900 415.950 ;
        RECT 533.100 414.150 534.900 415.950 ;
        RECT 523.950 412.050 526.050 414.150 ;
        RECT 532.950 412.050 535.050 414.150 ;
        RECT 537.000 411.150 538.050 418.350 ;
        RECT 551.100 417.150 552.900 418.950 ;
        RECT 553.950 418.050 556.050 420.150 ;
        RECT 557.250 417.150 559.050 418.950 ;
        RECT 539.100 414.150 540.900 415.950 ;
        RECT 550.950 415.050 553.050 417.150 ;
        RECT 556.950 415.050 559.050 417.150 ;
        RECT 560.700 415.950 561.750 424.200 ;
        RECT 575.550 417.150 576.750 425.400 ;
        RECT 592.650 419.400 594.450 431.250 ;
        RECT 595.650 419.400 597.450 431.250 ;
        RECT 608.400 425.400 610.200 431.250 ;
        RECT 611.700 419.400 613.500 431.250 ;
        RECT 615.900 419.400 617.700 431.250 ;
        RECT 626.550 425.400 628.350 431.250 ;
        RECT 629.550 425.400 631.350 431.250 ;
        RECT 632.550 425.400 634.350 431.250 ;
        RECT 538.950 412.050 541.050 414.150 ;
        RECT 559.950 413.850 562.050 415.950 ;
        RECT 571.950 413.850 574.050 415.950 ;
        RECT 574.950 415.050 577.050 417.150 ;
        RECT 535.950 409.050 538.050 411.150 ;
        RECT 560.400 409.650 561.600 413.850 ;
        RECT 572.100 412.050 573.900 413.850 ;
        RECT 517.950 407.100 525.450 408.300 ;
        RECT 517.950 406.500 519.750 407.100 ;
        RECT 514.650 404.100 517.950 405.600 ;
        RECT 516.150 399.750 517.950 404.100 ;
        RECT 519.150 399.750 520.950 405.600 ;
        RECT 523.650 399.750 525.450 407.100 ;
        RECT 537.000 402.600 538.050 409.050 ;
        RECT 533.550 399.750 535.350 402.600 ;
        RECT 536.550 399.750 538.350 402.600 ;
        RECT 539.550 399.750 541.350 402.600 ;
        RECT 551.700 399.750 553.500 408.600 ;
        RECT 557.100 408.000 561.600 409.650 ;
        RECT 557.100 399.750 558.900 408.000 ;
        RECT 575.550 407.700 576.750 415.050 ;
        RECT 577.950 413.850 580.050 415.950 ;
        RECT 593.400 414.150 594.600 419.400 ;
        RECT 608.250 417.150 610.050 418.950 ;
        RECT 607.950 415.050 610.050 417.150 ;
        RECT 611.850 414.150 613.050 419.400 ;
        RECT 629.550 417.150 630.750 425.400 ;
        RECT 644.550 419.400 646.350 431.250 ;
        RECT 647.550 419.400 649.350 431.250 ;
        RECT 659.550 425.400 661.350 431.250 ;
        RECT 662.550 425.400 664.350 431.250 ;
        RECT 617.100 414.150 618.900 415.950 ;
        RECT 578.100 412.050 579.900 413.850 ;
        RECT 592.950 412.050 595.050 414.150 ;
        RECT 575.550 406.800 579.150 407.700 ;
        RECT 572.850 399.750 574.650 405.600 ;
        RECT 577.350 399.750 579.150 406.800 ;
        RECT 593.400 405.600 594.600 412.050 ;
        RECT 595.950 410.850 598.050 412.950 ;
        RECT 610.950 412.050 613.050 414.150 ;
        RECT 596.100 409.050 597.900 410.850 ;
        RECT 610.950 408.750 612.150 412.050 ;
        RECT 613.950 410.850 616.050 412.950 ;
        RECT 616.950 412.050 619.050 414.150 ;
        RECT 625.950 413.850 628.050 415.950 ;
        RECT 628.950 415.050 631.050 417.150 ;
        RECT 626.100 412.050 627.900 413.850 ;
        RECT 614.100 409.050 615.900 410.850 ;
        RECT 608.250 407.700 612.000 408.750 ;
        RECT 629.550 407.700 630.750 415.050 ;
        RECT 631.950 413.850 634.050 415.950 ;
        RECT 647.400 414.150 648.600 419.400 ;
        RECT 632.100 412.050 633.900 413.850 ;
        RECT 643.950 410.850 646.050 412.950 ;
        RECT 646.950 412.050 649.050 414.150 ;
        RECT 662.400 412.950 663.600 425.400 ;
        RECT 668.550 419.400 670.350 431.250 ;
        RECT 671.550 428.400 673.350 431.250 ;
        RECT 676.050 425.400 677.850 431.250 ;
        RECT 680.250 425.400 682.050 431.250 ;
        RECT 673.950 423.300 677.850 425.400 ;
        RECT 684.150 424.500 685.950 431.250 ;
        RECT 687.150 425.400 688.950 431.250 ;
        RECT 691.950 425.400 693.750 431.250 ;
        RECT 697.050 425.400 698.850 431.250 ;
        RECT 692.250 424.500 693.450 425.400 ;
        RECT 682.950 422.700 689.850 424.500 ;
        RECT 692.250 422.400 697.050 424.500 ;
        RECT 675.150 420.600 677.850 422.400 ;
        RECT 678.750 421.800 680.550 422.400 ;
        RECT 678.750 420.900 685.050 421.800 ;
        RECT 692.250 421.500 693.450 422.400 ;
        RECT 678.750 420.600 680.550 420.900 ;
        RECT 676.950 419.700 677.850 420.600 ;
        RECT 644.100 409.050 645.900 410.850 ;
        RECT 608.250 405.600 609.450 407.700 ;
        RECT 629.550 406.800 633.150 407.700 ;
        RECT 592.650 399.750 594.450 405.600 ;
        RECT 595.650 399.750 597.450 405.600 ;
        RECT 607.650 399.750 609.450 405.600 ;
        RECT 610.650 404.700 618.450 406.050 ;
        RECT 610.650 399.750 612.450 404.700 ;
        RECT 613.650 399.750 615.450 403.800 ;
        RECT 616.650 399.750 618.450 404.700 ;
        RECT 626.850 399.750 628.650 405.600 ;
        RECT 631.350 399.750 633.150 406.800 ;
        RECT 647.400 405.600 648.600 412.050 ;
        RECT 659.100 411.150 660.900 412.950 ;
        RECT 658.950 409.050 661.050 411.150 ;
        RECT 661.950 410.850 664.050 412.950 ;
        RECT 644.550 399.750 646.350 405.600 ;
        RECT 647.550 399.750 649.350 405.600 ;
        RECT 662.400 402.600 663.600 410.850 ;
        RECT 668.550 409.950 669.750 419.400 ;
        RECT 673.950 418.800 676.050 419.700 ;
        RECT 676.950 418.800 682.950 419.700 ;
        RECT 671.850 417.600 676.050 418.800 ;
        RECT 670.950 415.800 672.750 417.600 ;
        RECT 682.050 414.150 682.950 418.800 ;
        RECT 684.150 418.800 685.050 420.900 ;
        RECT 685.950 420.300 693.450 421.500 ;
        RECT 685.950 419.700 687.750 420.300 ;
        RECT 700.050 419.400 701.850 431.250 ;
        RECT 690.750 418.800 701.850 419.400 ;
        RECT 684.150 418.200 701.850 418.800 ;
        RECT 684.150 417.900 692.550 418.200 ;
        RECT 690.750 417.600 692.550 417.900 ;
        RECT 682.050 412.050 685.050 414.150 ;
        RECT 688.950 413.100 691.050 414.150 ;
        RECT 688.950 412.050 696.900 413.100 ;
        RECT 670.950 411.750 673.050 412.050 ;
        RECT 670.950 409.950 674.850 411.750 ;
        RECT 668.550 407.850 673.050 409.950 ;
        RECT 682.050 408.000 682.950 412.050 ;
        RECT 695.100 411.300 696.900 412.050 ;
        RECT 698.100 411.150 699.900 412.950 ;
        RECT 692.100 410.400 693.900 411.000 ;
        RECT 698.100 410.400 699.000 411.150 ;
        RECT 692.100 409.200 699.000 410.400 ;
        RECT 692.100 408.000 693.150 409.200 ;
        RECT 668.550 405.600 669.750 407.850 ;
        RECT 682.050 407.100 693.150 408.000 ;
        RECT 682.050 406.800 682.950 407.100 ;
        RECT 659.550 399.750 661.350 402.600 ;
        RECT 662.550 399.750 664.350 402.600 ;
        RECT 668.550 399.750 670.350 405.600 ;
        RECT 673.950 404.700 676.050 405.600 ;
        RECT 681.150 405.000 682.950 406.800 ;
        RECT 692.100 406.200 693.150 407.100 ;
        RECT 688.350 405.450 690.150 406.200 ;
        RECT 673.950 403.500 677.700 404.700 ;
        RECT 676.650 402.600 677.700 403.500 ;
        RECT 685.200 404.400 690.150 405.450 ;
        RECT 691.650 404.400 693.450 406.200 ;
        RECT 700.950 405.600 701.850 418.200 ;
        RECT 685.200 402.600 686.250 404.400 ;
        RECT 694.950 403.500 697.050 405.600 ;
        RECT 694.950 402.600 696.000 403.500 ;
        RECT 671.850 399.750 673.650 402.600 ;
        RECT 676.350 399.750 678.150 402.600 ;
        RECT 680.550 399.750 682.350 402.600 ;
        RECT 684.450 399.750 686.250 402.600 ;
        RECT 687.750 399.750 689.550 402.600 ;
        RECT 692.250 401.700 696.000 402.600 ;
        RECT 692.250 399.750 694.050 401.700 ;
        RECT 697.050 399.750 698.850 402.600 ;
        RECT 700.050 399.750 701.850 405.600 ;
        RECT 705.150 419.400 706.950 431.250 ;
        RECT 708.150 425.400 709.950 431.250 ;
        RECT 713.250 425.400 715.050 431.250 ;
        RECT 718.050 425.400 719.850 431.250 ;
        RECT 713.550 424.500 714.750 425.400 ;
        RECT 721.050 424.500 722.850 431.250 ;
        RECT 724.950 425.400 726.750 431.250 ;
        RECT 729.150 425.400 730.950 431.250 ;
        RECT 733.650 428.400 735.450 431.250 ;
        RECT 709.950 422.400 714.750 424.500 ;
        RECT 717.150 422.700 724.050 424.500 ;
        RECT 729.150 423.300 733.050 425.400 ;
        RECT 713.550 421.500 714.750 422.400 ;
        RECT 726.450 421.800 728.250 422.400 ;
        RECT 713.550 420.300 721.050 421.500 ;
        RECT 719.250 419.700 721.050 420.300 ;
        RECT 721.950 420.900 728.250 421.800 ;
        RECT 705.150 418.800 716.250 419.400 ;
        RECT 721.950 418.800 722.850 420.900 ;
        RECT 726.450 420.600 728.250 420.900 ;
        RECT 729.150 420.600 731.850 422.400 ;
        RECT 729.150 419.700 730.050 420.600 ;
        RECT 705.150 418.200 722.850 418.800 ;
        RECT 705.150 405.600 706.050 418.200 ;
        RECT 714.450 417.900 722.850 418.200 ;
        RECT 724.050 418.800 730.050 419.700 ;
        RECT 730.950 418.800 733.050 419.700 ;
        RECT 736.650 419.400 738.450 431.250 ;
        RECT 750.300 419.400 752.100 431.250 ;
        RECT 754.500 419.400 756.300 431.250 ;
        RECT 757.800 425.400 759.600 431.250 ;
        RECT 770.550 425.400 772.350 431.250 ;
        RECT 773.550 425.400 775.350 431.250 ;
        RECT 776.550 425.400 778.350 431.250 ;
        RECT 714.450 417.600 716.250 417.900 ;
        RECT 724.050 414.150 724.950 418.800 ;
        RECT 730.950 417.600 735.150 418.800 ;
        RECT 734.250 415.800 736.050 417.600 ;
        RECT 715.950 413.100 718.050 414.150 ;
        RECT 707.100 411.150 708.900 412.950 ;
        RECT 710.100 412.050 718.050 413.100 ;
        RECT 721.950 412.050 724.950 414.150 ;
        RECT 710.100 411.300 711.900 412.050 ;
        RECT 708.000 410.400 708.900 411.150 ;
        RECT 713.100 410.400 714.900 411.000 ;
        RECT 708.000 409.200 714.900 410.400 ;
        RECT 713.850 408.000 714.900 409.200 ;
        RECT 724.050 408.000 724.950 412.050 ;
        RECT 733.950 411.750 736.050 412.050 ;
        RECT 732.150 409.950 736.050 411.750 ;
        RECT 737.250 409.950 738.450 419.400 ;
        RECT 749.100 414.150 750.900 415.950 ;
        RECT 754.950 414.150 756.150 419.400 ;
        RECT 757.950 417.150 759.750 418.950 ;
        RECT 773.550 417.150 774.750 425.400 ;
        RECT 788.550 419.400 790.350 431.250 ;
        RECT 791.550 419.400 793.350 431.250 ;
        RECT 794.550 419.400 796.350 431.250 ;
        RECT 800.550 419.400 802.350 431.250 ;
        RECT 803.550 428.400 805.350 431.250 ;
        RECT 808.050 425.400 809.850 431.250 ;
        RECT 812.250 425.400 814.050 431.250 ;
        RECT 805.950 423.300 809.850 425.400 ;
        RECT 816.150 424.500 817.950 431.250 ;
        RECT 819.150 425.400 820.950 431.250 ;
        RECT 823.950 425.400 825.750 431.250 ;
        RECT 829.050 425.400 830.850 431.250 ;
        RECT 824.250 424.500 825.450 425.400 ;
        RECT 814.950 422.700 821.850 424.500 ;
        RECT 824.250 422.400 829.050 424.500 ;
        RECT 807.150 420.600 809.850 422.400 ;
        RECT 810.750 421.800 812.550 422.400 ;
        RECT 810.750 420.900 817.050 421.800 ;
        RECT 824.250 421.500 825.450 422.400 ;
        RECT 810.750 420.600 812.550 420.900 ;
        RECT 808.950 419.700 809.850 420.600 ;
        RECT 757.950 415.050 760.050 417.150 ;
        RECT 748.950 412.050 751.050 414.150 ;
        RECT 751.950 410.850 754.050 412.950 ;
        RECT 754.950 412.050 757.050 414.150 ;
        RECT 769.950 413.850 772.050 415.950 ;
        RECT 772.950 415.050 775.050 417.150 ;
        RECT 770.100 412.050 771.900 413.850 ;
        RECT 713.850 407.100 724.950 408.000 ;
        RECT 733.950 407.850 738.450 409.950 ;
        RECT 752.100 409.050 753.900 410.850 ;
        RECT 755.850 408.750 757.050 412.050 ;
        RECT 713.850 406.200 714.900 407.100 ;
        RECT 724.050 406.800 724.950 407.100 ;
        RECT 705.150 399.750 706.950 405.600 ;
        RECT 709.950 403.500 712.050 405.600 ;
        RECT 713.550 404.400 715.350 406.200 ;
        RECT 716.850 405.450 718.650 406.200 ;
        RECT 716.850 404.400 721.800 405.450 ;
        RECT 724.050 405.000 725.850 406.800 ;
        RECT 737.250 405.600 738.450 407.850 ;
        RECT 756.000 407.700 759.750 408.750 ;
        RECT 730.950 404.700 733.050 405.600 ;
        RECT 711.000 402.600 712.050 403.500 ;
        RECT 720.750 402.600 721.800 404.400 ;
        RECT 729.300 403.500 733.050 404.700 ;
        RECT 729.300 402.600 730.350 403.500 ;
        RECT 708.150 399.750 709.950 402.600 ;
        RECT 711.000 401.700 714.750 402.600 ;
        RECT 712.950 399.750 714.750 401.700 ;
        RECT 717.450 399.750 719.250 402.600 ;
        RECT 720.750 399.750 722.550 402.600 ;
        RECT 724.650 399.750 726.450 402.600 ;
        RECT 728.850 399.750 730.650 402.600 ;
        RECT 733.350 399.750 735.150 402.600 ;
        RECT 736.650 399.750 738.450 405.600 ;
        RECT 749.550 404.700 757.350 406.050 ;
        RECT 749.550 399.750 751.350 404.700 ;
        RECT 752.550 399.750 754.350 403.800 ;
        RECT 755.550 399.750 757.350 404.700 ;
        RECT 758.550 405.600 759.750 407.700 ;
        RECT 773.550 407.700 774.750 415.050 ;
        RECT 775.950 413.850 778.050 415.950 ;
        RECT 776.100 412.050 777.900 413.850 ;
        RECT 791.850 412.950 793.200 419.400 ;
        RECT 787.950 410.850 790.050 412.950 ;
        RECT 791.850 410.850 796.050 412.950 ;
        RECT 788.100 409.050 789.900 410.850 ;
        RECT 773.550 406.800 777.150 407.700 ;
        RECT 758.550 399.750 760.350 405.600 ;
        RECT 770.850 399.750 772.650 405.600 ;
        RECT 775.350 399.750 777.150 406.800 ;
        RECT 791.850 405.600 793.200 410.850 ;
        RECT 800.550 409.950 801.750 419.400 ;
        RECT 805.950 418.800 808.050 419.700 ;
        RECT 808.950 418.800 814.950 419.700 ;
        RECT 803.850 417.600 808.050 418.800 ;
        RECT 802.950 415.800 804.750 417.600 ;
        RECT 814.050 414.150 814.950 418.800 ;
        RECT 816.150 418.800 817.050 420.900 ;
        RECT 817.950 420.300 825.450 421.500 ;
        RECT 817.950 419.700 819.750 420.300 ;
        RECT 832.050 419.400 833.850 431.250 ;
        RECT 843.300 419.400 845.100 431.250 ;
        RECT 847.500 419.400 849.300 431.250 ;
        RECT 850.800 425.400 852.600 431.250 ;
        RECT 822.750 418.800 833.850 419.400 ;
        RECT 816.150 418.200 833.850 418.800 ;
        RECT 816.150 417.900 824.550 418.200 ;
        RECT 822.750 417.600 824.550 417.900 ;
        RECT 814.050 412.050 817.050 414.150 ;
        RECT 820.950 413.100 823.050 414.150 ;
        RECT 820.950 412.050 828.900 413.100 ;
        RECT 802.950 411.750 805.050 412.050 ;
        RECT 802.950 409.950 806.850 411.750 ;
        RECT 800.550 407.850 805.050 409.950 ;
        RECT 814.050 408.000 814.950 412.050 ;
        RECT 827.100 411.300 828.900 412.050 ;
        RECT 830.100 411.150 831.900 412.950 ;
        RECT 824.100 410.400 825.900 411.000 ;
        RECT 830.100 410.400 831.000 411.150 ;
        RECT 824.100 409.200 831.000 410.400 ;
        RECT 824.100 408.000 825.150 409.200 ;
        RECT 800.550 405.600 801.750 407.850 ;
        RECT 814.050 407.100 825.150 408.000 ;
        RECT 814.050 406.800 814.950 407.100 ;
        RECT 788.550 399.750 790.350 405.600 ;
        RECT 791.550 399.750 793.350 405.600 ;
        RECT 794.550 399.750 796.350 405.600 ;
        RECT 800.550 399.750 802.350 405.600 ;
        RECT 805.950 404.700 808.050 405.600 ;
        RECT 813.150 405.000 814.950 406.800 ;
        RECT 824.100 406.200 825.150 407.100 ;
        RECT 820.350 405.450 822.150 406.200 ;
        RECT 805.950 403.500 809.700 404.700 ;
        RECT 808.650 402.600 809.700 403.500 ;
        RECT 817.200 404.400 822.150 405.450 ;
        RECT 823.650 404.400 825.450 406.200 ;
        RECT 832.950 405.600 833.850 418.200 ;
        RECT 842.100 414.150 843.900 415.950 ;
        RECT 847.950 414.150 849.150 419.400 ;
        RECT 850.950 417.150 852.750 418.950 ;
        RECT 850.950 415.050 853.050 417.150 ;
        RECT 841.950 412.050 844.050 414.150 ;
        RECT 844.950 410.850 847.050 412.950 ;
        RECT 847.950 412.050 850.050 414.150 ;
        RECT 845.100 409.050 846.900 410.850 ;
        RECT 848.850 408.750 850.050 412.050 ;
        RECT 849.000 407.700 852.750 408.750 ;
        RECT 817.200 402.600 818.250 404.400 ;
        RECT 826.950 403.500 829.050 405.600 ;
        RECT 826.950 402.600 828.000 403.500 ;
        RECT 803.850 399.750 805.650 402.600 ;
        RECT 808.350 399.750 810.150 402.600 ;
        RECT 812.550 399.750 814.350 402.600 ;
        RECT 816.450 399.750 818.250 402.600 ;
        RECT 819.750 399.750 821.550 402.600 ;
        RECT 824.250 401.700 828.000 402.600 ;
        RECT 824.250 399.750 826.050 401.700 ;
        RECT 829.050 399.750 830.850 402.600 ;
        RECT 832.050 399.750 833.850 405.600 ;
        RECT 842.550 404.700 850.350 406.050 ;
        RECT 842.550 399.750 844.350 404.700 ;
        RECT 845.550 399.750 847.350 403.800 ;
        RECT 848.550 399.750 850.350 404.700 ;
        RECT 851.550 405.600 852.750 407.700 ;
        RECT 851.550 399.750 853.350 405.600 ;
        RECT 10.650 392.400 12.450 395.250 ;
        RECT 13.650 392.400 15.450 395.250 ;
        RECT 23.550 392.400 25.350 395.250 ;
        RECT 26.550 392.400 28.350 395.250 ;
        RECT 41.700 392.400 43.500 395.250 ;
        RECT 11.400 384.150 12.600 392.400 ;
        RECT 10.950 382.050 13.050 384.150 ;
        RECT 13.950 383.850 16.050 385.950 ;
        RECT 22.950 383.850 25.050 385.950 ;
        RECT 26.400 384.150 27.600 392.400 ;
        RECT 45.000 391.050 46.800 395.250 ;
        RECT 41.100 389.400 46.800 391.050 ;
        RECT 49.200 389.400 51.000 395.250 ;
        RECT 14.100 382.050 15.900 383.850 ;
        RECT 23.100 382.050 24.900 383.850 ;
        RECT 25.950 382.050 28.050 384.150 ;
        RECT 41.100 382.950 42.300 389.400 ;
        RECT 59.700 386.400 61.500 395.250 ;
        RECT 65.100 387.000 66.900 395.250 ;
        RECT 80.550 392.400 82.350 395.250 ;
        RECT 83.550 392.400 85.350 395.250 ;
        RECT 95.550 392.400 97.350 395.250 ;
        RECT 98.550 392.400 100.350 395.250 ;
        RECT 101.550 392.400 103.350 395.250 ;
        RECT 44.100 384.150 45.900 385.950 ;
        RECT 11.400 369.600 12.600 382.050 ;
        RECT 26.400 369.600 27.600 382.050 ;
        RECT 40.950 380.850 43.050 382.950 ;
        RECT 43.950 382.050 46.050 384.150 ;
        RECT 46.950 383.850 49.050 385.950 ;
        RECT 50.100 384.150 51.900 385.950 ;
        RECT 65.100 385.350 69.600 387.000 ;
        RECT 47.100 382.050 48.900 383.850 ;
        RECT 49.950 382.050 52.050 384.150 ;
        RECT 68.400 381.150 69.600 385.350 ;
        RECT 79.950 383.850 82.050 385.950 ;
        RECT 83.400 384.150 84.600 392.400 ;
        RECT 99.000 385.950 100.050 392.400 ;
        RECT 113.550 390.300 115.350 395.250 ;
        RECT 116.550 391.200 118.350 395.250 ;
        RECT 119.550 390.300 121.350 395.250 ;
        RECT 113.550 388.950 121.350 390.300 ;
        RECT 122.550 389.400 124.350 395.250 ;
        RECT 138.000 389.400 139.800 395.250 ;
        RECT 142.200 391.050 144.000 395.250 ;
        RECT 145.500 392.400 147.300 395.250 ;
        RECT 142.200 389.400 147.900 391.050 ;
        RECT 160.650 389.400 162.450 395.250 ;
        RECT 122.550 387.300 123.750 389.400 ;
        RECT 120.000 386.250 123.750 387.300 ;
        RECT 80.100 382.050 81.900 383.850 ;
        RECT 82.950 382.050 85.050 384.150 ;
        RECT 97.950 383.850 100.050 385.950 ;
        RECT 116.100 384.150 117.900 385.950 ;
        RECT 41.100 375.600 42.300 380.850 ;
        RECT 58.950 377.850 61.050 379.950 ;
        RECT 64.950 377.850 67.050 379.950 ;
        RECT 67.950 379.050 70.050 381.150 ;
        RECT 59.100 376.050 60.900 377.850 ;
        RECT 10.650 363.750 12.450 369.600 ;
        RECT 13.650 363.750 15.450 369.600 ;
        RECT 23.550 363.750 25.350 369.600 ;
        RECT 26.550 363.750 28.350 369.600 ;
        RECT 40.650 363.750 42.450 375.600 ;
        RECT 43.650 374.700 51.450 375.600 ;
        RECT 61.950 374.850 64.050 376.950 ;
        RECT 65.250 376.050 67.050 377.850 ;
        RECT 43.650 363.750 45.450 374.700 ;
        RECT 46.650 363.750 48.450 373.800 ;
        RECT 49.650 363.750 51.450 374.700 ;
        RECT 62.100 373.050 63.900 374.850 ;
        RECT 68.700 370.800 69.750 379.050 ;
        RECT 62.700 369.900 69.750 370.800 ;
        RECT 62.700 369.600 64.350 369.900 ;
        RECT 59.550 363.750 61.350 369.600 ;
        RECT 62.550 363.750 64.350 369.600 ;
        RECT 68.550 369.600 69.750 369.900 ;
        RECT 83.400 369.600 84.600 382.050 ;
        RECT 94.950 380.850 97.050 382.950 ;
        RECT 95.100 379.050 96.900 380.850 ;
        RECT 99.000 376.650 100.050 383.850 ;
        RECT 100.950 380.850 103.050 382.950 ;
        RECT 112.950 380.850 115.050 382.950 ;
        RECT 115.950 382.050 118.050 384.150 ;
        RECT 119.850 382.950 121.050 386.250 ;
        RECT 137.100 384.150 138.900 385.950 ;
        RECT 118.950 380.850 121.050 382.950 ;
        RECT 136.950 382.050 139.050 384.150 ;
        RECT 139.950 383.850 142.050 385.950 ;
        RECT 143.100 384.150 144.900 385.950 ;
        RECT 140.100 382.050 141.900 383.850 ;
        RECT 142.950 382.050 145.050 384.150 ;
        RECT 146.700 382.950 147.900 389.400 ;
        RECT 161.250 387.300 162.450 389.400 ;
        RECT 163.650 390.300 165.450 395.250 ;
        RECT 166.650 391.200 168.450 395.250 ;
        RECT 169.650 390.300 171.450 395.250 ;
        RECT 163.650 388.950 171.450 390.300 ;
        RECT 182.850 388.200 184.650 395.250 ;
        RECT 187.350 389.400 189.150 395.250 ;
        RECT 182.850 387.300 186.450 388.200 ;
        RECT 161.250 386.250 165.000 387.300 ;
        RECT 163.950 382.950 165.150 386.250 ;
        RECT 167.100 384.150 168.900 385.950 ;
        RECT 145.950 380.850 148.050 382.950 ;
        RECT 163.950 380.850 166.050 382.950 ;
        RECT 166.950 382.050 169.050 384.150 ;
        RECT 169.950 380.850 172.050 382.950 ;
        RECT 182.100 381.150 183.900 382.950 ;
        RECT 101.100 379.050 102.900 380.850 ;
        RECT 113.100 379.050 114.900 380.850 ;
        RECT 99.000 375.600 101.550 376.650 ;
        RECT 118.950 375.600 120.150 380.850 ;
        RECT 121.950 377.850 124.050 379.950 ;
        RECT 121.950 376.050 123.750 377.850 ;
        RECT 146.700 375.600 147.900 380.850 ;
        RECT 160.950 377.850 163.050 379.950 ;
        RECT 161.250 376.050 163.050 377.850 ;
        RECT 164.850 375.600 166.050 380.850 ;
        RECT 170.100 379.050 171.900 380.850 ;
        RECT 181.950 379.050 184.050 381.150 ;
        RECT 185.250 379.950 186.450 387.300 ;
        RECT 197.550 387.900 199.350 395.250 ;
        RECT 202.050 389.400 203.850 395.250 ;
        RECT 205.050 390.900 206.850 395.250 ;
        RECT 205.050 389.400 208.350 390.900 ;
        RECT 203.250 387.900 205.050 388.500 ;
        RECT 197.550 386.700 205.050 387.900 ;
        RECT 188.100 381.150 189.900 382.950 ;
        RECT 184.950 377.850 187.050 379.950 ;
        RECT 187.950 379.050 190.050 381.150 ;
        RECT 196.950 380.850 199.050 382.950 ;
        RECT 197.100 379.050 198.900 380.850 ;
        RECT 65.550 363.750 67.350 369.000 ;
        RECT 68.550 363.750 70.350 369.600 ;
        RECT 80.550 363.750 82.350 369.600 ;
        RECT 83.550 363.750 85.350 369.600 ;
        RECT 95.550 363.750 97.350 375.600 ;
        RECT 99.750 363.750 101.550 375.600 ;
        RECT 114.300 363.750 116.100 375.600 ;
        RECT 118.500 363.750 120.300 375.600 ;
        RECT 137.550 374.700 145.350 375.600 ;
        RECT 121.800 363.750 123.600 369.600 ;
        RECT 137.550 363.750 139.350 374.700 ;
        RECT 140.550 363.750 142.350 373.800 ;
        RECT 143.550 363.750 145.350 374.700 ;
        RECT 146.550 363.750 148.350 375.600 ;
        RECT 161.400 363.750 163.200 369.600 ;
        RECT 164.700 363.750 166.500 375.600 ;
        RECT 168.900 363.750 170.700 375.600 ;
        RECT 185.250 369.600 186.450 377.850 ;
        RECT 200.700 369.600 201.900 386.700 ;
        RECT 207.150 382.950 208.350 389.400 ;
        RECT 224.100 387.000 225.900 395.250 ;
        RECT 203.100 381.150 204.900 382.950 ;
        RECT 202.950 379.050 205.050 381.150 ;
        RECT 205.950 380.850 208.350 382.950 ;
        RECT 221.400 385.350 225.900 387.000 ;
        RECT 229.500 386.400 231.300 395.250 ;
        RECT 239.550 392.400 241.350 395.250 ;
        RECT 242.550 392.400 244.350 395.250 ;
        RECT 221.400 381.150 222.600 385.350 ;
        RECT 238.950 383.850 241.050 385.950 ;
        RECT 242.400 384.150 243.600 392.400 ;
        RECT 254.550 390.300 256.350 395.250 ;
        RECT 257.550 391.200 259.350 395.250 ;
        RECT 260.550 390.300 262.350 395.250 ;
        RECT 254.550 388.950 262.350 390.300 ;
        RECT 263.550 389.400 265.350 395.250 ;
        RECT 277.650 389.400 279.450 395.250 ;
        RECT 263.550 387.300 264.750 389.400 ;
        RECT 261.000 386.250 264.750 387.300 ;
        RECT 278.250 387.300 279.450 389.400 ;
        RECT 280.650 390.300 282.450 395.250 ;
        RECT 283.650 391.200 285.450 395.250 ;
        RECT 286.650 390.300 288.450 395.250 ;
        RECT 280.650 388.950 288.450 390.300 ;
        RECT 296.550 390.300 298.350 395.250 ;
        RECT 299.550 391.200 301.350 395.250 ;
        RECT 302.550 390.300 304.350 395.250 ;
        RECT 296.550 388.950 304.350 390.300 ;
        RECT 305.550 389.400 307.350 395.250 ;
        RECT 305.550 387.300 306.750 389.400 ;
        RECT 278.250 386.250 282.000 387.300 ;
        RECT 303.000 386.250 306.750 387.300 ;
        RECT 323.100 387.000 324.900 395.250 ;
        RECT 257.100 384.150 258.900 385.950 ;
        RECT 239.100 382.050 240.900 383.850 ;
        RECT 241.950 382.050 244.050 384.150 ;
        RECT 207.150 375.600 208.350 380.850 ;
        RECT 220.950 379.050 223.050 381.150 ;
        RECT 181.650 363.750 183.450 369.600 ;
        RECT 184.650 363.750 186.450 369.600 ;
        RECT 187.650 363.750 189.450 369.600 ;
        RECT 197.550 363.750 199.350 369.600 ;
        RECT 200.550 363.750 202.350 369.600 ;
        RECT 204.150 363.750 205.950 375.600 ;
        RECT 207.150 363.750 208.950 375.600 ;
        RECT 221.250 370.800 222.300 379.050 ;
        RECT 223.950 377.850 226.050 379.950 ;
        RECT 229.950 377.850 232.050 379.950 ;
        RECT 223.950 376.050 225.750 377.850 ;
        RECT 226.950 374.850 229.050 376.950 ;
        RECT 230.100 376.050 231.900 377.850 ;
        RECT 227.100 373.050 228.900 374.850 ;
        RECT 221.250 369.900 228.300 370.800 ;
        RECT 221.250 369.600 222.450 369.900 ;
        RECT 220.650 363.750 222.450 369.600 ;
        RECT 226.650 369.600 228.300 369.900 ;
        RECT 242.400 369.600 243.600 382.050 ;
        RECT 253.950 380.850 256.050 382.950 ;
        RECT 256.950 382.050 259.050 384.150 ;
        RECT 260.850 382.950 262.050 386.250 ;
        RECT 268.950 382.950 271.050 385.050 ;
        RECT 280.950 382.950 282.150 386.250 ;
        RECT 284.100 384.150 285.900 385.950 ;
        RECT 299.100 384.150 300.900 385.950 ;
        RECT 259.950 380.850 262.050 382.950 ;
        RECT 254.100 379.050 255.900 380.850 ;
        RECT 259.950 375.600 261.150 380.850 ;
        RECT 262.950 377.850 265.050 379.950 ;
        RECT 262.950 376.050 264.750 377.850 ;
        RECT 223.650 363.750 225.450 369.000 ;
        RECT 226.650 363.750 228.450 369.600 ;
        RECT 229.650 363.750 231.450 369.600 ;
        RECT 239.550 363.750 241.350 369.600 ;
        RECT 242.550 363.750 244.350 369.600 ;
        RECT 255.300 363.750 257.100 375.600 ;
        RECT 259.500 363.750 261.300 375.600 ;
        RECT 269.550 375.450 270.450 382.950 ;
        RECT 280.950 380.850 283.050 382.950 ;
        RECT 283.950 382.050 286.050 384.150 ;
        RECT 286.950 380.850 289.050 382.950 ;
        RECT 295.950 380.850 298.050 382.950 ;
        RECT 298.950 382.050 301.050 384.150 ;
        RECT 302.850 382.950 304.050 386.250 ;
        RECT 301.950 380.850 304.050 382.950 ;
        RECT 320.400 385.350 324.900 387.000 ;
        RECT 328.500 386.400 330.300 395.250 ;
        RECT 341.700 392.400 343.500 395.250 ;
        RECT 345.000 391.050 346.800 395.250 ;
        RECT 341.100 389.400 346.800 391.050 ;
        RECT 349.200 389.400 351.000 395.250 ;
        RECT 359.850 389.400 361.650 395.250 ;
        RECT 320.400 381.150 321.600 385.350 ;
        RECT 341.100 382.950 342.300 389.400 ;
        RECT 364.350 388.200 366.150 395.250 ;
        RECT 382.650 389.400 384.450 395.250 ;
        RECT 362.550 387.300 366.150 388.200 ;
        RECT 383.250 387.300 384.450 389.400 ;
        RECT 385.650 390.300 387.450 395.250 ;
        RECT 388.650 391.200 390.450 395.250 ;
        RECT 391.650 390.300 393.450 395.250 ;
        RECT 385.650 388.950 393.450 390.300 ;
        RECT 401.550 390.300 403.350 395.250 ;
        RECT 404.550 391.200 406.350 395.250 ;
        RECT 407.550 390.300 409.350 395.250 ;
        RECT 401.550 388.950 409.350 390.300 ;
        RECT 410.550 389.400 412.350 395.250 ;
        RECT 425.700 392.400 427.500 395.250 ;
        RECT 429.000 391.050 430.800 395.250 ;
        RECT 410.550 387.300 411.750 389.400 ;
        RECT 421.950 388.950 424.050 391.050 ;
        RECT 425.100 389.400 430.800 391.050 ;
        RECT 433.200 389.400 435.000 395.250 ;
        RECT 445.650 392.400 447.450 395.250 ;
        RECT 448.650 392.400 450.450 395.250 ;
        RECT 344.100 384.150 345.900 385.950 ;
        RECT 277.950 377.850 280.050 379.950 ;
        RECT 278.250 376.050 280.050 377.850 ;
        RECT 281.850 375.600 283.050 380.850 ;
        RECT 287.100 379.050 288.900 380.850 ;
        RECT 296.100 379.050 297.900 380.850 ;
        RECT 301.950 375.600 303.150 380.850 ;
        RECT 304.950 377.850 307.050 379.950 ;
        RECT 319.950 379.050 322.050 381.150 ;
        RECT 340.950 380.850 343.050 382.950 ;
        RECT 343.950 382.050 346.050 384.150 ;
        RECT 346.950 383.850 349.050 385.950 ;
        RECT 350.100 384.150 351.900 385.950 ;
        RECT 347.100 382.050 348.900 383.850 ;
        RECT 349.950 382.050 352.050 384.150 ;
        RECT 359.100 381.150 360.900 382.950 ;
        RECT 304.950 376.050 306.750 377.850 ;
        RECT 269.550 374.550 276.450 375.450 ;
        RECT 262.950 372.450 265.050 373.050 ;
        RECT 271.950 372.450 274.050 373.050 ;
        RECT 262.950 371.550 274.050 372.450 ;
        RECT 262.950 370.950 265.050 371.550 ;
        RECT 271.950 370.950 274.050 371.550 ;
        RECT 262.800 363.750 264.600 369.600 ;
        RECT 271.950 369.450 274.050 370.050 ;
        RECT 275.550 369.450 276.450 374.550 ;
        RECT 271.950 368.550 276.450 369.450 ;
        RECT 271.950 367.950 274.050 368.550 ;
        RECT 278.400 363.750 280.200 369.600 ;
        RECT 281.700 363.750 283.500 375.600 ;
        RECT 285.900 363.750 287.700 375.600 ;
        RECT 297.300 363.750 299.100 375.600 ;
        RECT 301.500 363.750 303.300 375.600 ;
        RECT 320.250 370.800 321.300 379.050 ;
        RECT 322.950 377.850 325.050 379.950 ;
        RECT 328.950 377.850 331.050 379.950 ;
        RECT 322.950 376.050 324.750 377.850 ;
        RECT 325.950 374.850 328.050 376.950 ;
        RECT 329.100 376.050 330.900 377.850 ;
        RECT 341.100 375.600 342.300 380.850 ;
        RECT 358.950 379.050 361.050 381.150 ;
        RECT 362.550 379.950 363.750 387.300 ;
        RECT 383.250 386.250 387.000 387.300 ;
        RECT 408.000 386.250 411.750 387.300 ;
        RECT 385.950 382.950 387.150 386.250 ;
        RECT 389.100 384.150 390.900 385.950 ;
        RECT 404.100 384.150 405.900 385.950 ;
        RECT 365.100 381.150 366.900 382.950 ;
        RECT 361.950 377.850 364.050 379.950 ;
        RECT 364.950 379.050 367.050 381.150 ;
        RECT 385.950 380.850 388.050 382.950 ;
        RECT 388.950 382.050 391.050 384.150 ;
        RECT 391.950 380.850 394.050 382.950 ;
        RECT 400.950 380.850 403.050 382.950 ;
        RECT 403.950 382.050 406.050 384.150 ;
        RECT 407.850 382.950 409.050 386.250 ;
        RECT 406.950 380.850 409.050 382.950 ;
        RECT 382.950 377.850 385.050 379.950 ;
        RECT 326.100 373.050 327.900 374.850 ;
        RECT 320.250 369.900 327.300 370.800 ;
        RECT 320.250 369.600 321.450 369.900 ;
        RECT 304.800 363.750 306.600 369.600 ;
        RECT 319.650 363.750 321.450 369.600 ;
        RECT 325.650 369.600 327.300 369.900 ;
        RECT 322.650 363.750 324.450 369.000 ;
        RECT 325.650 363.750 327.450 369.600 ;
        RECT 328.650 363.750 330.450 369.600 ;
        RECT 340.650 363.750 342.450 375.600 ;
        RECT 343.650 374.700 351.450 375.600 ;
        RECT 343.650 363.750 345.450 374.700 ;
        RECT 346.650 363.750 348.450 373.800 ;
        RECT 349.650 363.750 351.450 374.700 ;
        RECT 362.550 369.600 363.750 377.850 ;
        RECT 383.250 376.050 385.050 377.850 ;
        RECT 386.850 375.600 388.050 380.850 ;
        RECT 392.100 379.050 393.900 380.850 ;
        RECT 401.100 379.050 402.900 380.850 ;
        RECT 406.950 375.600 408.150 380.850 ;
        RECT 409.950 377.850 412.050 379.950 ;
        RECT 422.550 379.050 423.450 388.950 ;
        RECT 425.100 382.950 426.300 389.400 ;
        RECT 428.100 384.150 429.900 385.950 ;
        RECT 424.950 380.850 427.050 382.950 ;
        RECT 427.950 382.050 430.050 384.150 ;
        RECT 430.950 383.850 433.050 385.950 ;
        RECT 434.100 384.150 435.900 385.950 ;
        RECT 446.400 384.150 447.600 392.400 ;
        RECT 458.550 390.300 460.350 395.250 ;
        RECT 461.550 391.200 463.350 395.250 ;
        RECT 464.550 390.300 466.350 395.250 ;
        RECT 458.550 388.950 466.350 390.300 ;
        RECT 467.550 389.400 469.350 395.250 ;
        RECT 482.850 389.400 484.650 395.250 ;
        RECT 467.550 387.300 468.750 389.400 ;
        RECT 487.350 388.200 489.150 395.250 ;
        RECT 465.000 386.250 468.750 387.300 ;
        RECT 475.950 387.450 478.050 388.050 ;
        RECT 481.950 387.450 484.050 388.050 ;
        RECT 475.950 386.550 484.050 387.450 ;
        RECT 431.100 382.050 432.900 383.850 ;
        RECT 433.950 382.050 436.050 384.150 ;
        RECT 445.950 382.050 448.050 384.150 ;
        RECT 448.950 383.850 451.050 385.950 ;
        RECT 461.100 384.150 462.900 385.950 ;
        RECT 449.100 382.050 450.900 383.850 ;
        RECT 409.950 376.050 411.750 377.850 ;
        RECT 421.950 376.950 424.050 379.050 ;
        RECT 425.100 375.600 426.300 380.850 ;
        RECT 359.550 363.750 361.350 369.600 ;
        RECT 362.550 363.750 364.350 369.600 ;
        RECT 365.550 363.750 367.350 369.600 ;
        RECT 383.400 363.750 385.200 369.600 ;
        RECT 386.700 363.750 388.500 375.600 ;
        RECT 390.900 363.750 392.700 375.600 ;
        RECT 402.300 363.750 404.100 375.600 ;
        RECT 406.500 363.750 408.300 375.600 ;
        RECT 409.800 363.750 411.600 369.600 ;
        RECT 424.650 363.750 426.450 375.600 ;
        RECT 427.650 374.700 435.450 375.600 ;
        RECT 427.650 363.750 429.450 374.700 ;
        RECT 430.650 363.750 432.450 373.800 ;
        RECT 433.650 363.750 435.450 374.700 ;
        RECT 446.400 369.600 447.600 382.050 ;
        RECT 457.950 380.850 460.050 382.950 ;
        RECT 460.950 382.050 463.050 384.150 ;
        RECT 464.850 382.950 466.050 386.250 ;
        RECT 475.950 385.950 478.050 386.550 ;
        RECT 481.950 385.950 484.050 386.550 ;
        RECT 485.550 387.300 489.150 388.200 ;
        RECT 466.950 384.450 469.050 385.050 ;
        RECT 466.950 383.550 471.450 384.450 ;
        RECT 466.950 382.950 469.050 383.550 ;
        RECT 463.950 380.850 466.050 382.950 ;
        RECT 470.550 381.450 471.450 383.550 ;
        RECT 478.950 381.450 481.050 382.050 ;
        RECT 458.100 379.050 459.900 380.850 ;
        RECT 463.950 375.600 465.150 380.850 ;
        RECT 470.550 380.550 481.050 381.450 ;
        RECT 482.100 381.150 483.900 382.950 ;
        RECT 478.950 379.950 481.050 380.550 ;
        RECT 466.950 377.850 469.050 379.950 ;
        RECT 481.950 379.050 484.050 381.150 ;
        RECT 485.550 379.950 486.750 387.300 ;
        RECT 506.100 387.000 507.900 395.250 ;
        RECT 503.400 385.350 507.900 387.000 ;
        RECT 511.500 386.400 513.300 395.250 ;
        RECT 521.550 387.900 523.350 395.250 ;
        RECT 526.050 389.400 527.850 395.250 ;
        RECT 529.050 390.900 530.850 395.250 ;
        RECT 529.050 389.400 532.350 390.900 ;
        RECT 542.850 389.400 544.650 395.250 ;
        RECT 527.250 387.900 529.050 388.500 ;
        RECT 521.550 386.700 529.050 387.900 ;
        RECT 488.100 381.150 489.900 382.950 ;
        RECT 503.400 381.150 504.600 385.350 ;
        RECT 484.950 377.850 487.050 379.950 ;
        RECT 487.950 379.050 490.050 381.150 ;
        RECT 502.950 379.050 505.050 381.150 ;
        RECT 520.950 380.850 523.050 382.950 ;
        RECT 466.950 376.050 468.750 377.850 ;
        RECT 445.650 363.750 447.450 369.600 ;
        RECT 448.650 363.750 450.450 369.600 ;
        RECT 459.300 363.750 461.100 375.600 ;
        RECT 463.500 363.750 465.300 375.600 ;
        RECT 485.550 369.600 486.750 377.850 ;
        RECT 503.250 370.800 504.300 379.050 ;
        RECT 505.950 377.850 508.050 379.950 ;
        RECT 511.950 377.850 514.050 379.950 ;
        RECT 521.100 379.050 522.900 380.850 ;
        RECT 505.950 376.050 507.750 377.850 ;
        RECT 508.950 374.850 511.050 376.950 ;
        RECT 512.100 376.050 513.900 377.850 ;
        RECT 509.100 373.050 510.900 374.850 ;
        RECT 503.250 369.900 510.300 370.800 ;
        RECT 503.250 369.600 504.450 369.900 ;
        RECT 466.800 363.750 468.600 369.600 ;
        RECT 482.550 363.750 484.350 369.600 ;
        RECT 485.550 363.750 487.350 369.600 ;
        RECT 488.550 363.750 490.350 369.600 ;
        RECT 502.650 363.750 504.450 369.600 ;
        RECT 508.650 369.600 510.300 369.900 ;
        RECT 524.700 369.600 525.900 386.700 ;
        RECT 531.150 382.950 532.350 389.400 ;
        RECT 547.350 388.200 549.150 395.250 ;
        RECT 561.000 389.400 562.800 395.250 ;
        RECT 565.200 389.400 567.000 395.250 ;
        RECT 569.400 389.400 571.200 395.250 ;
        RECT 584.550 392.400 586.350 395.250 ;
        RECT 587.550 392.400 589.350 395.250 ;
        RECT 590.550 392.400 592.350 395.250 ;
        RECT 597.750 392.400 599.550 395.250 ;
        RECT 600.750 392.400 602.550 395.250 ;
        RECT 545.550 387.300 549.150 388.200 ;
        RECT 527.100 381.150 528.900 382.950 ;
        RECT 526.950 379.050 529.050 381.150 ;
        RECT 529.950 380.850 532.350 382.950 ;
        RECT 542.100 381.150 543.900 382.950 ;
        RECT 531.150 375.600 532.350 380.850 ;
        RECT 541.950 379.050 544.050 381.150 ;
        RECT 545.550 379.950 546.750 387.300 ;
        RECT 563.250 384.150 565.050 385.950 ;
        RECT 548.100 381.150 549.900 382.950 ;
        RECT 544.950 377.850 547.050 379.950 ;
        RECT 547.950 379.050 550.050 381.150 ;
        RECT 559.950 380.850 562.050 382.950 ;
        RECT 562.950 382.050 565.050 384.150 ;
        RECT 565.950 382.950 567.000 389.400 ;
        RECT 588.000 385.950 589.050 392.400 ;
        RECT 568.950 384.150 570.750 385.950 ;
        RECT 565.950 380.850 568.050 382.950 ;
        RECT 568.950 382.050 571.050 384.150 ;
        RECT 586.950 383.850 589.050 385.950 ;
        RECT 601.050 384.150 602.550 392.400 ;
        RECT 571.950 380.850 574.050 382.950 ;
        RECT 583.950 380.850 586.050 382.950 ;
        RECT 560.250 379.050 562.050 380.850 ;
        RECT 505.650 363.750 507.450 369.000 ;
        RECT 508.650 363.750 510.450 369.600 ;
        RECT 511.650 363.750 513.450 369.600 ;
        RECT 521.550 363.750 523.350 369.600 ;
        RECT 524.550 363.750 526.350 369.600 ;
        RECT 528.150 363.750 529.950 375.600 ;
        RECT 531.150 363.750 532.950 375.600 ;
        RECT 545.550 369.600 546.750 377.850 ;
        RECT 567.150 377.400 568.050 380.850 ;
        RECT 572.100 379.050 573.900 380.850 ;
        RECT 584.100 379.050 585.900 380.850 ;
        RECT 567.150 376.500 571.200 377.400 ;
        RECT 569.400 375.600 571.200 376.500 ;
        RECT 588.000 376.650 589.050 383.850 ;
        RECT 589.950 380.850 592.050 382.950 ;
        RECT 598.950 382.050 602.550 384.150 ;
        RECT 590.100 379.050 591.900 380.850 ;
        RECT 588.000 375.600 590.550 376.650 ;
        RECT 560.550 374.400 568.350 375.300 ;
        RECT 542.550 363.750 544.350 369.600 ;
        RECT 545.550 363.750 547.350 369.600 ;
        RECT 548.550 363.750 550.350 369.600 ;
        RECT 560.550 363.750 562.350 374.400 ;
        RECT 563.550 363.750 565.350 373.500 ;
        RECT 566.550 364.500 568.350 374.400 ;
        RECT 569.550 365.400 571.350 375.600 ;
        RECT 572.550 364.500 574.350 375.600 ;
        RECT 566.550 363.750 574.350 364.500 ;
        RECT 584.550 363.750 586.350 375.600 ;
        RECT 588.750 363.750 590.550 375.600 ;
        RECT 601.050 369.600 602.550 382.050 ;
        RECT 604.650 389.400 606.450 395.250 ;
        RECT 610.050 389.400 611.850 395.250 ;
        RECT 615.600 390.600 617.400 395.250 ;
        RECT 620.250 391.500 622.050 395.250 ;
        RECT 623.250 391.500 625.050 395.250 ;
        RECT 626.250 391.500 628.050 395.250 ;
        RECT 613.200 389.400 617.400 390.600 ;
        RECT 619.950 389.400 622.050 391.500 ;
        RECT 622.950 389.400 625.050 391.500 ;
        RECT 625.950 389.400 628.050 391.500 ;
        RECT 630.000 391.500 631.800 395.250 ;
        RECT 633.000 392.400 634.800 395.250 ;
        RECT 636.000 391.500 637.800 395.250 ;
        RECT 640.500 392.400 642.300 395.250 ;
        RECT 643.500 392.400 645.300 395.250 ;
        RECT 646.500 392.400 648.300 395.250 ;
        RECT 649.500 392.400 651.300 395.250 ;
        RECT 630.000 389.700 632.850 391.500 ;
        RECT 630.750 389.400 632.850 389.700 ;
        RECT 634.950 389.700 637.800 391.500 ;
        RECT 638.700 390.750 640.500 391.200 ;
        RECT 643.950 391.050 645.300 392.400 ;
        RECT 646.950 391.050 648.300 392.400 ;
        RECT 649.950 391.050 651.300 392.400 ;
        RECT 634.950 389.400 637.050 389.700 ;
        RECT 638.700 389.400 642.750 390.750 ;
        RECT 604.650 374.550 605.850 389.400 ;
        RECT 613.200 385.800 614.700 389.400 ;
        RECT 619.350 386.700 626.100 388.500 ;
        RECT 627.000 386.700 633.900 388.500 ;
        RECT 641.850 388.050 642.750 389.400 ;
        RECT 643.950 388.950 646.050 391.050 ;
        RECT 646.950 388.950 649.050 391.050 ;
        RECT 649.950 388.950 652.050 391.050 ;
        RECT 641.850 387.900 646.950 388.050 ;
        RECT 641.850 387.150 649.500 387.900 ;
        RECT 645.150 386.700 649.500 387.150 ;
        RECT 627.000 385.800 628.050 386.700 ;
        RECT 645.150 386.250 646.950 386.700 ;
        RECT 606.900 384.000 614.700 385.800 ;
        RECT 618.150 384.750 628.050 385.800 ;
        RECT 618.150 382.950 619.200 384.750 ;
        RECT 628.950 384.450 636.600 385.800 ;
        RECT 628.950 383.700 629.850 384.450 ;
        RECT 610.950 381.900 619.200 382.950 ;
        RECT 620.250 382.650 629.850 383.700 ;
        RECT 610.950 377.850 613.050 381.900 ;
        RECT 620.250 381.000 621.150 382.650 ;
        RECT 630.750 381.750 634.650 383.550 ;
        RECT 635.550 382.950 636.600 384.450 ;
        RECT 637.950 385.650 640.050 385.950 ;
        RECT 637.950 383.850 641.850 385.650 ;
        RECT 648.450 383.250 649.500 386.700 ;
        RECT 651.000 385.800 652.050 388.950 ;
        RECT 653.700 389.400 655.500 395.250 ;
        RECT 659.100 389.400 660.900 395.250 ;
        RECT 664.500 389.400 666.300 395.250 ;
        RECT 653.700 388.500 655.200 389.400 ;
        RECT 653.700 387.300 662.100 388.500 ;
        RECT 660.300 386.700 662.100 387.300 ;
        RECT 665.100 385.800 666.300 389.400 ;
        RECT 651.000 384.900 666.300 385.800 ;
        RECT 635.550 382.050 647.550 382.950 ;
        RECT 614.100 379.200 621.150 381.000 ;
        RECT 622.500 379.950 624.300 381.750 ;
        RECT 630.750 381.450 632.850 381.750 ;
        RECT 634.950 380.550 637.050 380.850 ;
        RECT 643.800 380.550 645.600 381.150 ;
        RECT 634.950 379.950 645.600 380.550 ;
        RECT 622.500 379.350 645.600 379.950 ;
        RECT 646.500 380.550 647.550 382.050 ;
        RECT 648.450 381.450 650.250 383.250 ;
        RECT 652.050 382.950 663.900 384.000 ;
        RECT 652.050 380.550 653.250 382.950 ;
        RECT 662.100 381.150 663.900 382.950 ;
        RECT 646.500 379.650 653.250 380.550 ;
        RECT 655.950 379.650 658.050 379.950 ;
        RECT 622.500 378.750 637.050 379.350 ;
        RECT 654.150 378.450 658.050 379.650 ;
        RECT 661.950 379.050 664.050 381.150 ;
        RECT 644.100 377.850 658.050 378.450 ;
        RECT 618.000 377.550 657.750 377.850 ;
        RECT 606.750 376.650 608.550 377.250 ;
        RECT 618.000 376.650 646.050 377.550 ;
        RECT 606.750 375.450 619.050 376.650 ;
        RECT 646.950 376.050 649.050 376.350 ;
        RECT 656.700 376.050 658.500 376.650 ;
        RECT 619.950 374.550 622.050 375.750 ;
        RECT 604.650 373.650 622.050 374.550 ;
        RECT 625.950 374.400 646.050 375.750 ;
        RECT 625.950 373.650 628.050 374.400 ;
        RECT 607.500 369.600 608.700 373.650 ;
        RECT 609.600 371.700 611.400 372.300 ;
        RECT 616.350 372.150 618.150 372.300 ;
        RECT 609.600 370.500 615.300 371.700 ;
        RECT 616.350 370.950 625.050 372.150 ;
        RECT 616.350 370.500 618.150 370.950 ;
        RECT 597.750 363.750 599.550 369.600 ;
        RECT 600.750 363.750 602.550 369.600 ;
        RECT 604.500 363.750 606.300 369.600 ;
        RECT 607.500 363.750 609.300 369.600 ;
        RECT 610.500 363.750 612.300 369.600 ;
        RECT 613.500 363.750 615.300 370.500 ;
        RECT 622.950 370.050 625.050 370.950 ;
        RECT 616.500 363.750 618.300 369.600 ;
        RECT 619.800 367.800 621.900 369.900 ;
        RECT 620.400 366.600 621.900 367.800 ;
        RECT 620.250 363.750 622.050 366.600 ;
        RECT 623.250 363.750 625.050 370.050 ;
        RECT 626.550 366.600 627.900 373.650 ;
        RECT 644.100 373.350 646.050 374.400 ;
        RECT 646.950 374.850 658.500 376.050 ;
        RECT 646.950 374.250 649.050 374.850 ;
        RECT 660.000 373.350 661.800 374.100 ;
        RECT 629.100 370.800 633.000 372.600 ;
        RECT 630.000 370.500 633.000 370.800 ;
        RECT 634.950 372.150 637.050 372.600 ;
        RECT 644.100 372.300 661.800 373.350 ;
        RECT 634.950 370.500 637.350 372.150 ;
        RECT 626.250 363.750 628.050 366.600 ;
        RECT 630.000 363.750 631.800 370.500 ;
        RECT 636.000 369.600 637.350 370.500 ;
        RECT 643.950 369.600 646.050 370.050 ;
        RECT 633.000 363.750 634.800 369.600 ;
        RECT 636.000 363.750 637.800 369.600 ;
        RECT 639.750 363.750 641.550 369.600 ;
        RECT 643.500 367.950 646.050 369.600 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 643.500 366.600 644.700 367.950 ;
        RECT 646.950 366.600 647.850 367.950 ;
        RECT 649.950 366.600 651.150 367.950 ;
        RECT 642.750 363.750 644.700 366.600 ;
        RECT 645.750 363.750 647.850 366.600 ;
        RECT 648.750 363.750 651.150 366.600 ;
        RECT 652.500 363.750 654.300 367.050 ;
        RECT 655.500 363.750 657.300 372.300 ;
        RECT 665.100 371.400 666.300 384.900 ;
        RECT 662.250 370.500 666.300 371.400 ;
        RECT 668.700 389.400 670.500 395.250 ;
        RECT 674.100 389.400 675.900 395.250 ;
        RECT 679.500 389.400 681.300 395.250 ;
        RECT 683.700 392.400 685.500 395.250 ;
        RECT 686.700 392.400 688.500 395.250 ;
        RECT 689.700 392.400 691.500 395.250 ;
        RECT 692.700 392.400 694.500 395.250 ;
        RECT 683.700 391.050 685.050 392.400 ;
        RECT 686.700 391.050 688.050 392.400 ;
        RECT 689.700 391.050 691.050 392.400 ;
        RECT 697.200 391.500 699.000 395.250 ;
        RECT 700.200 392.400 702.000 395.250 ;
        RECT 703.200 391.500 705.000 395.250 ;
        RECT 668.700 385.800 669.900 389.400 ;
        RECT 679.800 388.500 681.300 389.400 ;
        RECT 672.900 387.300 681.300 388.500 ;
        RECT 682.950 388.950 685.050 391.050 ;
        RECT 685.950 388.950 688.050 391.050 ;
        RECT 688.950 388.950 691.050 391.050 ;
        RECT 694.500 390.750 696.300 391.200 ;
        RECT 692.250 389.400 696.300 390.750 ;
        RECT 697.200 389.700 700.050 391.500 ;
        RECT 697.950 389.400 700.050 389.700 ;
        RECT 702.150 389.700 705.000 391.500 ;
        RECT 706.950 391.500 708.750 395.250 ;
        RECT 709.950 391.500 711.750 395.250 ;
        RECT 712.950 391.500 714.750 395.250 ;
        RECT 702.150 389.400 704.250 389.700 ;
        RECT 706.950 389.400 709.050 391.500 ;
        RECT 709.950 389.400 712.050 391.500 ;
        RECT 712.950 389.400 715.050 391.500 ;
        RECT 717.600 390.600 719.400 395.250 ;
        RECT 717.600 389.400 721.800 390.600 ;
        RECT 723.150 389.400 724.950 395.250 ;
        RECT 728.550 389.400 730.350 395.250 ;
        RECT 672.900 386.700 674.700 387.300 ;
        RECT 682.950 385.800 684.000 388.950 ;
        RECT 692.250 388.050 693.150 389.400 ;
        RECT 688.050 387.900 693.150 388.050 ;
        RECT 668.700 384.900 684.000 385.800 ;
        RECT 685.500 387.150 693.150 387.900 ;
        RECT 685.500 386.700 689.850 387.150 ;
        RECT 701.100 386.700 708.000 388.500 ;
        RECT 708.900 386.700 715.650 388.500 ;
        RECT 668.700 371.400 669.900 384.900 ;
        RECT 671.100 382.950 682.950 384.000 ;
        RECT 685.500 383.250 686.550 386.700 ;
        RECT 688.050 386.250 689.850 386.700 ;
        RECT 694.950 385.650 697.050 385.950 ;
        RECT 706.950 385.800 708.000 386.700 ;
        RECT 720.300 385.800 721.800 389.400 ;
        RECT 693.150 383.850 697.050 385.650 ;
        RECT 698.400 384.450 706.050 385.800 ;
        RECT 706.950 384.750 716.850 385.800 ;
        RECT 671.100 381.150 672.900 382.950 ;
        RECT 670.950 379.050 673.050 381.150 ;
        RECT 681.750 380.550 682.950 382.950 ;
        RECT 684.750 381.450 686.550 383.250 ;
        RECT 698.400 382.950 699.450 384.450 ;
        RECT 705.150 383.700 706.050 384.450 ;
        RECT 687.450 382.050 699.450 382.950 ;
        RECT 687.450 380.550 688.500 382.050 ;
        RECT 700.350 381.750 704.250 383.550 ;
        RECT 705.150 382.650 714.750 383.700 ;
        RECT 702.150 381.450 704.250 381.750 ;
        RECT 676.950 379.650 679.050 379.950 ;
        RECT 681.750 379.650 688.500 380.550 ;
        RECT 689.400 380.550 691.200 381.150 ;
        RECT 697.950 380.550 700.050 380.850 ;
        RECT 689.400 379.950 700.050 380.550 ;
        RECT 710.700 379.950 712.500 381.750 ;
        RECT 676.950 378.450 680.850 379.650 ;
        RECT 689.400 379.350 712.500 379.950 ;
        RECT 697.950 378.750 712.500 379.350 ;
        RECT 713.850 381.000 714.750 382.650 ;
        RECT 715.800 382.950 716.850 384.750 ;
        RECT 720.300 384.000 728.100 385.800 ;
        RECT 715.800 381.900 724.050 382.950 ;
        RECT 713.850 379.200 720.900 381.000 ;
        RECT 676.950 377.850 690.900 378.450 ;
        RECT 721.950 377.850 724.050 381.900 ;
        RECT 677.250 377.550 717.000 377.850 ;
        RECT 688.950 376.650 717.000 377.550 ;
        RECT 726.450 376.650 728.250 377.250 ;
        RECT 676.500 376.050 678.300 376.650 ;
        RECT 685.950 376.050 688.050 376.350 ;
        RECT 676.500 374.850 688.050 376.050 ;
        RECT 685.950 374.250 688.050 374.850 ;
        RECT 688.950 374.400 709.050 375.750 ;
        RECT 673.200 373.350 675.000 374.100 ;
        RECT 688.950 373.350 690.900 374.400 ;
        RECT 706.950 373.650 709.050 374.400 ;
        RECT 712.950 374.550 715.050 375.750 ;
        RECT 715.950 375.450 728.250 376.650 ;
        RECT 729.150 374.550 730.350 389.400 ;
        RECT 712.950 373.650 730.350 374.550 ;
        RECT 732.450 392.400 734.250 395.250 ;
        RECT 735.450 392.400 737.250 395.250 ;
        RECT 732.450 384.150 733.950 392.400 ;
        RECT 741.150 389.400 742.950 395.250 ;
        RECT 744.150 392.400 745.950 395.250 ;
        RECT 748.950 393.300 750.750 395.250 ;
        RECT 747.000 392.400 750.750 393.300 ;
        RECT 753.450 392.400 755.250 395.250 ;
        RECT 756.750 392.400 758.550 395.250 ;
        RECT 760.650 392.400 762.450 395.250 ;
        RECT 764.850 392.400 766.650 395.250 ;
        RECT 769.350 392.400 771.150 395.250 ;
        RECT 747.000 391.500 748.050 392.400 ;
        RECT 745.950 389.400 748.050 391.500 ;
        RECT 756.750 390.600 757.800 392.400 ;
        RECT 732.450 382.050 736.050 384.150 ;
        RECT 673.200 372.300 690.900 373.350 ;
        RECT 668.700 370.500 672.750 371.400 ;
        RECT 662.250 369.600 663.300 370.500 ;
        RECT 671.700 369.600 672.750 370.500 ;
        RECT 658.500 363.750 660.300 369.600 ;
        RECT 661.500 363.750 663.300 369.600 ;
        RECT 664.500 363.750 666.300 369.600 ;
        RECT 668.700 363.750 670.500 369.600 ;
        RECT 671.700 363.750 673.500 369.600 ;
        RECT 674.700 363.750 676.500 369.600 ;
        RECT 677.700 363.750 679.500 372.300 ;
        RECT 697.950 372.150 700.050 372.600 ;
        RECT 697.650 370.500 700.050 372.150 ;
        RECT 702.000 370.800 705.900 372.600 ;
        RECT 702.000 370.500 705.000 370.800 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 369.600 691.050 370.050 ;
        RECT 697.650 369.600 699.000 370.500 ;
        RECT 688.950 367.950 691.500 369.600 ;
        RECT 680.700 363.750 682.500 367.050 ;
        RECT 683.850 366.600 685.050 367.950 ;
        RECT 687.150 366.600 688.050 367.950 ;
        RECT 690.300 366.600 691.500 367.950 ;
        RECT 683.850 363.750 686.250 366.600 ;
        RECT 687.150 363.750 689.250 366.600 ;
        RECT 690.300 363.750 692.250 366.600 ;
        RECT 693.450 363.750 695.250 369.600 ;
        RECT 697.200 363.750 699.000 369.600 ;
        RECT 700.200 363.750 702.000 369.600 ;
        RECT 703.200 363.750 705.000 370.500 ;
        RECT 707.100 366.600 708.450 373.650 ;
        RECT 716.850 372.150 718.650 372.300 ;
        RECT 709.950 370.950 718.650 372.150 ;
        RECT 723.600 371.700 725.400 372.300 ;
        RECT 709.950 370.050 712.050 370.950 ;
        RECT 716.850 370.500 718.650 370.950 ;
        RECT 719.700 370.500 725.400 371.700 ;
        RECT 706.950 363.750 708.750 366.600 ;
        RECT 709.950 363.750 711.750 370.050 ;
        RECT 713.100 367.800 715.200 369.900 ;
        RECT 713.100 366.600 714.600 367.800 ;
        RECT 712.950 363.750 714.750 366.600 ;
        RECT 716.700 363.750 718.500 369.600 ;
        RECT 719.700 363.750 721.500 370.500 ;
        RECT 726.300 369.600 727.500 373.650 ;
        RECT 732.450 369.600 733.950 382.050 ;
        RECT 741.150 376.800 742.050 389.400 ;
        RECT 749.550 388.800 751.350 390.600 ;
        RECT 752.850 389.550 757.800 390.600 ;
        RECT 765.300 391.500 766.350 392.400 ;
        RECT 765.300 390.300 769.050 391.500 ;
        RECT 752.850 388.800 754.650 389.550 ;
        RECT 749.850 387.900 750.900 388.800 ;
        RECT 760.050 388.200 761.850 390.000 ;
        RECT 766.950 389.400 769.050 390.300 ;
        RECT 772.650 389.400 774.450 395.250 ;
        RECT 784.650 389.400 786.450 395.250 ;
        RECT 787.650 389.400 789.450 395.250 ;
        RECT 790.650 389.400 792.450 395.250 ;
        RECT 793.650 389.400 795.450 395.250 ;
        RECT 796.650 389.400 798.450 395.250 ;
        RECT 760.050 387.900 760.950 388.200 ;
        RECT 749.850 387.000 760.950 387.900 ;
        RECT 773.250 387.150 774.450 389.400 ;
        RECT 787.800 388.500 789.600 389.400 ;
        RECT 793.800 388.500 795.600 389.400 ;
        RECT 799.650 388.500 801.450 395.250 ;
        RECT 802.650 389.400 804.450 395.250 ;
        RECT 805.650 389.400 807.450 395.250 ;
        RECT 808.650 389.400 810.450 395.250 ;
        RECT 821.550 389.400 823.350 395.250 ;
        RECT 824.550 389.400 826.350 395.250 ;
        RECT 827.550 389.400 829.350 395.250 ;
        RECT 805.800 388.500 807.600 389.400 ;
        RECT 786.900 388.350 789.600 388.500 ;
        RECT 749.850 385.800 750.900 387.000 ;
        RECT 744.000 384.600 750.900 385.800 ;
        RECT 744.000 383.850 744.900 384.600 ;
        RECT 749.100 384.000 750.900 384.600 ;
        RECT 743.100 382.050 744.900 383.850 ;
        RECT 746.100 382.950 747.900 383.700 ;
        RECT 760.050 382.950 760.950 387.000 ;
        RECT 769.950 385.050 774.450 387.150 ;
        RECT 768.150 383.250 772.050 385.050 ;
        RECT 769.950 382.950 772.050 383.250 ;
        RECT 746.100 381.900 754.050 382.950 ;
        RECT 751.950 380.850 754.050 381.900 ;
        RECT 757.950 380.850 760.950 382.950 ;
        RECT 750.450 377.100 752.250 377.400 ;
        RECT 750.450 376.800 758.850 377.100 ;
        RECT 741.150 376.200 758.850 376.800 ;
        RECT 741.150 375.600 752.250 376.200 ;
        RECT 722.700 363.750 724.500 369.600 ;
        RECT 725.700 363.750 727.500 369.600 ;
        RECT 728.700 363.750 730.500 369.600 ;
        RECT 732.450 363.750 734.250 369.600 ;
        RECT 735.450 363.750 737.250 369.600 ;
        RECT 741.150 363.750 742.950 375.600 ;
        RECT 755.250 374.700 757.050 375.300 ;
        RECT 749.550 373.500 757.050 374.700 ;
        RECT 757.950 374.100 758.850 376.200 ;
        RECT 760.050 376.200 760.950 380.850 ;
        RECT 770.250 377.400 772.050 379.200 ;
        RECT 766.950 376.200 771.150 377.400 ;
        RECT 760.050 375.300 766.050 376.200 ;
        RECT 766.950 375.300 769.050 376.200 ;
        RECT 773.250 375.600 774.450 385.050 ;
        RECT 786.750 387.300 789.600 388.350 ;
        RECT 791.700 387.300 795.600 388.500 ;
        RECT 797.700 387.300 801.450 388.500 ;
        RECT 803.550 387.300 807.600 388.500 ;
        RECT 824.400 388.500 826.200 389.400 ;
        RECT 830.550 388.500 832.350 395.250 ;
        RECT 833.550 389.400 835.350 395.250 ;
        RECT 836.550 389.400 838.350 395.250 ;
        RECT 839.550 389.400 841.350 395.250 ;
        RECT 842.550 389.400 844.350 395.250 ;
        RECT 845.550 389.400 847.350 395.250 ;
        RECT 857.550 389.400 859.350 395.250 ;
        RECT 860.550 389.400 862.350 395.250 ;
        RECT 836.400 388.500 838.200 389.400 ;
        RECT 842.400 388.500 844.200 389.400 ;
        RECT 824.400 387.300 828.450 388.500 ;
        RECT 830.550 387.300 834.300 388.500 ;
        RECT 836.400 387.300 840.300 388.500 ;
        RECT 842.400 388.350 845.100 388.500 ;
        RECT 842.400 387.300 845.250 388.350 ;
        RECT 786.750 384.150 787.800 387.300 ;
        RECT 791.700 386.400 792.900 387.300 ;
        RECT 797.700 386.400 798.900 387.300 ;
        RECT 803.550 386.400 804.750 387.300 ;
        RECT 788.700 384.600 792.900 386.400 ;
        RECT 794.700 384.600 798.900 386.400 ;
        RECT 800.700 384.600 804.750 386.400 ;
        RECT 827.250 386.400 828.450 387.300 ;
        RECT 833.100 386.400 834.300 387.300 ;
        RECT 839.100 386.400 840.300 387.300 ;
        RECT 784.950 382.050 787.800 384.150 ;
        RECT 786.750 377.700 787.800 382.050 ;
        RECT 791.700 377.700 792.900 384.600 ;
        RECT 797.700 377.700 798.900 384.600 ;
        RECT 803.550 377.700 804.750 384.600 ;
        RECT 806.100 384.150 807.900 385.950 ;
        RECT 824.100 384.150 825.900 385.950 ;
        RECT 827.250 384.600 831.300 386.400 ;
        RECT 833.100 384.600 837.300 386.400 ;
        RECT 839.100 384.600 843.300 386.400 ;
        RECT 805.950 382.050 808.050 384.150 ;
        RECT 823.950 382.050 826.050 384.150 ;
        RECT 827.250 377.700 828.450 384.600 ;
        RECT 833.100 377.700 834.300 384.600 ;
        RECT 839.100 377.700 840.300 384.600 ;
        RECT 844.200 384.150 845.250 387.300 ;
        RECT 857.100 384.150 858.900 385.950 ;
        RECT 844.200 382.050 847.050 384.150 ;
        RECT 856.950 382.050 859.050 384.150 ;
        RECT 860.400 382.950 861.600 389.400 ;
        RECT 844.200 377.700 845.250 382.050 ;
        RECT 859.950 380.850 862.050 382.950 ;
        RECT 786.750 376.500 789.450 377.700 ;
        RECT 791.700 376.500 795.450 377.700 ;
        RECT 797.700 376.500 801.450 377.700 ;
        RECT 803.550 376.500 807.450 377.700 ;
        RECT 765.150 374.400 766.050 375.300 ;
        RECT 762.450 374.100 764.250 374.400 ;
        RECT 749.550 372.600 750.750 373.500 ;
        RECT 757.950 373.200 764.250 374.100 ;
        RECT 762.450 372.600 764.250 373.200 ;
        RECT 765.150 372.600 767.850 374.400 ;
        RECT 745.950 370.500 750.750 372.600 ;
        RECT 753.150 370.500 760.050 372.300 ;
        RECT 749.550 369.600 750.750 370.500 ;
        RECT 744.150 363.750 745.950 369.600 ;
        RECT 749.250 363.750 751.050 369.600 ;
        RECT 754.050 363.750 755.850 369.600 ;
        RECT 757.050 363.750 758.850 370.500 ;
        RECT 765.150 369.600 769.050 371.700 ;
        RECT 760.950 363.750 762.750 369.600 ;
        RECT 765.150 363.750 766.950 369.600 ;
        RECT 769.650 363.750 771.450 366.600 ;
        RECT 772.650 363.750 774.450 375.600 ;
        RECT 784.650 363.750 786.450 375.600 ;
        RECT 787.650 363.750 789.450 376.500 ;
        RECT 790.650 363.750 792.450 375.600 ;
        RECT 793.650 363.750 795.450 376.500 ;
        RECT 796.650 363.750 798.450 375.600 ;
        RECT 799.650 363.750 801.450 376.500 ;
        RECT 802.650 363.750 804.450 375.600 ;
        RECT 805.650 363.750 807.450 376.500 ;
        RECT 824.550 376.500 828.450 377.700 ;
        RECT 830.550 376.500 834.300 377.700 ;
        RECT 836.550 376.500 840.300 377.700 ;
        RECT 842.550 376.500 845.250 377.700 ;
        RECT 808.650 363.750 810.450 375.600 ;
        RECT 821.550 363.750 823.350 375.600 ;
        RECT 824.550 363.750 826.350 376.500 ;
        RECT 827.550 363.750 829.350 375.600 ;
        RECT 830.550 363.750 832.350 376.500 ;
        RECT 833.550 363.750 835.350 375.600 ;
        RECT 836.550 363.750 838.350 376.500 ;
        RECT 839.550 363.750 841.350 375.600 ;
        RECT 842.550 363.750 844.350 376.500 ;
        RECT 860.400 375.600 861.600 380.850 ;
        RECT 845.550 363.750 847.350 375.600 ;
        RECT 857.550 363.750 859.350 375.600 ;
        RECT 860.550 363.750 862.350 375.600 ;
        RECT 10.350 347.400 12.150 359.250 ;
        RECT 13.350 347.400 15.150 359.250 ;
        RECT 16.650 353.400 18.450 359.250 ;
        RECT 28.650 353.400 30.450 359.250 ;
        RECT 31.650 354.000 33.450 359.250 ;
        RECT 10.650 342.150 11.850 347.400 ;
        RECT 17.250 346.500 18.450 353.400 ;
        RECT 12.750 345.600 18.450 346.500 ;
        RECT 29.250 353.100 30.450 353.400 ;
        RECT 34.650 353.400 36.450 359.250 ;
        RECT 37.650 353.400 39.450 359.250 ;
        RECT 47.550 353.400 49.350 359.250 ;
        RECT 50.550 353.400 52.350 359.250 ;
        RECT 53.550 353.400 55.350 359.250 ;
        RECT 34.650 353.100 36.300 353.400 ;
        RECT 29.250 352.200 36.300 353.100 ;
        RECT 12.750 344.700 15.000 345.600 ;
        RECT 10.650 340.050 13.050 342.150 ;
        RECT 10.650 333.600 11.850 340.050 ;
        RECT 13.950 336.300 15.000 344.700 ;
        RECT 29.250 343.950 30.300 352.200 ;
        RECT 35.100 348.150 36.900 349.950 ;
        RECT 31.950 345.150 33.750 346.950 ;
        RECT 34.950 346.050 37.050 348.150 ;
        RECT 38.100 345.150 39.900 346.950 ;
        RECT 50.550 345.150 51.750 353.400 ;
        RECT 66.300 347.400 68.100 359.250 ;
        RECT 70.500 347.400 72.300 359.250 ;
        RECT 73.800 353.400 75.600 359.250 ;
        RECT 89.400 353.400 91.200 359.250 ;
        RECT 92.700 347.400 94.500 359.250 ;
        RECT 96.900 347.400 98.700 359.250 ;
        RECT 112.650 353.400 114.450 359.250 ;
        RECT 115.650 354.000 117.450 359.250 ;
        RECT 113.250 353.100 114.450 353.400 ;
        RECT 118.650 353.400 120.450 359.250 ;
        RECT 121.650 353.400 123.450 359.250 ;
        RECT 133.650 353.400 135.450 359.250 ;
        RECT 136.650 353.400 138.450 359.250 ;
        RECT 139.650 353.400 141.450 359.250 ;
        RECT 118.650 353.100 120.300 353.400 ;
        RECT 113.250 352.200 120.300 353.100 ;
        RECT 17.100 342.150 18.900 343.950 ;
        RECT 16.950 340.050 19.050 342.150 ;
        RECT 28.950 341.850 31.050 343.950 ;
        RECT 31.950 343.050 34.050 345.150 ;
        RECT 37.950 343.050 40.050 345.150 ;
        RECT 46.950 341.850 49.050 343.950 ;
        RECT 49.950 343.050 52.050 345.150 ;
        RECT 12.750 335.400 15.000 336.300 ;
        RECT 29.400 337.650 30.600 341.850 ;
        RECT 47.100 340.050 48.900 341.850 ;
        RECT 29.400 336.000 33.900 337.650 ;
        RECT 12.750 334.500 17.850 335.400 ;
        RECT 10.350 327.750 12.150 333.600 ;
        RECT 13.350 327.750 15.150 333.600 ;
        RECT 16.650 330.600 17.850 334.500 ;
        RECT 16.650 327.750 18.450 330.600 ;
        RECT 32.100 327.750 33.900 336.000 ;
        RECT 37.500 327.750 39.300 336.600 ;
        RECT 50.550 335.700 51.750 343.050 ;
        RECT 52.950 341.850 55.050 343.950 ;
        RECT 65.100 342.150 66.900 343.950 ;
        RECT 70.950 342.150 72.150 347.400 ;
        RECT 73.950 345.150 75.750 346.950 ;
        RECT 89.250 345.150 91.050 346.950 ;
        RECT 73.950 343.050 76.050 345.150 ;
        RECT 88.950 343.050 91.050 345.150 ;
        RECT 92.850 342.150 94.050 347.400 ;
        RECT 113.250 343.950 114.300 352.200 ;
        RECT 119.100 348.150 120.900 349.950 ;
        RECT 115.950 345.150 117.750 346.950 ;
        RECT 118.950 346.050 121.050 348.150 ;
        RECT 122.100 345.150 123.900 346.950 ;
        RECT 137.250 345.150 138.450 353.400 ;
        RECT 153.150 348.900 154.950 359.250 ;
        RECT 152.550 347.550 154.950 348.900 ;
        RECT 156.150 347.550 157.950 359.250 ;
        RECT 98.100 342.150 99.900 343.950 ;
        RECT 53.100 340.050 54.900 341.850 ;
        RECT 64.950 340.050 67.050 342.150 ;
        RECT 67.950 338.850 70.050 340.950 ;
        RECT 70.950 340.050 73.050 342.150 ;
        RECT 68.100 337.050 69.900 338.850 ;
        RECT 71.850 336.750 73.050 340.050 ;
        RECT 91.950 340.050 94.050 342.150 ;
        RECT 91.950 336.750 93.150 340.050 ;
        RECT 94.950 338.850 97.050 340.950 ;
        RECT 97.950 340.050 100.050 342.150 ;
        RECT 112.950 341.850 115.050 343.950 ;
        RECT 115.950 343.050 118.050 345.150 ;
        RECT 121.950 343.050 124.050 345.150 ;
        RECT 133.950 341.850 136.050 343.950 ;
        RECT 136.950 343.050 139.050 345.150 ;
        RECT 95.100 337.050 96.900 338.850 ;
        RECT 113.400 337.650 114.600 341.850 ;
        RECT 134.100 340.050 135.900 341.850 ;
        RECT 72.000 335.700 75.750 336.750 ;
        RECT 50.550 334.800 54.150 335.700 ;
        RECT 47.850 327.750 49.650 333.600 ;
        RECT 52.350 327.750 54.150 334.800 ;
        RECT 65.550 332.700 73.350 334.050 ;
        RECT 65.550 327.750 67.350 332.700 ;
        RECT 68.550 327.750 70.350 331.800 ;
        RECT 71.550 327.750 73.350 332.700 ;
        RECT 74.550 333.600 75.750 335.700 ;
        RECT 89.250 335.700 93.000 336.750 ;
        RECT 113.400 336.000 117.900 337.650 ;
        RECT 89.250 333.600 90.450 335.700 ;
        RECT 74.550 327.750 76.350 333.600 ;
        RECT 88.650 327.750 90.450 333.600 ;
        RECT 91.650 332.700 99.450 334.050 ;
        RECT 91.650 327.750 93.450 332.700 ;
        RECT 94.650 327.750 96.450 331.800 ;
        RECT 97.650 327.750 99.450 332.700 ;
        RECT 116.100 327.750 117.900 336.000 ;
        RECT 121.500 327.750 123.300 336.600 ;
        RECT 137.250 335.700 138.450 343.050 ;
        RECT 139.950 341.850 142.050 343.950 ;
        RECT 140.100 340.050 141.900 341.850 ;
        RECT 152.550 340.950 153.900 347.550 ;
        RECT 160.650 347.400 162.450 359.250 ;
        RECT 170.550 347.400 172.350 359.250 ;
        RECT 173.550 347.400 175.350 359.250 ;
        RECT 187.650 353.400 189.450 359.250 ;
        RECT 190.650 354.000 192.450 359.250 ;
        RECT 188.250 353.100 189.450 353.400 ;
        RECT 193.650 353.400 195.450 359.250 ;
        RECT 196.650 353.400 198.450 359.250 ;
        RECT 193.650 353.100 195.300 353.400 ;
        RECT 188.250 352.200 195.300 353.100 ;
        RECT 155.250 346.200 157.050 346.650 ;
        RECT 161.250 346.200 162.450 347.400 ;
        RECT 155.250 345.000 162.450 346.200 ;
        RECT 155.250 344.850 157.050 345.000 ;
        RECT 134.850 334.800 138.450 335.700 ;
        RECT 151.950 338.850 154.050 340.950 ;
        RECT 134.850 327.750 136.650 334.800 ;
        RECT 151.950 333.600 153.000 338.850 ;
        RECT 155.400 336.600 156.300 344.850 ;
        RECT 158.100 342.150 159.900 343.950 ;
        RECT 173.400 342.150 174.600 347.400 ;
        RECT 188.250 343.950 189.300 352.200 ;
        RECT 194.100 348.150 195.900 349.950 ;
        RECT 190.950 345.150 192.750 346.950 ;
        RECT 193.950 346.050 196.050 348.150 ;
        RECT 208.650 347.400 210.450 359.250 ;
        RECT 211.650 348.300 213.450 359.250 ;
        RECT 214.650 349.200 216.450 359.250 ;
        RECT 217.650 348.300 219.450 359.250 ;
        RECT 233.400 353.400 235.200 359.250 ;
        RECT 211.650 347.400 219.450 348.300 ;
        RECT 236.700 347.400 238.500 359.250 ;
        RECT 240.900 347.400 242.700 359.250 ;
        RECT 253.650 347.400 255.450 359.250 ;
        RECT 256.650 348.300 258.450 359.250 ;
        RECT 259.650 349.200 261.450 359.250 ;
        RECT 262.650 348.300 264.450 359.250 ;
        RECT 274.650 353.400 276.450 359.250 ;
        RECT 277.650 354.000 279.450 359.250 ;
        RECT 256.650 347.400 264.450 348.300 ;
        RECT 275.250 353.100 276.450 353.400 ;
        RECT 280.650 353.400 282.450 359.250 ;
        RECT 283.650 353.400 285.450 359.250 ;
        RECT 295.650 353.400 297.450 359.250 ;
        RECT 298.650 354.000 300.450 359.250 ;
        RECT 280.650 353.100 282.300 353.400 ;
        RECT 275.250 352.200 282.300 353.100 ;
        RECT 296.250 353.100 297.450 353.400 ;
        RECT 301.650 353.400 303.450 359.250 ;
        RECT 304.650 353.400 306.450 359.250 ;
        RECT 309.750 353.400 311.550 359.250 ;
        RECT 312.750 353.400 314.550 359.250 ;
        RECT 316.500 353.400 318.300 359.250 ;
        RECT 319.500 353.400 321.300 359.250 ;
        RECT 322.500 353.400 324.300 359.250 ;
        RECT 301.650 353.100 303.300 353.400 ;
        RECT 296.250 352.200 303.300 353.100 ;
        RECT 197.100 345.150 198.900 346.950 ;
        RECT 157.950 340.050 160.050 342.150 ;
        RECT 161.100 339.150 162.900 340.950 ;
        RECT 160.950 337.050 163.050 339.150 ;
        RECT 169.950 338.850 172.050 340.950 ;
        RECT 172.950 340.050 175.050 342.150 ;
        RECT 187.950 341.850 190.050 343.950 ;
        RECT 190.950 343.050 193.050 345.150 ;
        RECT 196.950 343.050 199.050 345.150 ;
        RECT 209.100 342.150 210.300 347.400 ;
        RECT 233.250 345.150 235.050 346.950 ;
        RECT 232.950 343.050 235.050 345.150 ;
        RECT 236.850 342.150 238.050 347.400 ;
        RECT 242.100 342.150 243.900 343.950 ;
        RECT 254.100 342.150 255.300 347.400 ;
        RECT 275.250 343.950 276.300 352.200 ;
        RECT 281.100 348.150 282.900 349.950 ;
        RECT 277.950 345.150 279.750 346.950 ;
        RECT 280.950 346.050 283.050 348.150 ;
        RECT 284.100 345.150 285.900 346.950 ;
        RECT 170.100 337.050 171.900 338.850 ;
        RECT 155.250 335.700 157.050 336.600 ;
        RECT 155.250 334.800 158.550 335.700 ;
        RECT 139.350 327.750 141.150 333.600 ;
        RECT 151.650 327.750 153.450 333.600 ;
        RECT 157.650 330.600 158.550 334.800 ;
        RECT 173.400 333.600 174.600 340.050 ;
        RECT 188.400 337.650 189.600 341.850 ;
        RECT 208.950 340.050 211.050 342.150 ;
        RECT 188.400 336.000 192.900 337.650 ;
        RECT 154.650 327.750 156.450 330.600 ;
        RECT 157.650 327.750 159.450 330.600 ;
        RECT 160.650 327.750 162.450 330.600 ;
        RECT 170.550 327.750 172.350 333.600 ;
        RECT 173.550 327.750 175.350 333.600 ;
        RECT 191.100 327.750 192.900 336.000 ;
        RECT 196.500 327.750 198.300 336.600 ;
        RECT 209.100 333.600 210.300 340.050 ;
        RECT 211.950 338.850 214.050 340.950 ;
        RECT 215.100 339.150 216.900 340.950 ;
        RECT 212.100 337.050 213.900 338.850 ;
        RECT 214.950 337.050 217.050 339.150 ;
        RECT 217.950 338.850 220.050 340.950 ;
        RECT 235.950 340.050 238.050 342.150 ;
        RECT 218.100 337.050 219.900 338.850 ;
        RECT 235.950 336.750 237.150 340.050 ;
        RECT 238.950 338.850 241.050 340.950 ;
        RECT 241.950 340.050 244.050 342.150 ;
        RECT 253.950 340.050 256.050 342.150 ;
        RECT 274.950 341.850 277.050 343.950 ;
        RECT 277.950 343.050 280.050 345.150 ;
        RECT 283.950 343.050 286.050 345.150 ;
        RECT 296.250 343.950 297.300 352.200 ;
        RECT 302.100 348.150 303.900 349.950 ;
        RECT 298.950 345.150 300.750 346.950 ;
        RECT 301.950 346.050 304.050 348.150 ;
        RECT 305.100 345.150 306.900 346.950 ;
        RECT 295.950 341.850 298.050 343.950 ;
        RECT 298.950 343.050 301.050 345.150 ;
        RECT 304.950 343.050 307.050 345.150 ;
        RECT 239.100 337.050 240.900 338.850 ;
        RECT 233.250 335.700 237.000 336.750 ;
        RECT 233.250 333.600 234.450 335.700 ;
        RECT 209.100 331.950 214.800 333.600 ;
        RECT 209.700 327.750 211.500 330.600 ;
        RECT 213.000 327.750 214.800 331.950 ;
        RECT 217.200 327.750 219.000 333.600 ;
        RECT 232.650 327.750 234.450 333.600 ;
        RECT 235.650 332.700 243.450 334.050 ;
        RECT 235.650 327.750 237.450 332.700 ;
        RECT 238.650 327.750 240.450 331.800 ;
        RECT 241.650 327.750 243.450 332.700 ;
        RECT 254.100 333.600 255.300 340.050 ;
        RECT 256.950 338.850 259.050 340.950 ;
        RECT 260.100 339.150 261.900 340.950 ;
        RECT 257.100 337.050 258.900 338.850 ;
        RECT 259.950 337.050 262.050 339.150 ;
        RECT 262.950 338.850 265.050 340.950 ;
        RECT 263.100 337.050 264.900 338.850 ;
        RECT 275.400 337.650 276.600 341.850 ;
        RECT 296.400 337.650 297.600 341.850 ;
        RECT 313.050 340.950 314.550 353.400 ;
        RECT 319.500 349.350 320.700 353.400 ;
        RECT 325.500 352.500 327.300 359.250 ;
        RECT 328.500 353.400 330.300 359.250 ;
        RECT 332.250 356.400 334.050 359.250 ;
        RECT 332.400 355.200 333.900 356.400 ;
        RECT 331.800 353.100 333.900 355.200 ;
        RECT 335.250 352.950 337.050 359.250 ;
        RECT 338.250 356.400 340.050 359.250 ;
        RECT 321.600 351.300 327.300 352.500 ;
        RECT 328.350 352.050 330.150 352.500 ;
        RECT 334.950 352.050 337.050 352.950 ;
        RECT 321.600 350.700 323.400 351.300 ;
        RECT 328.350 350.850 337.050 352.050 ;
        RECT 328.350 350.700 330.150 350.850 ;
        RECT 338.550 349.350 339.900 356.400 ;
        RECT 342.000 352.500 343.800 359.250 ;
        RECT 345.000 353.400 346.800 359.250 ;
        RECT 348.000 353.400 349.800 359.250 ;
        RECT 351.750 353.400 353.550 359.250 ;
        RECT 354.750 356.400 356.700 359.250 ;
        RECT 357.750 356.400 359.850 359.250 ;
        RECT 360.750 356.400 363.150 359.250 ;
        RECT 355.500 355.050 356.700 356.400 ;
        RECT 358.950 355.050 359.850 356.400 ;
        RECT 361.950 355.050 363.150 356.400 ;
        RECT 364.500 355.950 366.300 359.250 ;
        RECT 355.500 353.400 358.050 355.050 ;
        RECT 348.000 352.500 349.350 353.400 ;
        RECT 355.950 352.950 358.050 353.400 ;
        RECT 358.950 352.950 361.050 355.050 ;
        RECT 361.950 352.950 364.050 355.050 ;
        RECT 342.000 352.200 345.000 352.500 ;
        RECT 341.100 350.400 345.000 352.200 ;
        RECT 346.950 350.850 349.350 352.500 ;
        RECT 346.950 350.400 349.050 350.850 ;
        RECT 367.500 350.700 369.300 359.250 ;
        RECT 370.500 353.400 372.300 359.250 ;
        RECT 373.500 353.400 375.300 359.250 ;
        RECT 376.500 353.400 378.300 359.250 ;
        RECT 374.250 352.500 375.300 353.400 ;
        RECT 374.250 351.600 378.300 352.500 ;
        RECT 356.100 349.650 373.800 350.700 ;
        RECT 310.950 338.850 314.550 340.950 ;
        RECT 275.400 336.000 279.900 337.650 ;
        RECT 254.100 331.950 259.800 333.600 ;
        RECT 254.700 327.750 256.500 330.600 ;
        RECT 258.000 327.750 259.800 331.950 ;
        RECT 262.200 327.750 264.000 333.600 ;
        RECT 278.100 327.750 279.900 336.000 ;
        RECT 283.500 327.750 285.300 336.600 ;
        RECT 296.400 336.000 300.900 337.650 ;
        RECT 299.100 327.750 300.900 336.000 ;
        RECT 304.500 327.750 306.300 336.600 ;
        RECT 313.050 330.600 314.550 338.850 ;
        RECT 309.750 327.750 311.550 330.600 ;
        RECT 312.750 327.750 314.550 330.600 ;
        RECT 316.650 348.450 334.050 349.350 ;
        RECT 316.650 333.600 317.850 348.450 ;
        RECT 318.750 346.350 331.050 347.550 ;
        RECT 331.950 347.250 334.050 348.450 ;
        RECT 337.950 348.600 340.050 349.350 ;
        RECT 356.100 348.600 358.050 349.650 ;
        RECT 372.000 348.900 373.800 349.650 ;
        RECT 337.950 347.250 358.050 348.600 ;
        RECT 358.950 348.150 361.050 348.750 ;
        RECT 358.950 346.950 370.500 348.150 ;
        RECT 358.950 346.650 361.050 346.950 ;
        RECT 368.700 346.350 370.500 346.950 ;
        RECT 318.750 345.750 320.550 346.350 ;
        RECT 330.000 345.450 358.050 346.350 ;
        RECT 330.000 345.150 369.750 345.450 ;
        RECT 322.950 341.100 325.050 345.150 ;
        RECT 356.100 344.550 370.050 345.150 ;
        RECT 326.100 342.000 333.150 343.800 ;
        RECT 322.950 340.050 331.200 341.100 ;
        RECT 318.900 337.200 326.700 339.000 ;
        RECT 330.150 338.250 331.200 340.050 ;
        RECT 332.250 340.350 333.150 342.000 ;
        RECT 334.500 343.650 349.050 344.250 ;
        RECT 334.500 343.050 357.600 343.650 ;
        RECT 366.150 343.350 370.050 344.550 ;
        RECT 334.500 341.250 336.300 343.050 ;
        RECT 346.950 342.450 357.600 343.050 ;
        RECT 346.950 342.150 349.050 342.450 ;
        RECT 355.800 341.850 357.600 342.450 ;
        RECT 358.500 342.450 365.250 343.350 ;
        RECT 367.950 343.050 370.050 343.350 ;
        RECT 342.750 341.250 344.850 341.550 ;
        RECT 332.250 339.300 341.850 340.350 ;
        RECT 342.750 339.450 346.650 341.250 ;
        RECT 358.500 340.950 359.550 342.450 ;
        RECT 347.550 340.050 359.550 340.950 ;
        RECT 340.950 338.550 341.850 339.300 ;
        RECT 347.550 338.550 348.600 340.050 ;
        RECT 360.450 339.750 362.250 341.550 ;
        RECT 364.050 340.050 365.250 342.450 ;
        RECT 373.950 341.850 376.050 343.950 ;
        RECT 374.100 340.050 375.900 341.850 ;
        RECT 330.150 337.200 340.050 338.250 ;
        RECT 340.950 337.200 348.600 338.550 ;
        RECT 349.950 337.350 353.850 339.150 ;
        RECT 325.200 333.600 326.700 337.200 ;
        RECT 339.000 336.300 340.050 337.200 ;
        RECT 349.950 337.050 352.050 337.350 ;
        RECT 357.150 336.300 358.950 336.750 ;
        RECT 360.450 336.300 361.500 339.750 ;
        RECT 364.050 339.000 375.900 340.050 ;
        RECT 377.100 338.100 378.300 351.600 ;
        RECT 388.350 347.400 390.150 359.250 ;
        RECT 391.350 347.400 393.150 359.250 ;
        RECT 394.650 353.400 396.450 359.250 ;
        RECT 331.350 334.500 338.100 336.300 ;
        RECT 339.000 334.500 345.900 336.300 ;
        RECT 357.150 335.850 361.500 336.300 ;
        RECT 353.850 335.100 361.500 335.850 ;
        RECT 363.000 337.200 378.300 338.100 ;
        RECT 353.850 334.950 358.950 335.100 ;
        RECT 353.850 333.600 354.750 334.950 ;
        RECT 363.000 334.050 364.050 337.200 ;
        RECT 372.300 335.700 374.100 336.300 ;
        RECT 316.650 327.750 318.450 333.600 ;
        RECT 322.050 327.750 323.850 333.600 ;
        RECT 325.200 332.400 329.400 333.600 ;
        RECT 327.600 327.750 329.400 332.400 ;
        RECT 331.950 331.500 334.050 333.600 ;
        RECT 334.950 331.500 337.050 333.600 ;
        RECT 337.950 331.500 340.050 333.600 ;
        RECT 342.750 333.300 344.850 333.600 ;
        RECT 332.250 327.750 334.050 331.500 ;
        RECT 335.250 327.750 337.050 331.500 ;
        RECT 338.250 327.750 340.050 331.500 ;
        RECT 342.000 331.500 344.850 333.300 ;
        RECT 346.950 333.300 349.050 333.600 ;
        RECT 346.950 331.500 349.800 333.300 ;
        RECT 350.700 332.250 354.750 333.600 ;
        RECT 350.700 331.800 352.500 332.250 ;
        RECT 355.950 331.950 358.050 334.050 ;
        RECT 358.950 331.950 361.050 334.050 ;
        RECT 361.950 331.950 364.050 334.050 ;
        RECT 365.700 334.500 374.100 335.700 ;
        RECT 365.700 333.600 367.200 334.500 ;
        RECT 377.100 333.600 378.300 337.200 ;
        RECT 388.650 342.150 389.850 347.400 ;
        RECT 395.250 346.500 396.450 353.400 ;
        RECT 408.300 347.400 410.100 359.250 ;
        RECT 412.500 347.400 414.300 359.250 ;
        RECT 415.800 353.400 417.600 359.250 ;
        RECT 429.300 347.400 431.100 359.250 ;
        RECT 433.500 347.400 435.300 359.250 ;
        RECT 436.800 353.400 438.600 359.250 ;
        RECT 451.650 353.400 453.450 359.250 ;
        RECT 454.650 353.400 456.450 359.250 ;
        RECT 457.650 353.400 459.450 359.250 ;
        RECT 470.550 353.400 472.350 359.250 ;
        RECT 473.550 353.400 475.350 359.250 ;
        RECT 476.550 353.400 478.350 359.250 ;
        RECT 390.750 345.600 396.450 346.500 ;
        RECT 390.750 344.700 393.000 345.600 ;
        RECT 388.650 340.050 391.050 342.150 ;
        RECT 388.650 333.600 389.850 340.050 ;
        RECT 391.950 336.300 393.000 344.700 ;
        RECT 395.100 342.150 396.900 343.950 ;
        RECT 407.100 342.150 408.900 343.950 ;
        RECT 412.950 342.150 414.150 347.400 ;
        RECT 415.950 345.150 417.750 346.950 ;
        RECT 415.950 343.050 418.050 345.150 ;
        RECT 428.100 342.150 429.900 343.950 ;
        RECT 433.950 342.150 435.150 347.400 ;
        RECT 436.950 345.150 438.750 346.950 ;
        RECT 455.250 345.150 456.450 353.400 ;
        RECT 473.550 345.150 474.750 353.400 ;
        RECT 490.650 347.400 492.450 359.250 ;
        RECT 493.650 348.300 495.450 359.250 ;
        RECT 496.650 349.200 498.450 359.250 ;
        RECT 499.650 348.300 501.450 359.250 ;
        RECT 493.650 347.400 501.450 348.300 ;
        RECT 436.950 343.050 439.050 345.150 ;
        RECT 394.950 340.050 397.050 342.150 ;
        RECT 406.950 340.050 409.050 342.150 ;
        RECT 409.950 338.850 412.050 340.950 ;
        RECT 412.950 340.050 415.050 342.150 ;
        RECT 427.950 340.050 430.050 342.150 ;
        RECT 410.100 337.050 411.900 338.850 ;
        RECT 413.850 336.750 415.050 340.050 ;
        RECT 430.950 338.850 433.050 340.950 ;
        RECT 433.950 340.050 436.050 342.150 ;
        RECT 451.950 341.850 454.050 343.950 ;
        RECT 454.950 343.050 457.050 345.150 ;
        RECT 452.100 340.050 453.900 341.850 ;
        RECT 431.100 337.050 432.900 338.850 ;
        RECT 434.850 336.750 436.050 340.050 ;
        RECT 390.750 335.400 393.000 336.300 ;
        RECT 414.000 335.700 417.750 336.750 ;
        RECT 435.000 335.700 438.750 336.750 ;
        RECT 455.250 335.700 456.450 343.050 ;
        RECT 457.950 341.850 460.050 343.950 ;
        RECT 469.950 341.850 472.050 343.950 ;
        RECT 472.950 343.050 475.050 345.150 ;
        RECT 487.950 343.950 490.050 346.050 ;
        RECT 458.100 340.050 459.900 341.850 ;
        RECT 470.100 340.050 471.900 341.850 ;
        RECT 390.750 334.500 395.850 335.400 ;
        RECT 342.000 327.750 343.800 331.500 ;
        RECT 345.000 327.750 346.800 330.600 ;
        RECT 348.000 327.750 349.800 331.500 ;
        RECT 355.950 330.600 357.300 331.950 ;
        RECT 358.950 330.600 360.300 331.950 ;
        RECT 361.950 330.600 363.300 331.950 ;
        RECT 352.500 327.750 354.300 330.600 ;
        RECT 355.500 327.750 357.300 330.600 ;
        RECT 358.500 327.750 360.300 330.600 ;
        RECT 361.500 327.750 363.300 330.600 ;
        RECT 365.700 327.750 367.500 333.600 ;
        RECT 371.100 327.750 372.900 333.600 ;
        RECT 376.500 327.750 378.300 333.600 ;
        RECT 388.350 327.750 390.150 333.600 ;
        RECT 391.350 327.750 393.150 333.600 ;
        RECT 394.650 330.600 395.850 334.500 ;
        RECT 407.550 332.700 415.350 334.050 ;
        RECT 394.650 327.750 396.450 330.600 ;
        RECT 407.550 327.750 409.350 332.700 ;
        RECT 410.550 327.750 412.350 331.800 ;
        RECT 413.550 327.750 415.350 332.700 ;
        RECT 416.550 333.600 417.750 335.700 ;
        RECT 416.550 327.750 418.350 333.600 ;
        RECT 428.550 332.700 436.350 334.050 ;
        RECT 428.550 327.750 430.350 332.700 ;
        RECT 431.550 327.750 433.350 331.800 ;
        RECT 434.550 327.750 436.350 332.700 ;
        RECT 437.550 333.600 438.750 335.700 ;
        RECT 452.850 334.800 456.450 335.700 ;
        RECT 473.550 335.700 474.750 343.050 ;
        RECT 475.950 341.850 478.050 343.950 ;
        RECT 476.100 340.050 477.900 341.850 ;
        RECT 481.950 336.450 484.050 337.050 ;
        RECT 488.550 336.450 489.450 343.950 ;
        RECT 491.100 342.150 492.300 347.400 ;
        RECT 505.950 346.950 508.050 349.050 ;
        RECT 509.550 347.400 511.350 359.250 ;
        RECT 513.750 347.400 515.550 359.250 ;
        RECT 517.950 357.450 520.050 358.050 ;
        RECT 526.950 357.450 529.050 358.050 ;
        RECT 517.950 356.550 529.050 357.450 ;
        RECT 517.950 355.950 520.050 356.550 ;
        RECT 526.950 355.950 529.050 356.550 ;
        RECT 531.300 347.400 533.100 359.250 ;
        RECT 535.500 347.400 537.300 359.250 ;
        RECT 538.800 353.400 540.600 359.250 ;
        RECT 551.550 353.400 553.350 359.250 ;
        RECT 554.550 353.400 556.350 359.250 ;
        RECT 557.550 353.400 559.350 359.250 ;
        RECT 569.550 353.400 571.350 359.250 ;
        RECT 493.950 345.450 496.050 346.050 ;
        RECT 506.550 345.450 507.450 346.950 ;
        RECT 493.950 344.550 507.450 345.450 ;
        RECT 513.000 346.350 515.550 347.400 ;
        RECT 493.950 343.950 496.050 344.550 ;
        RECT 509.100 342.150 510.900 343.950 ;
        RECT 490.950 340.050 493.050 342.150 ;
        RECT 473.550 334.800 477.150 335.700 ;
        RECT 481.950 335.550 489.450 336.450 ;
        RECT 481.950 334.950 484.050 335.550 ;
        RECT 437.550 327.750 439.350 333.600 ;
        RECT 452.850 327.750 454.650 334.800 ;
        RECT 457.350 327.750 459.150 333.600 ;
        RECT 470.850 327.750 472.650 333.600 ;
        RECT 475.350 327.750 477.150 334.800 ;
        RECT 491.100 333.600 492.300 340.050 ;
        RECT 493.950 338.850 496.050 340.950 ;
        RECT 497.100 339.150 498.900 340.950 ;
        RECT 494.100 337.050 495.900 338.850 ;
        RECT 496.950 337.050 499.050 339.150 ;
        RECT 499.950 338.850 502.050 340.950 ;
        RECT 508.950 340.050 511.050 342.150 ;
        RECT 513.000 339.150 514.050 346.350 ;
        RECT 515.100 342.150 516.900 343.950 ;
        RECT 530.100 342.150 531.900 343.950 ;
        RECT 535.950 342.150 537.150 347.400 ;
        RECT 538.950 345.150 540.750 346.950 ;
        RECT 554.550 345.150 555.750 353.400 ;
        RECT 569.550 346.500 570.750 353.400 ;
        RECT 572.850 347.400 574.650 359.250 ;
        RECT 575.850 347.400 577.650 359.250 ;
        RECT 582.750 353.400 584.550 359.250 ;
        RECT 585.750 353.400 587.550 359.250 ;
        RECT 589.500 353.400 591.300 359.250 ;
        RECT 592.500 353.400 594.300 359.250 ;
        RECT 595.500 353.400 597.300 359.250 ;
        RECT 569.550 345.600 575.250 346.500 ;
        RECT 538.950 343.050 541.050 345.150 ;
        RECT 514.950 340.050 517.050 342.150 ;
        RECT 529.950 340.050 532.050 342.150 ;
        RECT 500.100 337.050 501.900 338.850 ;
        RECT 511.950 337.050 514.050 339.150 ;
        RECT 532.950 338.850 535.050 340.950 ;
        RECT 535.950 340.050 538.050 342.150 ;
        RECT 550.950 341.850 553.050 343.950 ;
        RECT 553.950 343.050 556.050 345.150 ;
        RECT 573.000 344.700 575.250 345.600 ;
        RECT 551.100 340.050 552.900 341.850 ;
        RECT 533.100 337.050 534.900 338.850 ;
        RECT 491.100 331.950 496.800 333.600 ;
        RECT 491.700 327.750 493.500 330.600 ;
        RECT 495.000 327.750 496.800 331.950 ;
        RECT 499.200 327.750 501.000 333.600 ;
        RECT 513.000 330.600 514.050 337.050 ;
        RECT 536.850 336.750 538.050 340.050 ;
        RECT 537.000 335.700 540.750 336.750 ;
        RECT 530.550 332.700 538.350 334.050 ;
        RECT 509.550 327.750 511.350 330.600 ;
        RECT 512.550 327.750 514.350 330.600 ;
        RECT 515.550 327.750 517.350 330.600 ;
        RECT 530.550 327.750 532.350 332.700 ;
        RECT 533.550 327.750 535.350 331.800 ;
        RECT 536.550 327.750 538.350 332.700 ;
        RECT 539.550 333.600 540.750 335.700 ;
        RECT 554.550 335.700 555.750 343.050 ;
        RECT 556.950 341.850 559.050 343.950 ;
        RECT 569.100 342.150 570.900 343.950 ;
        RECT 557.100 340.050 558.900 341.850 ;
        RECT 568.950 340.050 571.050 342.150 ;
        RECT 573.000 336.300 574.050 344.700 ;
        RECT 576.150 342.150 577.350 347.400 ;
        RECT 574.950 340.050 577.350 342.150 ;
        RECT 586.050 340.950 587.550 353.400 ;
        RECT 592.500 349.350 593.700 353.400 ;
        RECT 598.500 352.500 600.300 359.250 ;
        RECT 601.500 353.400 603.300 359.250 ;
        RECT 605.250 356.400 607.050 359.250 ;
        RECT 605.400 355.200 606.900 356.400 ;
        RECT 604.800 353.100 606.900 355.200 ;
        RECT 608.250 352.950 610.050 359.250 ;
        RECT 611.250 356.400 613.050 359.250 ;
        RECT 594.600 351.300 600.300 352.500 ;
        RECT 601.350 352.050 603.150 352.500 ;
        RECT 607.950 352.050 610.050 352.950 ;
        RECT 594.600 350.700 596.400 351.300 ;
        RECT 601.350 350.850 610.050 352.050 ;
        RECT 601.350 350.700 603.150 350.850 ;
        RECT 611.550 349.350 612.900 356.400 ;
        RECT 615.000 352.500 616.800 359.250 ;
        RECT 618.000 353.400 619.800 359.250 ;
        RECT 621.000 353.400 622.800 359.250 ;
        RECT 624.750 353.400 626.550 359.250 ;
        RECT 627.750 356.400 629.700 359.250 ;
        RECT 630.750 356.400 632.850 359.250 ;
        RECT 633.750 356.400 636.150 359.250 ;
        RECT 628.500 355.050 629.700 356.400 ;
        RECT 631.950 355.050 632.850 356.400 ;
        RECT 634.950 355.050 636.150 356.400 ;
        RECT 637.500 355.950 639.300 359.250 ;
        RECT 628.500 353.400 631.050 355.050 ;
        RECT 621.000 352.500 622.350 353.400 ;
        RECT 628.950 352.950 631.050 353.400 ;
        RECT 631.950 352.950 634.050 355.050 ;
        RECT 634.950 352.950 637.050 355.050 ;
        RECT 615.000 352.200 618.000 352.500 ;
        RECT 614.100 350.400 618.000 352.200 ;
        RECT 619.950 350.850 622.350 352.500 ;
        RECT 619.950 350.400 622.050 350.850 ;
        RECT 640.500 350.700 642.300 359.250 ;
        RECT 643.500 353.400 645.300 359.250 ;
        RECT 646.500 353.400 648.300 359.250 ;
        RECT 649.500 353.400 651.300 359.250 ;
        RECT 659.550 353.400 661.350 359.250 ;
        RECT 662.550 353.400 664.350 359.250 ;
        RECT 647.250 352.500 648.300 353.400 ;
        RECT 647.250 351.600 651.300 352.500 ;
        RECT 629.100 349.650 646.800 350.700 ;
        RECT 554.550 334.800 558.150 335.700 ;
        RECT 573.000 335.400 575.250 336.300 ;
        RECT 539.550 327.750 541.350 333.600 ;
        RECT 551.850 327.750 553.650 333.600 ;
        RECT 556.350 327.750 558.150 334.800 ;
        RECT 570.150 334.500 575.250 335.400 ;
        RECT 570.150 330.600 571.350 334.500 ;
        RECT 576.150 333.600 577.350 340.050 ;
        RECT 583.950 338.850 587.550 340.950 ;
        RECT 569.550 327.750 571.350 330.600 ;
        RECT 572.850 327.750 574.650 333.600 ;
        RECT 575.850 327.750 577.650 333.600 ;
        RECT 586.050 330.600 587.550 338.850 ;
        RECT 582.750 327.750 584.550 330.600 ;
        RECT 585.750 327.750 587.550 330.600 ;
        RECT 589.650 348.450 607.050 349.350 ;
        RECT 589.650 333.600 590.850 348.450 ;
        RECT 591.750 346.350 604.050 347.550 ;
        RECT 604.950 347.250 607.050 348.450 ;
        RECT 610.950 348.600 613.050 349.350 ;
        RECT 629.100 348.600 631.050 349.650 ;
        RECT 645.000 348.900 646.800 349.650 ;
        RECT 610.950 347.250 631.050 348.600 ;
        RECT 631.950 348.150 634.050 348.750 ;
        RECT 631.950 346.950 643.500 348.150 ;
        RECT 631.950 346.650 634.050 346.950 ;
        RECT 641.700 346.350 643.500 346.950 ;
        RECT 591.750 345.750 593.550 346.350 ;
        RECT 603.000 345.450 631.050 346.350 ;
        RECT 603.000 345.150 642.750 345.450 ;
        RECT 595.950 341.100 598.050 345.150 ;
        RECT 629.100 344.550 643.050 345.150 ;
        RECT 599.100 342.000 606.150 343.800 ;
        RECT 595.950 340.050 604.200 341.100 ;
        RECT 591.900 337.200 599.700 339.000 ;
        RECT 603.150 338.250 604.200 340.050 ;
        RECT 605.250 340.350 606.150 342.000 ;
        RECT 607.500 343.650 622.050 344.250 ;
        RECT 607.500 343.050 630.600 343.650 ;
        RECT 639.150 343.350 643.050 344.550 ;
        RECT 607.500 341.250 609.300 343.050 ;
        RECT 619.950 342.450 630.600 343.050 ;
        RECT 619.950 342.150 622.050 342.450 ;
        RECT 628.800 341.850 630.600 342.450 ;
        RECT 631.500 342.450 638.250 343.350 ;
        RECT 640.950 343.050 643.050 343.350 ;
        RECT 615.750 341.250 617.850 341.550 ;
        RECT 605.250 339.300 614.850 340.350 ;
        RECT 615.750 339.450 619.650 341.250 ;
        RECT 631.500 340.950 632.550 342.450 ;
        RECT 620.550 340.050 632.550 340.950 ;
        RECT 613.950 338.550 614.850 339.300 ;
        RECT 620.550 338.550 621.600 340.050 ;
        RECT 633.450 339.750 635.250 341.550 ;
        RECT 637.050 340.050 638.250 342.450 ;
        RECT 646.950 341.850 649.050 343.950 ;
        RECT 647.100 340.050 648.900 341.850 ;
        RECT 603.150 337.200 613.050 338.250 ;
        RECT 613.950 337.200 621.600 338.550 ;
        RECT 622.950 337.350 626.850 339.150 ;
        RECT 598.200 333.600 599.700 337.200 ;
        RECT 612.000 336.300 613.050 337.200 ;
        RECT 622.950 337.050 625.050 337.350 ;
        RECT 630.150 336.300 631.950 336.750 ;
        RECT 633.450 336.300 634.500 339.750 ;
        RECT 637.050 339.000 648.900 340.050 ;
        RECT 650.100 338.100 651.300 351.600 ;
        RECT 659.100 342.150 660.900 343.950 ;
        RECT 658.950 340.050 661.050 342.150 ;
        RECT 604.350 334.500 611.100 336.300 ;
        RECT 612.000 334.500 618.900 336.300 ;
        RECT 630.150 335.850 634.500 336.300 ;
        RECT 626.850 335.100 634.500 335.850 ;
        RECT 636.000 337.200 651.300 338.100 ;
        RECT 626.850 334.950 631.950 335.100 ;
        RECT 626.850 333.600 627.750 334.950 ;
        RECT 636.000 334.050 637.050 337.200 ;
        RECT 645.300 335.700 647.100 336.300 ;
        RECT 589.650 327.750 591.450 333.600 ;
        RECT 595.050 327.750 596.850 333.600 ;
        RECT 598.200 332.400 602.400 333.600 ;
        RECT 600.600 327.750 602.400 332.400 ;
        RECT 604.950 331.500 607.050 333.600 ;
        RECT 607.950 331.500 610.050 333.600 ;
        RECT 610.950 331.500 613.050 333.600 ;
        RECT 615.750 333.300 617.850 333.600 ;
        RECT 605.250 327.750 607.050 331.500 ;
        RECT 608.250 327.750 610.050 331.500 ;
        RECT 611.250 327.750 613.050 331.500 ;
        RECT 615.000 331.500 617.850 333.300 ;
        RECT 619.950 333.300 622.050 333.600 ;
        RECT 619.950 331.500 622.800 333.300 ;
        RECT 623.700 332.250 627.750 333.600 ;
        RECT 623.700 331.800 625.500 332.250 ;
        RECT 628.950 331.950 631.050 334.050 ;
        RECT 631.950 331.950 634.050 334.050 ;
        RECT 634.950 331.950 637.050 334.050 ;
        RECT 638.700 334.500 647.100 335.700 ;
        RECT 638.700 333.600 640.200 334.500 ;
        RECT 650.100 333.600 651.300 337.200 ;
        RECT 662.700 336.300 663.900 353.400 ;
        RECT 666.150 347.400 667.950 359.250 ;
        RECT 669.150 347.400 670.950 359.250 ;
        RECT 680.550 348.600 682.350 359.250 ;
        RECT 683.550 349.500 685.350 359.250 ;
        RECT 686.550 358.500 694.350 359.250 ;
        RECT 686.550 348.600 688.350 358.500 ;
        RECT 680.550 347.700 688.350 348.600 ;
        RECT 689.550 347.400 691.350 357.600 ;
        RECT 692.550 347.400 694.350 358.500 ;
        RECT 704.550 353.400 706.350 359.250 ;
        RECT 707.550 353.400 709.350 359.250 ;
        RECT 710.550 353.400 712.350 359.250 ;
        RECT 664.950 341.850 667.050 343.950 ;
        RECT 669.150 342.150 670.350 347.400 ;
        RECT 689.400 346.500 691.200 347.400 ;
        RECT 687.150 345.600 691.200 346.500 ;
        RECT 680.250 342.150 682.050 343.950 ;
        RECT 687.150 342.150 688.050 345.600 ;
        RECT 707.550 345.150 708.750 353.400 ;
        RECT 724.350 347.400 726.150 359.250 ;
        RECT 727.350 347.400 729.150 359.250 ;
        RECT 730.650 353.400 732.450 359.250 ;
        RECT 740.550 353.400 742.350 359.250 ;
        RECT 743.550 353.400 745.350 359.250 ;
        RECT 692.100 342.150 693.900 343.950 ;
        RECT 665.100 340.050 666.900 341.850 ;
        RECT 667.950 340.050 670.350 342.150 ;
        RECT 679.950 340.050 682.050 342.150 ;
        RECT 615.000 327.750 616.800 331.500 ;
        RECT 618.000 327.750 619.800 330.600 ;
        RECT 621.000 327.750 622.800 331.500 ;
        RECT 628.950 330.600 630.300 331.950 ;
        RECT 631.950 330.600 633.300 331.950 ;
        RECT 634.950 330.600 636.300 331.950 ;
        RECT 625.500 327.750 627.300 330.600 ;
        RECT 628.500 327.750 630.300 330.600 ;
        RECT 631.500 327.750 633.300 330.600 ;
        RECT 634.500 327.750 636.300 330.600 ;
        RECT 638.700 327.750 640.500 333.600 ;
        RECT 644.100 327.750 645.900 333.600 ;
        RECT 649.500 327.750 651.300 333.600 ;
        RECT 659.550 335.100 667.050 336.300 ;
        RECT 659.550 327.750 661.350 335.100 ;
        RECT 665.250 334.500 667.050 335.100 ;
        RECT 669.150 333.600 670.350 340.050 ;
        RECT 682.950 338.850 685.050 340.950 ;
        RECT 683.250 337.050 685.050 338.850 ;
        RECT 685.950 340.050 688.050 342.150 ;
        RECT 685.950 333.600 687.000 340.050 ;
        RECT 688.950 338.850 691.050 340.950 ;
        RECT 691.950 340.050 694.050 342.150 ;
        RECT 703.950 341.850 706.050 343.950 ;
        RECT 706.950 343.050 709.050 345.150 ;
        RECT 704.100 340.050 705.900 341.850 ;
        RECT 688.950 337.050 690.750 338.850 ;
        RECT 707.550 335.700 708.750 343.050 ;
        RECT 709.950 341.850 712.050 343.950 ;
        RECT 724.650 342.150 725.850 347.400 ;
        RECT 731.250 346.500 732.450 353.400 ;
        RECT 726.750 345.600 732.450 346.500 ;
        RECT 726.750 344.700 729.000 345.600 ;
        RECT 710.100 340.050 711.900 341.850 ;
        RECT 724.650 340.050 727.050 342.150 ;
        RECT 707.550 334.800 711.150 335.700 ;
        RECT 664.050 327.750 665.850 333.600 ;
        RECT 667.050 332.100 670.350 333.600 ;
        RECT 667.050 327.750 668.850 332.100 ;
        RECT 681.000 327.750 682.800 333.600 ;
        RECT 685.200 327.750 687.000 333.600 ;
        RECT 689.400 327.750 691.200 333.600 ;
        RECT 704.850 327.750 706.650 333.600 ;
        RECT 709.350 327.750 711.150 334.800 ;
        RECT 724.650 333.600 725.850 340.050 ;
        RECT 727.950 336.300 729.000 344.700 ;
        RECT 731.100 342.150 732.900 343.950 ;
        RECT 730.950 340.050 733.050 342.150 ;
        RECT 743.400 340.950 744.600 353.400 ;
        RECT 755.550 348.600 757.350 359.250 ;
        RECT 758.550 349.500 760.350 359.250 ;
        RECT 761.550 358.500 769.350 359.250 ;
        RECT 761.550 348.600 763.350 358.500 ;
        RECT 755.550 347.700 763.350 348.600 ;
        RECT 764.550 347.400 766.350 357.600 ;
        RECT 767.550 347.400 769.350 358.500 ;
        RECT 779.550 353.400 781.350 359.250 ;
        RECT 782.550 353.400 784.350 359.250 ;
        RECT 785.550 353.400 787.350 359.250 ;
        RECT 772.950 348.450 775.050 349.050 ;
        RECT 778.950 348.450 781.050 349.050 ;
        RECT 772.950 347.550 781.050 348.450 ;
        RECT 764.400 346.500 766.200 347.400 ;
        RECT 772.950 346.950 775.050 347.550 ;
        RECT 778.950 346.950 781.050 347.550 ;
        RECT 762.150 345.600 766.200 346.500 ;
        RECT 755.250 342.150 757.050 343.950 ;
        RECT 762.150 342.150 763.050 345.600 ;
        RECT 782.550 345.150 783.750 353.400 ;
        RECT 797.550 347.400 799.350 359.250 ;
        RECT 800.550 347.400 802.350 359.250 ;
        RECT 812.550 353.400 814.350 359.250 ;
        RECT 815.550 353.400 817.350 359.250 ;
        RECT 818.550 353.400 820.350 359.250 ;
        RECT 830.550 353.400 832.350 359.250 ;
        RECT 833.550 353.400 835.350 359.250 ;
        RECT 787.950 345.450 790.050 346.050 ;
        RECT 796.950 345.450 799.050 346.050 ;
        RECT 767.100 342.150 768.900 343.950 ;
        RECT 740.100 339.150 741.900 340.950 ;
        RECT 739.950 337.050 742.050 339.150 ;
        RECT 742.950 338.850 745.050 340.950 ;
        RECT 754.950 340.050 757.050 342.150 ;
        RECT 757.950 338.850 760.050 340.950 ;
        RECT 726.750 335.400 729.000 336.300 ;
        RECT 726.750 334.500 731.850 335.400 ;
        RECT 724.350 327.750 726.150 333.600 ;
        RECT 727.350 327.750 729.150 333.600 ;
        RECT 730.650 330.600 731.850 334.500 ;
        RECT 743.400 330.600 744.600 338.850 ;
        RECT 758.250 337.050 760.050 338.850 ;
        RECT 760.950 340.050 763.050 342.150 ;
        RECT 760.950 333.600 762.000 340.050 ;
        RECT 763.950 338.850 766.050 340.950 ;
        RECT 766.950 340.050 769.050 342.150 ;
        RECT 778.950 341.850 781.050 343.950 ;
        RECT 781.950 343.050 784.050 345.150 ;
        RECT 787.950 344.550 799.050 345.450 ;
        RECT 787.950 343.950 790.050 344.550 ;
        RECT 796.950 343.950 799.050 344.550 ;
        RECT 779.100 340.050 780.900 341.850 ;
        RECT 763.950 337.050 765.750 338.850 ;
        RECT 782.550 335.700 783.750 343.050 ;
        RECT 784.950 341.850 787.050 343.950 ;
        RECT 800.400 342.150 801.600 347.400 ;
        RECT 815.550 345.150 816.750 353.400 ;
        RECT 785.100 340.050 786.900 341.850 ;
        RECT 796.950 338.850 799.050 340.950 ;
        RECT 799.950 340.050 802.050 342.150 ;
        RECT 811.950 341.850 814.050 343.950 ;
        RECT 814.950 343.050 817.050 345.150 ;
        RECT 812.100 340.050 813.900 341.850 ;
        RECT 797.100 337.050 798.900 338.850 ;
        RECT 782.550 334.800 786.150 335.700 ;
        RECT 730.650 327.750 732.450 330.600 ;
        RECT 740.550 327.750 742.350 330.600 ;
        RECT 743.550 327.750 745.350 330.600 ;
        RECT 756.000 327.750 757.800 333.600 ;
        RECT 760.200 327.750 762.000 333.600 ;
        RECT 764.400 327.750 766.200 333.600 ;
        RECT 779.850 327.750 781.650 333.600 ;
        RECT 784.350 327.750 786.150 334.800 ;
        RECT 800.400 333.600 801.600 340.050 ;
        RECT 815.550 335.700 816.750 343.050 ;
        RECT 817.950 341.850 820.050 343.950 ;
        RECT 818.100 340.050 819.900 341.850 ;
        RECT 833.400 340.950 834.600 353.400 ;
        RECT 845.550 352.200 847.350 358.200 ;
        RECT 848.550 352.200 850.350 359.250 ;
        RECT 846.450 347.100 847.350 352.200 ;
        RECT 853.050 348.900 854.850 358.200 ;
        RECT 853.050 348.000 855.150 348.900 ;
        RECT 846.450 346.200 852.600 347.100 ;
        RECT 848.250 342.150 850.050 343.950 ;
        RECT 830.100 339.150 831.900 340.950 ;
        RECT 829.950 337.050 832.050 339.150 ;
        RECT 832.950 338.850 835.050 340.950 ;
        RECT 844.950 338.850 847.050 340.950 ;
        RECT 847.950 340.050 850.050 342.150 ;
        RECT 851.250 343.500 852.600 346.200 ;
        RECT 851.250 341.700 853.050 343.500 ;
        RECT 815.550 334.800 819.150 335.700 ;
        RECT 797.550 327.750 799.350 333.600 ;
        RECT 800.550 327.750 802.350 333.600 ;
        RECT 812.850 327.750 814.650 333.600 ;
        RECT 817.350 327.750 819.150 334.800 ;
        RECT 833.400 330.600 834.600 338.850 ;
        RECT 845.250 337.050 847.050 338.850 ;
        RECT 851.250 336.000 852.600 341.700 ;
        RECT 854.250 340.950 855.150 348.000 ;
        RECT 857.550 347.400 859.350 359.250 ;
        RECT 857.100 342.150 858.900 343.950 ;
        RECT 853.950 338.850 856.050 340.950 ;
        RECT 856.950 340.050 859.050 342.150 ;
        RECT 846.300 335.100 852.600 336.000 ;
        RECT 846.300 331.800 847.350 335.100 ;
        RECT 854.250 334.200 855.150 338.850 ;
        RECT 853.050 333.300 855.150 334.200 ;
        RECT 830.550 327.750 832.350 330.600 ;
        RECT 833.550 327.750 835.350 330.600 ;
        RECT 845.550 328.800 847.350 331.800 ;
        RECT 848.550 327.750 850.350 331.800 ;
        RECT 853.050 328.800 854.850 333.300 ;
        RECT 857.550 327.750 859.350 334.800 ;
        RECT 13.350 317.400 15.150 323.250 ;
        RECT 16.350 317.400 18.150 323.250 ;
        RECT 19.650 320.400 21.450 323.250 ;
        RECT 13.650 310.950 14.850 317.400 ;
        RECT 19.650 316.500 20.850 320.400 ;
        RECT 15.750 315.600 20.850 316.500 ;
        RECT 15.750 314.700 18.000 315.600 ;
        RECT 38.100 315.000 39.900 323.250 ;
        RECT 13.650 308.850 16.050 310.950 ;
        RECT 13.650 303.600 14.850 308.850 ;
        RECT 16.950 306.300 18.000 314.700 ;
        RECT 35.400 313.350 39.900 315.000 ;
        RECT 43.500 314.400 45.300 323.250 ;
        RECT 54.000 317.400 55.800 323.250 ;
        RECT 58.200 319.050 60.000 323.250 ;
        RECT 61.500 320.400 63.300 323.250 ;
        RECT 76.650 320.400 78.450 323.250 ;
        RECT 79.650 320.400 81.450 323.250 ;
        RECT 58.200 317.400 63.900 319.050 ;
        RECT 19.950 308.850 22.050 310.950 ;
        RECT 35.400 309.150 36.600 313.350 ;
        RECT 40.950 312.450 43.050 313.050 ;
        RECT 49.950 312.450 52.050 313.050 ;
        RECT 40.950 311.550 52.050 312.450 ;
        RECT 53.100 312.150 54.900 313.950 ;
        RECT 40.950 310.950 43.050 311.550 ;
        RECT 49.950 310.950 52.050 311.550 ;
        RECT 52.950 310.050 55.050 312.150 ;
        RECT 55.950 311.850 58.050 313.950 ;
        RECT 59.100 312.150 60.900 313.950 ;
        RECT 56.100 310.050 57.900 311.850 ;
        RECT 58.950 310.050 61.050 312.150 ;
        RECT 62.700 310.950 63.900 317.400 ;
        RECT 77.400 312.150 78.600 320.400 ;
        RECT 91.650 317.400 93.450 323.250 ;
        RECT 92.250 315.300 93.450 317.400 ;
        RECT 94.650 318.300 96.450 323.250 ;
        RECT 97.650 319.200 99.450 323.250 ;
        RECT 100.650 318.300 102.450 323.250 ;
        RECT 113.700 320.400 115.500 323.250 ;
        RECT 117.000 319.050 118.800 323.250 ;
        RECT 94.650 316.950 102.450 318.300 ;
        RECT 113.100 317.400 118.800 319.050 ;
        RECT 121.200 317.400 123.000 323.250 ;
        RECT 92.250 314.250 96.000 315.300 ;
        RECT 20.100 307.050 21.900 308.850 ;
        RECT 34.950 307.050 37.050 309.150 ;
        RECT 61.950 308.850 64.050 310.950 ;
        RECT 76.950 310.050 79.050 312.150 ;
        RECT 79.950 311.850 82.050 313.950 ;
        RECT 80.100 310.050 81.900 311.850 ;
        RECT 94.950 310.950 96.150 314.250 ;
        RECT 98.100 312.150 99.900 313.950 ;
        RECT 15.750 305.400 18.000 306.300 ;
        RECT 15.750 304.500 21.450 305.400 ;
        RECT 13.350 291.750 15.150 303.600 ;
        RECT 16.350 291.750 18.150 303.600 ;
        RECT 20.250 297.600 21.450 304.500 ;
        RECT 35.250 298.800 36.300 307.050 ;
        RECT 37.950 305.850 40.050 307.950 ;
        RECT 43.950 305.850 46.050 307.950 ;
        RECT 37.950 304.050 39.750 305.850 ;
        RECT 40.950 302.850 43.050 304.950 ;
        RECT 44.100 304.050 45.900 305.850 ;
        RECT 62.700 303.600 63.900 308.850 ;
        RECT 41.100 301.050 42.900 302.850 ;
        RECT 53.550 302.700 61.350 303.600 ;
        RECT 35.250 297.900 42.300 298.800 ;
        RECT 35.250 297.600 36.450 297.900 ;
        RECT 19.650 291.750 21.450 297.600 ;
        RECT 34.650 291.750 36.450 297.600 ;
        RECT 40.650 297.600 42.300 297.900 ;
        RECT 37.650 291.750 39.450 297.000 ;
        RECT 40.650 291.750 42.450 297.600 ;
        RECT 43.650 291.750 45.450 297.600 ;
        RECT 53.550 291.750 55.350 302.700 ;
        RECT 56.550 291.750 58.350 301.800 ;
        RECT 59.550 291.750 61.350 302.700 ;
        RECT 62.550 291.750 64.350 303.600 ;
        RECT 77.400 297.600 78.600 310.050 ;
        RECT 94.950 308.850 97.050 310.950 ;
        RECT 97.950 310.050 100.050 312.150 ;
        RECT 113.100 310.950 114.300 317.400 ;
        RECT 131.700 314.400 133.500 323.250 ;
        RECT 137.100 315.000 138.900 323.250 ;
        RECT 161.100 315.000 162.900 323.250 ;
        RECT 116.100 312.150 117.900 313.950 ;
        RECT 100.950 308.850 103.050 310.950 ;
        RECT 112.950 308.850 115.050 310.950 ;
        RECT 115.950 310.050 118.050 312.150 ;
        RECT 118.950 311.850 121.050 313.950 ;
        RECT 122.100 312.150 123.900 313.950 ;
        RECT 137.100 313.350 141.600 315.000 ;
        RECT 119.100 310.050 120.900 311.850 ;
        RECT 121.950 310.050 124.050 312.150 ;
        RECT 127.950 310.950 130.050 313.050 ;
        RECT 91.950 305.850 94.050 307.950 ;
        RECT 92.250 304.050 94.050 305.850 ;
        RECT 95.850 303.600 97.050 308.850 ;
        RECT 101.100 307.050 102.900 308.850 ;
        RECT 113.100 303.600 114.300 308.850 ;
        RECT 121.950 306.450 124.050 307.050 ;
        RECT 128.550 306.450 129.450 310.950 ;
        RECT 140.400 309.150 141.600 313.350 ;
        RECT 158.400 313.350 162.900 315.000 ;
        RECT 166.500 314.400 168.300 323.250 ;
        RECT 178.650 317.400 180.450 323.250 ;
        RECT 179.250 315.300 180.450 317.400 ;
        RECT 181.650 318.300 183.450 323.250 ;
        RECT 184.650 319.200 186.450 323.250 ;
        RECT 187.650 318.300 189.450 323.250 ;
        RECT 181.650 316.950 189.450 318.300 ;
        RECT 199.650 317.400 201.450 323.250 ;
        RECT 200.250 315.300 201.450 317.400 ;
        RECT 202.650 318.300 204.450 323.250 ;
        RECT 205.650 319.200 207.450 323.250 ;
        RECT 208.650 318.300 210.450 323.250 ;
        RECT 221.700 320.400 223.500 323.250 ;
        RECT 225.000 319.050 226.800 323.250 ;
        RECT 202.650 316.950 210.450 318.300 ;
        RECT 221.100 317.400 226.800 319.050 ;
        RECT 229.200 317.400 231.000 323.250 ;
        RECT 179.250 314.250 183.000 315.300 ;
        RECT 200.250 314.250 204.000 315.300 ;
        RECT 158.400 309.150 159.600 313.350 ;
        RECT 181.950 310.950 183.150 314.250 ;
        RECT 185.100 312.150 186.900 313.950 ;
        RECT 121.950 305.550 129.450 306.450 ;
        RECT 130.950 305.850 133.050 307.950 ;
        RECT 136.950 305.850 139.050 307.950 ;
        RECT 139.950 307.050 142.050 309.150 ;
        RECT 157.950 307.050 160.050 309.150 ;
        RECT 181.950 308.850 184.050 310.950 ;
        RECT 184.950 310.050 187.050 312.150 ;
        RECT 202.950 310.950 204.150 314.250 ;
        RECT 206.100 312.150 207.900 313.950 ;
        RECT 187.950 308.850 190.050 310.950 ;
        RECT 202.950 308.850 205.050 310.950 ;
        RECT 205.950 310.050 208.050 312.150 ;
        RECT 221.100 310.950 222.300 317.400 ;
        RECT 245.100 315.000 246.900 323.250 ;
        RECT 224.100 312.150 225.900 313.950 ;
        RECT 208.950 308.850 211.050 310.950 ;
        RECT 220.950 308.850 223.050 310.950 ;
        RECT 223.950 310.050 226.050 312.150 ;
        RECT 226.950 311.850 229.050 313.950 ;
        RECT 230.100 312.150 231.900 313.950 ;
        RECT 242.400 313.350 246.900 315.000 ;
        RECT 250.500 314.400 252.300 323.250 ;
        RECT 260.550 318.300 262.350 323.250 ;
        RECT 263.550 319.200 265.350 323.250 ;
        RECT 266.550 318.300 268.350 323.250 ;
        RECT 260.550 316.950 268.350 318.300 ;
        RECT 269.550 317.400 271.350 323.250 ;
        RECT 282.000 317.400 283.800 323.250 ;
        RECT 286.200 319.050 288.000 323.250 ;
        RECT 289.500 320.400 291.300 323.250 ;
        RECT 313.650 320.400 315.450 323.250 ;
        RECT 316.650 320.400 318.450 323.250 ;
        RECT 319.650 320.400 321.450 323.250 ;
        RECT 322.650 320.400 324.750 323.250 ;
        RECT 313.650 319.500 314.700 320.400 ;
        RECT 319.650 319.500 320.700 320.400 ;
        RECT 286.200 317.400 291.900 319.050 ;
        RECT 269.550 315.300 270.750 317.400 ;
        RECT 267.000 314.250 270.750 315.300 ;
        RECT 227.100 310.050 228.900 311.850 ;
        RECT 229.950 310.050 232.050 312.150 ;
        RECT 242.400 309.150 243.600 313.350 ;
        RECT 263.100 312.150 264.900 313.950 ;
        RECT 121.950 304.950 124.050 305.550 ;
        RECT 131.100 304.050 132.900 305.850 ;
        RECT 76.650 291.750 78.450 297.600 ;
        RECT 79.650 291.750 81.450 297.600 ;
        RECT 92.400 291.750 94.200 297.600 ;
        RECT 95.700 291.750 97.500 303.600 ;
        RECT 99.900 291.750 101.700 303.600 ;
        RECT 112.650 291.750 114.450 303.600 ;
        RECT 115.650 302.700 123.450 303.600 ;
        RECT 133.950 302.850 136.050 304.950 ;
        RECT 137.250 304.050 139.050 305.850 ;
        RECT 115.650 291.750 117.450 302.700 ;
        RECT 118.650 291.750 120.450 301.800 ;
        RECT 121.650 291.750 123.450 302.700 ;
        RECT 134.100 301.050 135.900 302.850 ;
        RECT 140.700 298.800 141.750 307.050 ;
        RECT 134.700 297.900 141.750 298.800 ;
        RECT 134.700 297.600 136.350 297.900 ;
        RECT 131.550 291.750 133.350 297.600 ;
        RECT 134.550 291.750 136.350 297.600 ;
        RECT 140.550 297.600 141.750 297.900 ;
        RECT 158.250 298.800 159.300 307.050 ;
        RECT 160.950 305.850 163.050 307.950 ;
        RECT 166.950 305.850 169.050 307.950 ;
        RECT 178.950 305.850 181.050 307.950 ;
        RECT 160.950 304.050 162.750 305.850 ;
        RECT 163.950 302.850 166.050 304.950 ;
        RECT 167.100 304.050 168.900 305.850 ;
        RECT 179.250 304.050 181.050 305.850 ;
        RECT 182.850 303.600 184.050 308.850 ;
        RECT 188.100 307.050 189.900 308.850 ;
        RECT 199.950 305.850 202.050 307.950 ;
        RECT 200.250 304.050 202.050 305.850 ;
        RECT 203.850 303.600 205.050 308.850 ;
        RECT 209.100 307.050 210.900 308.850 ;
        RECT 221.100 303.600 222.300 308.850 ;
        RECT 241.950 307.050 244.050 309.150 ;
        RECT 259.950 308.850 262.050 310.950 ;
        RECT 262.950 310.050 265.050 312.150 ;
        RECT 266.850 310.950 268.050 314.250 ;
        RECT 281.100 312.150 282.900 313.950 ;
        RECT 265.950 308.850 268.050 310.950 ;
        RECT 280.950 310.050 283.050 312.150 ;
        RECT 283.950 311.850 286.050 313.950 ;
        RECT 287.100 312.150 288.900 313.950 ;
        RECT 284.100 310.050 285.900 311.850 ;
        RECT 286.950 310.050 289.050 312.150 ;
        RECT 290.700 310.950 291.900 317.400 ;
        RECT 309.900 318.600 320.700 319.500 ;
        RECT 309.900 312.150 311.100 318.600 ;
        RECT 341.100 315.000 342.900 323.250 ;
        RECT 317.100 312.150 318.900 313.950 ;
        RECT 338.400 313.350 342.900 315.000 ;
        RECT 346.500 314.400 348.300 323.250 ;
        RECT 351.750 320.400 353.550 323.250 ;
        RECT 354.750 320.400 356.550 323.250 ;
        RECT 289.950 308.850 292.050 310.950 ;
        RECT 307.950 310.050 311.100 312.150 ;
        RECT 164.100 301.050 165.900 302.850 ;
        RECT 158.250 297.900 165.300 298.800 ;
        RECT 158.250 297.600 159.450 297.900 ;
        RECT 137.550 291.750 139.350 297.000 ;
        RECT 140.550 291.750 142.350 297.600 ;
        RECT 157.650 291.750 159.450 297.600 ;
        RECT 163.650 297.600 165.300 297.900 ;
        RECT 160.650 291.750 162.450 297.000 ;
        RECT 163.650 291.750 165.450 297.600 ;
        RECT 166.650 291.750 168.450 297.600 ;
        RECT 179.400 291.750 181.200 297.600 ;
        RECT 182.700 291.750 184.500 303.600 ;
        RECT 186.900 291.750 188.700 303.600 ;
        RECT 200.400 291.750 202.200 297.600 ;
        RECT 203.700 291.750 205.500 303.600 ;
        RECT 207.900 291.750 209.700 303.600 ;
        RECT 220.650 291.750 222.450 303.600 ;
        RECT 223.650 302.700 231.450 303.600 ;
        RECT 223.650 291.750 225.450 302.700 ;
        RECT 226.650 291.750 228.450 301.800 ;
        RECT 229.650 291.750 231.450 302.700 ;
        RECT 242.250 298.800 243.300 307.050 ;
        RECT 244.950 305.850 247.050 307.950 ;
        RECT 250.950 305.850 253.050 307.950 ;
        RECT 260.100 307.050 261.900 308.850 ;
        RECT 244.950 304.050 246.750 305.850 ;
        RECT 247.950 302.850 250.050 304.950 ;
        RECT 251.100 304.050 252.900 305.850 ;
        RECT 265.950 303.600 267.150 308.850 ;
        RECT 268.950 305.850 271.050 307.950 ;
        RECT 268.950 304.050 270.750 305.850 ;
        RECT 290.700 303.600 291.900 308.850 ;
        RECT 309.900 304.800 311.100 310.050 ;
        RECT 313.950 308.850 316.050 310.950 ;
        RECT 316.950 310.050 319.050 312.150 ;
        RECT 322.950 308.850 325.050 310.950 ;
        RECT 338.400 309.150 339.600 313.350 ;
        RECT 355.050 312.150 356.550 320.400 ;
        RECT 352.950 310.050 356.550 312.150 ;
        RECT 314.100 307.050 315.900 308.850 ;
        RECT 323.100 307.050 324.900 308.850 ;
        RECT 337.950 307.050 340.050 309.150 ;
        RECT 307.650 303.600 311.100 304.800 ;
        RECT 248.100 301.050 249.900 302.850 ;
        RECT 242.250 297.900 249.300 298.800 ;
        RECT 242.250 297.600 243.450 297.900 ;
        RECT 241.650 291.750 243.450 297.600 ;
        RECT 247.650 297.600 249.300 297.900 ;
        RECT 244.650 291.750 246.450 297.000 ;
        RECT 247.650 291.750 249.450 297.600 ;
        RECT 250.650 291.750 252.450 297.600 ;
        RECT 261.300 291.750 263.100 303.600 ;
        RECT 265.500 291.750 267.300 303.600 ;
        RECT 281.550 302.700 289.350 303.600 ;
        RECT 268.800 291.750 270.600 297.600 ;
        RECT 281.550 291.750 283.350 302.700 ;
        RECT 284.550 291.750 286.350 301.800 ;
        RECT 287.550 291.750 289.350 302.700 ;
        RECT 290.550 291.750 292.350 303.600 ;
        RECT 304.050 292.500 305.850 301.800 ;
        RECT 307.650 301.200 308.850 303.600 ;
        RECT 307.050 293.400 308.850 301.200 ;
        RECT 310.050 301.200 318.450 302.100 ;
        RECT 310.050 292.500 311.850 301.200 ;
        RECT 304.050 291.750 311.850 292.500 ;
        RECT 313.650 292.500 315.450 300.300 ;
        RECT 316.650 293.400 318.450 301.200 ;
        RECT 319.650 301.500 327.450 302.400 ;
        RECT 319.650 292.500 321.450 301.500 ;
        RECT 313.650 291.750 321.450 292.500 ;
        RECT 322.650 291.750 324.450 300.600 ;
        RECT 325.650 291.750 327.450 301.500 ;
        RECT 338.250 298.800 339.300 307.050 ;
        RECT 340.950 305.850 343.050 307.950 ;
        RECT 346.950 305.850 349.050 307.950 ;
        RECT 340.950 304.050 342.750 305.850 ;
        RECT 343.950 302.850 346.050 304.950 ;
        RECT 347.100 304.050 348.900 305.850 ;
        RECT 344.100 301.050 345.900 302.850 ;
        RECT 338.250 297.900 345.300 298.800 ;
        RECT 338.250 297.600 339.450 297.900 ;
        RECT 337.650 291.750 339.450 297.600 ;
        RECT 343.650 297.600 345.300 297.900 ;
        RECT 355.050 297.600 356.550 310.050 ;
        RECT 358.650 317.400 360.450 323.250 ;
        RECT 364.050 317.400 365.850 323.250 ;
        RECT 369.600 318.600 371.400 323.250 ;
        RECT 374.250 319.500 376.050 323.250 ;
        RECT 377.250 319.500 379.050 323.250 ;
        RECT 380.250 319.500 382.050 323.250 ;
        RECT 367.200 317.400 371.400 318.600 ;
        RECT 373.950 317.400 376.050 319.500 ;
        RECT 376.950 317.400 379.050 319.500 ;
        RECT 379.950 317.400 382.050 319.500 ;
        RECT 384.000 319.500 385.800 323.250 ;
        RECT 387.000 320.400 388.800 323.250 ;
        RECT 390.000 319.500 391.800 323.250 ;
        RECT 394.500 320.400 396.300 323.250 ;
        RECT 397.500 320.400 399.300 323.250 ;
        RECT 400.500 320.400 402.300 323.250 ;
        RECT 403.500 320.400 405.300 323.250 ;
        RECT 384.000 317.700 386.850 319.500 ;
        RECT 384.750 317.400 386.850 317.700 ;
        RECT 388.950 317.700 391.800 319.500 ;
        RECT 392.700 318.750 394.500 319.200 ;
        RECT 397.950 319.050 399.300 320.400 ;
        RECT 400.950 319.050 402.300 320.400 ;
        RECT 403.950 319.050 405.300 320.400 ;
        RECT 388.950 317.400 391.050 317.700 ;
        RECT 392.700 317.400 396.750 318.750 ;
        RECT 358.650 302.550 359.850 317.400 ;
        RECT 367.200 313.800 368.700 317.400 ;
        RECT 373.350 314.700 380.100 316.500 ;
        RECT 381.000 314.700 387.900 316.500 ;
        RECT 395.850 316.050 396.750 317.400 ;
        RECT 397.950 316.950 400.050 319.050 ;
        RECT 400.950 316.950 403.050 319.050 ;
        RECT 403.950 316.950 406.050 319.050 ;
        RECT 395.850 315.900 400.950 316.050 ;
        RECT 395.850 315.150 403.500 315.900 ;
        RECT 399.150 314.700 403.500 315.150 ;
        RECT 381.000 313.800 382.050 314.700 ;
        RECT 399.150 314.250 400.950 314.700 ;
        RECT 360.900 312.000 368.700 313.800 ;
        RECT 372.150 312.750 382.050 313.800 ;
        RECT 372.150 310.950 373.200 312.750 ;
        RECT 382.950 312.450 390.600 313.800 ;
        RECT 382.950 311.700 383.850 312.450 ;
        RECT 364.950 309.900 373.200 310.950 ;
        RECT 374.250 310.650 383.850 311.700 ;
        RECT 364.950 305.850 367.050 309.900 ;
        RECT 374.250 309.000 375.150 310.650 ;
        RECT 384.750 309.750 388.650 311.550 ;
        RECT 389.550 310.950 390.600 312.450 ;
        RECT 391.950 313.650 394.050 313.950 ;
        RECT 391.950 311.850 395.850 313.650 ;
        RECT 402.450 311.250 403.500 314.700 ;
        RECT 405.000 313.800 406.050 316.950 ;
        RECT 407.700 317.400 409.500 323.250 ;
        RECT 413.100 317.400 414.900 323.250 ;
        RECT 418.500 317.400 420.300 323.250 ;
        RECT 407.700 316.500 409.200 317.400 ;
        RECT 407.700 315.300 416.100 316.500 ;
        RECT 414.300 314.700 416.100 315.300 ;
        RECT 419.100 313.800 420.300 317.400 ;
        RECT 428.550 318.300 430.350 323.250 ;
        RECT 431.550 319.200 433.350 323.250 ;
        RECT 434.550 318.300 436.350 323.250 ;
        RECT 428.550 316.950 436.350 318.300 ;
        RECT 437.550 317.400 439.350 323.250 ;
        RECT 437.550 315.300 438.750 317.400 ;
        RECT 452.850 316.200 454.650 323.250 ;
        RECT 457.350 317.400 459.150 323.250 ;
        RECT 467.850 317.400 469.650 323.250 ;
        RECT 472.350 316.200 474.150 323.250 ;
        RECT 488.550 320.400 490.350 323.250 ;
        RECT 491.550 320.400 493.350 323.250 ;
        RECT 494.550 320.400 496.350 323.250 ;
        RECT 452.850 315.300 456.450 316.200 ;
        RECT 435.000 314.250 438.750 315.300 ;
        RECT 405.000 312.900 420.300 313.800 ;
        RECT 389.550 310.050 401.550 310.950 ;
        RECT 368.100 307.200 375.150 309.000 ;
        RECT 376.500 307.950 378.300 309.750 ;
        RECT 384.750 309.450 386.850 309.750 ;
        RECT 388.950 308.550 391.050 308.850 ;
        RECT 397.800 308.550 399.600 309.150 ;
        RECT 388.950 307.950 399.600 308.550 ;
        RECT 376.500 307.350 399.600 307.950 ;
        RECT 400.500 308.550 401.550 310.050 ;
        RECT 402.450 309.450 404.250 311.250 ;
        RECT 406.050 310.950 417.900 312.000 ;
        RECT 406.050 308.550 407.250 310.950 ;
        RECT 416.100 309.150 417.900 310.950 ;
        RECT 400.500 307.650 407.250 308.550 ;
        RECT 409.950 307.650 412.050 307.950 ;
        RECT 376.500 306.750 391.050 307.350 ;
        RECT 408.150 306.450 412.050 307.650 ;
        RECT 415.950 307.050 418.050 309.150 ;
        RECT 398.100 305.850 412.050 306.450 ;
        RECT 372.000 305.550 411.750 305.850 ;
        RECT 360.750 304.650 362.550 305.250 ;
        RECT 372.000 304.650 400.050 305.550 ;
        RECT 360.750 303.450 373.050 304.650 ;
        RECT 400.950 304.050 403.050 304.350 ;
        RECT 410.700 304.050 412.500 304.650 ;
        RECT 373.950 302.550 376.050 303.750 ;
        RECT 358.650 301.650 376.050 302.550 ;
        RECT 379.950 302.400 400.050 303.750 ;
        RECT 379.950 301.650 382.050 302.400 ;
        RECT 361.500 297.600 362.700 301.650 ;
        RECT 363.600 299.700 365.400 300.300 ;
        RECT 370.350 300.150 372.150 300.300 ;
        RECT 363.600 298.500 369.300 299.700 ;
        RECT 370.350 298.950 379.050 300.150 ;
        RECT 370.350 298.500 372.150 298.950 ;
        RECT 340.650 291.750 342.450 297.000 ;
        RECT 343.650 291.750 345.450 297.600 ;
        RECT 346.650 291.750 348.450 297.600 ;
        RECT 351.750 291.750 353.550 297.600 ;
        RECT 354.750 291.750 356.550 297.600 ;
        RECT 358.500 291.750 360.300 297.600 ;
        RECT 361.500 291.750 363.300 297.600 ;
        RECT 364.500 291.750 366.300 297.600 ;
        RECT 367.500 291.750 369.300 298.500 ;
        RECT 376.950 298.050 379.050 298.950 ;
        RECT 370.500 291.750 372.300 297.600 ;
        RECT 373.800 295.800 375.900 297.900 ;
        RECT 374.400 294.600 375.900 295.800 ;
        RECT 374.250 291.750 376.050 294.600 ;
        RECT 377.250 291.750 379.050 298.050 ;
        RECT 380.550 294.600 381.900 301.650 ;
        RECT 398.100 301.350 400.050 302.400 ;
        RECT 400.950 302.850 412.500 304.050 ;
        RECT 400.950 302.250 403.050 302.850 ;
        RECT 414.000 301.350 415.800 302.100 ;
        RECT 383.100 298.800 387.000 300.600 ;
        RECT 384.000 298.500 387.000 298.800 ;
        RECT 388.950 300.150 391.050 300.600 ;
        RECT 398.100 300.300 415.800 301.350 ;
        RECT 388.950 298.500 391.350 300.150 ;
        RECT 380.250 291.750 382.050 294.600 ;
        RECT 384.000 291.750 385.800 298.500 ;
        RECT 390.000 297.600 391.350 298.500 ;
        RECT 397.950 297.600 400.050 298.050 ;
        RECT 387.000 291.750 388.800 297.600 ;
        RECT 390.000 291.750 391.800 297.600 ;
        RECT 393.750 291.750 395.550 297.600 ;
        RECT 397.500 295.950 400.050 297.600 ;
        RECT 400.950 295.950 403.050 298.050 ;
        RECT 403.950 295.950 406.050 298.050 ;
        RECT 397.500 294.600 398.700 295.950 ;
        RECT 400.950 294.600 401.850 295.950 ;
        RECT 403.950 294.600 405.150 295.950 ;
        RECT 396.750 291.750 398.700 294.600 ;
        RECT 399.750 291.750 401.850 294.600 ;
        RECT 402.750 291.750 405.150 294.600 ;
        RECT 406.500 291.750 408.300 295.050 ;
        RECT 409.500 291.750 411.300 300.300 ;
        RECT 419.100 299.400 420.300 312.900 ;
        RECT 431.100 312.150 432.900 313.950 ;
        RECT 427.950 308.850 430.050 310.950 ;
        RECT 430.950 310.050 433.050 312.150 ;
        RECT 434.850 310.950 436.050 314.250 ;
        RECT 433.950 308.850 436.050 310.950 ;
        RECT 452.100 309.150 453.900 310.950 ;
        RECT 428.100 307.050 429.900 308.850 ;
        RECT 433.950 303.600 435.150 308.850 ;
        RECT 436.950 305.850 439.050 307.950 ;
        RECT 451.950 307.050 454.050 309.150 ;
        RECT 455.250 307.950 456.450 315.300 ;
        RECT 470.550 315.300 474.150 316.200 ;
        RECT 458.100 309.150 459.900 310.950 ;
        RECT 467.100 309.150 468.900 310.950 ;
        RECT 454.950 305.850 457.050 307.950 ;
        RECT 457.950 307.050 460.050 309.150 ;
        RECT 466.950 307.050 469.050 309.150 ;
        RECT 470.550 307.950 471.750 315.300 ;
        RECT 492.000 313.950 493.050 320.400 ;
        RECT 510.150 318.900 511.950 323.250 ;
        RECT 490.950 311.850 493.050 313.950 ;
        RECT 473.100 309.150 474.900 310.950 ;
        RECT 469.950 305.850 472.050 307.950 ;
        RECT 472.950 307.050 475.050 309.150 ;
        RECT 487.950 308.850 490.050 310.950 ;
        RECT 488.100 307.050 489.900 308.850 ;
        RECT 436.950 304.050 438.750 305.850 ;
        RECT 416.250 298.500 420.300 299.400 ;
        RECT 416.250 297.600 417.300 298.500 ;
        RECT 412.500 291.750 414.300 297.600 ;
        RECT 415.500 291.750 417.300 297.600 ;
        RECT 418.500 291.750 420.300 297.600 ;
        RECT 429.300 291.750 431.100 303.600 ;
        RECT 433.500 291.750 435.300 303.600 ;
        RECT 436.950 300.450 439.050 301.050 ;
        RECT 448.950 300.450 451.050 301.050 ;
        RECT 436.950 299.550 451.050 300.450 ;
        RECT 436.950 298.950 439.050 299.550 ;
        RECT 448.950 298.950 451.050 299.550 ;
        RECT 455.250 297.600 456.450 305.850 ;
        RECT 470.550 297.600 471.750 305.850 ;
        RECT 492.000 304.650 493.050 311.850 ;
        RECT 508.650 317.400 511.950 318.900 ;
        RECT 513.150 317.400 514.950 323.250 ;
        RECT 508.650 310.950 509.850 317.400 ;
        RECT 511.950 315.900 513.750 316.500 ;
        RECT 517.650 315.900 519.450 323.250 ;
        RECT 528.000 317.400 529.800 323.250 ;
        RECT 532.200 319.050 534.000 323.250 ;
        RECT 535.500 320.400 537.300 323.250 ;
        RECT 532.200 317.400 537.900 319.050 ;
        RECT 553.650 317.400 555.450 323.250 ;
        RECT 556.650 317.400 558.450 323.250 ;
        RECT 511.950 314.700 519.450 315.900 ;
        RECT 493.950 308.850 496.050 310.950 ;
        RECT 508.650 308.850 511.050 310.950 ;
        RECT 512.100 309.150 513.900 310.950 ;
        RECT 494.100 307.050 495.900 308.850 ;
        RECT 492.000 303.600 494.550 304.650 ;
        RECT 508.650 303.600 509.850 308.850 ;
        RECT 511.950 307.050 514.050 309.150 ;
        RECT 436.800 291.750 438.600 297.600 ;
        RECT 451.650 291.750 453.450 297.600 ;
        RECT 454.650 291.750 456.450 297.600 ;
        RECT 457.650 291.750 459.450 297.600 ;
        RECT 467.550 291.750 469.350 297.600 ;
        RECT 470.550 291.750 472.350 297.600 ;
        RECT 473.550 291.750 475.350 297.600 ;
        RECT 488.550 291.750 490.350 303.600 ;
        RECT 492.750 291.750 494.550 303.600 ;
        RECT 508.050 291.750 509.850 303.600 ;
        RECT 511.050 291.750 512.850 303.600 ;
        RECT 515.100 297.600 516.300 314.700 ;
        RECT 527.100 312.150 528.900 313.950 ;
        RECT 517.950 308.850 520.050 310.950 ;
        RECT 526.950 310.050 529.050 312.150 ;
        RECT 529.950 311.850 532.050 313.950 ;
        RECT 533.100 312.150 534.900 313.950 ;
        RECT 530.100 310.050 531.900 311.850 ;
        RECT 532.950 310.050 535.050 312.150 ;
        RECT 536.700 310.950 537.900 317.400 ;
        RECT 554.400 310.950 555.600 317.400 ;
        RECT 569.700 314.400 571.500 323.250 ;
        RECT 575.100 315.000 576.900 323.250 ;
        RECT 593.550 317.400 595.350 323.250 ;
        RECT 596.550 317.400 598.350 323.250 ;
        RECT 615.150 318.900 616.950 323.250 ;
        RECT 613.650 317.400 616.950 318.900 ;
        RECT 618.150 317.400 619.950 323.250 ;
        RECT 557.100 312.150 558.900 313.950 ;
        RECT 575.100 313.350 579.600 315.000 ;
        RECT 535.950 308.850 538.050 310.950 ;
        RECT 553.950 308.850 556.050 310.950 ;
        RECT 556.950 310.050 559.050 312.150 ;
        RECT 578.400 309.150 579.600 313.350 ;
        RECT 593.100 312.150 594.900 313.950 ;
        RECT 592.950 310.050 595.050 312.150 ;
        RECT 596.400 310.950 597.600 317.400 ;
        RECT 613.650 310.950 614.850 317.400 ;
        RECT 616.950 315.900 618.750 316.500 ;
        RECT 622.650 315.900 624.450 323.250 ;
        RECT 616.950 314.700 624.450 315.900 ;
        RECT 635.850 316.200 637.650 323.250 ;
        RECT 640.350 317.400 642.150 323.250 ;
        RECT 652.650 317.400 654.450 323.250 ;
        RECT 635.850 315.300 639.450 316.200 ;
        RECT 518.100 307.050 519.900 308.850 ;
        RECT 536.700 303.600 537.900 308.850 ;
        RECT 554.400 303.600 555.600 308.850 ;
        RECT 556.950 306.450 559.050 307.050 ;
        RECT 565.950 306.450 568.050 307.050 ;
        RECT 556.950 305.550 568.050 306.450 ;
        RECT 568.950 305.850 571.050 307.950 ;
        RECT 574.950 305.850 577.050 307.950 ;
        RECT 577.950 307.050 580.050 309.150 ;
        RECT 595.950 308.850 598.050 310.950 ;
        RECT 613.650 308.850 616.050 310.950 ;
        RECT 617.100 309.150 618.900 310.950 ;
        RECT 556.950 304.950 559.050 305.550 ;
        RECT 565.950 304.950 568.050 305.550 ;
        RECT 569.100 304.050 570.900 305.850 ;
        RECT 527.550 302.700 535.350 303.600 ;
        RECT 514.650 291.750 516.450 297.600 ;
        RECT 517.650 291.750 519.450 297.600 ;
        RECT 527.550 291.750 529.350 302.700 ;
        RECT 530.550 291.750 532.350 301.800 ;
        RECT 533.550 291.750 535.350 302.700 ;
        RECT 536.550 291.750 538.350 303.600 ;
        RECT 553.650 291.750 555.450 303.600 ;
        RECT 556.650 291.750 558.450 303.600 ;
        RECT 571.950 302.850 574.050 304.950 ;
        RECT 575.250 304.050 577.050 305.850 ;
        RECT 572.100 301.050 573.900 302.850 ;
        RECT 578.700 298.800 579.750 307.050 ;
        RECT 596.400 303.600 597.600 308.850 ;
        RECT 613.650 303.600 614.850 308.850 ;
        RECT 616.950 307.050 619.050 309.150 ;
        RECT 572.700 297.900 579.750 298.800 ;
        RECT 572.700 297.600 574.350 297.900 ;
        RECT 569.550 291.750 571.350 297.600 ;
        RECT 572.550 291.750 574.350 297.600 ;
        RECT 578.550 297.600 579.750 297.900 ;
        RECT 575.550 291.750 577.350 297.000 ;
        RECT 578.550 291.750 580.350 297.600 ;
        RECT 593.550 291.750 595.350 303.600 ;
        RECT 596.550 291.750 598.350 303.600 ;
        RECT 613.050 291.750 614.850 303.600 ;
        RECT 616.050 291.750 617.850 303.600 ;
        RECT 620.100 297.600 621.300 314.700 ;
        RECT 622.950 308.850 625.050 310.950 ;
        RECT 635.100 309.150 636.900 310.950 ;
        RECT 623.100 307.050 624.900 308.850 ;
        RECT 634.950 307.050 637.050 309.150 ;
        RECT 638.250 307.950 639.450 315.300 ;
        RECT 653.250 315.300 654.450 317.400 ;
        RECT 655.650 318.300 657.450 323.250 ;
        RECT 658.650 319.200 660.450 323.250 ;
        RECT 661.650 318.300 663.450 323.250 ;
        RECT 655.650 316.950 663.450 318.300 ;
        RECT 671.550 318.300 673.350 323.250 ;
        RECT 674.550 319.200 676.350 323.250 ;
        RECT 677.550 318.300 679.350 323.250 ;
        RECT 671.550 316.950 679.350 318.300 ;
        RECT 680.550 317.400 682.350 323.250 ;
        RECT 692.850 317.400 694.650 323.250 ;
        RECT 680.550 315.300 681.750 317.400 ;
        RECT 697.350 316.200 699.150 323.250 ;
        RECT 710.850 317.400 712.650 323.250 ;
        RECT 715.350 316.200 717.150 323.250 ;
        RECT 733.650 317.400 735.450 323.250 ;
        RECT 653.250 314.250 657.000 315.300 ;
        RECT 678.000 314.250 681.750 315.300 ;
        RECT 695.550 315.300 699.150 316.200 ;
        RECT 713.550 315.300 717.150 316.200 ;
        RECT 734.250 315.300 735.450 317.400 ;
        RECT 736.650 318.300 738.450 323.250 ;
        RECT 739.650 319.200 741.450 323.250 ;
        RECT 742.650 318.300 744.450 323.250 ;
        RECT 736.650 316.950 744.450 318.300 ;
        RECT 754.650 317.400 756.450 323.250 ;
        RECT 755.250 315.300 756.450 317.400 ;
        RECT 757.650 318.300 759.450 323.250 ;
        RECT 760.650 319.200 762.450 323.250 ;
        RECT 763.650 318.300 765.450 323.250 ;
        RECT 773.550 320.400 775.350 323.250 ;
        RECT 776.550 320.400 778.350 323.250 ;
        RECT 788.550 320.400 790.350 323.250 ;
        RECT 791.550 320.400 793.350 323.250 ;
        RECT 794.550 320.400 796.350 323.250 ;
        RECT 757.650 316.950 765.450 318.300 ;
        RECT 655.950 310.950 657.150 314.250 ;
        RECT 659.100 312.150 660.900 313.950 ;
        RECT 674.100 312.150 675.900 313.950 ;
        RECT 641.100 309.150 642.900 310.950 ;
        RECT 637.950 305.850 640.050 307.950 ;
        RECT 640.950 307.050 643.050 309.150 ;
        RECT 655.950 308.850 658.050 310.950 ;
        RECT 658.950 310.050 661.050 312.150 ;
        RECT 661.950 308.850 664.050 310.950 ;
        RECT 670.950 308.850 673.050 310.950 ;
        RECT 673.950 310.050 676.050 312.150 ;
        RECT 677.850 310.950 679.050 314.250 ;
        RECT 676.950 308.850 679.050 310.950 ;
        RECT 692.100 309.150 693.900 310.950 ;
        RECT 652.950 305.850 655.050 307.950 ;
        RECT 638.250 297.600 639.450 305.850 ;
        RECT 653.250 304.050 655.050 305.850 ;
        RECT 656.850 303.600 658.050 308.850 ;
        RECT 662.100 307.050 663.900 308.850 ;
        RECT 671.100 307.050 672.900 308.850 ;
        RECT 676.950 303.600 678.150 308.850 ;
        RECT 679.950 305.850 682.050 307.950 ;
        RECT 691.950 307.050 694.050 309.150 ;
        RECT 695.550 307.950 696.750 315.300 ;
        RECT 698.100 309.150 699.900 310.950 ;
        RECT 710.100 309.150 711.900 310.950 ;
        RECT 694.950 305.850 697.050 307.950 ;
        RECT 697.950 307.050 700.050 309.150 ;
        RECT 709.950 307.050 712.050 309.150 ;
        RECT 713.550 307.950 714.750 315.300 ;
        RECT 734.250 314.250 738.000 315.300 ;
        RECT 755.250 314.250 759.000 315.300 ;
        RECT 736.950 310.950 738.150 314.250 ;
        RECT 740.100 312.150 741.900 313.950 ;
        RECT 716.100 309.150 717.900 310.950 ;
        RECT 712.950 305.850 715.050 307.950 ;
        RECT 715.950 307.050 718.050 309.150 ;
        RECT 736.950 308.850 739.050 310.950 ;
        RECT 739.950 310.050 742.050 312.150 ;
        RECT 757.950 310.950 759.150 314.250 ;
        RECT 761.100 312.150 762.900 313.950 ;
        RECT 742.950 308.850 745.050 310.950 ;
        RECT 757.950 308.850 760.050 310.950 ;
        RECT 760.950 310.050 763.050 312.150 ;
        RECT 772.950 311.850 775.050 313.950 ;
        RECT 776.400 312.150 777.600 320.400 ;
        RECT 792.000 313.950 793.050 320.400 ;
        RECT 806.850 317.400 808.650 323.250 ;
        RECT 811.350 316.200 813.150 323.250 ;
        RECT 824.550 320.400 826.350 323.250 ;
        RECT 827.550 320.400 829.350 323.250 ;
        RECT 841.650 320.400 843.450 323.250 ;
        RECT 844.650 320.400 846.450 323.250 ;
        RECT 763.950 308.850 766.050 310.950 ;
        RECT 773.100 310.050 774.900 311.850 ;
        RECT 775.950 310.050 778.050 312.150 ;
        RECT 790.950 311.850 793.050 313.950 ;
        RECT 733.950 305.850 736.050 307.950 ;
        RECT 679.950 304.050 681.750 305.850 ;
        RECT 619.650 291.750 621.450 297.600 ;
        RECT 622.650 291.750 624.450 297.600 ;
        RECT 634.650 291.750 636.450 297.600 ;
        RECT 637.650 291.750 639.450 297.600 ;
        RECT 640.650 291.750 642.450 297.600 ;
        RECT 653.400 291.750 655.200 297.600 ;
        RECT 656.700 291.750 658.500 303.600 ;
        RECT 660.900 291.750 662.700 303.600 ;
        RECT 672.300 291.750 674.100 303.600 ;
        RECT 676.500 291.750 678.300 303.600 ;
        RECT 695.550 297.600 696.750 305.850 ;
        RECT 713.550 297.600 714.750 305.850 ;
        RECT 734.250 304.050 736.050 305.850 ;
        RECT 737.850 303.600 739.050 308.850 ;
        RECT 743.100 307.050 744.900 308.850 ;
        RECT 754.950 305.850 757.050 307.950 ;
        RECT 755.250 304.050 757.050 305.850 ;
        RECT 758.850 303.600 760.050 308.850 ;
        RECT 764.100 307.050 765.900 308.850 ;
        RECT 679.800 291.750 681.600 297.600 ;
        RECT 692.550 291.750 694.350 297.600 ;
        RECT 695.550 291.750 697.350 297.600 ;
        RECT 698.550 291.750 700.350 297.600 ;
        RECT 710.550 291.750 712.350 297.600 ;
        RECT 713.550 291.750 715.350 297.600 ;
        RECT 716.550 291.750 718.350 297.600 ;
        RECT 734.400 291.750 736.200 297.600 ;
        RECT 737.700 291.750 739.500 303.600 ;
        RECT 741.900 291.750 743.700 303.600 ;
        RECT 755.400 291.750 757.200 297.600 ;
        RECT 758.700 291.750 760.500 303.600 ;
        RECT 762.900 291.750 764.700 303.600 ;
        RECT 776.400 297.600 777.600 310.050 ;
        RECT 787.950 308.850 790.050 310.950 ;
        RECT 788.100 307.050 789.900 308.850 ;
        RECT 792.000 304.650 793.050 311.850 ;
        RECT 809.550 315.300 813.150 316.200 ;
        RECT 793.950 308.850 796.050 310.950 ;
        RECT 806.100 309.150 807.900 310.950 ;
        RECT 794.100 307.050 795.900 308.850 ;
        RECT 805.950 307.050 808.050 309.150 ;
        RECT 809.550 307.950 810.750 315.300 ;
        RECT 823.950 311.850 826.050 313.950 ;
        RECT 827.400 312.150 828.600 320.400 ;
        RECT 842.400 312.150 843.600 320.400 ;
        RECT 854.550 318.300 856.350 323.250 ;
        RECT 857.550 319.200 859.350 323.250 ;
        RECT 860.550 318.300 862.350 323.250 ;
        RECT 854.550 316.950 862.350 318.300 ;
        RECT 863.550 317.400 865.350 323.250 ;
        RECT 863.550 315.300 864.750 317.400 ;
        RECT 861.000 314.250 864.750 315.300 ;
        RECT 812.100 309.150 813.900 310.950 ;
        RECT 824.100 310.050 825.900 311.850 ;
        RECT 826.950 310.050 829.050 312.150 ;
        RECT 841.950 310.050 844.050 312.150 ;
        RECT 844.950 311.850 847.050 313.950 ;
        RECT 857.100 312.150 858.900 313.950 ;
        RECT 845.100 310.050 846.900 311.850 ;
        RECT 808.950 305.850 811.050 307.950 ;
        RECT 811.950 307.050 814.050 309.150 ;
        RECT 792.000 303.600 794.550 304.650 ;
        RECT 773.550 291.750 775.350 297.600 ;
        RECT 776.550 291.750 778.350 297.600 ;
        RECT 788.550 291.750 790.350 303.600 ;
        RECT 792.750 291.750 794.550 303.600 ;
        RECT 809.550 297.600 810.750 305.850 ;
        RECT 827.400 297.600 828.600 310.050 ;
        RECT 842.400 297.600 843.600 310.050 ;
        RECT 853.950 308.850 856.050 310.950 ;
        RECT 856.950 310.050 859.050 312.150 ;
        RECT 860.850 310.950 862.050 314.250 ;
        RECT 859.950 308.850 862.050 310.950 ;
        RECT 854.100 307.050 855.900 308.850 ;
        RECT 859.950 303.600 861.150 308.850 ;
        RECT 862.950 305.850 865.050 307.950 ;
        RECT 862.950 304.050 864.750 305.850 ;
        RECT 806.550 291.750 808.350 297.600 ;
        RECT 809.550 291.750 811.350 297.600 ;
        RECT 812.550 291.750 814.350 297.600 ;
        RECT 824.550 291.750 826.350 297.600 ;
        RECT 827.550 291.750 829.350 297.600 ;
        RECT 841.650 291.750 843.450 297.600 ;
        RECT 844.650 291.750 846.450 297.600 ;
        RECT 855.300 291.750 857.100 303.600 ;
        RECT 859.500 291.750 861.300 303.600 ;
        RECT 862.800 291.750 864.600 297.600 ;
        RECT 10.650 281.400 12.450 287.250 ;
        RECT 13.650 282.000 15.450 287.250 ;
        RECT 11.250 281.100 12.450 281.400 ;
        RECT 16.650 281.400 18.450 287.250 ;
        RECT 19.650 281.400 21.450 287.250 ;
        RECT 16.650 281.100 18.300 281.400 ;
        RECT 11.250 280.200 18.300 281.100 ;
        RECT 11.250 271.950 12.300 280.200 ;
        RECT 17.100 276.150 18.900 277.950 ;
        RECT 29.550 276.300 31.350 287.250 ;
        RECT 32.550 277.200 34.350 287.250 ;
        RECT 35.550 276.300 37.350 287.250 ;
        RECT 13.950 273.150 15.750 274.950 ;
        RECT 16.950 274.050 19.050 276.150 ;
        RECT 29.550 275.400 37.350 276.300 ;
        RECT 38.550 275.400 40.350 287.250 ;
        RECT 53.400 281.400 55.200 287.250 ;
        RECT 56.700 275.400 58.500 287.250 ;
        RECT 60.900 275.400 62.700 287.250 ;
        RECT 73.650 281.400 75.450 287.250 ;
        RECT 76.650 282.000 78.450 287.250 ;
        RECT 74.250 281.100 75.450 281.400 ;
        RECT 79.650 281.400 81.450 287.250 ;
        RECT 82.650 281.400 84.450 287.250 ;
        RECT 79.650 281.100 81.300 281.400 ;
        RECT 74.250 280.200 81.300 281.100 ;
        RECT 20.100 273.150 21.900 274.950 ;
        RECT 10.950 269.850 13.050 271.950 ;
        RECT 13.950 271.050 16.050 273.150 ;
        RECT 19.950 271.050 22.050 273.150 ;
        RECT 38.700 270.150 39.900 275.400 ;
        RECT 53.250 273.150 55.050 274.950 ;
        RECT 52.950 271.050 55.050 273.150 ;
        RECT 56.850 270.150 58.050 275.400 ;
        RECT 74.250 271.950 75.300 280.200 ;
        RECT 80.100 276.150 81.900 277.950 ;
        RECT 76.950 273.150 78.750 274.950 ;
        RECT 79.950 274.050 82.050 276.150 ;
        RECT 99.450 275.400 101.250 287.250 ;
        RECT 103.650 275.400 105.450 287.250 ;
        RECT 113.550 276.300 115.350 287.250 ;
        RECT 116.550 277.200 118.350 287.250 ;
        RECT 119.550 276.300 121.350 287.250 ;
        RECT 113.550 275.400 121.350 276.300 ;
        RECT 122.550 275.400 124.350 287.250 ;
        RECT 139.650 281.400 141.450 287.250 ;
        RECT 142.650 281.400 144.450 287.250 ;
        RECT 158.400 281.400 160.200 287.250 ;
        RECT 83.100 273.150 84.900 274.950 ;
        RECT 99.450 274.350 102.000 275.400 ;
        RECT 62.100 270.150 63.900 271.950 ;
        RECT 11.400 265.650 12.600 269.850 ;
        RECT 28.950 266.850 31.050 268.950 ;
        RECT 32.100 267.150 33.900 268.950 ;
        RECT 11.400 264.000 15.900 265.650 ;
        RECT 29.100 265.050 30.900 266.850 ;
        RECT 31.950 265.050 34.050 267.150 ;
        RECT 34.950 266.850 37.050 268.950 ;
        RECT 37.950 268.050 40.050 270.150 ;
        RECT 55.950 268.050 58.050 270.150 ;
        RECT 35.100 265.050 36.900 266.850 ;
        RECT 14.100 255.750 15.900 264.000 ;
        RECT 19.500 255.750 21.300 264.600 ;
        RECT 38.700 261.600 39.900 268.050 ;
        RECT 55.950 264.750 57.150 268.050 ;
        RECT 58.950 266.850 61.050 268.950 ;
        RECT 61.950 268.050 64.050 270.150 ;
        RECT 73.950 269.850 76.050 271.950 ;
        RECT 76.950 271.050 79.050 273.150 ;
        RECT 82.950 271.050 85.050 273.150 ;
        RECT 98.100 270.150 99.900 271.950 ;
        RECT 59.100 265.050 60.900 266.850 ;
        RECT 74.400 265.650 75.600 269.850 ;
        RECT 97.950 268.050 100.050 270.150 ;
        RECT 100.950 267.150 102.000 274.350 ;
        RECT 118.950 273.450 121.050 274.050 ;
        RECT 110.550 272.550 121.050 273.450 ;
        RECT 104.100 270.150 105.900 271.950 ;
        RECT 103.950 268.050 106.050 270.150 ;
        RECT 53.250 263.700 57.000 264.750 ;
        RECT 74.400 264.000 78.900 265.650 ;
        RECT 100.950 265.050 103.050 267.150 ;
        RECT 53.250 261.600 54.450 263.700 ;
        RECT 30.000 255.750 31.800 261.600 ;
        RECT 34.200 259.950 39.900 261.600 ;
        RECT 34.200 255.750 36.000 259.950 ;
        RECT 37.500 255.750 39.300 258.600 ;
        RECT 52.650 255.750 54.450 261.600 ;
        RECT 55.650 260.700 63.450 262.050 ;
        RECT 55.650 255.750 57.450 260.700 ;
        RECT 58.650 255.750 60.450 259.800 ;
        RECT 61.650 255.750 63.450 260.700 ;
        RECT 77.100 255.750 78.900 264.000 ;
        RECT 82.500 255.750 84.300 264.600 ;
        RECT 100.950 258.600 102.000 265.050 ;
        RECT 103.950 264.450 106.050 265.050 ;
        RECT 110.550 264.450 111.450 272.550 ;
        RECT 118.950 271.950 121.050 272.550 ;
        RECT 122.700 270.150 123.900 275.400 ;
        RECT 112.950 266.850 115.050 268.950 ;
        RECT 116.100 267.150 117.900 268.950 ;
        RECT 113.100 265.050 114.900 266.850 ;
        RECT 115.950 265.050 118.050 267.150 ;
        RECT 118.950 266.850 121.050 268.950 ;
        RECT 121.950 268.050 124.050 270.150 ;
        RECT 140.400 268.950 141.600 281.400 ;
        RECT 161.700 275.400 163.500 287.250 ;
        RECT 165.900 275.400 167.700 287.250 ;
        RECT 179.400 281.400 181.200 287.250 ;
        RECT 182.700 275.400 184.500 287.250 ;
        RECT 186.900 275.400 188.700 287.250 ;
        RECT 199.650 281.400 201.450 287.250 ;
        RECT 202.650 281.400 204.450 287.250 ;
        RECT 215.400 281.400 217.200 287.250 ;
        RECT 158.250 273.150 160.050 274.950 ;
        RECT 157.950 271.050 160.050 273.150 ;
        RECT 161.850 270.150 163.050 275.400 ;
        RECT 179.250 273.150 181.050 274.950 ;
        RECT 167.100 270.150 168.900 271.950 ;
        RECT 178.950 271.050 181.050 273.150 ;
        RECT 182.850 270.150 184.050 275.400 ;
        RECT 188.100 270.150 189.900 271.950 ;
        RECT 119.100 265.050 120.900 266.850 ;
        RECT 103.950 263.550 111.450 264.450 ;
        RECT 103.950 262.950 106.050 263.550 ;
        RECT 122.700 261.600 123.900 268.050 ;
        RECT 139.950 266.850 142.050 268.950 ;
        RECT 143.100 267.150 144.900 268.950 ;
        RECT 160.950 268.050 163.050 270.150 ;
        RECT 97.650 255.750 99.450 258.600 ;
        RECT 100.650 255.750 102.450 258.600 ;
        RECT 103.650 255.750 105.450 258.600 ;
        RECT 114.000 255.750 115.800 261.600 ;
        RECT 118.200 259.950 123.900 261.600 ;
        RECT 118.200 255.750 120.000 259.950 ;
        RECT 140.400 258.600 141.600 266.850 ;
        RECT 142.950 265.050 145.050 267.150 ;
        RECT 160.950 264.750 162.150 268.050 ;
        RECT 163.950 266.850 166.050 268.950 ;
        RECT 166.950 268.050 169.050 270.150 ;
        RECT 181.950 268.050 184.050 270.150 ;
        RECT 164.100 265.050 165.900 266.850 ;
        RECT 181.950 264.750 183.150 268.050 ;
        RECT 184.950 266.850 187.050 268.950 ;
        RECT 187.950 268.050 190.050 270.150 ;
        RECT 200.400 268.950 201.600 281.400 ;
        RECT 218.700 275.400 220.500 287.250 ;
        RECT 222.900 275.400 224.700 287.250 ;
        RECT 234.300 275.400 236.100 287.250 ;
        RECT 238.500 275.400 240.300 287.250 ;
        RECT 241.800 281.400 243.600 287.250 ;
        RECT 257.400 281.400 259.200 287.250 ;
        RECT 260.700 275.400 262.500 287.250 ;
        RECT 264.900 275.400 266.700 287.250 ;
        RECT 277.650 281.400 279.450 287.250 ;
        RECT 280.650 281.400 282.450 287.250 ;
        RECT 283.650 281.400 285.450 287.250 ;
        RECT 295.650 281.400 297.450 287.250 ;
        RECT 298.650 281.400 300.450 287.250 ;
        RECT 301.650 281.400 303.450 287.250 ;
        RECT 215.250 273.150 217.050 274.950 ;
        RECT 214.950 271.050 217.050 273.150 ;
        RECT 218.850 270.150 220.050 275.400 ;
        RECT 224.100 270.150 225.900 271.950 ;
        RECT 233.100 270.150 234.900 271.950 ;
        RECT 238.950 270.150 240.150 275.400 ;
        RECT 241.950 273.150 243.750 274.950 ;
        RECT 257.250 273.150 259.050 274.950 ;
        RECT 241.950 271.050 244.050 273.150 ;
        RECT 256.950 271.050 259.050 273.150 ;
        RECT 260.850 270.150 262.050 275.400 ;
        RECT 281.250 273.150 282.450 281.400 ;
        RECT 299.250 273.150 300.450 281.400 ;
        RECT 316.650 275.400 318.450 287.250 ;
        RECT 319.650 275.400 321.450 287.250 ;
        RECT 322.650 275.400 324.450 287.250 ;
        RECT 327.750 281.400 329.550 287.250 ;
        RECT 330.750 281.400 332.550 287.250 ;
        RECT 334.500 281.400 336.300 287.250 ;
        RECT 337.500 281.400 339.300 287.250 ;
        RECT 340.500 281.400 342.300 287.250 ;
        RECT 266.100 270.150 267.900 271.950 ;
        RECT 199.950 266.850 202.050 268.950 ;
        RECT 203.100 267.150 204.900 268.950 ;
        RECT 217.950 268.050 220.050 270.150 ;
        RECT 185.100 265.050 186.900 266.850 ;
        RECT 158.250 263.700 162.000 264.750 ;
        RECT 179.250 263.700 183.000 264.750 ;
        RECT 158.250 261.600 159.450 263.700 ;
        RECT 121.500 255.750 123.300 258.600 ;
        RECT 139.650 255.750 141.450 258.600 ;
        RECT 142.650 255.750 144.450 258.600 ;
        RECT 157.650 255.750 159.450 261.600 ;
        RECT 160.650 260.700 168.450 262.050 ;
        RECT 179.250 261.600 180.450 263.700 ;
        RECT 160.650 255.750 162.450 260.700 ;
        RECT 163.650 255.750 165.450 259.800 ;
        RECT 166.650 255.750 168.450 260.700 ;
        RECT 178.650 255.750 180.450 261.600 ;
        RECT 181.650 260.700 189.450 262.050 ;
        RECT 181.650 255.750 183.450 260.700 ;
        RECT 184.650 255.750 186.450 259.800 ;
        RECT 187.650 255.750 189.450 260.700 ;
        RECT 200.400 258.600 201.600 266.850 ;
        RECT 202.950 265.050 205.050 267.150 ;
        RECT 217.950 264.750 219.150 268.050 ;
        RECT 220.950 266.850 223.050 268.950 ;
        RECT 223.950 268.050 226.050 270.150 ;
        RECT 232.950 268.050 235.050 270.150 ;
        RECT 235.950 266.850 238.050 268.950 ;
        RECT 238.950 268.050 241.050 270.150 ;
        RECT 221.100 265.050 222.900 266.850 ;
        RECT 236.100 265.050 237.900 266.850 ;
        RECT 239.850 264.750 241.050 268.050 ;
        RECT 259.950 268.050 262.050 270.150 ;
        RECT 259.950 264.750 261.150 268.050 ;
        RECT 262.950 266.850 265.050 268.950 ;
        RECT 265.950 268.050 268.050 270.150 ;
        RECT 277.950 269.850 280.050 271.950 ;
        RECT 280.950 271.050 283.050 273.150 ;
        RECT 278.100 268.050 279.900 269.850 ;
        RECT 263.100 265.050 264.900 266.850 ;
        RECT 215.250 263.700 219.000 264.750 ;
        RECT 240.000 263.700 243.750 264.750 ;
        RECT 215.250 261.600 216.450 263.700 ;
        RECT 199.650 255.750 201.450 258.600 ;
        RECT 202.650 255.750 204.450 258.600 ;
        RECT 214.650 255.750 216.450 261.600 ;
        RECT 217.650 260.700 225.450 262.050 ;
        RECT 217.650 255.750 219.450 260.700 ;
        RECT 220.650 255.750 222.450 259.800 ;
        RECT 223.650 255.750 225.450 260.700 ;
        RECT 233.550 260.700 241.350 262.050 ;
        RECT 233.550 255.750 235.350 260.700 ;
        RECT 236.550 255.750 238.350 259.800 ;
        RECT 239.550 255.750 241.350 260.700 ;
        RECT 242.550 261.600 243.750 263.700 ;
        RECT 257.250 263.700 261.000 264.750 ;
        RECT 281.250 263.700 282.450 271.050 ;
        RECT 283.950 269.850 286.050 271.950 ;
        RECT 295.950 269.850 298.050 271.950 ;
        RECT 298.950 271.050 301.050 273.150 ;
        RECT 284.100 268.050 285.900 269.850 ;
        RECT 296.100 268.050 297.900 269.850 ;
        RECT 299.250 263.700 300.450 271.050 ;
        RECT 301.950 269.850 304.050 271.950 ;
        RECT 302.100 268.050 303.900 269.850 ;
        RECT 319.800 268.950 321.150 275.400 ;
        RECT 331.050 268.950 332.550 281.400 ;
        RECT 337.500 277.350 338.700 281.400 ;
        RECT 343.500 280.500 345.300 287.250 ;
        RECT 346.500 281.400 348.300 287.250 ;
        RECT 350.250 284.400 352.050 287.250 ;
        RECT 350.400 283.200 351.900 284.400 ;
        RECT 349.800 281.100 351.900 283.200 ;
        RECT 353.250 280.950 355.050 287.250 ;
        RECT 356.250 284.400 358.050 287.250 ;
        RECT 339.600 279.300 345.300 280.500 ;
        RECT 346.350 280.050 348.150 280.500 ;
        RECT 352.950 280.050 355.050 280.950 ;
        RECT 339.600 278.700 341.400 279.300 ;
        RECT 346.350 278.850 355.050 280.050 ;
        RECT 346.350 278.700 348.150 278.850 ;
        RECT 356.550 277.350 357.900 284.400 ;
        RECT 360.000 280.500 361.800 287.250 ;
        RECT 363.000 281.400 364.800 287.250 ;
        RECT 366.000 281.400 367.800 287.250 ;
        RECT 369.750 281.400 371.550 287.250 ;
        RECT 372.750 284.400 374.700 287.250 ;
        RECT 375.750 284.400 377.850 287.250 ;
        RECT 378.750 284.400 381.150 287.250 ;
        RECT 373.500 283.050 374.700 284.400 ;
        RECT 376.950 283.050 377.850 284.400 ;
        RECT 379.950 283.050 381.150 284.400 ;
        RECT 382.500 283.950 384.300 287.250 ;
        RECT 373.500 281.400 376.050 283.050 ;
        RECT 366.000 280.500 367.350 281.400 ;
        RECT 373.950 280.950 376.050 281.400 ;
        RECT 376.950 280.950 379.050 283.050 ;
        RECT 379.950 280.950 382.050 283.050 ;
        RECT 360.000 280.200 363.000 280.500 ;
        RECT 359.100 278.400 363.000 280.200 ;
        RECT 364.950 278.850 367.350 280.500 ;
        RECT 364.950 278.400 367.050 278.850 ;
        RECT 385.500 278.700 387.300 287.250 ;
        RECT 388.500 281.400 390.300 287.250 ;
        RECT 391.500 281.400 393.300 287.250 ;
        RECT 394.500 281.400 396.300 287.250 ;
        RECT 404.550 281.400 406.350 287.250 ;
        RECT 407.550 281.400 409.350 287.250 ;
        RECT 410.550 281.400 412.350 287.250 ;
        RECT 424.650 281.400 426.450 287.250 ;
        RECT 427.650 282.000 429.450 287.250 ;
        RECT 392.250 280.500 393.300 281.400 ;
        RECT 392.250 279.600 396.300 280.500 ;
        RECT 374.100 277.650 391.800 278.700 ;
        RECT 316.950 266.850 321.150 268.950 ;
        RECT 322.950 266.850 325.050 268.950 ;
        RECT 328.950 266.850 332.550 268.950 ;
        RECT 257.250 261.600 258.450 263.700 ;
        RECT 278.850 262.800 282.450 263.700 ;
        RECT 296.850 262.800 300.450 263.700 ;
        RECT 242.550 255.750 244.350 261.600 ;
        RECT 256.650 255.750 258.450 261.600 ;
        RECT 259.650 260.700 267.450 262.050 ;
        RECT 259.650 255.750 261.450 260.700 ;
        RECT 262.650 255.750 264.450 259.800 ;
        RECT 265.650 255.750 267.450 260.700 ;
        RECT 278.850 255.750 280.650 262.800 ;
        RECT 283.350 255.750 285.150 261.600 ;
        RECT 296.850 255.750 298.650 262.800 ;
        RECT 319.800 261.600 321.150 266.850 ;
        RECT 323.100 265.050 324.900 266.850 ;
        RECT 301.350 255.750 303.150 261.600 ;
        RECT 316.650 255.750 318.450 261.600 ;
        RECT 319.650 255.750 321.450 261.600 ;
        RECT 322.650 255.750 324.450 261.600 ;
        RECT 331.050 258.600 332.550 266.850 ;
        RECT 327.750 255.750 329.550 258.600 ;
        RECT 330.750 255.750 332.550 258.600 ;
        RECT 334.650 276.450 352.050 277.350 ;
        RECT 334.650 261.600 335.850 276.450 ;
        RECT 336.750 274.350 349.050 275.550 ;
        RECT 349.950 275.250 352.050 276.450 ;
        RECT 355.950 276.600 358.050 277.350 ;
        RECT 374.100 276.600 376.050 277.650 ;
        RECT 390.000 276.900 391.800 277.650 ;
        RECT 355.950 275.250 376.050 276.600 ;
        RECT 376.950 276.150 379.050 276.750 ;
        RECT 376.950 274.950 388.500 276.150 ;
        RECT 376.950 274.650 379.050 274.950 ;
        RECT 386.700 274.350 388.500 274.950 ;
        RECT 336.750 273.750 338.550 274.350 ;
        RECT 348.000 273.450 376.050 274.350 ;
        RECT 348.000 273.150 387.750 273.450 ;
        RECT 340.950 269.100 343.050 273.150 ;
        RECT 374.100 272.550 388.050 273.150 ;
        RECT 344.100 270.000 351.150 271.800 ;
        RECT 340.950 268.050 349.200 269.100 ;
        RECT 336.900 265.200 344.700 267.000 ;
        RECT 348.150 266.250 349.200 268.050 ;
        RECT 350.250 268.350 351.150 270.000 ;
        RECT 352.500 271.650 367.050 272.250 ;
        RECT 352.500 271.050 375.600 271.650 ;
        RECT 384.150 271.350 388.050 272.550 ;
        RECT 352.500 269.250 354.300 271.050 ;
        RECT 364.950 270.450 375.600 271.050 ;
        RECT 364.950 270.150 367.050 270.450 ;
        RECT 373.800 269.850 375.600 270.450 ;
        RECT 376.500 270.450 383.250 271.350 ;
        RECT 385.950 271.050 388.050 271.350 ;
        RECT 360.750 269.250 362.850 269.550 ;
        RECT 350.250 267.300 359.850 268.350 ;
        RECT 360.750 267.450 364.650 269.250 ;
        RECT 376.500 268.950 377.550 270.450 ;
        RECT 365.550 268.050 377.550 268.950 ;
        RECT 358.950 266.550 359.850 267.300 ;
        RECT 365.550 266.550 366.600 268.050 ;
        RECT 378.450 267.750 380.250 269.550 ;
        RECT 382.050 268.050 383.250 270.450 ;
        RECT 391.950 269.850 394.050 271.950 ;
        RECT 392.100 268.050 393.900 269.850 ;
        RECT 348.150 265.200 358.050 266.250 ;
        RECT 358.950 265.200 366.600 266.550 ;
        RECT 367.950 265.350 371.850 267.150 ;
        RECT 343.200 261.600 344.700 265.200 ;
        RECT 357.000 264.300 358.050 265.200 ;
        RECT 367.950 265.050 370.050 265.350 ;
        RECT 375.150 264.300 376.950 264.750 ;
        RECT 378.450 264.300 379.500 267.750 ;
        RECT 382.050 267.000 393.900 268.050 ;
        RECT 395.100 266.100 396.300 279.600 ;
        RECT 407.550 273.150 408.750 281.400 ;
        RECT 425.250 281.100 426.450 281.400 ;
        RECT 430.650 281.400 432.450 287.250 ;
        RECT 433.650 281.400 435.450 287.250 ;
        RECT 446.400 281.400 448.200 287.250 ;
        RECT 430.650 281.100 432.300 281.400 ;
        RECT 425.250 280.200 432.300 281.100 ;
        RECT 403.950 269.850 406.050 271.950 ;
        RECT 406.950 271.050 409.050 273.150 ;
        RECT 425.250 271.950 426.300 280.200 ;
        RECT 431.100 276.150 432.900 277.950 ;
        RECT 427.950 273.150 429.750 274.950 ;
        RECT 430.950 274.050 433.050 276.150 ;
        RECT 449.700 275.400 451.500 287.250 ;
        RECT 453.900 275.400 455.700 287.250 ;
        RECT 464.550 275.400 466.350 287.250 ;
        RECT 468.750 275.400 470.550 287.250 ;
        RECT 482.550 280.200 484.350 286.200 ;
        RECT 485.550 280.200 487.350 287.250 ;
        RECT 434.100 273.150 435.900 274.950 ;
        RECT 446.250 273.150 448.050 274.950 ;
        RECT 404.100 268.050 405.900 269.850 ;
        RECT 349.350 262.500 356.100 264.300 ;
        RECT 357.000 262.500 363.900 264.300 ;
        RECT 375.150 263.850 379.500 264.300 ;
        RECT 371.850 263.100 379.500 263.850 ;
        RECT 381.000 265.200 396.300 266.100 ;
        RECT 371.850 262.950 376.950 263.100 ;
        RECT 371.850 261.600 372.750 262.950 ;
        RECT 381.000 262.050 382.050 265.200 ;
        RECT 390.300 263.700 392.100 264.300 ;
        RECT 334.650 255.750 336.450 261.600 ;
        RECT 340.050 255.750 341.850 261.600 ;
        RECT 343.200 260.400 347.400 261.600 ;
        RECT 345.600 255.750 347.400 260.400 ;
        RECT 349.950 259.500 352.050 261.600 ;
        RECT 352.950 259.500 355.050 261.600 ;
        RECT 355.950 259.500 358.050 261.600 ;
        RECT 360.750 261.300 362.850 261.600 ;
        RECT 350.250 255.750 352.050 259.500 ;
        RECT 353.250 255.750 355.050 259.500 ;
        RECT 356.250 255.750 358.050 259.500 ;
        RECT 360.000 259.500 362.850 261.300 ;
        RECT 364.950 261.300 367.050 261.600 ;
        RECT 364.950 259.500 367.800 261.300 ;
        RECT 368.700 260.250 372.750 261.600 ;
        RECT 368.700 259.800 370.500 260.250 ;
        RECT 373.950 259.950 376.050 262.050 ;
        RECT 376.950 259.950 379.050 262.050 ;
        RECT 379.950 259.950 382.050 262.050 ;
        RECT 383.700 262.500 392.100 263.700 ;
        RECT 383.700 261.600 385.200 262.500 ;
        RECT 395.100 261.600 396.300 265.200 ;
        RECT 407.550 263.700 408.750 271.050 ;
        RECT 409.950 269.850 412.050 271.950 ;
        RECT 424.950 269.850 427.050 271.950 ;
        RECT 427.950 271.050 430.050 273.150 ;
        RECT 433.950 271.050 436.050 273.150 ;
        RECT 445.950 271.050 448.050 273.150 ;
        RECT 449.850 270.150 451.050 275.400 ;
        RECT 468.000 274.350 470.550 275.400 ;
        RECT 483.450 275.100 484.350 280.200 ;
        RECT 490.050 276.900 491.850 286.200 ;
        RECT 490.050 276.000 492.150 276.900 ;
        RECT 455.100 270.150 456.900 271.950 ;
        RECT 464.100 270.150 465.900 271.950 ;
        RECT 410.100 268.050 411.900 269.850 ;
        RECT 425.400 265.650 426.600 269.850 ;
        RECT 448.950 268.050 451.050 270.150 ;
        RECT 425.400 264.000 429.900 265.650 ;
        RECT 448.950 264.750 450.150 268.050 ;
        RECT 451.950 266.850 454.050 268.950 ;
        RECT 454.950 268.050 457.050 270.150 ;
        RECT 463.950 268.050 466.050 270.150 ;
        RECT 468.000 267.150 469.050 274.350 ;
        RECT 483.450 274.200 489.600 275.100 ;
        RECT 470.100 270.150 471.900 271.950 ;
        RECT 485.250 270.150 487.050 271.950 ;
        RECT 469.950 268.050 472.050 270.150 ;
        RECT 452.100 265.050 453.900 266.850 ;
        RECT 466.950 265.050 469.050 267.150 ;
        RECT 481.950 266.850 484.050 268.950 ;
        RECT 484.950 268.050 487.050 270.150 ;
        RECT 488.250 271.500 489.600 274.200 ;
        RECT 488.250 269.700 490.050 271.500 ;
        RECT 482.250 265.050 484.050 266.850 ;
        RECT 407.550 262.800 411.150 263.700 ;
        RECT 360.000 255.750 361.800 259.500 ;
        RECT 363.000 255.750 364.800 258.600 ;
        RECT 366.000 255.750 367.800 259.500 ;
        RECT 373.950 258.600 375.300 259.950 ;
        RECT 376.950 258.600 378.300 259.950 ;
        RECT 379.950 258.600 381.300 259.950 ;
        RECT 370.500 255.750 372.300 258.600 ;
        RECT 373.500 255.750 375.300 258.600 ;
        RECT 376.500 255.750 378.300 258.600 ;
        RECT 379.500 255.750 381.300 258.600 ;
        RECT 383.700 255.750 385.500 261.600 ;
        RECT 389.100 255.750 390.900 261.600 ;
        RECT 394.500 255.750 396.300 261.600 ;
        RECT 404.850 255.750 406.650 261.600 ;
        RECT 409.350 255.750 411.150 262.800 ;
        RECT 428.100 255.750 429.900 264.000 ;
        RECT 433.500 255.750 435.300 264.600 ;
        RECT 446.250 263.700 450.000 264.750 ;
        RECT 446.250 261.600 447.450 263.700 ;
        RECT 445.650 255.750 447.450 261.600 ;
        RECT 448.650 260.700 456.450 262.050 ;
        RECT 448.650 255.750 450.450 260.700 ;
        RECT 451.650 255.750 453.450 259.800 ;
        RECT 454.650 255.750 456.450 260.700 ;
        RECT 468.000 258.600 469.050 265.050 ;
        RECT 488.250 264.000 489.600 269.700 ;
        RECT 491.250 268.950 492.150 276.000 ;
        RECT 494.550 275.400 496.350 287.250 ;
        RECT 508.650 281.400 510.450 287.250 ;
        RECT 511.650 281.400 513.450 287.250 ;
        RECT 494.100 270.150 495.900 271.950 ;
        RECT 490.950 266.850 493.050 268.950 ;
        RECT 493.950 268.050 496.050 270.150 ;
        RECT 509.400 268.950 510.600 281.400 ;
        RECT 521.550 275.400 523.350 287.250 ;
        RECT 526.050 275.400 529.350 287.250 ;
        RECT 532.050 275.400 533.850 287.250 ;
        RECT 548.400 281.400 550.200 287.250 ;
        RECT 551.700 275.400 553.500 287.250 ;
        RECT 555.900 275.400 557.700 287.250 ;
        RECT 572.400 281.400 574.200 287.250 ;
        RECT 575.700 275.400 577.500 287.250 ;
        RECT 579.900 275.400 581.700 287.250 ;
        RECT 591.300 275.400 593.100 287.250 ;
        RECT 595.500 275.400 597.300 287.250 ;
        RECT 598.800 281.400 600.600 287.250 ;
        RECT 613.650 281.400 615.450 287.250 ;
        RECT 616.650 281.400 618.450 287.250 ;
        RECT 619.650 281.400 621.450 287.250 ;
        RECT 631.650 286.500 639.450 287.250 ;
        RECT 521.100 270.150 522.900 271.950 ;
        RECT 527.550 270.150 528.750 275.400 ;
        RECT 548.250 273.150 550.050 274.950 ;
        RECT 532.950 270.150 534.750 271.950 ;
        RECT 547.950 271.050 550.050 273.150 ;
        RECT 551.850 270.150 553.050 275.400 ;
        RECT 572.250 273.150 574.050 274.950 ;
        RECT 557.100 270.150 558.900 271.950 ;
        RECT 571.950 271.050 574.050 273.150 ;
        RECT 575.850 270.150 577.050 275.400 ;
        RECT 586.950 271.950 589.050 274.050 ;
        RECT 581.100 270.150 582.900 271.950 ;
        RECT 508.950 266.850 511.050 268.950 ;
        RECT 512.100 267.150 513.900 268.950 ;
        RECT 520.950 268.050 523.050 270.150 ;
        RECT 483.300 263.100 489.600 264.000 ;
        RECT 483.300 259.800 484.350 263.100 ;
        RECT 491.250 262.200 492.150 266.850 ;
        RECT 490.050 261.300 492.150 262.200 ;
        RECT 464.550 255.750 466.350 258.600 ;
        RECT 467.550 255.750 469.350 258.600 ;
        RECT 470.550 255.750 472.350 258.600 ;
        RECT 482.550 256.800 484.350 259.800 ;
        RECT 485.550 255.750 487.350 259.800 ;
        RECT 490.050 256.800 491.850 261.300 ;
        RECT 494.550 255.750 496.350 262.800 ;
        RECT 509.400 258.600 510.600 266.850 ;
        RECT 511.950 265.050 514.050 267.150 ;
        RECT 523.950 266.850 526.050 268.950 ;
        RECT 526.950 268.050 529.050 270.150 ;
        RECT 524.100 265.050 525.900 266.850 ;
        RECT 527.400 264.150 528.600 268.050 ;
        RECT 529.950 266.850 532.050 268.950 ;
        RECT 532.950 268.050 535.050 270.150 ;
        RECT 550.950 268.050 553.050 270.150 ;
        RECT 529.500 265.050 531.300 266.850 ;
        RECT 550.950 264.750 552.150 268.050 ;
        RECT 553.950 266.850 556.050 268.950 ;
        RECT 556.950 268.050 559.050 270.150 ;
        RECT 574.950 268.050 577.050 270.150 ;
        RECT 554.100 265.050 555.900 266.850 ;
        RECT 574.950 264.750 576.150 268.050 ;
        RECT 577.950 266.850 580.050 268.950 ;
        RECT 580.950 268.050 583.050 270.150 ;
        RECT 578.100 265.050 579.900 266.850 ;
        RECT 527.400 263.100 531.750 264.150 ;
        RECT 521.550 261.000 529.350 261.900 ;
        RECT 530.850 261.600 531.750 263.100 ;
        RECT 548.250 263.700 552.000 264.750 ;
        RECT 572.250 263.700 576.000 264.750 ;
        RECT 580.950 264.450 583.050 265.050 ;
        RECT 587.550 264.450 588.450 271.950 ;
        RECT 590.100 270.150 591.900 271.950 ;
        RECT 595.950 270.150 597.150 275.400 ;
        RECT 598.950 273.150 600.750 274.950 ;
        RECT 617.250 273.150 618.450 281.400 ;
        RECT 631.650 275.400 633.450 286.500 ;
        RECT 634.650 275.400 636.450 285.600 ;
        RECT 637.650 276.600 639.450 286.500 ;
        RECT 640.650 277.500 642.450 287.250 ;
        RECT 643.650 276.600 645.450 287.250 ;
        RECT 655.650 281.400 657.450 287.250 ;
        RECT 658.650 281.400 660.450 287.250 ;
        RECT 661.650 281.400 663.450 287.250 ;
        RECT 637.650 275.700 645.450 276.600 ;
        RECT 655.950 276.450 658.050 277.050 ;
        RECT 653.550 275.550 658.050 276.450 ;
        RECT 634.800 274.500 636.600 275.400 ;
        RECT 634.800 273.600 638.850 274.500 ;
        RECT 598.950 271.050 601.050 273.150 ;
        RECT 589.950 268.050 592.050 270.150 ;
        RECT 592.950 266.850 595.050 268.950 ;
        RECT 595.950 268.050 598.050 270.150 ;
        RECT 613.950 269.850 616.050 271.950 ;
        RECT 616.950 271.050 619.050 273.150 ;
        RECT 614.100 268.050 615.900 269.850 ;
        RECT 593.100 265.050 594.900 266.850 ;
        RECT 596.850 264.750 598.050 268.050 ;
        RECT 548.250 261.600 549.450 263.700 ;
        RECT 508.650 255.750 510.450 258.600 ;
        RECT 511.650 255.750 513.450 258.600 ;
        RECT 521.550 255.750 523.350 261.000 ;
        RECT 524.550 255.750 526.350 260.100 ;
        RECT 527.550 256.500 529.350 261.000 ;
        RECT 530.550 257.400 532.350 261.600 ;
        RECT 533.550 256.500 535.350 261.600 ;
        RECT 527.550 255.750 535.350 256.500 ;
        RECT 547.650 255.750 549.450 261.600 ;
        RECT 550.650 260.700 558.450 262.050 ;
        RECT 572.250 261.600 573.450 263.700 ;
        RECT 580.950 263.550 588.450 264.450 ;
        RECT 597.000 263.700 600.750 264.750 ;
        RECT 617.250 263.700 618.450 271.050 ;
        RECT 619.950 269.850 622.050 271.950 ;
        RECT 632.100 270.150 633.900 271.950 ;
        RECT 637.950 270.150 638.850 273.600 ;
        RECT 653.550 273.450 654.450 275.550 ;
        RECT 655.950 274.950 658.050 275.550 ;
        RECT 650.550 272.550 654.450 273.450 ;
        RECT 659.250 273.150 660.450 281.400 ;
        RECT 672.300 275.400 674.100 287.250 ;
        RECT 676.500 275.400 678.300 287.250 ;
        RECT 679.800 281.400 681.600 287.250 ;
        RECT 694.050 275.400 695.850 287.250 ;
        RECT 697.050 275.400 698.850 287.250 ;
        RECT 700.650 281.400 702.450 287.250 ;
        RECT 703.650 281.400 705.450 287.250 ;
        RECT 643.950 270.150 645.750 271.950 ;
        RECT 620.100 268.050 621.900 269.850 ;
        RECT 631.950 268.050 634.050 270.150 ;
        RECT 634.950 266.850 637.050 268.950 ;
        RECT 637.950 268.050 640.050 270.150 ;
        RECT 635.250 265.050 637.050 266.850 ;
        RECT 580.950 262.950 583.050 263.550 ;
        RECT 550.650 255.750 552.450 260.700 ;
        RECT 553.650 255.750 555.450 259.800 ;
        RECT 556.650 255.750 558.450 260.700 ;
        RECT 571.650 255.750 573.450 261.600 ;
        RECT 574.650 260.700 582.450 262.050 ;
        RECT 574.650 255.750 576.450 260.700 ;
        RECT 577.650 255.750 579.450 259.800 ;
        RECT 580.650 255.750 582.450 260.700 ;
        RECT 590.550 260.700 598.350 262.050 ;
        RECT 590.550 255.750 592.350 260.700 ;
        RECT 593.550 255.750 595.350 259.800 ;
        RECT 596.550 255.750 598.350 260.700 ;
        RECT 599.550 261.600 600.750 263.700 ;
        RECT 614.850 262.800 618.450 263.700 ;
        RECT 599.550 255.750 601.350 261.600 ;
        RECT 614.850 255.750 616.650 262.800 ;
        RECT 639.000 261.600 640.050 268.050 ;
        RECT 640.950 266.850 643.050 268.950 ;
        RECT 643.950 268.050 646.050 270.150 ;
        RECT 640.950 265.050 642.750 266.850 ;
        RECT 619.350 255.750 621.150 261.600 ;
        RECT 634.800 255.750 636.600 261.600 ;
        RECT 639.000 255.750 640.800 261.600 ;
        RECT 643.200 255.750 645.000 261.600 ;
        RECT 650.550 259.050 651.450 272.550 ;
        RECT 655.950 269.850 658.050 271.950 ;
        RECT 658.950 271.050 661.050 273.150 ;
        RECT 656.100 268.050 657.900 269.850 ;
        RECT 659.250 263.700 660.450 271.050 ;
        RECT 661.950 269.850 664.050 271.950 ;
        RECT 671.100 270.150 672.900 271.950 ;
        RECT 676.950 270.150 678.150 275.400 ;
        RECT 679.950 273.150 681.750 274.950 ;
        RECT 679.950 271.050 682.050 273.150 ;
        RECT 694.650 270.150 695.850 275.400 ;
        RECT 662.100 268.050 663.900 269.850 ;
        RECT 670.950 268.050 673.050 270.150 ;
        RECT 673.950 266.850 676.050 268.950 ;
        RECT 676.950 268.050 679.050 270.150 ;
        RECT 674.100 265.050 675.900 266.850 ;
        RECT 677.850 264.750 679.050 268.050 ;
        RECT 694.650 268.050 697.050 270.150 ;
        RECT 697.950 269.850 700.050 271.950 ;
        RECT 698.100 268.050 699.900 269.850 ;
        RECT 678.000 263.700 681.750 264.750 ;
        RECT 656.850 262.800 660.450 263.700 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 656.850 255.750 658.650 262.800 ;
        RECT 661.350 255.750 663.150 261.600 ;
        RECT 671.550 260.700 679.350 262.050 ;
        RECT 671.550 255.750 673.350 260.700 ;
        RECT 674.550 255.750 676.350 259.800 ;
        RECT 677.550 255.750 679.350 260.700 ;
        RECT 680.550 261.600 681.750 263.700 ;
        RECT 694.650 261.600 695.850 268.050 ;
        RECT 701.100 264.300 702.300 281.400 ;
        RECT 717.450 275.400 719.250 287.250 ;
        RECT 721.650 275.400 723.450 287.250 ;
        RECT 733.650 281.400 735.450 287.250 ;
        RECT 736.650 281.400 738.450 287.250 ;
        RECT 739.650 281.400 741.450 287.250 ;
        RECT 751.650 286.500 759.450 287.250 ;
        RECT 717.450 274.350 720.000 275.400 ;
        RECT 704.100 270.150 705.900 271.950 ;
        RECT 716.100 270.150 717.900 271.950 ;
        RECT 703.950 268.050 706.050 270.150 ;
        RECT 715.950 268.050 718.050 270.150 ;
        RECT 718.950 267.150 720.000 274.350 ;
        RECT 737.250 273.150 738.450 281.400 ;
        RECT 751.650 275.400 753.450 286.500 ;
        RECT 754.650 275.400 756.450 285.600 ;
        RECT 757.650 276.600 759.450 286.500 ;
        RECT 760.650 277.500 762.450 287.250 ;
        RECT 763.650 276.600 765.450 287.250 ;
        RECT 775.650 281.400 777.450 287.250 ;
        RECT 778.650 281.400 780.450 287.250 ;
        RECT 757.650 275.700 765.450 276.600 ;
        RECT 754.800 274.500 756.600 275.400 ;
        RECT 754.800 273.600 758.850 274.500 ;
        RECT 722.100 270.150 723.900 271.950 ;
        RECT 721.950 268.050 724.050 270.150 ;
        RECT 733.950 269.850 736.050 271.950 ;
        RECT 736.950 271.050 739.050 273.150 ;
        RECT 734.100 268.050 735.900 269.850 ;
        RECT 718.950 265.050 721.050 267.150 ;
        RECT 697.950 263.100 705.450 264.300 ;
        RECT 697.950 262.500 699.750 263.100 ;
        RECT 680.550 255.750 682.350 261.600 ;
        RECT 694.650 260.100 697.950 261.600 ;
        RECT 696.150 255.750 697.950 260.100 ;
        RECT 699.150 255.750 700.950 261.600 ;
        RECT 703.650 255.750 705.450 263.100 ;
        RECT 718.950 258.600 720.000 265.050 ;
        RECT 737.250 263.700 738.450 271.050 ;
        RECT 739.950 269.850 742.050 271.950 ;
        RECT 752.100 270.150 753.900 271.950 ;
        RECT 757.950 270.150 758.850 273.600 ;
        RECT 763.950 270.150 765.750 271.950 ;
        RECT 740.100 268.050 741.900 269.850 ;
        RECT 751.950 268.050 754.050 270.150 ;
        RECT 754.950 266.850 757.050 268.950 ;
        RECT 757.950 268.050 760.050 270.150 ;
        RECT 755.250 265.050 757.050 266.850 ;
        RECT 734.850 262.800 738.450 263.700 ;
        RECT 715.650 255.750 717.450 258.600 ;
        RECT 718.650 255.750 720.450 258.600 ;
        RECT 721.650 255.750 723.450 258.600 ;
        RECT 734.850 255.750 736.650 262.800 ;
        RECT 759.000 261.600 760.050 268.050 ;
        RECT 760.950 266.850 763.050 268.950 ;
        RECT 763.950 268.050 766.050 270.150 ;
        RECT 776.400 268.950 777.600 281.400 ;
        RECT 792.450 275.400 794.250 287.250 ;
        RECT 796.650 275.400 798.450 287.250 ;
        RECT 792.450 274.350 795.000 275.400 ;
        RECT 802.950 274.950 805.050 277.050 ;
        RECT 807.300 275.400 809.100 287.250 ;
        RECT 811.500 275.400 813.300 287.250 ;
        RECT 814.800 281.400 816.600 287.250 ;
        RECT 830.400 281.400 832.200 287.250 ;
        RECT 833.700 275.400 835.500 287.250 ;
        RECT 837.900 275.400 839.700 287.250 ;
        RECT 848.550 275.400 850.350 287.250 ;
        RECT 851.550 275.400 853.350 287.250 ;
        RECT 854.550 275.400 856.350 287.250 ;
        RECT 791.100 270.150 792.900 271.950 ;
        RECT 775.950 266.850 778.050 268.950 ;
        RECT 779.100 267.150 780.900 268.950 ;
        RECT 790.950 268.050 793.050 270.150 ;
        RECT 793.950 267.150 795.000 274.350 ;
        RECT 797.100 270.150 798.900 271.950 ;
        RECT 796.950 268.050 799.050 270.150 ;
        RECT 760.950 265.050 762.750 266.850 ;
        RECT 739.350 255.750 741.150 261.600 ;
        RECT 754.800 255.750 756.600 261.600 ;
        RECT 759.000 255.750 760.800 261.600 ;
        RECT 763.200 255.750 765.000 261.600 ;
        RECT 776.400 258.600 777.600 266.850 ;
        RECT 778.950 265.050 781.050 267.150 ;
        RECT 793.950 265.050 796.050 267.150 ;
        RECT 793.950 258.600 795.000 265.050 ;
        RECT 796.950 261.450 799.050 262.050 ;
        RECT 803.550 261.450 804.450 274.950 ;
        RECT 806.100 270.150 807.900 271.950 ;
        RECT 811.950 270.150 813.150 275.400 ;
        RECT 814.950 273.150 816.750 274.950 ;
        RECT 830.250 273.150 832.050 274.950 ;
        RECT 814.950 271.050 817.050 273.150 ;
        RECT 829.950 271.050 832.050 273.150 ;
        RECT 833.850 270.150 835.050 275.400 ;
        RECT 839.100 270.150 840.900 271.950 ;
        RECT 805.950 268.050 808.050 270.150 ;
        RECT 808.950 266.850 811.050 268.950 ;
        RECT 811.950 268.050 814.050 270.150 ;
        RECT 809.100 265.050 810.900 266.850 ;
        RECT 812.850 264.750 814.050 268.050 ;
        RECT 832.950 268.050 835.050 270.150 ;
        RECT 832.950 264.750 834.150 268.050 ;
        RECT 835.950 266.850 838.050 268.950 ;
        RECT 838.950 268.050 841.050 270.150 ;
        RECT 851.850 268.950 853.200 275.400 ;
        RECT 847.950 266.850 850.050 268.950 ;
        RECT 851.850 266.850 856.050 268.950 ;
        RECT 836.100 265.050 837.900 266.850 ;
        RECT 848.100 265.050 849.900 266.850 ;
        RECT 813.000 263.700 816.750 264.750 ;
        RECT 796.950 260.550 804.450 261.450 ;
        RECT 806.550 260.700 814.350 262.050 ;
        RECT 796.950 259.950 799.050 260.550 ;
        RECT 775.650 255.750 777.450 258.600 ;
        RECT 778.650 255.750 780.450 258.600 ;
        RECT 790.650 255.750 792.450 258.600 ;
        RECT 793.650 255.750 795.450 258.600 ;
        RECT 796.650 255.750 798.450 258.600 ;
        RECT 806.550 255.750 808.350 260.700 ;
        RECT 809.550 255.750 811.350 259.800 ;
        RECT 812.550 255.750 814.350 260.700 ;
        RECT 815.550 261.600 816.750 263.700 ;
        RECT 830.250 263.700 834.000 264.750 ;
        RECT 830.250 261.600 831.450 263.700 ;
        RECT 815.550 255.750 817.350 261.600 ;
        RECT 829.650 255.750 831.450 261.600 ;
        RECT 832.650 260.700 840.450 262.050 ;
        RECT 851.850 261.600 853.200 266.850 ;
        RECT 832.650 255.750 834.450 260.700 ;
        RECT 835.650 255.750 837.450 259.800 ;
        RECT 838.650 255.750 840.450 260.700 ;
        RECT 848.550 255.750 850.350 261.600 ;
        RECT 851.550 255.750 853.350 261.600 ;
        RECT 854.550 255.750 856.350 261.600 ;
        RECT 11.700 242.400 13.500 251.250 ;
        RECT 17.100 243.000 18.900 251.250 ;
        RECT 38.100 243.000 39.900 251.250 ;
        RECT 17.100 241.350 21.600 243.000 ;
        RECT 20.400 237.150 21.600 241.350 ;
        RECT 35.400 241.350 39.900 243.000 ;
        RECT 43.500 242.400 45.300 251.250 ;
        RECT 54.000 245.400 55.800 251.250 ;
        RECT 58.200 247.050 60.000 251.250 ;
        RECT 61.500 248.400 63.300 251.250 ;
        RECT 77.700 248.400 79.500 251.250 ;
        RECT 81.000 247.050 82.800 251.250 ;
        RECT 58.200 245.400 63.900 247.050 ;
        RECT 35.400 237.150 36.600 241.350 ;
        RECT 53.100 240.150 54.900 241.950 ;
        RECT 52.950 238.050 55.050 240.150 ;
        RECT 55.950 239.850 58.050 241.950 ;
        RECT 59.100 240.150 60.900 241.950 ;
        RECT 56.100 238.050 57.900 239.850 ;
        RECT 58.950 238.050 61.050 240.150 ;
        RECT 62.700 238.950 63.900 245.400 ;
        RECT 77.100 245.400 82.800 247.050 ;
        RECT 85.200 245.400 87.000 251.250 ;
        RECT 95.850 245.400 97.650 251.250 ;
        RECT 77.100 238.950 78.300 245.400 ;
        RECT 100.350 244.200 102.150 251.250 ;
        RECT 113.550 248.400 115.350 251.250 ;
        RECT 116.550 248.400 118.350 251.250 ;
        RECT 98.550 243.300 102.150 244.200 ;
        RECT 80.100 240.150 81.900 241.950 ;
        RECT 10.950 233.850 13.050 235.950 ;
        RECT 16.950 233.850 19.050 235.950 ;
        RECT 19.950 235.050 22.050 237.150 ;
        RECT 34.950 235.050 37.050 237.150 ;
        RECT 61.950 236.850 64.050 238.950 ;
        RECT 76.950 236.850 79.050 238.950 ;
        RECT 79.950 238.050 82.050 240.150 ;
        RECT 82.950 239.850 85.050 241.950 ;
        RECT 86.100 240.150 87.900 241.950 ;
        RECT 83.100 238.050 84.900 239.850 ;
        RECT 85.950 238.050 88.050 240.150 ;
        RECT 95.100 237.150 96.900 238.950 ;
        RECT 11.100 232.050 12.900 233.850 ;
        RECT 13.950 230.850 16.050 232.950 ;
        RECT 17.250 232.050 19.050 233.850 ;
        RECT 14.100 229.050 15.900 230.850 ;
        RECT 20.700 226.800 21.750 235.050 ;
        RECT 14.700 225.900 21.750 226.800 ;
        RECT 14.700 225.600 16.350 225.900 ;
        RECT 11.550 219.750 13.350 225.600 ;
        RECT 14.550 219.750 16.350 225.600 ;
        RECT 20.550 225.600 21.750 225.900 ;
        RECT 35.250 226.800 36.300 235.050 ;
        RECT 37.950 233.850 40.050 235.950 ;
        RECT 43.950 233.850 46.050 235.950 ;
        RECT 37.950 232.050 39.750 233.850 ;
        RECT 40.950 230.850 43.050 232.950 ;
        RECT 44.100 232.050 45.900 233.850 ;
        RECT 62.700 231.600 63.900 236.850 ;
        RECT 77.100 231.600 78.300 236.850 ;
        RECT 94.950 235.050 97.050 237.150 ;
        RECT 98.550 235.950 99.750 243.300 ;
        RECT 112.950 239.850 115.050 241.950 ;
        RECT 116.400 240.150 117.600 248.400 ;
        RECT 130.650 245.400 132.450 251.250 ;
        RECT 131.250 243.300 132.450 245.400 ;
        RECT 133.650 246.300 135.450 251.250 ;
        RECT 136.650 247.200 138.450 251.250 ;
        RECT 139.650 246.300 141.450 251.250 ;
        RECT 133.650 244.950 141.450 246.300 ;
        RECT 131.250 242.250 135.000 243.300 ;
        RECT 155.100 243.000 156.900 251.250 ;
        RECT 101.100 237.150 102.900 238.950 ;
        RECT 113.100 238.050 114.900 239.850 ;
        RECT 115.950 238.050 118.050 240.150 ;
        RECT 133.950 238.950 135.150 242.250 ;
        RECT 137.100 240.150 138.900 241.950 ;
        RECT 152.400 241.350 156.900 243.000 ;
        RECT 160.500 242.400 162.300 251.250 ;
        RECT 173.850 244.200 175.650 251.250 ;
        RECT 178.350 245.400 180.150 251.250 ;
        RECT 191.550 248.400 193.350 251.250 ;
        RECT 194.550 248.400 196.350 251.250 ;
        RECT 197.550 248.400 199.350 251.250 ;
        RECT 173.850 243.300 177.450 244.200 ;
        RECT 97.950 233.850 100.050 235.950 ;
        RECT 100.950 235.050 103.050 237.150 ;
        RECT 41.100 229.050 42.900 230.850 ;
        RECT 53.550 230.700 61.350 231.600 ;
        RECT 35.250 225.900 42.300 226.800 ;
        RECT 35.250 225.600 36.450 225.900 ;
        RECT 17.550 219.750 19.350 225.000 ;
        RECT 20.550 219.750 22.350 225.600 ;
        RECT 34.650 219.750 36.450 225.600 ;
        RECT 40.650 225.600 42.300 225.900 ;
        RECT 37.650 219.750 39.450 225.000 ;
        RECT 40.650 219.750 42.450 225.600 ;
        RECT 43.650 219.750 45.450 225.600 ;
        RECT 53.550 219.750 55.350 230.700 ;
        RECT 56.550 219.750 58.350 229.800 ;
        RECT 59.550 219.750 61.350 230.700 ;
        RECT 62.550 219.750 64.350 231.600 ;
        RECT 76.650 219.750 78.450 231.600 ;
        RECT 79.650 230.700 87.450 231.600 ;
        RECT 79.650 219.750 81.450 230.700 ;
        RECT 82.650 219.750 84.450 229.800 ;
        RECT 85.650 219.750 87.450 230.700 ;
        RECT 98.550 225.600 99.750 233.850 ;
        RECT 116.400 225.600 117.600 238.050 ;
        RECT 133.950 236.850 136.050 238.950 ;
        RECT 136.950 238.050 139.050 240.150 ;
        RECT 139.950 236.850 142.050 238.950 ;
        RECT 152.400 237.150 153.600 241.350 ;
        RECT 173.100 237.150 174.900 238.950 ;
        RECT 130.950 233.850 133.050 235.950 ;
        RECT 131.250 232.050 133.050 233.850 ;
        RECT 134.850 231.600 136.050 236.850 ;
        RECT 140.100 235.050 141.900 236.850 ;
        RECT 151.950 235.050 154.050 237.150 ;
        RECT 95.550 219.750 97.350 225.600 ;
        RECT 98.550 219.750 100.350 225.600 ;
        RECT 101.550 219.750 103.350 225.600 ;
        RECT 113.550 219.750 115.350 225.600 ;
        RECT 116.550 219.750 118.350 225.600 ;
        RECT 131.400 219.750 133.200 225.600 ;
        RECT 134.700 219.750 136.500 231.600 ;
        RECT 138.900 219.750 140.700 231.600 ;
        RECT 152.250 226.800 153.300 235.050 ;
        RECT 154.950 233.850 157.050 235.950 ;
        RECT 160.950 233.850 163.050 235.950 ;
        RECT 172.950 235.050 175.050 237.150 ;
        RECT 176.250 235.950 177.450 243.300 ;
        RECT 195.000 241.950 196.050 248.400 ;
        RECT 211.350 245.400 213.150 251.250 ;
        RECT 214.350 245.400 216.150 251.250 ;
        RECT 217.650 248.400 219.450 251.250 ;
        RECT 232.650 248.400 234.450 251.250 ;
        RECT 235.650 248.400 237.450 251.250 ;
        RECT 193.950 239.850 196.050 241.950 ;
        RECT 179.100 237.150 180.900 238.950 ;
        RECT 175.950 233.850 178.050 235.950 ;
        RECT 178.950 235.050 181.050 237.150 ;
        RECT 190.950 236.850 193.050 238.950 ;
        RECT 191.100 235.050 192.900 236.850 ;
        RECT 154.950 232.050 156.750 233.850 ;
        RECT 157.950 230.850 160.050 232.950 ;
        RECT 161.100 232.050 162.900 233.850 ;
        RECT 158.100 229.050 159.900 230.850 ;
        RECT 152.250 225.900 159.300 226.800 ;
        RECT 152.250 225.600 153.450 225.900 ;
        RECT 151.650 219.750 153.450 225.600 ;
        RECT 157.650 225.600 159.300 225.900 ;
        RECT 176.250 225.600 177.450 233.850 ;
        RECT 195.000 232.650 196.050 239.850 ;
        RECT 211.650 238.950 212.850 245.400 ;
        RECT 217.650 244.500 218.850 248.400 ;
        RECT 213.750 243.600 218.850 244.500 ;
        RECT 213.750 242.700 216.000 243.600 ;
        RECT 196.950 236.850 199.050 238.950 ;
        RECT 211.650 236.850 214.050 238.950 ;
        RECT 197.100 235.050 198.900 236.850 ;
        RECT 195.000 231.600 197.550 232.650 ;
        RECT 211.650 231.600 212.850 236.850 ;
        RECT 214.950 234.300 216.000 242.700 ;
        RECT 233.400 240.150 234.600 248.400 ;
        RECT 246.000 245.400 247.800 251.250 ;
        RECT 250.200 245.400 252.000 251.250 ;
        RECT 254.400 245.400 256.200 251.250 ;
        RECT 264.750 248.400 266.550 251.250 ;
        RECT 267.750 248.400 269.550 251.250 ;
        RECT 217.950 236.850 220.050 238.950 ;
        RECT 232.950 238.050 235.050 240.150 ;
        RECT 235.950 239.850 238.050 241.950 ;
        RECT 248.250 240.150 250.050 241.950 ;
        RECT 236.100 238.050 237.900 239.850 ;
        RECT 218.100 235.050 219.900 236.850 ;
        RECT 213.750 233.400 216.000 234.300 ;
        RECT 213.750 232.500 219.450 233.400 ;
        RECT 154.650 219.750 156.450 225.000 ;
        RECT 157.650 219.750 159.450 225.600 ;
        RECT 160.650 219.750 162.450 225.600 ;
        RECT 172.650 219.750 174.450 225.600 ;
        RECT 175.650 219.750 177.450 225.600 ;
        RECT 178.650 219.750 180.450 225.600 ;
        RECT 191.550 219.750 193.350 231.600 ;
        RECT 195.750 219.750 197.550 231.600 ;
        RECT 211.350 219.750 213.150 231.600 ;
        RECT 214.350 219.750 216.150 231.600 ;
        RECT 218.250 225.600 219.450 232.500 ;
        RECT 233.400 225.600 234.600 238.050 ;
        RECT 244.950 236.850 247.050 238.950 ;
        RECT 247.950 238.050 250.050 240.150 ;
        RECT 250.950 238.950 252.000 245.400 ;
        RECT 253.950 240.150 255.750 241.950 ;
        RECT 268.050 240.150 269.550 248.400 ;
        RECT 250.950 236.850 253.050 238.950 ;
        RECT 253.950 238.050 256.050 240.150 ;
        RECT 256.950 236.850 259.050 238.950 ;
        RECT 265.950 238.050 269.550 240.150 ;
        RECT 245.250 235.050 247.050 236.850 ;
        RECT 252.150 233.400 253.050 236.850 ;
        RECT 257.100 235.050 258.900 236.850 ;
        RECT 252.150 232.500 256.200 233.400 ;
        RECT 254.400 231.600 256.200 232.500 ;
        RECT 245.550 230.400 253.350 231.300 ;
        RECT 217.650 219.750 219.450 225.600 ;
        RECT 232.650 219.750 234.450 225.600 ;
        RECT 235.650 219.750 237.450 225.600 ;
        RECT 245.550 219.750 247.350 230.400 ;
        RECT 248.550 219.750 250.350 229.500 ;
        RECT 251.550 220.500 253.350 230.400 ;
        RECT 254.550 221.400 256.350 231.600 ;
        RECT 257.550 220.500 259.350 231.600 ;
        RECT 268.050 225.600 269.550 238.050 ;
        RECT 271.650 245.400 273.450 251.250 ;
        RECT 277.050 245.400 278.850 251.250 ;
        RECT 282.600 246.600 284.400 251.250 ;
        RECT 287.250 247.500 289.050 251.250 ;
        RECT 290.250 247.500 292.050 251.250 ;
        RECT 293.250 247.500 295.050 251.250 ;
        RECT 280.200 245.400 284.400 246.600 ;
        RECT 286.950 245.400 289.050 247.500 ;
        RECT 289.950 245.400 292.050 247.500 ;
        RECT 292.950 245.400 295.050 247.500 ;
        RECT 297.000 247.500 298.800 251.250 ;
        RECT 300.000 248.400 301.800 251.250 ;
        RECT 303.000 247.500 304.800 251.250 ;
        RECT 307.500 248.400 309.300 251.250 ;
        RECT 310.500 248.400 312.300 251.250 ;
        RECT 313.500 248.400 315.300 251.250 ;
        RECT 316.500 248.400 318.300 251.250 ;
        RECT 297.000 245.700 299.850 247.500 ;
        RECT 297.750 245.400 299.850 245.700 ;
        RECT 301.950 245.700 304.800 247.500 ;
        RECT 305.700 246.750 307.500 247.200 ;
        RECT 310.950 247.050 312.300 248.400 ;
        RECT 313.950 247.050 315.300 248.400 ;
        RECT 316.950 247.050 318.300 248.400 ;
        RECT 301.950 245.400 304.050 245.700 ;
        RECT 305.700 245.400 309.750 246.750 ;
        RECT 271.650 230.550 272.850 245.400 ;
        RECT 280.200 241.800 281.700 245.400 ;
        RECT 286.350 242.700 293.100 244.500 ;
        RECT 294.000 242.700 300.900 244.500 ;
        RECT 308.850 244.050 309.750 245.400 ;
        RECT 310.950 244.950 313.050 247.050 ;
        RECT 313.950 244.950 316.050 247.050 ;
        RECT 316.950 244.950 319.050 247.050 ;
        RECT 308.850 243.900 313.950 244.050 ;
        RECT 308.850 243.150 316.500 243.900 ;
        RECT 312.150 242.700 316.500 243.150 ;
        RECT 294.000 241.800 295.050 242.700 ;
        RECT 312.150 242.250 313.950 242.700 ;
        RECT 273.900 240.000 281.700 241.800 ;
        RECT 285.150 240.750 295.050 241.800 ;
        RECT 285.150 238.950 286.200 240.750 ;
        RECT 295.950 240.450 303.600 241.800 ;
        RECT 295.950 239.700 296.850 240.450 ;
        RECT 277.950 237.900 286.200 238.950 ;
        RECT 287.250 238.650 296.850 239.700 ;
        RECT 277.950 233.850 280.050 237.900 ;
        RECT 287.250 237.000 288.150 238.650 ;
        RECT 297.750 237.750 301.650 239.550 ;
        RECT 302.550 238.950 303.600 240.450 ;
        RECT 304.950 241.650 307.050 241.950 ;
        RECT 304.950 239.850 308.850 241.650 ;
        RECT 315.450 239.250 316.500 242.700 ;
        RECT 318.000 241.800 319.050 244.950 ;
        RECT 320.700 245.400 322.500 251.250 ;
        RECT 326.100 245.400 327.900 251.250 ;
        RECT 331.500 245.400 333.300 251.250 ;
        RECT 320.700 244.500 322.200 245.400 ;
        RECT 320.700 243.300 329.100 244.500 ;
        RECT 327.300 242.700 329.100 243.300 ;
        RECT 332.100 241.800 333.300 245.400 ;
        RECT 344.550 246.300 346.350 251.250 ;
        RECT 347.550 247.200 349.350 251.250 ;
        RECT 350.550 246.300 352.350 251.250 ;
        RECT 344.550 244.950 352.350 246.300 ;
        RECT 353.550 245.400 355.350 251.250 ;
        RECT 365.850 245.400 367.650 251.250 ;
        RECT 353.550 243.300 354.750 245.400 ;
        RECT 370.350 244.200 372.150 251.250 ;
        RECT 385.650 245.400 387.450 251.250 ;
        RECT 351.000 242.250 354.750 243.300 ;
        RECT 368.550 243.300 372.150 244.200 ;
        RECT 386.250 243.300 387.450 245.400 ;
        RECT 388.650 246.300 390.450 251.250 ;
        RECT 391.650 247.200 393.450 251.250 ;
        RECT 394.650 246.300 396.450 251.250 ;
        RECT 388.650 244.950 396.450 246.300 ;
        RECT 407.850 244.200 409.650 251.250 ;
        RECT 412.350 245.400 414.150 251.250 ;
        RECT 424.650 245.400 426.450 251.250 ;
        RECT 407.850 243.300 411.450 244.200 ;
        RECT 318.000 240.900 333.300 241.800 ;
        RECT 302.550 238.050 314.550 238.950 ;
        RECT 281.100 235.200 288.150 237.000 ;
        RECT 289.500 235.950 291.300 237.750 ;
        RECT 297.750 237.450 299.850 237.750 ;
        RECT 301.950 236.550 304.050 236.850 ;
        RECT 310.800 236.550 312.600 237.150 ;
        RECT 301.950 235.950 312.600 236.550 ;
        RECT 289.500 235.350 312.600 235.950 ;
        RECT 313.500 236.550 314.550 238.050 ;
        RECT 315.450 237.450 317.250 239.250 ;
        RECT 319.050 238.950 330.900 240.000 ;
        RECT 319.050 236.550 320.250 238.950 ;
        RECT 329.100 237.150 330.900 238.950 ;
        RECT 313.500 235.650 320.250 236.550 ;
        RECT 322.950 235.650 325.050 235.950 ;
        RECT 289.500 234.750 304.050 235.350 ;
        RECT 321.150 234.450 325.050 235.650 ;
        RECT 328.950 235.050 331.050 237.150 ;
        RECT 311.100 233.850 325.050 234.450 ;
        RECT 285.000 233.550 324.750 233.850 ;
        RECT 273.750 232.650 275.550 233.250 ;
        RECT 285.000 232.650 313.050 233.550 ;
        RECT 273.750 231.450 286.050 232.650 ;
        RECT 313.950 232.050 316.050 232.350 ;
        RECT 323.700 232.050 325.500 232.650 ;
        RECT 286.950 230.550 289.050 231.750 ;
        RECT 271.650 229.650 289.050 230.550 ;
        RECT 292.950 230.400 313.050 231.750 ;
        RECT 292.950 229.650 295.050 230.400 ;
        RECT 274.500 225.600 275.700 229.650 ;
        RECT 276.600 227.700 278.400 228.300 ;
        RECT 283.350 228.150 285.150 228.300 ;
        RECT 276.600 226.500 282.300 227.700 ;
        RECT 283.350 226.950 292.050 228.150 ;
        RECT 283.350 226.500 285.150 226.950 ;
        RECT 251.550 219.750 259.350 220.500 ;
        RECT 264.750 219.750 266.550 225.600 ;
        RECT 267.750 219.750 269.550 225.600 ;
        RECT 271.500 219.750 273.300 225.600 ;
        RECT 274.500 219.750 276.300 225.600 ;
        RECT 277.500 219.750 279.300 225.600 ;
        RECT 280.500 219.750 282.300 226.500 ;
        RECT 289.950 226.050 292.050 226.950 ;
        RECT 283.500 219.750 285.300 225.600 ;
        RECT 286.800 223.800 288.900 225.900 ;
        RECT 287.400 222.600 288.900 223.800 ;
        RECT 287.250 219.750 289.050 222.600 ;
        RECT 290.250 219.750 292.050 226.050 ;
        RECT 293.550 222.600 294.900 229.650 ;
        RECT 311.100 229.350 313.050 230.400 ;
        RECT 313.950 230.850 325.500 232.050 ;
        RECT 313.950 230.250 316.050 230.850 ;
        RECT 327.000 229.350 328.800 230.100 ;
        RECT 296.100 226.800 300.000 228.600 ;
        RECT 297.000 226.500 300.000 226.800 ;
        RECT 301.950 228.150 304.050 228.600 ;
        RECT 311.100 228.300 328.800 229.350 ;
        RECT 301.950 226.500 304.350 228.150 ;
        RECT 293.250 219.750 295.050 222.600 ;
        RECT 297.000 219.750 298.800 226.500 ;
        RECT 303.000 225.600 304.350 226.500 ;
        RECT 310.950 225.600 313.050 226.050 ;
        RECT 300.000 219.750 301.800 225.600 ;
        RECT 303.000 219.750 304.800 225.600 ;
        RECT 306.750 219.750 308.550 225.600 ;
        RECT 310.500 223.950 313.050 225.600 ;
        RECT 313.950 223.950 316.050 226.050 ;
        RECT 316.950 223.950 319.050 226.050 ;
        RECT 310.500 222.600 311.700 223.950 ;
        RECT 313.950 222.600 314.850 223.950 ;
        RECT 316.950 222.600 318.150 223.950 ;
        RECT 309.750 219.750 311.700 222.600 ;
        RECT 312.750 219.750 314.850 222.600 ;
        RECT 315.750 219.750 318.150 222.600 ;
        RECT 319.500 219.750 321.300 223.050 ;
        RECT 322.500 219.750 324.300 228.300 ;
        RECT 332.100 227.400 333.300 240.900 ;
        RECT 347.100 240.150 348.900 241.950 ;
        RECT 343.950 236.850 346.050 238.950 ;
        RECT 346.950 238.050 349.050 240.150 ;
        RECT 350.850 238.950 352.050 242.250 ;
        RECT 349.950 236.850 352.050 238.950 ;
        RECT 365.100 237.150 366.900 238.950 ;
        RECT 344.100 235.050 345.900 236.850 ;
        RECT 349.950 231.600 351.150 236.850 ;
        RECT 352.950 233.850 355.050 235.950 ;
        RECT 364.950 235.050 367.050 237.150 ;
        RECT 368.550 235.950 369.750 243.300 ;
        RECT 386.250 242.250 390.000 243.300 ;
        RECT 388.950 238.950 390.150 242.250 ;
        RECT 392.100 240.150 393.900 241.950 ;
        RECT 371.100 237.150 372.900 238.950 ;
        RECT 367.950 233.850 370.050 235.950 ;
        RECT 370.950 235.050 373.050 237.150 ;
        RECT 388.950 236.850 391.050 238.950 ;
        RECT 391.950 238.050 394.050 240.150 ;
        RECT 394.950 236.850 397.050 238.950 ;
        RECT 407.100 237.150 408.900 238.950 ;
        RECT 385.950 233.850 388.050 235.950 ;
        RECT 352.950 232.050 354.750 233.850 ;
        RECT 329.250 226.500 333.300 227.400 ;
        RECT 329.250 225.600 330.300 226.500 ;
        RECT 325.500 219.750 327.300 225.600 ;
        RECT 328.500 219.750 330.300 225.600 ;
        RECT 331.500 219.750 333.300 225.600 ;
        RECT 345.300 219.750 347.100 231.600 ;
        RECT 349.500 219.750 351.300 231.600 ;
        RECT 368.550 225.600 369.750 233.850 ;
        RECT 386.250 232.050 388.050 233.850 ;
        RECT 389.850 231.600 391.050 236.850 ;
        RECT 395.100 235.050 396.900 236.850 ;
        RECT 406.950 235.050 409.050 237.150 ;
        RECT 410.250 235.950 411.450 243.300 ;
        RECT 425.250 243.300 426.450 245.400 ;
        RECT 427.650 246.300 429.450 251.250 ;
        RECT 430.650 247.200 432.450 251.250 ;
        RECT 433.650 246.300 435.450 251.250 ;
        RECT 427.650 244.950 435.450 246.300 ;
        RECT 445.650 245.400 447.450 251.250 ;
        RECT 446.250 243.300 447.450 245.400 ;
        RECT 448.650 246.300 450.450 251.250 ;
        RECT 451.650 247.200 453.450 251.250 ;
        RECT 454.650 246.300 456.450 251.250 ;
        RECT 448.650 244.950 456.450 246.300 ;
        RECT 458.700 245.400 460.500 251.250 ;
        RECT 464.100 245.400 465.900 251.250 ;
        RECT 469.500 245.400 471.300 251.250 ;
        RECT 473.700 248.400 475.500 251.250 ;
        RECT 476.700 248.400 478.500 251.250 ;
        RECT 479.700 248.400 481.500 251.250 ;
        RECT 482.700 248.400 484.500 251.250 ;
        RECT 473.700 247.050 475.050 248.400 ;
        RECT 476.700 247.050 478.050 248.400 ;
        RECT 479.700 247.050 481.050 248.400 ;
        RECT 487.200 247.500 489.000 251.250 ;
        RECT 490.200 248.400 492.000 251.250 ;
        RECT 493.200 247.500 495.000 251.250 ;
        RECT 425.250 242.250 429.000 243.300 ;
        RECT 446.250 242.250 450.000 243.300 ;
        RECT 415.950 240.450 418.050 241.050 ;
        RECT 424.950 240.450 427.050 241.050 ;
        RECT 415.950 239.550 427.050 240.450 ;
        RECT 415.950 238.950 418.050 239.550 ;
        RECT 424.950 238.950 427.050 239.550 ;
        RECT 427.950 238.950 429.150 242.250 ;
        RECT 431.100 240.150 432.900 241.950 ;
        RECT 413.100 237.150 414.900 238.950 ;
        RECT 409.950 233.850 412.050 235.950 ;
        RECT 412.950 235.050 415.050 237.150 ;
        RECT 427.950 236.850 430.050 238.950 ;
        RECT 430.950 238.050 433.050 240.150 ;
        RECT 448.950 238.950 450.150 242.250 ;
        RECT 452.100 240.150 453.900 241.950 ;
        RECT 458.700 241.800 459.900 245.400 ;
        RECT 469.800 244.500 471.300 245.400 ;
        RECT 462.900 243.300 471.300 244.500 ;
        RECT 472.950 244.950 475.050 247.050 ;
        RECT 475.950 244.950 478.050 247.050 ;
        RECT 478.950 244.950 481.050 247.050 ;
        RECT 484.500 246.750 486.300 247.200 ;
        RECT 482.250 245.400 486.300 246.750 ;
        RECT 487.200 245.700 490.050 247.500 ;
        RECT 487.950 245.400 490.050 245.700 ;
        RECT 492.150 245.700 495.000 247.500 ;
        RECT 496.950 247.500 498.750 251.250 ;
        RECT 499.950 247.500 501.750 251.250 ;
        RECT 502.950 247.500 504.750 251.250 ;
        RECT 492.150 245.400 494.250 245.700 ;
        RECT 496.950 245.400 499.050 247.500 ;
        RECT 499.950 245.400 502.050 247.500 ;
        RECT 502.950 245.400 505.050 247.500 ;
        RECT 507.600 246.600 509.400 251.250 ;
        RECT 507.600 245.400 511.800 246.600 ;
        RECT 513.150 245.400 514.950 251.250 ;
        RECT 518.550 245.400 520.350 251.250 ;
        RECT 462.900 242.700 464.700 243.300 ;
        RECT 472.950 241.800 474.000 244.950 ;
        RECT 482.250 244.050 483.150 245.400 ;
        RECT 478.050 243.900 483.150 244.050 ;
        RECT 458.700 240.900 474.000 241.800 ;
        RECT 475.500 243.150 483.150 243.900 ;
        RECT 475.500 242.700 479.850 243.150 ;
        RECT 491.100 242.700 498.000 244.500 ;
        RECT 498.900 242.700 505.650 244.500 ;
        RECT 433.950 236.850 436.050 238.950 ;
        RECT 448.950 236.850 451.050 238.950 ;
        RECT 451.950 238.050 454.050 240.150 ;
        RECT 454.950 236.850 457.050 238.950 ;
        RECT 424.950 233.850 427.050 235.950 ;
        RECT 352.800 219.750 354.600 225.600 ;
        RECT 365.550 219.750 367.350 225.600 ;
        RECT 368.550 219.750 370.350 225.600 ;
        RECT 371.550 219.750 373.350 225.600 ;
        RECT 386.400 219.750 388.200 225.600 ;
        RECT 389.700 219.750 391.500 231.600 ;
        RECT 393.900 219.750 395.700 231.600 ;
        RECT 410.250 225.600 411.450 233.850 ;
        RECT 425.250 232.050 427.050 233.850 ;
        RECT 428.850 231.600 430.050 236.850 ;
        RECT 434.100 235.050 435.900 236.850 ;
        RECT 445.950 233.850 448.050 235.950 ;
        RECT 446.250 232.050 448.050 233.850 ;
        RECT 449.850 231.600 451.050 236.850 ;
        RECT 455.100 235.050 456.900 236.850 ;
        RECT 406.650 219.750 408.450 225.600 ;
        RECT 409.650 219.750 411.450 225.600 ;
        RECT 412.650 219.750 414.450 225.600 ;
        RECT 425.400 219.750 427.200 225.600 ;
        RECT 428.700 219.750 430.500 231.600 ;
        RECT 432.900 219.750 434.700 231.600 ;
        RECT 446.400 219.750 448.200 225.600 ;
        RECT 449.700 219.750 451.500 231.600 ;
        RECT 453.900 219.750 455.700 231.600 ;
        RECT 458.700 227.400 459.900 240.900 ;
        RECT 461.100 238.950 472.950 240.000 ;
        RECT 475.500 239.250 476.550 242.700 ;
        RECT 478.050 242.250 479.850 242.700 ;
        RECT 484.950 241.650 487.050 241.950 ;
        RECT 496.950 241.800 498.000 242.700 ;
        RECT 510.300 241.800 511.800 245.400 ;
        RECT 483.150 239.850 487.050 241.650 ;
        RECT 488.400 240.450 496.050 241.800 ;
        RECT 496.950 240.750 506.850 241.800 ;
        RECT 461.100 237.150 462.900 238.950 ;
        RECT 460.950 235.050 463.050 237.150 ;
        RECT 471.750 236.550 472.950 238.950 ;
        RECT 474.750 237.450 476.550 239.250 ;
        RECT 488.400 238.950 489.450 240.450 ;
        RECT 495.150 239.700 496.050 240.450 ;
        RECT 477.450 238.050 489.450 238.950 ;
        RECT 477.450 236.550 478.500 238.050 ;
        RECT 490.350 237.750 494.250 239.550 ;
        RECT 495.150 238.650 504.750 239.700 ;
        RECT 492.150 237.450 494.250 237.750 ;
        RECT 466.950 235.650 469.050 235.950 ;
        RECT 471.750 235.650 478.500 236.550 ;
        RECT 479.400 236.550 481.200 237.150 ;
        RECT 487.950 236.550 490.050 236.850 ;
        RECT 479.400 235.950 490.050 236.550 ;
        RECT 500.700 235.950 502.500 237.750 ;
        RECT 466.950 234.450 470.850 235.650 ;
        RECT 479.400 235.350 502.500 235.950 ;
        RECT 487.950 234.750 502.500 235.350 ;
        RECT 503.850 237.000 504.750 238.650 ;
        RECT 505.800 238.950 506.850 240.750 ;
        RECT 510.300 240.000 518.100 241.800 ;
        RECT 505.800 237.900 514.050 238.950 ;
        RECT 503.850 235.200 510.900 237.000 ;
        RECT 466.950 233.850 480.900 234.450 ;
        RECT 511.950 233.850 514.050 237.900 ;
        RECT 467.250 233.550 507.000 233.850 ;
        RECT 478.950 232.650 507.000 233.550 ;
        RECT 516.450 232.650 518.250 233.250 ;
        RECT 466.500 232.050 468.300 232.650 ;
        RECT 475.950 232.050 478.050 232.350 ;
        RECT 466.500 230.850 478.050 232.050 ;
        RECT 475.950 230.250 478.050 230.850 ;
        RECT 478.950 230.400 499.050 231.750 ;
        RECT 463.200 229.350 465.000 230.100 ;
        RECT 478.950 229.350 480.900 230.400 ;
        RECT 496.950 229.650 499.050 230.400 ;
        RECT 502.950 230.550 505.050 231.750 ;
        RECT 505.950 231.450 518.250 232.650 ;
        RECT 519.150 230.550 520.350 245.400 ;
        RECT 502.950 229.650 520.350 230.550 ;
        RECT 522.450 248.400 524.250 251.250 ;
        RECT 525.450 248.400 527.250 251.250 ;
        RECT 539.700 248.400 541.500 251.250 ;
        RECT 522.450 240.150 523.950 248.400 ;
        RECT 543.000 247.050 544.800 251.250 ;
        RECT 539.100 245.400 544.800 247.050 ;
        RECT 547.200 245.400 549.000 251.250 ;
        RECT 557.550 246.300 559.350 251.250 ;
        RECT 560.550 247.200 562.350 251.250 ;
        RECT 563.550 246.300 565.350 251.250 ;
        RECT 522.450 238.050 526.050 240.150 ;
        RECT 539.100 238.950 540.300 245.400 ;
        RECT 557.550 244.950 565.350 246.300 ;
        RECT 566.550 245.400 568.350 251.250 ;
        RECT 580.350 245.400 582.150 251.250 ;
        RECT 583.350 245.400 585.150 251.250 ;
        RECT 586.650 248.400 588.450 251.250 ;
        RECT 566.550 243.300 567.750 245.400 ;
        RECT 564.000 242.250 567.750 243.300 ;
        RECT 542.100 240.150 543.900 241.950 ;
        RECT 463.200 228.300 480.900 229.350 ;
        RECT 458.700 226.500 462.750 227.400 ;
        RECT 461.700 225.600 462.750 226.500 ;
        RECT 458.700 219.750 460.500 225.600 ;
        RECT 461.700 219.750 463.500 225.600 ;
        RECT 464.700 219.750 466.500 225.600 ;
        RECT 467.700 219.750 469.500 228.300 ;
        RECT 487.950 228.150 490.050 228.600 ;
        RECT 487.650 226.500 490.050 228.150 ;
        RECT 492.000 226.800 495.900 228.600 ;
        RECT 492.000 226.500 495.000 226.800 ;
        RECT 472.950 223.950 475.050 226.050 ;
        RECT 475.950 223.950 478.050 226.050 ;
        RECT 478.950 225.600 481.050 226.050 ;
        RECT 487.650 225.600 489.000 226.500 ;
        RECT 478.950 223.950 481.500 225.600 ;
        RECT 470.700 219.750 472.500 223.050 ;
        RECT 473.850 222.600 475.050 223.950 ;
        RECT 477.150 222.600 478.050 223.950 ;
        RECT 480.300 222.600 481.500 223.950 ;
        RECT 473.850 219.750 476.250 222.600 ;
        RECT 477.150 219.750 479.250 222.600 ;
        RECT 480.300 219.750 482.250 222.600 ;
        RECT 483.450 219.750 485.250 225.600 ;
        RECT 487.200 219.750 489.000 225.600 ;
        RECT 490.200 219.750 492.000 225.600 ;
        RECT 493.200 219.750 495.000 226.500 ;
        RECT 497.100 222.600 498.450 229.650 ;
        RECT 506.850 228.150 508.650 228.300 ;
        RECT 499.950 226.950 508.650 228.150 ;
        RECT 513.600 227.700 515.400 228.300 ;
        RECT 499.950 226.050 502.050 226.950 ;
        RECT 506.850 226.500 508.650 226.950 ;
        RECT 509.700 226.500 515.400 227.700 ;
        RECT 496.950 219.750 498.750 222.600 ;
        RECT 499.950 219.750 501.750 226.050 ;
        RECT 503.100 223.800 505.200 225.900 ;
        RECT 503.100 222.600 504.600 223.800 ;
        RECT 502.950 219.750 504.750 222.600 ;
        RECT 506.700 219.750 508.500 225.600 ;
        RECT 509.700 219.750 511.500 226.500 ;
        RECT 516.300 225.600 517.500 229.650 ;
        RECT 522.450 225.600 523.950 238.050 ;
        RECT 538.950 236.850 541.050 238.950 ;
        RECT 541.950 238.050 544.050 240.150 ;
        RECT 544.950 239.850 547.050 241.950 ;
        RECT 548.100 240.150 549.900 241.950 ;
        RECT 560.100 240.150 561.900 241.950 ;
        RECT 545.100 238.050 546.900 239.850 ;
        RECT 547.950 238.050 550.050 240.150 ;
        RECT 556.950 236.850 559.050 238.950 ;
        RECT 559.950 238.050 562.050 240.150 ;
        RECT 563.850 238.950 565.050 242.250 ;
        RECT 562.950 236.850 565.050 238.950 ;
        RECT 580.650 238.950 581.850 245.400 ;
        RECT 586.650 244.500 587.850 248.400 ;
        RECT 600.150 246.900 601.950 251.250 ;
        RECT 582.750 243.600 587.850 244.500 ;
        RECT 598.650 245.400 601.950 246.900 ;
        RECT 603.150 245.400 604.950 251.250 ;
        RECT 582.750 242.700 585.000 243.600 ;
        RECT 580.650 236.850 583.050 238.950 ;
        RECT 539.100 231.600 540.300 236.850 ;
        RECT 557.100 235.050 558.900 236.850 ;
        RECT 562.950 231.600 564.150 236.850 ;
        RECT 565.950 233.850 568.050 235.950 ;
        RECT 565.950 232.050 567.750 233.850 ;
        RECT 580.650 231.600 581.850 236.850 ;
        RECT 583.950 234.300 585.000 242.700 ;
        RECT 598.650 238.950 599.850 245.400 ;
        RECT 601.950 243.900 603.750 244.500 ;
        RECT 607.650 243.900 609.450 251.250 ;
        RECT 617.850 245.400 619.650 251.250 ;
        RECT 622.350 244.200 624.150 251.250 ;
        RECT 640.800 245.400 642.600 251.250 ;
        RECT 645.000 245.400 646.800 251.250 ;
        RECT 649.200 245.400 651.000 251.250 ;
        RECT 664.800 245.400 666.600 251.250 ;
        RECT 669.000 245.400 670.800 251.250 ;
        RECT 673.200 245.400 675.000 251.250 ;
        RECT 687.000 245.400 688.800 251.250 ;
        RECT 691.200 245.400 693.000 251.250 ;
        RECT 695.400 245.400 697.200 251.250 ;
        RECT 710.850 245.400 712.650 251.250 ;
        RECT 601.950 242.700 609.450 243.900 ;
        RECT 620.550 243.300 624.150 244.200 ;
        RECT 586.950 236.850 589.050 238.950 ;
        RECT 598.650 236.850 601.050 238.950 ;
        RECT 602.100 237.150 603.900 238.950 ;
        RECT 587.100 235.050 588.900 236.850 ;
        RECT 582.750 233.400 585.000 234.300 ;
        RECT 582.750 232.500 588.450 233.400 ;
        RECT 512.700 219.750 514.500 225.600 ;
        RECT 515.700 219.750 517.500 225.600 ;
        RECT 518.700 219.750 520.500 225.600 ;
        RECT 522.450 219.750 524.250 225.600 ;
        RECT 525.450 219.750 527.250 225.600 ;
        RECT 538.650 219.750 540.450 231.600 ;
        RECT 541.650 230.700 549.450 231.600 ;
        RECT 541.650 219.750 543.450 230.700 ;
        RECT 544.650 219.750 546.450 229.800 ;
        RECT 547.650 219.750 549.450 230.700 ;
        RECT 558.300 219.750 560.100 231.600 ;
        RECT 562.500 219.750 564.300 231.600 ;
        RECT 565.800 219.750 567.600 225.600 ;
        RECT 580.350 219.750 582.150 231.600 ;
        RECT 583.350 219.750 585.150 231.600 ;
        RECT 587.250 225.600 588.450 232.500 ;
        RECT 598.650 231.600 599.850 236.850 ;
        RECT 601.950 235.050 604.050 237.150 ;
        RECT 586.650 219.750 588.450 225.600 ;
        RECT 598.050 219.750 599.850 231.600 ;
        RECT 601.050 219.750 602.850 231.600 ;
        RECT 605.100 225.600 606.300 242.700 ;
        RECT 607.950 236.850 610.050 238.950 ;
        RECT 617.100 237.150 618.900 238.950 ;
        RECT 608.100 235.050 609.900 236.850 ;
        RECT 616.950 235.050 619.050 237.150 ;
        RECT 620.550 235.950 621.750 243.300 ;
        RECT 641.250 240.150 643.050 241.950 ;
        RECT 623.100 237.150 624.900 238.950 ;
        RECT 619.950 233.850 622.050 235.950 ;
        RECT 622.950 235.050 625.050 237.150 ;
        RECT 637.950 236.850 640.050 238.950 ;
        RECT 640.950 238.050 643.050 240.150 ;
        RECT 645.000 238.950 646.050 245.400 ;
        RECT 643.950 236.850 646.050 238.950 ;
        RECT 646.950 240.150 648.750 241.950 ;
        RECT 665.250 240.150 667.050 241.950 ;
        RECT 646.950 238.050 649.050 240.150 ;
        RECT 649.950 236.850 652.050 238.950 ;
        RECT 661.950 236.850 664.050 238.950 ;
        RECT 664.950 238.050 667.050 240.150 ;
        RECT 669.000 238.950 670.050 245.400 ;
        RECT 673.950 243.450 676.050 244.050 ;
        RECT 673.950 242.550 684.450 243.450 ;
        RECT 673.950 241.950 676.050 242.550 ;
        RECT 667.950 236.850 670.050 238.950 ;
        RECT 670.950 240.150 672.750 241.950 ;
        RECT 670.950 238.050 673.050 240.150 ;
        RECT 673.950 236.850 676.050 238.950 ;
        RECT 638.100 235.050 639.900 236.850 ;
        RECT 620.550 225.600 621.750 233.850 ;
        RECT 643.950 233.400 644.850 236.850 ;
        RECT 649.950 235.050 651.750 236.850 ;
        RECT 662.100 235.050 663.900 236.850 ;
        RECT 667.950 233.400 668.850 236.850 ;
        RECT 673.950 235.050 675.750 236.850 ;
        RECT 683.550 235.050 684.450 242.550 ;
        RECT 689.250 240.150 691.050 241.950 ;
        RECT 685.950 236.850 688.050 238.950 ;
        RECT 688.950 238.050 691.050 240.150 ;
        RECT 691.950 238.950 693.000 245.400 ;
        RECT 715.350 244.200 717.150 251.250 ;
        RECT 728.550 246.300 730.350 251.250 ;
        RECT 731.550 247.200 733.350 251.250 ;
        RECT 734.550 246.300 736.350 251.250 ;
        RECT 728.550 244.950 736.350 246.300 ;
        RECT 737.550 245.400 739.350 251.250 ;
        RECT 753.150 246.900 754.950 251.250 ;
        RECT 751.650 245.400 754.950 246.900 ;
        RECT 756.150 245.400 757.950 251.250 ;
        RECT 713.550 243.300 717.150 244.200 ;
        RECT 737.550 243.300 738.750 245.400 ;
        RECT 694.950 240.150 696.750 241.950 ;
        RECT 691.950 236.850 694.050 238.950 ;
        RECT 694.950 238.050 697.050 240.150 ;
        RECT 697.950 236.850 700.050 238.950 ;
        RECT 710.100 237.150 711.900 238.950 ;
        RECT 686.250 235.050 688.050 236.850 ;
        RECT 640.800 232.500 644.850 233.400 ;
        RECT 664.800 232.500 668.850 233.400 ;
        RECT 682.950 232.950 685.050 235.050 ;
        RECT 693.150 233.400 694.050 236.850 ;
        RECT 698.100 235.050 699.900 236.850 ;
        RECT 709.950 235.050 712.050 237.150 ;
        RECT 713.550 235.950 714.750 243.300 ;
        RECT 735.000 242.250 738.750 243.300 ;
        RECT 731.100 240.150 732.900 241.950 ;
        RECT 716.100 237.150 717.900 238.950 ;
        RECT 712.950 233.850 715.050 235.950 ;
        RECT 715.950 235.050 718.050 237.150 ;
        RECT 727.950 236.850 730.050 238.950 ;
        RECT 730.950 238.050 733.050 240.150 ;
        RECT 734.850 238.950 736.050 242.250 ;
        RECT 733.950 236.850 736.050 238.950 ;
        RECT 751.650 238.950 752.850 245.400 ;
        RECT 754.950 243.900 756.750 244.500 ;
        RECT 760.650 243.900 762.450 251.250 ;
        RECT 754.950 242.700 762.450 243.900 ;
        RECT 751.650 236.850 754.050 238.950 ;
        RECT 755.100 237.150 756.900 238.950 ;
        RECT 728.100 235.050 729.900 236.850 ;
        RECT 693.150 232.500 697.200 233.400 ;
        RECT 640.800 231.600 642.600 232.500 ;
        RECT 664.800 231.600 666.600 232.500 ;
        RECT 695.400 231.600 697.200 232.500 ;
        RECT 604.650 219.750 606.450 225.600 ;
        RECT 607.650 219.750 609.450 225.600 ;
        RECT 617.550 219.750 619.350 225.600 ;
        RECT 620.550 219.750 622.350 225.600 ;
        RECT 623.550 219.750 625.350 225.600 ;
        RECT 637.650 220.500 639.450 231.600 ;
        RECT 640.650 221.400 642.450 231.600 ;
        RECT 643.650 230.400 651.450 231.300 ;
        RECT 643.650 220.500 645.450 230.400 ;
        RECT 637.650 219.750 645.450 220.500 ;
        RECT 646.650 219.750 648.450 229.500 ;
        RECT 649.650 219.750 651.450 230.400 ;
        RECT 661.650 220.500 663.450 231.600 ;
        RECT 664.650 221.400 666.450 231.600 ;
        RECT 667.650 230.400 675.450 231.300 ;
        RECT 667.650 220.500 669.450 230.400 ;
        RECT 661.650 219.750 669.450 220.500 ;
        RECT 670.650 219.750 672.450 229.500 ;
        RECT 673.650 219.750 675.450 230.400 ;
        RECT 686.550 230.400 694.350 231.300 ;
        RECT 686.550 219.750 688.350 230.400 ;
        RECT 689.550 219.750 691.350 229.500 ;
        RECT 692.550 220.500 694.350 230.400 ;
        RECT 695.550 221.400 697.350 231.600 ;
        RECT 698.550 220.500 700.350 231.600 ;
        RECT 713.550 225.600 714.750 233.850 ;
        RECT 733.950 231.600 735.150 236.850 ;
        RECT 736.950 233.850 739.050 235.950 ;
        RECT 736.950 232.050 738.750 233.850 ;
        RECT 751.650 231.600 752.850 236.850 ;
        RECT 754.950 235.050 757.050 237.150 ;
        RECT 692.550 219.750 700.350 220.500 ;
        RECT 710.550 219.750 712.350 225.600 ;
        RECT 713.550 219.750 715.350 225.600 ;
        RECT 716.550 219.750 718.350 225.600 ;
        RECT 729.300 219.750 731.100 231.600 ;
        RECT 733.500 219.750 735.300 231.600 ;
        RECT 736.800 219.750 738.600 225.600 ;
        RECT 751.050 219.750 752.850 231.600 ;
        RECT 754.050 219.750 755.850 231.600 ;
        RECT 758.100 225.600 759.300 242.700 ;
        RECT 773.700 242.400 775.500 251.250 ;
        RECT 779.100 243.000 780.900 251.250 ;
        RECT 781.950 246.450 784.050 247.050 ;
        RECT 787.950 246.450 790.050 247.050 ;
        RECT 781.950 245.550 790.050 246.450 ;
        RECT 781.950 244.950 784.050 245.550 ;
        RECT 787.950 244.950 790.050 245.550 ;
        RECT 795.000 245.400 796.800 251.250 ;
        RECT 799.200 245.400 801.000 251.250 ;
        RECT 803.400 245.400 805.200 251.250 ;
        RECT 818.850 245.400 820.650 251.250 ;
        RECT 790.950 243.450 793.050 244.050 ;
        RECT 779.100 241.350 783.600 243.000 ;
        RECT 772.950 240.450 775.050 241.050 ;
        RECT 770.550 239.550 775.050 240.450 ;
        RECT 760.950 236.850 763.050 238.950 ;
        RECT 761.100 235.050 762.900 236.850 ;
        RECT 770.550 228.450 771.450 239.550 ;
        RECT 772.950 238.950 775.050 239.550 ;
        RECT 782.400 237.150 783.600 241.350 ;
        RECT 788.550 242.550 793.050 243.450 ;
        RECT 772.950 233.850 775.050 235.950 ;
        RECT 778.950 233.850 781.050 235.950 ;
        RECT 781.950 235.050 784.050 237.150 ;
        RECT 773.100 232.050 774.900 233.850 ;
        RECT 775.950 230.850 778.050 232.950 ;
        RECT 779.250 232.050 781.050 233.850 ;
        RECT 776.100 229.050 777.900 230.850 ;
        RECT 772.950 228.450 775.050 229.050 ;
        RECT 770.550 227.550 775.050 228.450 ;
        RECT 772.950 226.950 775.050 227.550 ;
        RECT 782.700 226.800 783.750 235.050 ;
        RECT 788.550 229.050 789.450 242.550 ;
        RECT 790.950 241.950 793.050 242.550 ;
        RECT 797.250 240.150 799.050 241.950 ;
        RECT 793.950 236.850 796.050 238.950 ;
        RECT 796.950 238.050 799.050 240.150 ;
        RECT 799.950 238.950 801.000 245.400 ;
        RECT 823.350 244.200 825.150 251.250 ;
        RECT 821.550 243.300 825.150 244.200 ;
        RECT 829.950 243.450 832.050 244.050 ;
        RECT 802.950 240.150 804.750 241.950 ;
        RECT 799.950 236.850 802.050 238.950 ;
        RECT 802.950 238.050 805.050 240.150 ;
        RECT 805.950 236.850 808.050 238.950 ;
        RECT 818.100 237.150 819.900 238.950 ;
        RECT 794.250 235.050 796.050 236.850 ;
        RECT 801.150 233.400 802.050 236.850 ;
        RECT 806.100 235.050 807.900 236.850 ;
        RECT 817.950 235.050 820.050 237.150 ;
        RECT 821.550 235.950 822.750 243.300 ;
        RECT 827.550 242.550 832.050 243.450 ;
        RECT 824.100 237.150 825.900 238.950 ;
        RECT 820.950 233.850 823.050 235.950 ;
        RECT 823.950 235.050 826.050 237.150 ;
        RECT 801.150 232.500 805.200 233.400 ;
        RECT 803.400 231.600 805.200 232.500 ;
        RECT 794.550 230.400 802.350 231.300 ;
        RECT 787.950 226.950 790.050 229.050 ;
        RECT 776.700 225.900 783.750 226.800 ;
        RECT 776.700 225.600 778.350 225.900 ;
        RECT 757.650 219.750 759.450 225.600 ;
        RECT 760.650 219.750 762.450 225.600 ;
        RECT 773.550 219.750 775.350 225.600 ;
        RECT 776.550 219.750 778.350 225.600 ;
        RECT 782.550 225.600 783.750 225.900 ;
        RECT 779.550 219.750 781.350 225.000 ;
        RECT 782.550 219.750 784.350 225.600 ;
        RECT 794.550 219.750 796.350 230.400 ;
        RECT 797.550 219.750 799.350 229.500 ;
        RECT 800.550 220.500 802.350 230.400 ;
        RECT 803.550 221.400 805.350 231.600 ;
        RECT 806.550 220.500 808.350 231.600 ;
        RECT 821.550 225.600 822.750 233.850 ;
        RECT 823.950 231.450 826.050 232.050 ;
        RECT 827.550 231.450 828.450 242.550 ;
        RECT 829.950 241.950 832.050 242.550 ;
        RECT 836.700 242.400 838.500 251.250 ;
        RECT 842.100 243.000 843.900 251.250 ;
        RECT 862.650 245.400 864.450 251.250 ;
        RECT 865.650 245.400 867.450 251.250 ;
        RECT 842.100 241.350 846.600 243.000 ;
        RECT 845.400 237.150 846.600 241.350 ;
        RECT 863.400 238.950 864.600 245.400 ;
        RECT 866.100 240.150 867.900 241.950 ;
        RECT 835.950 233.850 838.050 235.950 ;
        RECT 841.950 233.850 844.050 235.950 ;
        RECT 844.950 235.050 847.050 237.150 ;
        RECT 862.950 236.850 865.050 238.950 ;
        RECT 865.950 238.050 868.050 240.150 ;
        RECT 836.100 232.050 837.900 233.850 ;
        RECT 823.950 230.550 828.450 231.450 ;
        RECT 838.950 230.850 841.050 232.950 ;
        RECT 842.250 232.050 844.050 233.850 ;
        RECT 823.950 229.950 826.050 230.550 ;
        RECT 839.100 229.050 840.900 230.850 ;
        RECT 845.700 226.800 846.750 235.050 ;
        RECT 863.400 231.600 864.600 236.850 ;
        RECT 839.700 225.900 846.750 226.800 ;
        RECT 839.700 225.600 841.350 225.900 ;
        RECT 800.550 219.750 808.350 220.500 ;
        RECT 818.550 219.750 820.350 225.600 ;
        RECT 821.550 219.750 823.350 225.600 ;
        RECT 824.550 219.750 826.350 225.600 ;
        RECT 836.550 219.750 838.350 225.600 ;
        RECT 839.550 219.750 841.350 225.600 ;
        RECT 845.550 225.600 846.750 225.900 ;
        RECT 842.550 219.750 844.350 225.000 ;
        RECT 845.550 219.750 847.350 225.600 ;
        RECT 862.650 219.750 864.450 231.600 ;
        RECT 865.650 219.750 867.450 231.600 ;
        RECT 10.650 209.400 12.450 215.250 ;
        RECT 13.650 210.000 15.450 215.250 ;
        RECT 11.250 209.100 12.450 209.400 ;
        RECT 16.650 209.400 18.450 215.250 ;
        RECT 19.650 209.400 21.450 215.250 ;
        RECT 16.650 209.100 18.300 209.400 ;
        RECT 11.250 208.200 18.300 209.100 ;
        RECT 11.250 199.950 12.300 208.200 ;
        RECT 17.100 204.150 18.900 205.950 ;
        RECT 29.550 204.300 31.350 215.250 ;
        RECT 32.550 205.200 34.350 215.250 ;
        RECT 35.550 204.300 37.350 215.250 ;
        RECT 13.950 201.150 15.750 202.950 ;
        RECT 16.950 202.050 19.050 204.150 ;
        RECT 29.550 203.400 37.350 204.300 ;
        RECT 38.550 203.400 40.350 215.250 ;
        RECT 52.650 209.400 54.450 215.250 ;
        RECT 55.650 210.000 57.450 215.250 ;
        RECT 53.250 209.100 54.450 209.400 ;
        RECT 58.650 209.400 60.450 215.250 ;
        RECT 61.650 209.400 63.450 215.250 ;
        RECT 74.400 209.400 76.200 215.250 ;
        RECT 58.650 209.100 60.300 209.400 ;
        RECT 53.250 208.200 60.300 209.100 ;
        RECT 20.100 201.150 21.900 202.950 ;
        RECT 10.950 197.850 13.050 199.950 ;
        RECT 13.950 199.050 16.050 201.150 ;
        RECT 19.950 199.050 22.050 201.150 ;
        RECT 38.700 198.150 39.900 203.400 ;
        RECT 53.250 199.950 54.300 208.200 ;
        RECT 59.100 204.150 60.900 205.950 ;
        RECT 55.950 201.150 57.750 202.950 ;
        RECT 58.950 202.050 61.050 204.150 ;
        RECT 77.700 203.400 79.500 215.250 ;
        RECT 81.900 203.400 83.700 215.250 ;
        RECT 95.400 209.400 97.200 215.250 ;
        RECT 98.700 203.400 100.500 215.250 ;
        RECT 102.900 203.400 104.700 215.250 ;
        RECT 118.050 203.400 119.850 215.250 ;
        RECT 121.050 203.400 122.850 215.250 ;
        RECT 124.650 209.400 126.450 215.250 ;
        RECT 127.650 209.400 129.450 215.250 ;
        RECT 137.550 209.400 139.350 215.250 ;
        RECT 140.550 209.400 142.350 215.250 ;
        RECT 143.550 209.400 145.350 215.250 ;
        RECT 157.650 209.400 159.450 215.250 ;
        RECT 160.650 209.400 162.450 215.250 ;
        RECT 170.550 209.400 172.350 215.250 ;
        RECT 173.550 209.400 175.350 215.250 ;
        RECT 176.550 210.000 178.350 215.250 ;
        RECT 62.100 201.150 63.900 202.950 ;
        RECT 74.250 201.150 76.050 202.950 ;
        RECT 11.400 193.650 12.600 197.850 ;
        RECT 28.950 194.850 31.050 196.950 ;
        RECT 32.100 195.150 33.900 196.950 ;
        RECT 11.400 192.000 15.900 193.650 ;
        RECT 29.100 193.050 30.900 194.850 ;
        RECT 31.950 193.050 34.050 195.150 ;
        RECT 34.950 194.850 37.050 196.950 ;
        RECT 37.950 196.050 40.050 198.150 ;
        RECT 52.950 197.850 55.050 199.950 ;
        RECT 55.950 199.050 58.050 201.150 ;
        RECT 61.950 199.050 64.050 201.150 ;
        RECT 73.950 199.050 76.050 201.150 ;
        RECT 77.850 198.150 79.050 203.400 ;
        RECT 95.250 201.150 97.050 202.950 ;
        RECT 83.100 198.150 84.900 199.950 ;
        RECT 94.950 199.050 97.050 201.150 ;
        RECT 98.850 198.150 100.050 203.400 ;
        RECT 104.100 198.150 105.900 199.950 ;
        RECT 118.650 198.150 119.850 203.400 ;
        RECT 35.100 193.050 36.900 194.850 ;
        RECT 14.100 183.750 15.900 192.000 ;
        RECT 19.500 183.750 21.300 192.600 ;
        RECT 38.700 189.600 39.900 196.050 ;
        RECT 53.400 193.650 54.600 197.850 ;
        RECT 76.950 196.050 79.050 198.150 ;
        RECT 53.400 192.000 57.900 193.650 ;
        RECT 76.950 192.750 78.150 196.050 ;
        RECT 79.950 194.850 82.050 196.950 ;
        RECT 82.950 196.050 85.050 198.150 ;
        RECT 97.950 196.050 100.050 198.150 ;
        RECT 80.100 193.050 81.900 194.850 ;
        RECT 97.950 192.750 99.150 196.050 ;
        RECT 100.950 194.850 103.050 196.950 ;
        RECT 103.950 196.050 106.050 198.150 ;
        RECT 118.650 196.050 121.050 198.150 ;
        RECT 121.950 197.850 124.050 199.950 ;
        RECT 122.100 196.050 123.900 197.850 ;
        RECT 101.100 193.050 102.900 194.850 ;
        RECT 30.000 183.750 31.800 189.600 ;
        RECT 34.200 187.950 39.900 189.600 ;
        RECT 34.200 183.750 36.000 187.950 ;
        RECT 37.500 183.750 39.300 186.600 ;
        RECT 56.100 183.750 57.900 192.000 ;
        RECT 61.500 183.750 63.300 192.600 ;
        RECT 74.250 191.700 78.000 192.750 ;
        RECT 95.250 191.700 99.000 192.750 ;
        RECT 74.250 189.600 75.450 191.700 ;
        RECT 73.650 183.750 75.450 189.600 ;
        RECT 76.650 188.700 84.450 190.050 ;
        RECT 95.250 189.600 96.450 191.700 ;
        RECT 76.650 183.750 78.450 188.700 ;
        RECT 79.650 183.750 81.450 187.800 ;
        RECT 82.650 183.750 84.450 188.700 ;
        RECT 94.650 183.750 96.450 189.600 ;
        RECT 97.650 188.700 105.450 190.050 ;
        RECT 97.650 183.750 99.450 188.700 ;
        RECT 100.650 183.750 102.450 187.800 ;
        RECT 103.650 183.750 105.450 188.700 ;
        RECT 118.650 189.600 119.850 196.050 ;
        RECT 125.100 192.300 126.300 209.400 ;
        RECT 140.550 201.150 141.750 209.400 ;
        RECT 128.100 198.150 129.900 199.950 ;
        RECT 127.950 196.050 130.050 198.150 ;
        RECT 136.950 197.850 139.050 199.950 ;
        RECT 139.950 199.050 142.050 201.150 ;
        RECT 137.100 196.050 138.900 197.850 ;
        RECT 121.950 191.100 129.450 192.300 ;
        RECT 121.950 190.500 123.750 191.100 ;
        RECT 118.650 188.100 121.950 189.600 ;
        RECT 120.150 183.750 121.950 188.100 ;
        RECT 123.150 183.750 124.950 189.600 ;
        RECT 127.650 183.750 129.450 191.100 ;
        RECT 140.550 191.700 141.750 199.050 ;
        RECT 142.950 197.850 145.050 199.950 ;
        RECT 143.100 196.050 144.900 197.850 ;
        RECT 158.400 196.950 159.600 209.400 ;
        RECT 173.700 209.100 175.350 209.400 ;
        RECT 179.550 209.400 181.350 215.250 ;
        RECT 191.550 209.400 193.350 215.250 ;
        RECT 194.550 209.400 196.350 215.250 ;
        RECT 197.550 209.400 199.350 215.250 ;
        RECT 211.650 209.400 213.450 215.250 ;
        RECT 214.650 209.400 216.450 215.250 ;
        RECT 217.650 209.400 219.450 215.250 ;
        RECT 229.650 209.400 231.450 215.250 ;
        RECT 232.650 209.400 234.450 215.250 ;
        RECT 235.650 209.400 237.450 215.250 ;
        RECT 250.650 209.400 252.450 215.250 ;
        RECT 253.650 210.000 255.450 215.250 ;
        RECT 179.550 209.100 180.750 209.400 ;
        RECT 173.700 208.200 180.750 209.100 ;
        RECT 173.100 204.150 174.900 205.950 ;
        RECT 170.100 201.150 171.900 202.950 ;
        RECT 172.950 202.050 175.050 204.150 ;
        RECT 176.250 201.150 178.050 202.950 ;
        RECT 169.950 199.050 172.050 201.150 ;
        RECT 175.950 199.050 178.050 201.150 ;
        RECT 179.700 199.950 180.750 208.200 ;
        RECT 194.550 201.150 195.750 209.400 ;
        RECT 215.250 201.150 216.450 209.400 ;
        RECT 233.250 201.150 234.450 209.400 ;
        RECT 251.250 209.100 252.450 209.400 ;
        RECT 256.650 209.400 258.450 215.250 ;
        RECT 259.650 209.400 261.450 215.250 ;
        RECT 269.550 209.400 271.350 215.250 ;
        RECT 272.550 209.400 274.350 215.250 ;
        RECT 275.550 209.400 277.350 215.250 ;
        RECT 289.650 209.400 291.450 215.250 ;
        RECT 292.650 210.000 294.450 215.250 ;
        RECT 256.650 209.100 258.300 209.400 ;
        RECT 251.250 208.200 258.300 209.100 ;
        RECT 178.950 197.850 181.050 199.950 ;
        RECT 190.950 197.850 193.050 199.950 ;
        RECT 193.950 199.050 196.050 201.150 ;
        RECT 157.950 194.850 160.050 196.950 ;
        RECT 161.100 195.150 162.900 196.950 ;
        RECT 140.550 190.800 144.150 191.700 ;
        RECT 137.850 183.750 139.650 189.600 ;
        RECT 142.350 183.750 144.150 190.800 ;
        RECT 158.400 186.600 159.600 194.850 ;
        RECT 160.950 193.050 163.050 195.150 ;
        RECT 179.400 193.650 180.600 197.850 ;
        RECT 191.100 196.050 192.900 197.850 ;
        RECT 157.650 183.750 159.450 186.600 ;
        RECT 160.650 183.750 162.450 186.600 ;
        RECT 170.700 183.750 172.500 192.600 ;
        RECT 176.100 192.000 180.600 193.650 ;
        RECT 176.100 183.750 177.900 192.000 ;
        RECT 194.550 191.700 195.750 199.050 ;
        RECT 196.950 197.850 199.050 199.950 ;
        RECT 211.950 197.850 214.050 199.950 ;
        RECT 214.950 199.050 217.050 201.150 ;
        RECT 197.100 196.050 198.900 197.850 ;
        RECT 212.100 196.050 213.900 197.850 ;
        RECT 215.250 191.700 216.450 199.050 ;
        RECT 217.950 197.850 220.050 199.950 ;
        RECT 229.950 197.850 232.050 199.950 ;
        RECT 232.950 199.050 235.050 201.150 ;
        RECT 251.250 199.950 252.300 208.200 ;
        RECT 257.100 204.150 258.900 205.950 ;
        RECT 253.950 201.150 255.750 202.950 ;
        RECT 256.950 202.050 259.050 204.150 ;
        RECT 260.100 201.150 261.900 202.950 ;
        RECT 272.550 201.150 273.750 209.400 ;
        RECT 290.250 209.100 291.450 209.400 ;
        RECT 295.650 209.400 297.450 215.250 ;
        RECT 298.650 209.400 300.450 215.250 ;
        RECT 310.650 209.400 312.450 215.250 ;
        RECT 313.650 209.400 315.450 215.250 ;
        RECT 328.650 209.400 330.450 215.250 ;
        RECT 331.650 210.000 333.450 215.250 ;
        RECT 295.650 209.100 297.300 209.400 ;
        RECT 290.250 208.200 297.300 209.100 ;
        RECT 218.100 196.050 219.900 197.850 ;
        RECT 230.100 196.050 231.900 197.850 ;
        RECT 233.250 191.700 234.450 199.050 ;
        RECT 235.950 197.850 238.050 199.950 ;
        RECT 250.950 197.850 253.050 199.950 ;
        RECT 253.950 199.050 256.050 201.150 ;
        RECT 259.950 199.050 262.050 201.150 ;
        RECT 268.950 197.850 271.050 199.950 ;
        RECT 271.950 199.050 274.050 201.150 ;
        RECT 290.250 199.950 291.300 208.200 ;
        RECT 296.100 204.150 297.900 205.950 ;
        RECT 292.950 201.150 294.750 202.950 ;
        RECT 295.950 202.050 298.050 204.150 ;
        RECT 299.100 201.150 300.900 202.950 ;
        RECT 236.100 196.050 237.900 197.850 ;
        RECT 251.400 193.650 252.600 197.850 ;
        RECT 269.100 196.050 270.900 197.850 ;
        RECT 251.400 192.000 255.900 193.650 ;
        RECT 194.550 190.800 198.150 191.700 ;
        RECT 191.850 183.750 193.650 189.600 ;
        RECT 196.350 183.750 198.150 190.800 ;
        RECT 212.850 190.800 216.450 191.700 ;
        RECT 230.850 190.800 234.450 191.700 ;
        RECT 212.850 183.750 214.650 190.800 ;
        RECT 217.350 183.750 219.150 189.600 ;
        RECT 230.850 183.750 232.650 190.800 ;
        RECT 235.350 183.750 237.150 189.600 ;
        RECT 254.100 183.750 255.900 192.000 ;
        RECT 259.500 183.750 261.300 192.600 ;
        RECT 272.550 191.700 273.750 199.050 ;
        RECT 274.950 197.850 277.050 199.950 ;
        RECT 289.950 197.850 292.050 199.950 ;
        RECT 292.950 199.050 295.050 201.150 ;
        RECT 298.950 199.050 301.050 201.150 ;
        RECT 275.100 196.050 276.900 197.850 ;
        RECT 290.400 193.650 291.600 197.850 ;
        RECT 311.400 196.950 312.600 209.400 ;
        RECT 329.250 209.100 330.450 209.400 ;
        RECT 334.650 209.400 336.450 215.250 ;
        RECT 337.650 209.400 339.450 215.250 ;
        RECT 349.650 209.400 351.450 215.250 ;
        RECT 352.650 210.000 354.450 215.250 ;
        RECT 334.650 209.100 336.300 209.400 ;
        RECT 329.250 208.200 336.300 209.100 ;
        RECT 350.250 209.100 351.450 209.400 ;
        RECT 355.650 209.400 357.450 215.250 ;
        RECT 358.650 209.400 360.450 215.250 ;
        RECT 368.550 209.400 370.350 215.250 ;
        RECT 371.550 209.400 373.350 215.250 ;
        RECT 389.400 209.400 391.200 215.250 ;
        RECT 355.650 209.100 357.300 209.400 ;
        RECT 350.250 208.200 357.300 209.100 ;
        RECT 329.250 199.950 330.300 208.200 ;
        RECT 335.100 204.150 336.900 205.950 ;
        RECT 331.950 201.150 333.750 202.950 ;
        RECT 334.950 202.050 337.050 204.150 ;
        RECT 338.100 201.150 339.900 202.950 ;
        RECT 328.950 197.850 331.050 199.950 ;
        RECT 331.950 199.050 334.050 201.150 ;
        RECT 337.950 199.050 340.050 201.150 ;
        RECT 350.250 199.950 351.300 208.200 ;
        RECT 356.100 204.150 357.900 205.950 ;
        RECT 352.950 201.150 354.750 202.950 ;
        RECT 355.950 202.050 358.050 204.150 ;
        RECT 359.100 201.150 360.900 202.950 ;
        RECT 349.950 197.850 352.050 199.950 ;
        RECT 352.950 199.050 355.050 201.150 ;
        RECT 358.950 199.050 361.050 201.150 ;
        RECT 310.950 194.850 313.050 196.950 ;
        RECT 314.100 195.150 315.900 196.950 ;
        RECT 290.400 192.000 294.900 193.650 ;
        RECT 272.550 190.800 276.150 191.700 ;
        RECT 269.850 183.750 271.650 189.600 ;
        RECT 274.350 183.750 276.150 190.800 ;
        RECT 293.100 183.750 294.900 192.000 ;
        RECT 298.500 183.750 300.300 192.600 ;
        RECT 311.400 186.600 312.600 194.850 ;
        RECT 313.950 193.050 316.050 195.150 ;
        RECT 329.400 193.650 330.600 197.850 ;
        RECT 350.400 193.650 351.600 197.850 ;
        RECT 371.400 196.950 372.600 209.400 ;
        RECT 392.700 203.400 394.500 215.250 ;
        RECT 396.900 203.400 398.700 215.250 ;
        RECT 407.550 204.300 409.350 215.250 ;
        RECT 410.550 205.200 412.350 215.250 ;
        RECT 413.550 204.300 415.350 215.250 ;
        RECT 407.550 203.400 415.350 204.300 ;
        RECT 416.550 203.400 418.350 215.250 ;
        RECT 431.400 209.400 433.200 215.250 ;
        RECT 427.950 205.950 430.050 208.050 ;
        RECT 389.250 201.150 391.050 202.950 ;
        RECT 388.950 199.050 391.050 201.150 ;
        RECT 392.850 198.150 394.050 203.400 ;
        RECT 398.100 198.150 399.900 199.950 ;
        RECT 416.700 198.150 417.900 203.400 ;
        RECT 368.100 195.150 369.900 196.950 ;
        RECT 329.400 192.000 333.900 193.650 ;
        RECT 310.650 183.750 312.450 186.600 ;
        RECT 313.650 183.750 315.450 186.600 ;
        RECT 332.100 183.750 333.900 192.000 ;
        RECT 337.500 183.750 339.300 192.600 ;
        RECT 350.400 192.000 354.900 193.650 ;
        RECT 367.950 193.050 370.050 195.150 ;
        RECT 370.950 194.850 373.050 196.950 ;
        RECT 391.950 196.050 394.050 198.150 ;
        RECT 353.100 183.750 354.900 192.000 ;
        RECT 358.500 183.750 360.300 192.600 ;
        RECT 371.400 186.600 372.600 194.850 ;
        RECT 391.950 192.750 393.150 196.050 ;
        RECT 394.950 194.850 397.050 196.950 ;
        RECT 397.950 196.050 400.050 198.150 ;
        RECT 406.950 194.850 409.050 196.950 ;
        RECT 410.100 195.150 411.900 196.950 ;
        RECT 395.100 193.050 396.900 194.850 ;
        RECT 407.100 193.050 408.900 194.850 ;
        RECT 409.950 193.050 412.050 195.150 ;
        RECT 412.950 194.850 415.050 196.950 ;
        RECT 415.950 196.050 418.050 198.150 ;
        RECT 413.100 193.050 414.900 194.850 ;
        RECT 389.250 191.700 393.000 192.750 ;
        RECT 389.250 189.600 390.450 191.700 ;
        RECT 368.550 183.750 370.350 186.600 ;
        RECT 371.550 183.750 373.350 186.600 ;
        RECT 388.650 183.750 390.450 189.600 ;
        RECT 391.650 188.700 399.450 190.050 ;
        RECT 416.700 189.600 417.900 196.050 ;
        RECT 424.950 192.450 427.050 193.050 ;
        RECT 428.550 192.450 429.450 205.950 ;
        RECT 434.700 203.400 436.500 215.250 ;
        RECT 438.900 203.400 440.700 215.250 ;
        RECT 452.400 209.400 454.200 215.250 ;
        RECT 455.700 203.400 457.500 215.250 ;
        RECT 459.900 203.400 461.700 215.250 ;
        RECT 473.400 209.400 475.200 215.250 ;
        RECT 476.700 203.400 478.500 215.250 ;
        RECT 480.900 203.400 482.700 215.250 ;
        RECT 493.650 209.400 495.450 215.250 ;
        RECT 496.650 209.400 498.450 215.250 ;
        RECT 506.550 209.400 508.350 215.250 ;
        RECT 509.550 209.400 511.350 215.250 ;
        RECT 431.250 201.150 433.050 202.950 ;
        RECT 430.950 199.050 433.050 201.150 ;
        RECT 434.850 198.150 436.050 203.400 ;
        RECT 452.250 201.150 454.050 202.950 ;
        RECT 440.100 198.150 441.900 199.950 ;
        RECT 451.950 199.050 454.050 201.150 ;
        RECT 455.850 198.150 457.050 203.400 ;
        RECT 473.250 201.150 475.050 202.950 ;
        RECT 461.100 198.150 462.900 199.950 ;
        RECT 472.950 199.050 475.050 201.150 ;
        RECT 476.850 198.150 478.050 203.400 ;
        RECT 482.100 198.150 483.900 199.950 ;
        RECT 433.950 196.050 436.050 198.150 ;
        RECT 433.950 192.750 435.150 196.050 ;
        RECT 436.950 194.850 439.050 196.950 ;
        RECT 439.950 196.050 442.050 198.150 ;
        RECT 454.950 196.050 457.050 198.150 ;
        RECT 437.100 193.050 438.900 194.850 ;
        RECT 454.950 192.750 456.150 196.050 ;
        RECT 457.950 194.850 460.050 196.950 ;
        RECT 460.950 196.050 463.050 198.150 ;
        RECT 475.950 196.050 478.050 198.150 ;
        RECT 458.100 193.050 459.900 194.850 ;
        RECT 475.950 192.750 477.150 196.050 ;
        RECT 478.950 194.850 481.050 196.950 ;
        RECT 481.950 196.050 484.050 198.150 ;
        RECT 494.400 196.950 495.600 209.400 ;
        RECT 509.400 196.950 510.600 209.400 ;
        RECT 523.350 203.400 525.150 215.250 ;
        RECT 526.350 203.400 528.150 215.250 ;
        RECT 529.650 209.400 531.450 215.250 ;
        RECT 523.650 198.150 524.850 203.400 ;
        RECT 530.250 202.500 531.450 209.400 ;
        RECT 544.650 203.400 546.450 215.250 ;
        RECT 547.650 204.300 549.450 215.250 ;
        RECT 550.650 205.200 552.450 215.250 ;
        RECT 553.650 204.300 555.450 215.250 ;
        RECT 547.650 203.400 555.450 204.300 ;
        RECT 564.300 203.400 566.100 215.250 ;
        RECT 568.500 203.400 570.300 215.250 ;
        RECT 571.800 209.400 573.600 215.250 ;
        RECT 586.650 209.400 588.450 215.250 ;
        RECT 589.650 209.400 591.450 215.250 ;
        RECT 602.400 209.400 604.200 215.250 ;
        RECT 525.750 201.600 531.450 202.500 ;
        RECT 525.750 200.700 528.000 201.600 ;
        RECT 493.950 194.850 496.050 196.950 ;
        RECT 497.100 195.150 498.900 196.950 ;
        RECT 506.100 195.150 507.900 196.950 ;
        RECT 479.100 193.050 480.900 194.850 ;
        RECT 424.950 191.550 429.450 192.450 ;
        RECT 431.250 191.700 435.000 192.750 ;
        RECT 452.250 191.700 456.000 192.750 ;
        RECT 473.250 191.700 477.000 192.750 ;
        RECT 424.950 190.950 427.050 191.550 ;
        RECT 431.250 189.600 432.450 191.700 ;
        RECT 391.650 183.750 393.450 188.700 ;
        RECT 394.650 183.750 396.450 187.800 ;
        RECT 397.650 183.750 399.450 188.700 ;
        RECT 408.000 183.750 409.800 189.600 ;
        RECT 412.200 187.950 417.900 189.600 ;
        RECT 412.200 183.750 414.000 187.950 ;
        RECT 415.500 183.750 417.300 186.600 ;
        RECT 430.650 183.750 432.450 189.600 ;
        RECT 433.650 188.700 441.450 190.050 ;
        RECT 452.250 189.600 453.450 191.700 ;
        RECT 433.650 183.750 435.450 188.700 ;
        RECT 436.650 183.750 438.450 187.800 ;
        RECT 439.650 183.750 441.450 188.700 ;
        RECT 451.650 183.750 453.450 189.600 ;
        RECT 454.650 188.700 462.450 190.050 ;
        RECT 473.250 189.600 474.450 191.700 ;
        RECT 454.650 183.750 456.450 188.700 ;
        RECT 457.650 183.750 459.450 187.800 ;
        RECT 460.650 183.750 462.450 188.700 ;
        RECT 472.650 183.750 474.450 189.600 ;
        RECT 475.650 188.700 483.450 190.050 ;
        RECT 475.650 183.750 477.450 188.700 ;
        RECT 478.650 183.750 480.450 187.800 ;
        RECT 481.650 183.750 483.450 188.700 ;
        RECT 494.400 186.600 495.600 194.850 ;
        RECT 496.950 193.050 499.050 195.150 ;
        RECT 505.950 193.050 508.050 195.150 ;
        RECT 508.950 194.850 511.050 196.950 ;
        RECT 523.650 196.050 526.050 198.150 ;
        RECT 509.400 186.600 510.600 194.850 ;
        RECT 523.650 189.600 524.850 196.050 ;
        RECT 526.950 192.300 528.000 200.700 ;
        RECT 530.100 198.150 531.900 199.950 ;
        RECT 545.100 198.150 546.300 203.400 ;
        RECT 547.950 201.450 550.050 202.050 ;
        RECT 556.950 201.450 559.050 202.050 ;
        RECT 547.950 200.550 559.050 201.450 ;
        RECT 547.950 199.950 550.050 200.550 ;
        RECT 556.950 199.950 559.050 200.550 ;
        RECT 563.100 198.150 564.900 199.950 ;
        RECT 568.950 198.150 570.150 203.400 ;
        RECT 571.950 201.150 573.750 202.950 ;
        RECT 571.950 199.050 574.050 201.150 ;
        RECT 529.950 196.050 532.050 198.150 ;
        RECT 544.950 196.050 547.050 198.150 ;
        RECT 525.750 191.400 528.000 192.300 ;
        RECT 525.750 190.500 530.850 191.400 ;
        RECT 493.650 183.750 495.450 186.600 ;
        RECT 496.650 183.750 498.450 186.600 ;
        RECT 506.550 183.750 508.350 186.600 ;
        RECT 509.550 183.750 511.350 186.600 ;
        RECT 523.350 183.750 525.150 189.600 ;
        RECT 526.350 183.750 528.150 189.600 ;
        RECT 529.650 186.600 530.850 190.500 ;
        RECT 545.100 189.600 546.300 196.050 ;
        RECT 547.950 194.850 550.050 196.950 ;
        RECT 551.100 195.150 552.900 196.950 ;
        RECT 548.100 193.050 549.900 194.850 ;
        RECT 550.950 193.050 553.050 195.150 ;
        RECT 553.950 194.850 556.050 196.950 ;
        RECT 562.950 196.050 565.050 198.150 ;
        RECT 565.950 194.850 568.050 196.950 ;
        RECT 568.950 196.050 571.050 198.150 ;
        RECT 587.400 196.950 588.600 209.400 ;
        RECT 605.700 203.400 607.500 215.250 ;
        RECT 609.900 203.400 611.700 215.250 ;
        RECT 623.400 209.400 625.200 215.250 ;
        RECT 626.700 203.400 628.500 215.250 ;
        RECT 630.900 203.400 632.700 215.250 ;
        RECT 643.650 203.400 645.450 215.250 ;
        RECT 646.650 204.300 648.450 215.250 ;
        RECT 649.650 205.200 651.450 215.250 ;
        RECT 652.650 204.300 654.450 215.250 ;
        RECT 665.400 209.400 667.200 215.250 ;
        RECT 646.650 203.400 654.450 204.300 ;
        RECT 668.700 203.400 670.500 215.250 ;
        RECT 672.900 203.400 674.700 215.250 ;
        RECT 687.300 203.400 689.100 215.250 ;
        RECT 691.500 203.400 693.300 215.250 ;
        RECT 694.800 209.400 696.600 215.250 ;
        RECT 707.550 209.400 709.350 215.250 ;
        RECT 710.550 209.400 712.350 215.250 ;
        RECT 713.550 209.400 715.350 215.250 ;
        RECT 602.250 201.150 604.050 202.950 ;
        RECT 601.950 199.050 604.050 201.150 ;
        RECT 605.850 198.150 607.050 203.400 ;
        RECT 623.250 201.150 625.050 202.950 ;
        RECT 611.100 198.150 612.900 199.950 ;
        RECT 622.950 199.050 625.050 201.150 ;
        RECT 626.850 198.150 628.050 203.400 ;
        RECT 632.100 198.150 633.900 199.950 ;
        RECT 644.100 198.150 645.300 203.400 ;
        RECT 665.250 201.150 667.050 202.950 ;
        RECT 664.950 199.050 667.050 201.150 ;
        RECT 668.850 198.150 670.050 203.400 ;
        RECT 674.100 198.150 675.900 199.950 ;
        RECT 686.100 198.150 687.900 199.950 ;
        RECT 691.950 198.150 693.150 203.400 ;
        RECT 694.950 201.150 696.750 202.950 ;
        RECT 710.550 201.150 711.750 209.400 ;
        RECT 726.300 203.400 728.100 215.250 ;
        RECT 730.500 203.400 732.300 215.250 ;
        RECT 733.800 209.400 735.600 215.250 ;
        RECT 746.550 203.400 748.350 215.250 ;
        RECT 750.750 203.400 752.550 215.250 ;
        RECT 764.550 209.400 766.350 215.250 ;
        RECT 767.550 209.400 769.350 215.250 ;
        RECT 770.550 209.400 772.350 215.250 ;
        RECT 784.650 209.400 786.450 215.250 ;
        RECT 787.650 209.400 789.450 215.250 ;
        RECT 790.650 209.400 792.450 215.250 ;
        RECT 803.400 209.400 805.200 215.250 ;
        RECT 694.950 199.050 697.050 201.150 ;
        RECT 554.100 193.050 555.900 194.850 ;
        RECT 566.100 193.050 567.900 194.850 ;
        RECT 569.850 192.750 571.050 196.050 ;
        RECT 586.950 194.850 589.050 196.950 ;
        RECT 590.100 195.150 591.900 196.950 ;
        RECT 604.950 196.050 607.050 198.150 ;
        RECT 570.000 191.700 573.750 192.750 ;
        RECT 545.100 187.950 550.800 189.600 ;
        RECT 529.650 183.750 531.450 186.600 ;
        RECT 545.700 183.750 547.500 186.600 ;
        RECT 549.000 183.750 550.800 187.950 ;
        RECT 553.200 183.750 555.000 189.600 ;
        RECT 563.550 188.700 571.350 190.050 ;
        RECT 563.550 183.750 565.350 188.700 ;
        RECT 566.550 183.750 568.350 187.800 ;
        RECT 569.550 183.750 571.350 188.700 ;
        RECT 572.550 189.600 573.750 191.700 ;
        RECT 572.550 183.750 574.350 189.600 ;
        RECT 587.400 186.600 588.600 194.850 ;
        RECT 589.950 193.050 592.050 195.150 ;
        RECT 604.950 192.750 606.150 196.050 ;
        RECT 607.950 194.850 610.050 196.950 ;
        RECT 610.950 196.050 613.050 198.150 ;
        RECT 625.950 196.050 628.050 198.150 ;
        RECT 608.100 193.050 609.900 194.850 ;
        RECT 625.950 192.750 627.150 196.050 ;
        RECT 628.950 194.850 631.050 196.950 ;
        RECT 631.950 196.050 634.050 198.150 ;
        RECT 643.950 196.050 646.050 198.150 ;
        RECT 629.100 193.050 630.900 194.850 ;
        RECT 602.250 191.700 606.000 192.750 ;
        RECT 623.250 191.700 627.000 192.750 ;
        RECT 602.250 189.600 603.450 191.700 ;
        RECT 586.650 183.750 588.450 186.600 ;
        RECT 589.650 183.750 591.450 186.600 ;
        RECT 601.650 183.750 603.450 189.600 ;
        RECT 604.650 188.700 612.450 190.050 ;
        RECT 623.250 189.600 624.450 191.700 ;
        RECT 604.650 183.750 606.450 188.700 ;
        RECT 607.650 183.750 609.450 187.800 ;
        RECT 610.650 183.750 612.450 188.700 ;
        RECT 622.650 183.750 624.450 189.600 ;
        RECT 625.650 188.700 633.450 190.050 ;
        RECT 625.650 183.750 627.450 188.700 ;
        RECT 628.650 183.750 630.450 187.800 ;
        RECT 631.650 183.750 633.450 188.700 ;
        RECT 644.100 189.600 645.300 196.050 ;
        RECT 646.950 194.850 649.050 196.950 ;
        RECT 650.100 195.150 651.900 196.950 ;
        RECT 647.100 193.050 648.900 194.850 ;
        RECT 649.950 193.050 652.050 195.150 ;
        RECT 652.950 194.850 655.050 196.950 ;
        RECT 667.950 196.050 670.050 198.150 ;
        RECT 653.100 193.050 654.900 194.850 ;
        RECT 667.950 192.750 669.150 196.050 ;
        RECT 670.950 194.850 673.050 196.950 ;
        RECT 673.950 196.050 676.050 198.150 ;
        RECT 685.950 196.050 688.050 198.150 ;
        RECT 688.950 194.850 691.050 196.950 ;
        RECT 691.950 196.050 694.050 198.150 ;
        RECT 706.950 197.850 709.050 199.950 ;
        RECT 709.950 199.050 712.050 201.150 ;
        RECT 707.100 196.050 708.900 197.850 ;
        RECT 671.100 193.050 672.900 194.850 ;
        RECT 689.100 193.050 690.900 194.850 ;
        RECT 692.850 192.750 694.050 196.050 ;
        RECT 665.250 191.700 669.000 192.750 ;
        RECT 693.000 191.700 696.750 192.750 ;
        RECT 665.250 189.600 666.450 191.700 ;
        RECT 644.100 187.950 649.800 189.600 ;
        RECT 644.700 183.750 646.500 186.600 ;
        RECT 648.000 183.750 649.800 187.950 ;
        RECT 652.200 183.750 654.000 189.600 ;
        RECT 664.650 183.750 666.450 189.600 ;
        RECT 667.650 188.700 675.450 190.050 ;
        RECT 667.650 183.750 669.450 188.700 ;
        RECT 670.650 183.750 672.450 187.800 ;
        RECT 673.650 183.750 675.450 188.700 ;
        RECT 686.550 188.700 694.350 190.050 ;
        RECT 686.550 183.750 688.350 188.700 ;
        RECT 689.550 183.750 691.350 187.800 ;
        RECT 692.550 183.750 694.350 188.700 ;
        RECT 695.550 189.600 696.750 191.700 ;
        RECT 710.550 191.700 711.750 199.050 ;
        RECT 712.950 197.850 715.050 199.950 ;
        RECT 725.100 198.150 726.900 199.950 ;
        RECT 730.950 198.150 732.150 203.400 ;
        RECT 733.950 201.150 735.750 202.950 ;
        RECT 750.000 202.350 752.550 203.400 ;
        RECT 733.950 199.050 736.050 201.150 ;
        RECT 746.100 198.150 747.900 199.950 ;
        RECT 713.100 196.050 714.900 197.850 ;
        RECT 724.950 196.050 727.050 198.150 ;
        RECT 727.950 194.850 730.050 196.950 ;
        RECT 730.950 196.050 733.050 198.150 ;
        RECT 745.950 196.050 748.050 198.150 ;
        RECT 728.100 193.050 729.900 194.850 ;
        RECT 731.850 192.750 733.050 196.050 ;
        RECT 750.000 195.150 751.050 202.350 ;
        RECT 767.550 201.150 768.750 209.400 ;
        RECT 788.250 201.150 789.450 209.400 ;
        RECT 806.700 203.400 808.500 215.250 ;
        RECT 810.900 203.400 812.700 215.250 ;
        RECT 822.300 203.400 824.100 215.250 ;
        RECT 826.500 203.400 828.300 215.250 ;
        RECT 829.800 209.400 831.600 215.250 ;
        RECT 846.300 203.400 848.100 215.250 ;
        RECT 850.500 203.400 852.300 215.250 ;
        RECT 853.800 209.400 855.600 215.250 ;
        RECT 803.250 201.150 805.050 202.950 ;
        RECT 752.100 198.150 753.900 199.950 ;
        RECT 751.950 196.050 754.050 198.150 ;
        RECT 763.950 197.850 766.050 199.950 ;
        RECT 766.950 199.050 769.050 201.150 ;
        RECT 764.100 196.050 765.900 197.850 ;
        RECT 748.950 193.050 751.050 195.150 ;
        RECT 732.000 191.700 735.750 192.750 ;
        RECT 710.550 190.800 714.150 191.700 ;
        RECT 695.550 183.750 697.350 189.600 ;
        RECT 707.850 183.750 709.650 189.600 ;
        RECT 712.350 183.750 714.150 190.800 ;
        RECT 725.550 188.700 733.350 190.050 ;
        RECT 725.550 183.750 727.350 188.700 ;
        RECT 728.550 183.750 730.350 187.800 ;
        RECT 731.550 183.750 733.350 188.700 ;
        RECT 734.550 189.600 735.750 191.700 ;
        RECT 734.550 183.750 736.350 189.600 ;
        RECT 750.000 186.600 751.050 193.050 ;
        RECT 767.550 191.700 768.750 199.050 ;
        RECT 769.950 197.850 772.050 199.950 ;
        RECT 784.950 197.850 787.050 199.950 ;
        RECT 787.950 199.050 790.050 201.150 ;
        RECT 770.100 196.050 771.900 197.850 ;
        RECT 785.100 196.050 786.900 197.850 ;
        RECT 788.250 191.700 789.450 199.050 ;
        RECT 790.950 197.850 793.050 199.950 ;
        RECT 802.950 199.050 805.050 201.150 ;
        RECT 806.850 198.150 808.050 203.400 ;
        RECT 812.100 198.150 813.900 199.950 ;
        RECT 821.100 198.150 822.900 199.950 ;
        RECT 826.950 198.150 828.150 203.400 ;
        RECT 829.950 201.150 831.750 202.950 ;
        RECT 829.950 199.050 832.050 201.150 ;
        RECT 845.100 198.150 846.900 199.950 ;
        RECT 850.950 198.150 852.150 203.400 ;
        RECT 853.950 201.150 855.750 202.950 ;
        RECT 853.950 199.050 856.050 201.150 ;
        RECT 791.100 196.050 792.900 197.850 ;
        RECT 805.950 196.050 808.050 198.150 ;
        RECT 805.950 192.750 807.150 196.050 ;
        RECT 808.950 194.850 811.050 196.950 ;
        RECT 811.950 196.050 814.050 198.150 ;
        RECT 820.950 196.050 823.050 198.150 ;
        RECT 823.950 194.850 826.050 196.950 ;
        RECT 826.950 196.050 829.050 198.150 ;
        RECT 844.950 196.050 847.050 198.150 ;
        RECT 809.100 193.050 810.900 194.850 ;
        RECT 824.100 193.050 825.900 194.850 ;
        RECT 827.850 192.750 829.050 196.050 ;
        RECT 847.950 194.850 850.050 196.950 ;
        RECT 850.950 196.050 853.050 198.150 ;
        RECT 848.100 193.050 849.900 194.850 ;
        RECT 851.850 192.750 853.050 196.050 ;
        RECT 767.550 190.800 771.150 191.700 ;
        RECT 746.550 183.750 748.350 186.600 ;
        RECT 749.550 183.750 751.350 186.600 ;
        RECT 752.550 183.750 754.350 186.600 ;
        RECT 764.850 183.750 766.650 189.600 ;
        RECT 769.350 183.750 771.150 190.800 ;
        RECT 785.850 190.800 789.450 191.700 ;
        RECT 803.250 191.700 807.000 192.750 ;
        RECT 828.000 191.700 831.750 192.750 ;
        RECT 852.000 191.700 855.750 192.750 ;
        RECT 785.850 183.750 787.650 190.800 ;
        RECT 803.250 189.600 804.450 191.700 ;
        RECT 790.350 183.750 792.150 189.600 ;
        RECT 802.650 183.750 804.450 189.600 ;
        RECT 805.650 188.700 813.450 190.050 ;
        RECT 805.650 183.750 807.450 188.700 ;
        RECT 808.650 183.750 810.450 187.800 ;
        RECT 811.650 183.750 813.450 188.700 ;
        RECT 821.550 188.700 829.350 190.050 ;
        RECT 821.550 183.750 823.350 188.700 ;
        RECT 824.550 183.750 826.350 187.800 ;
        RECT 827.550 183.750 829.350 188.700 ;
        RECT 830.550 189.600 831.750 191.700 ;
        RECT 830.550 183.750 832.350 189.600 ;
        RECT 845.550 188.700 853.350 190.050 ;
        RECT 845.550 183.750 847.350 188.700 ;
        RECT 848.550 183.750 850.350 187.800 ;
        RECT 851.550 183.750 853.350 188.700 ;
        RECT 854.550 189.600 855.750 191.700 ;
        RECT 854.550 183.750 856.350 189.600 ;
        RECT 10.650 176.400 12.450 179.250 ;
        RECT 13.650 176.400 15.450 179.250 ;
        RECT 11.400 168.150 12.600 176.400 ;
        RECT 24.000 173.400 25.800 179.250 ;
        RECT 28.200 175.050 30.000 179.250 ;
        RECT 31.500 176.400 33.300 179.250 ;
        RECT 28.200 173.400 33.900 175.050 ;
        RECT 10.950 166.050 13.050 168.150 ;
        RECT 13.950 167.850 16.050 169.950 ;
        RECT 23.100 168.150 24.900 169.950 ;
        RECT 14.100 166.050 15.900 167.850 ;
        RECT 22.950 166.050 25.050 168.150 ;
        RECT 25.950 167.850 28.050 169.950 ;
        RECT 29.100 168.150 30.900 169.950 ;
        RECT 26.100 166.050 27.900 167.850 ;
        RECT 28.950 166.050 31.050 168.150 ;
        RECT 32.700 166.950 33.900 173.400 ;
        RECT 44.550 174.300 46.350 179.250 ;
        RECT 47.550 175.200 49.350 179.250 ;
        RECT 50.550 174.300 52.350 179.250 ;
        RECT 44.550 172.950 52.350 174.300 ;
        RECT 53.550 173.400 55.350 179.250 ;
        RECT 65.550 174.300 67.350 179.250 ;
        RECT 68.550 175.200 70.350 179.250 ;
        RECT 71.550 174.300 73.350 179.250 ;
        RECT 53.550 171.300 54.750 173.400 ;
        RECT 65.550 172.950 73.350 174.300 ;
        RECT 74.550 173.400 76.350 179.250 ;
        RECT 74.550 171.300 75.750 173.400 ;
        RECT 51.000 170.250 54.750 171.300 ;
        RECT 72.000 170.250 75.750 171.300 ;
        RECT 92.100 171.000 93.900 179.250 ;
        RECT 47.100 168.150 48.900 169.950 ;
        RECT 11.400 153.600 12.600 166.050 ;
        RECT 31.950 164.850 34.050 166.950 ;
        RECT 43.950 164.850 46.050 166.950 ;
        RECT 46.950 166.050 49.050 168.150 ;
        RECT 50.850 166.950 52.050 170.250 ;
        RECT 68.100 168.150 69.900 169.950 ;
        RECT 49.950 164.850 52.050 166.950 ;
        RECT 64.950 164.850 67.050 166.950 ;
        RECT 67.950 166.050 70.050 168.150 ;
        RECT 71.850 166.950 73.050 170.250 ;
        RECT 70.950 164.850 73.050 166.950 ;
        RECT 89.400 169.350 93.900 171.000 ;
        RECT 97.500 170.400 99.300 179.250 ;
        RECT 107.550 174.300 109.350 179.250 ;
        RECT 110.550 175.200 112.350 179.250 ;
        RECT 113.550 174.300 115.350 179.250 ;
        RECT 107.550 172.950 115.350 174.300 ;
        RECT 116.550 173.400 118.350 179.250 ;
        RECT 132.000 173.400 133.800 179.250 ;
        RECT 136.200 175.050 138.000 179.250 ;
        RECT 139.500 176.400 141.300 179.250 ;
        RECT 136.200 173.400 141.900 175.050 ;
        RECT 154.650 173.400 156.450 179.250 ;
        RECT 116.550 171.300 117.750 173.400 ;
        RECT 114.000 170.250 117.750 171.300 ;
        RECT 89.400 165.150 90.600 169.350 ;
        RECT 110.100 168.150 111.900 169.950 ;
        RECT 32.700 159.600 33.900 164.850 ;
        RECT 44.100 163.050 45.900 164.850 ;
        RECT 49.950 159.600 51.150 164.850 ;
        RECT 52.950 161.850 55.050 163.950 ;
        RECT 65.100 163.050 66.900 164.850 ;
        RECT 52.950 160.050 54.750 161.850 ;
        RECT 70.950 159.600 72.150 164.850 ;
        RECT 73.950 161.850 76.050 163.950 ;
        RECT 88.950 163.050 91.050 165.150 ;
        RECT 106.950 164.850 109.050 166.950 ;
        RECT 109.950 166.050 112.050 168.150 ;
        RECT 113.850 166.950 115.050 170.250 ;
        RECT 131.100 168.150 132.900 169.950 ;
        RECT 112.950 164.850 115.050 166.950 ;
        RECT 130.950 166.050 133.050 168.150 ;
        RECT 133.950 167.850 136.050 169.950 ;
        RECT 137.100 168.150 138.900 169.950 ;
        RECT 134.100 166.050 135.900 167.850 ;
        RECT 136.950 166.050 139.050 168.150 ;
        RECT 140.700 166.950 141.900 173.400 ;
        RECT 155.250 171.300 156.450 173.400 ;
        RECT 157.650 174.300 159.450 179.250 ;
        RECT 160.650 175.200 162.450 179.250 ;
        RECT 163.650 174.300 165.450 179.250 ;
        RECT 175.650 176.400 177.450 179.250 ;
        RECT 178.650 176.400 180.450 179.250 ;
        RECT 157.650 172.950 165.450 174.300 ;
        RECT 155.250 170.250 159.000 171.300 ;
        RECT 157.950 166.950 159.150 170.250 ;
        RECT 161.100 168.150 162.900 169.950 ;
        RECT 176.400 168.150 177.600 176.400 ;
        RECT 189.000 173.400 190.800 179.250 ;
        RECT 193.200 175.050 195.000 179.250 ;
        RECT 196.500 176.400 198.300 179.250 ;
        RECT 211.650 176.400 213.450 179.250 ;
        RECT 214.650 176.400 216.450 179.250 ;
        RECT 226.650 176.400 228.450 179.250 ;
        RECT 229.650 176.400 231.450 179.250 ;
        RECT 232.650 176.400 234.450 179.250 ;
        RECT 245.550 176.400 247.350 179.250 ;
        RECT 248.550 176.400 250.350 179.250 ;
        RECT 193.200 173.400 198.900 175.050 ;
        RECT 139.950 164.850 142.050 166.950 ;
        RECT 157.950 164.850 160.050 166.950 ;
        RECT 160.950 166.050 163.050 168.150 ;
        RECT 163.950 164.850 166.050 166.950 ;
        RECT 175.950 166.050 178.050 168.150 ;
        RECT 178.950 167.850 181.050 169.950 ;
        RECT 188.100 168.150 189.900 169.950 ;
        RECT 179.100 166.050 180.900 167.850 ;
        RECT 187.950 166.050 190.050 168.150 ;
        RECT 190.950 167.850 193.050 169.950 ;
        RECT 194.100 168.150 195.900 169.950 ;
        RECT 191.100 166.050 192.900 167.850 ;
        RECT 193.950 166.050 196.050 168.150 ;
        RECT 197.700 166.950 198.900 173.400 ;
        RECT 212.400 168.150 213.600 176.400 ;
        RECT 229.950 169.950 231.000 176.400 ;
        RECT 73.950 160.050 75.750 161.850 ;
        RECT 23.550 158.700 31.350 159.600 ;
        RECT 10.650 147.750 12.450 153.600 ;
        RECT 13.650 147.750 15.450 153.600 ;
        RECT 23.550 147.750 25.350 158.700 ;
        RECT 26.550 147.750 28.350 157.800 ;
        RECT 29.550 147.750 31.350 158.700 ;
        RECT 32.550 147.750 34.350 159.600 ;
        RECT 45.300 147.750 47.100 159.600 ;
        RECT 49.500 147.750 51.300 159.600 ;
        RECT 52.800 147.750 54.600 153.600 ;
        RECT 66.300 147.750 68.100 159.600 ;
        RECT 70.500 147.750 72.300 159.600 ;
        RECT 89.250 154.800 90.300 163.050 ;
        RECT 91.950 161.850 94.050 163.950 ;
        RECT 97.950 161.850 100.050 163.950 ;
        RECT 107.100 163.050 108.900 164.850 ;
        RECT 91.950 160.050 93.750 161.850 ;
        RECT 94.950 158.850 97.050 160.950 ;
        RECT 98.100 160.050 99.900 161.850 ;
        RECT 112.950 159.600 114.150 164.850 ;
        RECT 115.950 161.850 118.050 163.950 ;
        RECT 115.950 160.050 117.750 161.850 ;
        RECT 140.700 159.600 141.900 164.850 ;
        RECT 154.950 161.850 157.050 163.950 ;
        RECT 155.250 160.050 157.050 161.850 ;
        RECT 158.850 159.600 160.050 164.850 ;
        RECT 164.100 163.050 165.900 164.850 ;
        RECT 166.950 162.450 169.050 163.050 ;
        RECT 172.950 162.450 175.050 163.050 ;
        RECT 166.950 161.550 175.050 162.450 ;
        RECT 166.950 160.950 169.050 161.550 ;
        RECT 172.950 160.950 175.050 161.550 ;
        RECT 95.100 157.050 96.900 158.850 ;
        RECT 89.250 153.900 96.300 154.800 ;
        RECT 89.250 153.600 90.450 153.900 ;
        RECT 73.800 147.750 75.600 153.600 ;
        RECT 88.650 147.750 90.450 153.600 ;
        RECT 94.650 153.600 96.300 153.900 ;
        RECT 91.650 147.750 93.450 153.000 ;
        RECT 94.650 147.750 96.450 153.600 ;
        RECT 97.650 147.750 99.450 153.600 ;
        RECT 108.300 147.750 110.100 159.600 ;
        RECT 112.500 147.750 114.300 159.600 ;
        RECT 131.550 158.700 139.350 159.600 ;
        RECT 115.800 147.750 117.600 153.600 ;
        RECT 131.550 147.750 133.350 158.700 ;
        RECT 134.550 147.750 136.350 157.800 ;
        RECT 137.550 147.750 139.350 158.700 ;
        RECT 140.550 147.750 142.350 159.600 ;
        RECT 155.400 147.750 157.200 153.600 ;
        RECT 158.700 147.750 160.500 159.600 ;
        RECT 162.900 147.750 164.700 159.600 ;
        RECT 176.400 153.600 177.600 166.050 ;
        RECT 196.950 164.850 199.050 166.950 ;
        RECT 211.950 166.050 214.050 168.150 ;
        RECT 214.950 167.850 217.050 169.950 ;
        RECT 229.950 167.850 232.050 169.950 ;
        RECT 244.950 167.850 247.050 169.950 ;
        RECT 248.400 168.150 249.600 176.400 ;
        RECT 266.100 171.000 267.900 179.250 ;
        RECT 263.400 169.350 267.900 171.000 ;
        RECT 271.500 170.400 273.300 179.250 ;
        RECT 284.850 172.200 286.650 179.250 ;
        RECT 289.350 173.400 291.150 179.250 ;
        RECT 301.650 173.400 303.450 179.250 ;
        RECT 284.850 171.300 288.450 172.200 ;
        RECT 215.100 166.050 216.900 167.850 ;
        RECT 197.700 159.600 198.900 164.850 ;
        RECT 188.550 158.700 196.350 159.600 ;
        RECT 175.650 147.750 177.450 153.600 ;
        RECT 178.650 147.750 180.450 153.600 ;
        RECT 188.550 147.750 190.350 158.700 ;
        RECT 191.550 147.750 193.350 157.800 ;
        RECT 194.550 147.750 196.350 158.700 ;
        RECT 197.550 147.750 199.350 159.600 ;
        RECT 212.400 153.600 213.600 166.050 ;
        RECT 226.950 164.850 229.050 166.950 ;
        RECT 227.100 163.050 228.900 164.850 ;
        RECT 229.950 160.650 231.000 167.850 ;
        RECT 232.950 164.850 235.050 166.950 ;
        RECT 245.100 166.050 246.900 167.850 ;
        RECT 247.950 166.050 250.050 168.150 ;
        RECT 233.100 163.050 234.900 164.850 ;
        RECT 228.450 159.600 231.000 160.650 ;
        RECT 211.650 147.750 213.450 153.600 ;
        RECT 214.650 147.750 216.450 153.600 ;
        RECT 228.450 147.750 230.250 159.600 ;
        RECT 232.650 147.750 234.450 159.600 ;
        RECT 248.400 153.600 249.600 166.050 ;
        RECT 263.400 165.150 264.600 169.350 ;
        RECT 271.950 168.450 274.050 169.050 ;
        RECT 277.950 168.450 280.050 169.050 ;
        RECT 271.950 167.550 280.050 168.450 ;
        RECT 271.950 166.950 274.050 167.550 ;
        RECT 277.950 166.950 280.050 167.550 ;
        RECT 284.100 165.150 285.900 166.950 ;
        RECT 262.950 163.050 265.050 165.150 ;
        RECT 263.250 154.800 264.300 163.050 ;
        RECT 265.950 161.850 268.050 163.950 ;
        RECT 271.950 161.850 274.050 163.950 ;
        RECT 283.950 163.050 286.050 165.150 ;
        RECT 287.250 163.950 288.450 171.300 ;
        RECT 302.250 171.300 303.450 173.400 ;
        RECT 304.650 174.300 306.450 179.250 ;
        RECT 307.650 175.200 309.450 179.250 ;
        RECT 310.650 174.300 312.450 179.250 ;
        RECT 304.650 172.950 312.450 174.300 ;
        RECT 302.250 170.250 306.000 171.300 ;
        RECT 326.100 171.000 327.900 179.250 ;
        RECT 304.950 166.950 306.150 170.250 ;
        RECT 308.100 168.150 309.900 169.950 ;
        RECT 323.400 169.350 327.900 171.000 ;
        RECT 331.500 170.400 333.300 179.250 ;
        RECT 347.100 171.000 348.900 179.250 ;
        RECT 344.400 169.350 348.900 171.000 ;
        RECT 352.500 170.400 354.300 179.250 ;
        RECT 364.650 173.400 366.450 179.250 ;
        RECT 365.250 171.300 366.450 173.400 ;
        RECT 367.650 174.300 369.450 179.250 ;
        RECT 370.650 175.200 372.450 179.250 ;
        RECT 373.650 174.300 375.450 179.250 ;
        RECT 367.650 172.950 375.450 174.300 ;
        RECT 365.250 170.250 369.000 171.300 ;
        RECT 389.100 171.000 390.900 179.250 ;
        RECT 290.100 165.150 291.900 166.950 ;
        RECT 286.950 161.850 289.050 163.950 ;
        RECT 289.950 163.050 292.050 165.150 ;
        RECT 304.950 164.850 307.050 166.950 ;
        RECT 307.950 166.050 310.050 168.150 ;
        RECT 310.950 164.850 313.050 166.950 ;
        RECT 323.400 165.150 324.600 169.350 ;
        RECT 344.400 165.150 345.600 169.350 ;
        RECT 367.950 166.950 369.150 170.250 ;
        RECT 371.100 168.150 372.900 169.950 ;
        RECT 386.400 169.350 390.900 171.000 ;
        RECT 394.500 170.400 396.300 179.250 ;
        RECT 407.550 176.400 409.350 179.250 ;
        RECT 410.550 176.400 412.350 179.250 ;
        RECT 422.550 176.400 424.350 179.250 ;
        RECT 425.550 176.400 427.350 179.250 ;
        RECT 428.550 176.400 430.350 179.250 ;
        RECT 440.550 176.400 442.350 179.250 ;
        RECT 443.550 176.400 445.350 179.250 ;
        RECT 446.550 176.400 448.350 179.250 ;
        RECT 301.950 161.850 304.050 163.950 ;
        RECT 265.950 160.050 267.750 161.850 ;
        RECT 268.950 158.850 271.050 160.950 ;
        RECT 272.100 160.050 273.900 161.850 ;
        RECT 269.100 157.050 270.900 158.850 ;
        RECT 263.250 153.900 270.300 154.800 ;
        RECT 263.250 153.600 264.450 153.900 ;
        RECT 245.550 147.750 247.350 153.600 ;
        RECT 248.550 147.750 250.350 153.600 ;
        RECT 262.650 147.750 264.450 153.600 ;
        RECT 268.650 153.600 270.300 153.900 ;
        RECT 287.250 153.600 288.450 161.850 ;
        RECT 302.250 160.050 304.050 161.850 ;
        RECT 305.850 159.600 307.050 164.850 ;
        RECT 311.100 163.050 312.900 164.850 ;
        RECT 322.950 163.050 325.050 165.150 ;
        RECT 265.650 147.750 267.450 153.000 ;
        RECT 268.650 147.750 270.450 153.600 ;
        RECT 271.650 147.750 273.450 153.600 ;
        RECT 283.650 147.750 285.450 153.600 ;
        RECT 286.650 147.750 288.450 153.600 ;
        RECT 289.650 147.750 291.450 153.600 ;
        RECT 302.400 147.750 304.200 153.600 ;
        RECT 305.700 147.750 307.500 159.600 ;
        RECT 309.900 147.750 311.700 159.600 ;
        RECT 323.250 154.800 324.300 163.050 ;
        RECT 325.950 161.850 328.050 163.950 ;
        RECT 331.950 161.850 334.050 163.950 ;
        RECT 343.950 163.050 346.050 165.150 ;
        RECT 367.950 164.850 370.050 166.950 ;
        RECT 370.950 166.050 373.050 168.150 ;
        RECT 373.950 164.850 376.050 166.950 ;
        RECT 386.400 165.150 387.600 169.350 ;
        RECT 406.950 167.850 409.050 169.950 ;
        RECT 410.400 168.150 411.600 176.400 ;
        RECT 426.000 169.950 427.050 176.400 ;
        RECT 444.000 169.950 445.050 176.400 ;
        RECT 458.550 171.900 460.350 179.250 ;
        RECT 463.050 173.400 464.850 179.250 ;
        RECT 466.050 174.900 467.850 179.250 ;
        RECT 481.650 176.400 483.450 179.250 ;
        RECT 484.650 176.400 486.450 179.250 ;
        RECT 487.650 176.400 489.450 179.250 ;
        RECT 502.650 176.400 504.450 179.250 ;
        RECT 505.650 176.400 507.450 179.250 ;
        RECT 508.650 176.400 510.450 179.250 ;
        RECT 520.650 176.400 522.450 179.250 ;
        RECT 523.650 176.400 525.450 179.250 ;
        RECT 466.050 173.400 469.350 174.900 ;
        RECT 464.250 171.900 466.050 172.500 ;
        RECT 458.550 170.700 466.050 171.900 ;
        RECT 407.100 166.050 408.900 167.850 ;
        RECT 409.950 166.050 412.050 168.150 ;
        RECT 424.950 167.850 427.050 169.950 ;
        RECT 442.950 167.850 445.050 169.950 ;
        RECT 325.950 160.050 327.750 161.850 ;
        RECT 328.950 158.850 331.050 160.950 ;
        RECT 332.100 160.050 333.900 161.850 ;
        RECT 329.100 157.050 330.900 158.850 ;
        RECT 344.250 154.800 345.300 163.050 ;
        RECT 346.950 161.850 349.050 163.950 ;
        RECT 352.950 161.850 355.050 163.950 ;
        RECT 364.950 161.850 367.050 163.950 ;
        RECT 346.950 160.050 348.750 161.850 ;
        RECT 349.950 158.850 352.050 160.950 ;
        RECT 353.100 160.050 354.900 161.850 ;
        RECT 365.250 160.050 367.050 161.850 ;
        RECT 368.850 159.600 370.050 164.850 ;
        RECT 374.100 163.050 375.900 164.850 ;
        RECT 385.950 163.050 388.050 165.150 ;
        RECT 350.100 157.050 351.900 158.850 ;
        RECT 323.250 153.900 330.300 154.800 ;
        RECT 323.250 153.600 324.450 153.900 ;
        RECT 322.650 147.750 324.450 153.600 ;
        RECT 328.650 153.600 330.300 153.900 ;
        RECT 344.250 153.900 351.300 154.800 ;
        RECT 344.250 153.600 345.450 153.900 ;
        RECT 325.650 147.750 327.450 153.000 ;
        RECT 328.650 147.750 330.450 153.600 ;
        RECT 331.650 147.750 333.450 153.600 ;
        RECT 343.650 147.750 345.450 153.600 ;
        RECT 349.650 153.600 351.300 153.900 ;
        RECT 346.650 147.750 348.450 153.000 ;
        RECT 349.650 147.750 351.450 153.600 ;
        RECT 352.650 147.750 354.450 153.600 ;
        RECT 365.400 147.750 367.200 153.600 ;
        RECT 368.700 147.750 370.500 159.600 ;
        RECT 372.900 147.750 374.700 159.600 ;
        RECT 386.250 154.800 387.300 163.050 ;
        RECT 388.950 161.850 391.050 163.950 ;
        RECT 394.950 161.850 397.050 163.950 ;
        RECT 388.950 160.050 390.750 161.850 ;
        RECT 391.950 158.850 394.050 160.950 ;
        RECT 395.100 160.050 396.900 161.850 ;
        RECT 392.100 157.050 393.900 158.850 ;
        RECT 386.250 153.900 393.300 154.800 ;
        RECT 386.250 153.600 387.450 153.900 ;
        RECT 385.650 147.750 387.450 153.600 ;
        RECT 391.650 153.600 393.300 153.900 ;
        RECT 410.400 153.600 411.600 166.050 ;
        RECT 421.950 164.850 424.050 166.950 ;
        RECT 422.100 163.050 423.900 164.850 ;
        RECT 426.000 160.650 427.050 167.850 ;
        RECT 427.950 164.850 430.050 166.950 ;
        RECT 439.950 164.850 442.050 166.950 ;
        RECT 428.100 163.050 429.900 164.850 ;
        RECT 440.100 163.050 441.900 164.850 ;
        RECT 444.000 160.650 445.050 167.850 ;
        RECT 445.950 164.850 448.050 166.950 ;
        RECT 457.950 164.850 460.050 166.950 ;
        RECT 446.100 163.050 447.900 164.850 ;
        RECT 458.100 163.050 459.900 164.850 ;
        RECT 426.000 159.600 428.550 160.650 ;
        RECT 444.000 159.600 446.550 160.650 ;
        RECT 388.650 147.750 390.450 153.000 ;
        RECT 391.650 147.750 393.450 153.600 ;
        RECT 394.650 147.750 396.450 153.600 ;
        RECT 407.550 147.750 409.350 153.600 ;
        RECT 410.550 147.750 412.350 153.600 ;
        RECT 422.550 147.750 424.350 159.600 ;
        RECT 426.750 147.750 428.550 159.600 ;
        RECT 440.550 147.750 442.350 159.600 ;
        RECT 444.750 147.750 446.550 159.600 ;
        RECT 461.700 153.600 462.900 170.700 ;
        RECT 468.150 166.950 469.350 173.400 ;
        RECT 484.950 169.950 486.000 176.400 ;
        RECT 505.950 169.950 507.000 176.400 ;
        RECT 484.950 167.850 487.050 169.950 ;
        RECT 505.950 167.850 508.050 169.950 ;
        RECT 521.400 168.150 522.600 176.400 ;
        RECT 535.650 173.400 537.450 179.250 ;
        RECT 536.250 171.300 537.450 173.400 ;
        RECT 538.650 174.300 540.450 179.250 ;
        RECT 541.650 175.200 543.450 179.250 ;
        RECT 544.650 174.300 546.450 179.250 ;
        RECT 538.650 172.950 546.450 174.300 ;
        RECT 556.650 173.400 558.450 179.250 ;
        RECT 557.250 171.300 558.450 173.400 ;
        RECT 559.650 174.300 561.450 179.250 ;
        RECT 562.650 175.200 564.450 179.250 ;
        RECT 565.650 174.300 567.450 179.250 ;
        RECT 559.650 172.950 567.450 174.300 ;
        RECT 575.850 173.400 577.650 179.250 ;
        RECT 580.350 172.200 582.150 179.250 ;
        RECT 593.850 173.400 595.650 179.250 ;
        RECT 598.350 172.200 600.150 179.250 ;
        RECT 611.550 176.400 613.350 179.250 ;
        RECT 614.550 176.400 616.350 179.250 ;
        RECT 617.550 176.400 619.350 179.250 ;
        RECT 629.550 176.400 631.350 179.250 ;
        RECT 632.550 176.400 634.350 179.250 ;
        RECT 647.700 176.400 649.500 179.250 ;
        RECT 578.550 171.300 582.150 172.200 ;
        RECT 596.550 171.300 600.150 172.200 ;
        RECT 536.250 170.250 540.000 171.300 ;
        RECT 557.250 170.250 561.000 171.300 ;
        RECT 464.100 165.150 465.900 166.950 ;
        RECT 463.950 163.050 466.050 165.150 ;
        RECT 466.950 164.850 469.350 166.950 ;
        RECT 481.950 164.850 484.050 166.950 ;
        RECT 468.150 159.600 469.350 164.850 ;
        RECT 482.100 163.050 483.900 164.850 ;
        RECT 484.950 160.650 486.000 167.850 ;
        RECT 487.950 164.850 490.050 166.950 ;
        RECT 502.950 164.850 505.050 166.950 ;
        RECT 488.100 163.050 489.900 164.850 ;
        RECT 503.100 163.050 504.900 164.850 ;
        RECT 505.950 160.650 507.000 167.850 ;
        RECT 508.950 164.850 511.050 166.950 ;
        RECT 520.950 166.050 523.050 168.150 ;
        RECT 523.950 167.850 526.050 169.950 ;
        RECT 524.100 166.050 525.900 167.850 ;
        RECT 538.950 166.950 540.150 170.250 ;
        RECT 542.100 168.150 543.900 169.950 ;
        RECT 509.100 163.050 510.900 164.850 ;
        RECT 483.450 159.600 486.000 160.650 ;
        RECT 504.450 159.600 507.000 160.650 ;
        RECT 458.550 147.750 460.350 153.600 ;
        RECT 461.550 147.750 463.350 153.600 ;
        RECT 465.150 147.750 466.950 159.600 ;
        RECT 468.150 147.750 469.950 159.600 ;
        RECT 483.450 147.750 485.250 159.600 ;
        RECT 487.650 147.750 489.450 159.600 ;
        RECT 504.450 147.750 506.250 159.600 ;
        RECT 508.650 147.750 510.450 159.600 ;
        RECT 521.400 153.600 522.600 166.050 ;
        RECT 538.950 164.850 541.050 166.950 ;
        RECT 541.950 166.050 544.050 168.150 ;
        RECT 559.950 166.950 561.150 170.250 ;
        RECT 563.100 168.150 564.900 169.950 ;
        RECT 544.950 164.850 547.050 166.950 ;
        RECT 559.950 164.850 562.050 166.950 ;
        RECT 562.950 166.050 565.050 168.150 ;
        RECT 565.950 164.850 568.050 166.950 ;
        RECT 575.100 165.150 576.900 166.950 ;
        RECT 535.950 161.850 538.050 163.950 ;
        RECT 536.250 160.050 538.050 161.850 ;
        RECT 539.850 159.600 541.050 164.850 ;
        RECT 545.100 163.050 546.900 164.850 ;
        RECT 556.950 161.850 559.050 163.950 ;
        RECT 557.250 160.050 559.050 161.850 ;
        RECT 560.850 159.600 562.050 164.850 ;
        RECT 566.100 163.050 567.900 164.850 ;
        RECT 574.950 163.050 577.050 165.150 ;
        RECT 578.550 163.950 579.750 171.300 ;
        RECT 581.100 165.150 582.900 166.950 ;
        RECT 593.100 165.150 594.900 166.950 ;
        RECT 577.950 161.850 580.050 163.950 ;
        RECT 580.950 163.050 583.050 165.150 ;
        RECT 592.950 163.050 595.050 165.150 ;
        RECT 596.550 163.950 597.750 171.300 ;
        RECT 615.000 169.950 616.050 176.400 ;
        RECT 613.950 167.850 616.050 169.950 ;
        RECT 628.950 167.850 631.050 169.950 ;
        RECT 632.400 168.150 633.600 176.400 ;
        RECT 651.000 175.050 652.800 179.250 ;
        RECT 647.100 173.400 652.800 175.050 ;
        RECT 655.200 173.400 657.000 179.250 ;
        RECT 670.650 173.400 672.450 179.250 ;
        RECT 599.100 165.150 600.900 166.950 ;
        RECT 595.950 161.850 598.050 163.950 ;
        RECT 598.950 163.050 601.050 165.150 ;
        RECT 610.950 164.850 613.050 166.950 ;
        RECT 611.100 163.050 612.900 164.850 ;
        RECT 520.650 147.750 522.450 153.600 ;
        RECT 523.650 147.750 525.450 153.600 ;
        RECT 536.400 147.750 538.200 153.600 ;
        RECT 539.700 147.750 541.500 159.600 ;
        RECT 543.900 147.750 545.700 159.600 ;
        RECT 557.400 147.750 559.200 153.600 ;
        RECT 560.700 147.750 562.500 159.600 ;
        RECT 564.900 147.750 566.700 159.600 ;
        RECT 578.550 153.600 579.750 161.850 ;
        RECT 596.550 153.600 597.750 161.850 ;
        RECT 615.000 160.650 616.050 167.850 ;
        RECT 616.950 164.850 619.050 166.950 ;
        RECT 629.100 166.050 630.900 167.850 ;
        RECT 631.950 166.050 634.050 168.150 ;
        RECT 647.100 166.950 648.300 173.400 ;
        RECT 671.250 171.300 672.450 173.400 ;
        RECT 673.650 174.300 675.450 179.250 ;
        RECT 676.650 175.200 678.450 179.250 ;
        RECT 679.650 174.300 681.450 179.250 ;
        RECT 692.700 176.400 694.500 179.250 ;
        RECT 696.000 175.050 697.800 179.250 ;
        RECT 673.650 172.950 681.450 174.300 ;
        RECT 692.100 173.400 697.800 175.050 ;
        RECT 700.200 173.400 702.000 179.250 ;
        RECT 710.550 174.300 712.350 179.250 ;
        RECT 713.550 175.200 715.350 179.250 ;
        RECT 716.550 174.300 718.350 179.250 ;
        RECT 671.250 170.250 675.000 171.300 ;
        RECT 650.100 168.150 651.900 169.950 ;
        RECT 617.100 163.050 618.900 164.850 ;
        RECT 615.000 159.600 617.550 160.650 ;
        RECT 575.550 147.750 577.350 153.600 ;
        RECT 578.550 147.750 580.350 153.600 ;
        RECT 581.550 147.750 583.350 153.600 ;
        RECT 593.550 147.750 595.350 153.600 ;
        RECT 596.550 147.750 598.350 153.600 ;
        RECT 599.550 147.750 601.350 153.600 ;
        RECT 611.550 147.750 613.350 159.600 ;
        RECT 615.750 147.750 617.550 159.600 ;
        RECT 632.400 153.600 633.600 166.050 ;
        RECT 646.950 164.850 649.050 166.950 ;
        RECT 649.950 166.050 652.050 168.150 ;
        RECT 652.950 167.850 655.050 169.950 ;
        RECT 656.100 168.150 657.900 169.950 ;
        RECT 653.100 166.050 654.900 167.850 ;
        RECT 655.950 166.050 658.050 168.150 ;
        RECT 673.950 166.950 675.150 170.250 ;
        RECT 677.100 168.150 678.900 169.950 ;
        RECT 673.950 164.850 676.050 166.950 ;
        RECT 676.950 166.050 679.050 168.150 ;
        RECT 692.100 166.950 693.300 173.400 ;
        RECT 710.550 172.950 718.350 174.300 ;
        RECT 719.550 173.400 721.350 179.250 ;
        RECT 731.550 176.400 733.350 179.250 ;
        RECT 719.550 171.300 720.750 173.400 ;
        RECT 732.150 172.500 733.350 176.400 ;
        RECT 734.850 173.400 736.650 179.250 ;
        RECT 737.850 173.400 739.650 179.250 ;
        RECT 749.550 176.400 751.350 179.250 ;
        RECT 752.550 176.400 754.350 179.250 ;
        RECT 764.550 176.400 766.350 179.250 ;
        RECT 767.550 176.400 769.350 179.250 ;
        RECT 732.150 171.600 737.250 172.500 ;
        RECT 717.000 170.250 720.750 171.300 ;
        RECT 735.000 170.700 737.250 171.600 ;
        RECT 695.100 168.150 696.900 169.950 ;
        RECT 679.950 164.850 682.050 166.950 ;
        RECT 691.950 164.850 694.050 166.950 ;
        RECT 694.950 166.050 697.050 168.150 ;
        RECT 697.950 167.850 700.050 169.950 ;
        RECT 701.100 168.150 702.900 169.950 ;
        RECT 713.100 168.150 714.900 169.950 ;
        RECT 698.100 166.050 699.900 167.850 ;
        RECT 700.950 166.050 703.050 168.150 ;
        RECT 709.950 164.850 712.050 166.950 ;
        RECT 712.950 166.050 715.050 168.150 ;
        RECT 716.850 166.950 718.050 170.250 ;
        RECT 715.950 164.850 718.050 166.950 ;
        RECT 730.950 164.850 733.050 166.950 ;
        RECT 647.100 159.600 648.300 164.850 ;
        RECT 670.950 161.850 673.050 163.950 ;
        RECT 671.250 160.050 673.050 161.850 ;
        RECT 674.850 159.600 676.050 164.850 ;
        RECT 680.100 163.050 681.900 164.850 ;
        RECT 692.100 159.600 693.300 164.850 ;
        RECT 710.100 163.050 711.900 164.850 ;
        RECT 694.950 162.450 697.050 163.050 ;
        RECT 706.950 162.450 709.050 163.050 ;
        RECT 694.950 161.550 709.050 162.450 ;
        RECT 694.950 160.950 697.050 161.550 ;
        RECT 706.950 160.950 709.050 161.550 ;
        RECT 715.950 159.600 717.150 164.850 ;
        RECT 718.950 161.850 721.050 163.950 ;
        RECT 731.100 163.050 732.900 164.850 ;
        RECT 735.000 162.300 736.050 170.700 ;
        RECT 738.150 166.950 739.350 173.400 ;
        RECT 748.950 167.850 751.050 169.950 ;
        RECT 752.400 168.150 753.600 176.400 ;
        RECT 736.950 164.850 739.350 166.950 ;
        RECT 749.100 166.050 750.900 167.850 ;
        RECT 751.950 166.050 754.050 168.150 ;
        RECT 763.950 167.850 766.050 169.950 ;
        RECT 767.400 168.150 768.600 176.400 ;
        RECT 782.850 172.200 784.650 179.250 ;
        RECT 787.350 173.400 789.150 179.250 ;
        RECT 802.650 173.400 804.450 179.250 ;
        RECT 782.850 171.300 786.450 172.200 ;
        RECT 764.100 166.050 765.900 167.850 ;
        RECT 766.950 166.050 769.050 168.150 ;
        RECT 718.950 160.050 720.750 161.850 ;
        RECT 735.000 161.400 737.250 162.300 ;
        RECT 731.550 160.500 737.250 161.400 ;
        RECT 629.550 147.750 631.350 153.600 ;
        RECT 632.550 147.750 634.350 153.600 ;
        RECT 646.650 147.750 648.450 159.600 ;
        RECT 649.650 158.700 657.450 159.600 ;
        RECT 649.650 147.750 651.450 158.700 ;
        RECT 652.650 147.750 654.450 157.800 ;
        RECT 655.650 147.750 657.450 158.700 ;
        RECT 671.400 147.750 673.200 153.600 ;
        RECT 674.700 147.750 676.500 159.600 ;
        RECT 678.900 147.750 680.700 159.600 ;
        RECT 691.650 147.750 693.450 159.600 ;
        RECT 694.650 158.700 702.450 159.600 ;
        RECT 694.650 147.750 696.450 158.700 ;
        RECT 697.650 147.750 699.450 157.800 ;
        RECT 700.650 147.750 702.450 158.700 ;
        RECT 711.300 147.750 713.100 159.600 ;
        RECT 715.500 147.750 717.300 159.600 ;
        RECT 731.550 153.600 732.750 160.500 ;
        RECT 738.150 159.600 739.350 164.850 ;
        RECT 718.800 147.750 720.600 153.600 ;
        RECT 731.550 147.750 733.350 153.600 ;
        RECT 734.850 147.750 736.650 159.600 ;
        RECT 737.850 147.750 739.650 159.600 ;
        RECT 752.400 153.600 753.600 166.050 ;
        RECT 767.400 153.600 768.600 166.050 ;
        RECT 782.100 165.150 783.900 166.950 ;
        RECT 781.950 163.050 784.050 165.150 ;
        RECT 785.250 163.950 786.450 171.300 ;
        RECT 803.250 171.300 804.450 173.400 ;
        RECT 805.650 174.300 807.450 179.250 ;
        RECT 808.650 175.200 810.450 179.250 ;
        RECT 811.650 174.300 813.450 179.250 ;
        RECT 821.550 176.400 823.350 179.250 ;
        RECT 824.550 176.400 826.350 179.250 ;
        RECT 827.550 176.400 829.350 179.250 ;
        RECT 805.650 172.950 813.450 174.300 ;
        RECT 803.250 170.250 807.000 171.300 ;
        RECT 805.950 166.950 807.150 170.250 ;
        RECT 825.000 169.950 826.050 176.400 ;
        RECT 845.100 171.000 846.900 179.250 ;
        RECT 809.100 168.150 810.900 169.950 ;
        RECT 788.100 165.150 789.900 166.950 ;
        RECT 784.950 161.850 787.050 163.950 ;
        RECT 787.950 163.050 790.050 165.150 ;
        RECT 805.950 164.850 808.050 166.950 ;
        RECT 808.950 166.050 811.050 168.150 ;
        RECT 823.950 167.850 826.050 169.950 ;
        RECT 811.950 164.850 814.050 166.950 ;
        RECT 820.950 164.850 823.050 166.950 ;
        RECT 802.950 161.850 805.050 163.950 ;
        RECT 785.250 153.600 786.450 161.850 ;
        RECT 803.250 160.050 805.050 161.850 ;
        RECT 806.850 159.600 808.050 164.850 ;
        RECT 812.100 163.050 813.900 164.850 ;
        RECT 821.100 163.050 822.900 164.850 ;
        RECT 825.000 160.650 826.050 167.850 ;
        RECT 842.400 169.350 846.900 171.000 ;
        RECT 850.500 170.400 852.300 179.250 ;
        RECT 862.650 176.400 864.450 179.250 ;
        RECT 865.650 176.400 867.450 179.250 ;
        RECT 826.950 164.850 829.050 166.950 ;
        RECT 842.400 165.150 843.600 169.350 ;
        RECT 850.950 168.450 853.050 169.050 ;
        RECT 850.950 167.550 855.450 168.450 ;
        RECT 863.400 168.150 864.600 176.400 ;
        RECT 850.950 166.950 853.050 167.550 ;
        RECT 827.100 163.050 828.900 164.850 ;
        RECT 841.950 163.050 844.050 165.150 ;
        RECT 825.000 159.600 827.550 160.650 ;
        RECT 749.550 147.750 751.350 153.600 ;
        RECT 752.550 147.750 754.350 153.600 ;
        RECT 764.550 147.750 766.350 153.600 ;
        RECT 767.550 147.750 769.350 153.600 ;
        RECT 781.650 147.750 783.450 153.600 ;
        RECT 784.650 147.750 786.450 153.600 ;
        RECT 787.650 147.750 789.450 153.600 ;
        RECT 803.400 147.750 805.200 153.600 ;
        RECT 806.700 147.750 808.500 159.600 ;
        RECT 810.900 147.750 812.700 159.600 ;
        RECT 821.550 147.750 823.350 159.600 ;
        RECT 825.750 147.750 827.550 159.600 ;
        RECT 842.250 154.800 843.300 163.050 ;
        RECT 844.950 161.850 847.050 163.950 ;
        RECT 850.950 161.850 853.050 163.950 ;
        RECT 854.550 163.050 855.450 167.550 ;
        RECT 862.950 166.050 865.050 168.150 ;
        RECT 865.950 167.850 868.050 169.950 ;
        RECT 866.100 166.050 867.900 167.850 ;
        RECT 844.950 160.050 846.750 161.850 ;
        RECT 847.950 158.850 850.050 160.950 ;
        RECT 851.100 160.050 852.900 161.850 ;
        RECT 853.950 160.950 856.050 163.050 ;
        RECT 848.100 157.050 849.900 158.850 ;
        RECT 842.250 153.900 849.300 154.800 ;
        RECT 842.250 153.600 843.450 153.900 ;
        RECT 841.650 147.750 843.450 153.600 ;
        RECT 847.650 153.600 849.300 153.900 ;
        RECT 863.400 153.600 864.600 166.050 ;
        RECT 844.650 147.750 846.450 153.000 ;
        RECT 847.650 147.750 849.450 153.600 ;
        RECT 850.650 147.750 852.450 153.600 ;
        RECT 862.650 147.750 864.450 153.600 ;
        RECT 865.650 147.750 867.450 153.600 ;
        RECT 10.650 137.400 12.450 143.250 ;
        RECT 13.650 138.000 15.450 143.250 ;
        RECT 11.250 137.100 12.450 137.400 ;
        RECT 16.650 137.400 18.450 143.250 ;
        RECT 19.650 137.400 21.450 143.250 ;
        RECT 16.650 137.100 18.300 137.400 ;
        RECT 11.250 136.200 18.300 137.100 ;
        RECT 11.250 127.950 12.300 136.200 ;
        RECT 17.100 132.150 18.900 133.950 ;
        RECT 29.550 132.300 31.350 143.250 ;
        RECT 32.550 133.200 34.350 143.250 ;
        RECT 35.550 132.300 37.350 143.250 ;
        RECT 13.950 129.150 15.750 130.950 ;
        RECT 16.950 130.050 19.050 132.150 ;
        RECT 29.550 131.400 37.350 132.300 ;
        RECT 38.550 131.400 40.350 143.250 ;
        RECT 52.650 137.400 54.450 143.250 ;
        RECT 55.650 138.000 57.450 143.250 ;
        RECT 53.250 137.100 54.450 137.400 ;
        RECT 58.650 137.400 60.450 143.250 ;
        RECT 61.650 137.400 63.450 143.250 ;
        RECT 58.650 137.100 60.300 137.400 ;
        RECT 53.250 136.200 60.300 137.100 ;
        RECT 20.100 129.150 21.900 130.950 ;
        RECT 10.950 125.850 13.050 127.950 ;
        RECT 13.950 127.050 16.050 129.150 ;
        RECT 19.950 127.050 22.050 129.150 ;
        RECT 38.700 126.150 39.900 131.400 ;
        RECT 53.250 127.950 54.300 136.200 ;
        RECT 59.100 132.150 60.900 133.950 ;
        RECT 55.950 129.150 57.750 130.950 ;
        RECT 58.950 130.050 61.050 132.150 ;
        RECT 73.650 131.400 75.450 143.250 ;
        RECT 76.650 132.300 78.450 143.250 ;
        RECT 79.650 133.200 81.450 143.250 ;
        RECT 82.650 132.300 84.450 143.250 ;
        RECT 94.650 137.400 96.450 143.250 ;
        RECT 97.650 138.000 99.450 143.250 ;
        RECT 76.650 131.400 84.450 132.300 ;
        RECT 95.250 137.100 96.450 137.400 ;
        RECT 100.650 137.400 102.450 143.250 ;
        RECT 103.650 137.400 105.450 143.250 ;
        RECT 100.650 137.100 102.300 137.400 ;
        RECT 95.250 136.200 102.300 137.100 ;
        RECT 62.100 129.150 63.900 130.950 ;
        RECT 11.400 121.650 12.600 125.850 ;
        RECT 28.950 122.850 31.050 124.950 ;
        RECT 32.100 123.150 33.900 124.950 ;
        RECT 11.400 120.000 15.900 121.650 ;
        RECT 29.100 121.050 30.900 122.850 ;
        RECT 31.950 121.050 34.050 123.150 ;
        RECT 34.950 122.850 37.050 124.950 ;
        RECT 37.950 124.050 40.050 126.150 ;
        RECT 52.950 125.850 55.050 127.950 ;
        RECT 55.950 127.050 58.050 129.150 ;
        RECT 61.950 127.050 64.050 129.150 ;
        RECT 74.100 126.150 75.300 131.400 ;
        RECT 95.250 127.950 96.300 136.200 ;
        RECT 101.100 132.150 102.900 133.950 ;
        RECT 113.550 132.300 115.350 143.250 ;
        RECT 116.550 133.200 118.350 143.250 ;
        RECT 119.550 132.300 121.350 143.250 ;
        RECT 97.950 129.150 99.750 130.950 ;
        RECT 100.950 130.050 103.050 132.150 ;
        RECT 113.550 131.400 121.350 132.300 ;
        RECT 122.550 131.400 124.350 143.250 ;
        RECT 137.400 137.400 139.200 143.250 ;
        RECT 140.700 131.400 142.500 143.250 ;
        RECT 144.900 131.400 146.700 143.250 ;
        RECT 157.650 137.400 159.450 143.250 ;
        RECT 160.650 138.000 162.450 143.250 ;
        RECT 158.250 137.100 159.450 137.400 ;
        RECT 163.650 137.400 165.450 143.250 ;
        RECT 166.650 137.400 168.450 143.250 ;
        RECT 163.650 137.100 165.300 137.400 ;
        RECT 158.250 136.200 165.300 137.100 ;
        RECT 104.100 129.150 105.900 130.950 ;
        RECT 35.100 121.050 36.900 122.850 ;
        RECT 14.100 111.750 15.900 120.000 ;
        RECT 19.500 111.750 21.300 120.600 ;
        RECT 38.700 117.600 39.900 124.050 ;
        RECT 53.400 121.650 54.600 125.850 ;
        RECT 73.950 124.050 76.050 126.150 ;
        RECT 94.950 125.850 97.050 127.950 ;
        RECT 97.950 127.050 100.050 129.150 ;
        RECT 103.950 127.050 106.050 129.150 ;
        RECT 122.700 126.150 123.900 131.400 ;
        RECT 137.250 129.150 139.050 130.950 ;
        RECT 136.950 127.050 139.050 129.150 ;
        RECT 140.850 126.150 142.050 131.400 ;
        RECT 158.250 127.950 159.300 136.200 ;
        RECT 164.100 132.150 165.900 133.950 ;
        RECT 160.950 129.150 162.750 130.950 ;
        RECT 163.950 130.050 166.050 132.150 ;
        RECT 177.300 131.400 179.100 143.250 ;
        RECT 181.500 131.400 183.300 143.250 ;
        RECT 184.800 137.400 186.600 143.250 ;
        RECT 199.650 137.400 201.450 143.250 ;
        RECT 202.650 138.000 204.450 143.250 ;
        RECT 200.250 137.100 201.450 137.400 ;
        RECT 205.650 137.400 207.450 143.250 ;
        RECT 208.650 137.400 210.450 143.250 ;
        RECT 218.550 137.400 220.350 143.250 ;
        RECT 221.550 137.400 223.350 143.250 ;
        RECT 233.550 137.400 235.350 143.250 ;
        RECT 236.550 137.400 238.350 143.250 ;
        RECT 239.550 137.400 241.350 143.250 ;
        RECT 256.650 137.400 258.450 143.250 ;
        RECT 259.650 138.000 261.450 143.250 ;
        RECT 205.650 137.100 207.300 137.400 ;
        RECT 200.250 136.200 207.300 137.100 ;
        RECT 167.100 129.150 168.900 130.950 ;
        RECT 146.100 126.150 147.900 127.950 ;
        RECT 53.400 120.000 57.900 121.650 ;
        RECT 30.000 111.750 31.800 117.600 ;
        RECT 34.200 115.950 39.900 117.600 ;
        RECT 34.200 111.750 36.000 115.950 ;
        RECT 37.500 111.750 39.300 114.600 ;
        RECT 56.100 111.750 57.900 120.000 ;
        RECT 61.500 111.750 63.300 120.600 ;
        RECT 74.100 117.600 75.300 124.050 ;
        RECT 76.950 122.850 79.050 124.950 ;
        RECT 80.100 123.150 81.900 124.950 ;
        RECT 77.100 121.050 78.900 122.850 ;
        RECT 79.950 121.050 82.050 123.150 ;
        RECT 82.950 122.850 85.050 124.950 ;
        RECT 83.100 121.050 84.900 122.850 ;
        RECT 95.400 121.650 96.600 125.850 ;
        RECT 112.950 122.850 115.050 124.950 ;
        RECT 116.100 123.150 117.900 124.950 ;
        RECT 95.400 120.000 99.900 121.650 ;
        RECT 113.100 121.050 114.900 122.850 ;
        RECT 115.950 121.050 118.050 123.150 ;
        RECT 118.950 122.850 121.050 124.950 ;
        RECT 121.950 124.050 124.050 126.150 ;
        RECT 139.950 124.050 142.050 126.150 ;
        RECT 119.100 121.050 120.900 122.850 ;
        RECT 74.100 115.950 79.800 117.600 ;
        RECT 74.700 111.750 76.500 114.600 ;
        RECT 78.000 111.750 79.800 115.950 ;
        RECT 82.200 111.750 84.000 117.600 ;
        RECT 98.100 111.750 99.900 120.000 ;
        RECT 103.500 111.750 105.300 120.600 ;
        RECT 122.700 117.600 123.900 124.050 ;
        RECT 139.950 120.750 141.150 124.050 ;
        RECT 142.950 122.850 145.050 124.950 ;
        RECT 145.950 124.050 148.050 126.150 ;
        RECT 157.950 125.850 160.050 127.950 ;
        RECT 160.950 127.050 163.050 129.150 ;
        RECT 166.950 127.050 169.050 129.150 ;
        RECT 176.100 126.150 177.900 127.950 ;
        RECT 181.950 126.150 183.150 131.400 ;
        RECT 184.950 129.150 186.750 130.950 ;
        RECT 184.950 127.050 187.050 129.150 ;
        RECT 200.250 127.950 201.300 136.200 ;
        RECT 206.100 132.150 207.900 133.950 ;
        RECT 202.950 129.150 204.750 130.950 ;
        RECT 205.950 130.050 208.050 132.150 ;
        RECT 209.100 129.150 210.900 130.950 ;
        RECT 143.100 121.050 144.900 122.850 ;
        RECT 158.400 121.650 159.600 125.850 ;
        RECT 175.950 124.050 178.050 126.150 ;
        RECT 178.950 122.850 181.050 124.950 ;
        RECT 181.950 124.050 184.050 126.150 ;
        RECT 199.950 125.850 202.050 127.950 ;
        RECT 202.950 127.050 205.050 129.150 ;
        RECT 208.950 127.050 211.050 129.150 ;
        RECT 137.250 119.700 141.000 120.750 ;
        RECT 158.400 120.000 162.900 121.650 ;
        RECT 179.100 121.050 180.900 122.850 ;
        RECT 137.250 117.600 138.450 119.700 ;
        RECT 114.000 111.750 115.800 117.600 ;
        RECT 118.200 115.950 123.900 117.600 ;
        RECT 118.200 111.750 120.000 115.950 ;
        RECT 121.500 111.750 123.300 114.600 ;
        RECT 136.650 111.750 138.450 117.600 ;
        RECT 139.650 116.700 147.450 118.050 ;
        RECT 139.650 111.750 141.450 116.700 ;
        RECT 142.650 111.750 144.450 115.800 ;
        RECT 145.650 111.750 147.450 116.700 ;
        RECT 161.100 111.750 162.900 120.000 ;
        RECT 166.500 111.750 168.300 120.600 ;
        RECT 169.950 120.450 172.050 121.050 ;
        RECT 175.950 120.450 178.050 121.050 ;
        RECT 182.850 120.750 184.050 124.050 ;
        RECT 200.400 121.650 201.600 125.850 ;
        RECT 221.400 124.950 222.600 137.400 ;
        RECT 236.550 129.150 237.750 137.400 ;
        RECT 257.250 137.100 258.450 137.400 ;
        RECT 262.650 137.400 264.450 143.250 ;
        RECT 265.650 137.400 267.450 143.250 ;
        RECT 277.650 137.400 279.450 143.250 ;
        RECT 280.650 138.000 282.450 143.250 ;
        RECT 262.650 137.100 264.300 137.400 ;
        RECT 257.250 136.200 264.300 137.100 ;
        RECT 278.250 137.100 279.450 137.400 ;
        RECT 283.650 137.400 285.450 143.250 ;
        RECT 286.650 137.400 288.450 143.250 ;
        RECT 296.550 137.400 298.350 143.250 ;
        RECT 299.550 137.400 301.350 143.250 ;
        RECT 302.550 138.000 304.350 143.250 ;
        RECT 283.650 137.100 285.300 137.400 ;
        RECT 278.250 136.200 285.300 137.100 ;
        RECT 299.700 137.100 301.350 137.400 ;
        RECT 305.550 137.400 307.350 143.250 ;
        RECT 305.550 137.100 306.750 137.400 ;
        RECT 299.700 136.200 306.750 137.100 ;
        RECT 238.950 132.450 241.050 133.050 ;
        RECT 247.950 132.450 250.050 133.050 ;
        RECT 238.950 131.550 250.050 132.450 ;
        RECT 238.950 130.950 241.050 131.550 ;
        RECT 247.950 130.950 250.050 131.550 ;
        RECT 232.950 125.850 235.050 127.950 ;
        RECT 235.950 127.050 238.050 129.150 ;
        RECT 257.250 127.950 258.300 136.200 ;
        RECT 263.100 132.150 264.900 133.950 ;
        RECT 259.950 129.150 261.750 130.950 ;
        RECT 262.950 130.050 265.050 132.150 ;
        RECT 266.100 129.150 267.900 130.950 ;
        RECT 218.100 123.150 219.900 124.950 ;
        RECT 169.950 119.550 178.050 120.450 ;
        RECT 183.000 119.700 186.750 120.750 ;
        RECT 200.400 120.000 204.900 121.650 ;
        RECT 217.950 121.050 220.050 123.150 ;
        RECT 220.950 122.850 223.050 124.950 ;
        RECT 233.100 124.050 234.900 125.850 ;
        RECT 169.950 118.950 172.050 119.550 ;
        RECT 175.950 118.950 178.050 119.550 ;
        RECT 176.550 116.700 184.350 118.050 ;
        RECT 176.550 111.750 178.350 116.700 ;
        RECT 179.550 111.750 181.350 115.800 ;
        RECT 182.550 111.750 184.350 116.700 ;
        RECT 185.550 117.600 186.750 119.700 ;
        RECT 185.550 111.750 187.350 117.600 ;
        RECT 203.100 111.750 204.900 120.000 ;
        RECT 208.500 111.750 210.300 120.600 ;
        RECT 221.400 114.600 222.600 122.850 ;
        RECT 236.550 119.700 237.750 127.050 ;
        RECT 238.950 125.850 241.050 127.950 ;
        RECT 256.950 125.850 259.050 127.950 ;
        RECT 259.950 127.050 262.050 129.150 ;
        RECT 265.950 127.050 268.050 129.150 ;
        RECT 278.250 127.950 279.300 136.200 ;
        RECT 284.100 132.150 285.900 133.950 ;
        RECT 299.100 132.150 300.900 133.950 ;
        RECT 280.950 129.150 282.750 130.950 ;
        RECT 283.950 130.050 286.050 132.150 ;
        RECT 287.100 129.150 288.900 130.950 ;
        RECT 296.100 129.150 297.900 130.950 ;
        RECT 298.950 130.050 301.050 132.150 ;
        RECT 302.250 129.150 304.050 130.950 ;
        RECT 277.950 125.850 280.050 127.950 ;
        RECT 280.950 127.050 283.050 129.150 ;
        RECT 286.950 127.050 289.050 129.150 ;
        RECT 295.950 127.050 298.050 129.150 ;
        RECT 301.950 127.050 304.050 129.150 ;
        RECT 305.700 127.950 306.750 136.200 ;
        RECT 318.300 131.400 320.100 143.250 ;
        RECT 322.500 131.400 324.300 143.250 ;
        RECT 325.800 137.400 327.600 143.250 ;
        RECT 338.550 137.400 340.350 143.250 ;
        RECT 341.550 137.400 343.350 143.250 ;
        RECT 304.950 125.850 307.050 127.950 ;
        RECT 317.100 126.150 318.900 127.950 ;
        RECT 322.950 126.150 324.150 131.400 ;
        RECT 325.950 129.150 327.750 130.950 ;
        RECT 325.950 127.050 328.050 129.150 ;
        RECT 338.100 126.150 339.900 127.950 ;
        RECT 239.100 124.050 240.900 125.850 ;
        RECT 257.400 121.650 258.600 125.850 ;
        RECT 278.400 121.650 279.600 125.850 ;
        RECT 305.400 121.650 306.600 125.850 ;
        RECT 316.950 124.050 319.050 126.150 ;
        RECT 319.950 122.850 322.050 124.950 ;
        RECT 322.950 124.050 325.050 126.150 ;
        RECT 337.950 124.050 340.050 126.150 ;
        RECT 257.400 120.000 261.900 121.650 ;
        RECT 236.550 118.800 240.150 119.700 ;
        RECT 218.550 111.750 220.350 114.600 ;
        RECT 221.550 111.750 223.350 114.600 ;
        RECT 233.850 111.750 235.650 117.600 ;
        RECT 238.350 111.750 240.150 118.800 ;
        RECT 260.100 111.750 261.900 120.000 ;
        RECT 265.500 111.750 267.300 120.600 ;
        RECT 278.400 120.000 282.900 121.650 ;
        RECT 281.100 111.750 282.900 120.000 ;
        RECT 286.500 111.750 288.300 120.600 ;
        RECT 296.700 111.750 298.500 120.600 ;
        RECT 302.100 120.000 306.600 121.650 ;
        RECT 320.100 121.050 321.900 122.850 ;
        RECT 323.850 120.750 325.050 124.050 ;
        RECT 302.100 111.750 303.900 120.000 ;
        RECT 324.000 119.700 327.750 120.750 ;
        RECT 341.700 120.300 342.900 137.400 ;
        RECT 345.150 131.400 346.950 143.250 ;
        RECT 348.150 131.400 349.950 143.250 ;
        RECT 359.550 137.400 361.350 143.250 ;
        RECT 362.550 137.400 364.350 143.250 ;
        RECT 376.650 137.400 378.450 143.250 ;
        RECT 379.650 137.400 381.450 143.250 ;
        RECT 382.650 137.400 384.450 143.250 ;
        RECT 343.950 125.850 346.050 127.950 ;
        RECT 348.150 126.150 349.350 131.400 ;
        RECT 344.100 124.050 345.900 125.850 ;
        RECT 346.950 124.050 349.350 126.150 ;
        RECT 362.400 124.950 363.600 137.400 ;
        RECT 380.250 129.150 381.450 137.400 ;
        RECT 396.150 132.900 397.950 143.250 ;
        RECT 395.550 131.550 397.950 132.900 ;
        RECT 399.150 131.550 400.950 143.250 ;
        RECT 376.950 125.850 379.050 127.950 ;
        RECT 379.950 127.050 382.050 129.150 ;
        RECT 317.550 116.700 325.350 118.050 ;
        RECT 317.550 111.750 319.350 116.700 ;
        RECT 320.550 111.750 322.350 115.800 ;
        RECT 323.550 111.750 325.350 116.700 ;
        RECT 326.550 117.600 327.750 119.700 ;
        RECT 338.550 119.100 346.050 120.300 ;
        RECT 326.550 111.750 328.350 117.600 ;
        RECT 338.550 111.750 340.350 119.100 ;
        RECT 344.250 118.500 346.050 119.100 ;
        RECT 348.150 117.600 349.350 124.050 ;
        RECT 359.100 123.150 360.900 124.950 ;
        RECT 358.950 121.050 361.050 123.150 ;
        RECT 361.950 122.850 364.050 124.950 ;
        RECT 377.100 124.050 378.900 125.850 ;
        RECT 343.050 111.750 344.850 117.600 ;
        RECT 346.050 116.100 349.350 117.600 ;
        RECT 346.050 111.750 347.850 116.100 ;
        RECT 362.400 114.600 363.600 122.850 ;
        RECT 380.250 119.700 381.450 127.050 ;
        RECT 382.950 125.850 385.050 127.950 ;
        RECT 383.100 124.050 384.900 125.850 ;
        RECT 395.550 124.950 396.900 131.550 ;
        RECT 403.650 131.400 405.450 143.250 ;
        RECT 413.550 137.400 415.350 143.250 ;
        RECT 416.550 137.400 418.350 143.250 ;
        RECT 419.550 137.400 421.350 143.250 ;
        RECT 433.650 137.400 435.450 143.250 ;
        RECT 436.650 137.400 438.450 143.250 ;
        RECT 439.650 137.400 441.450 143.250 ;
        RECT 452.550 137.400 454.350 143.250 ;
        RECT 455.550 137.400 457.350 143.250 ;
        RECT 469.650 137.400 471.450 143.250 ;
        RECT 472.650 137.400 474.450 143.250 ;
        RECT 487.650 137.400 489.450 143.250 ;
        RECT 490.650 137.400 492.450 143.250 ;
        RECT 493.650 137.400 495.450 143.250 ;
        RECT 398.250 130.200 400.050 130.650 ;
        RECT 404.250 130.200 405.450 131.400 ;
        RECT 398.250 129.000 405.450 130.200 ;
        RECT 416.550 129.150 417.750 137.400 ;
        RECT 437.250 129.150 438.450 137.400 ;
        RECT 398.250 128.850 400.050 129.000 ;
        RECT 377.850 118.800 381.450 119.700 ;
        RECT 394.950 122.850 397.050 124.950 ;
        RECT 359.550 111.750 361.350 114.600 ;
        RECT 362.550 111.750 364.350 114.600 ;
        RECT 377.850 111.750 379.650 118.800 ;
        RECT 394.950 117.600 396.000 122.850 ;
        RECT 398.400 120.600 399.300 128.850 ;
        RECT 401.100 126.150 402.900 127.950 ;
        RECT 400.950 124.050 403.050 126.150 ;
        RECT 412.950 125.850 415.050 127.950 ;
        RECT 415.950 127.050 418.050 129.150 ;
        RECT 404.100 123.150 405.900 124.950 ;
        RECT 413.100 124.050 414.900 125.850 ;
        RECT 403.950 121.050 406.050 123.150 ;
        RECT 398.250 119.700 400.050 120.600 ;
        RECT 416.550 119.700 417.750 127.050 ;
        RECT 418.950 125.850 421.050 127.950 ;
        RECT 433.950 125.850 436.050 127.950 ;
        RECT 436.950 127.050 439.050 129.150 ;
        RECT 419.100 124.050 420.900 125.850 ;
        RECT 434.100 124.050 435.900 125.850 ;
        RECT 437.250 119.700 438.450 127.050 ;
        RECT 439.950 125.850 442.050 127.950 ;
        RECT 440.100 124.050 441.900 125.850 ;
        RECT 455.400 124.950 456.600 137.400 ;
        RECT 470.400 124.950 471.600 137.400 ;
        RECT 491.250 129.150 492.450 137.400 ;
        RECT 510.450 131.400 512.250 143.250 ;
        RECT 514.650 131.400 516.450 143.250 ;
        RECT 528.450 131.400 530.250 143.250 ;
        RECT 532.650 131.400 534.450 143.250 ;
        RECT 544.650 131.400 546.450 143.250 ;
        RECT 547.650 132.300 549.450 143.250 ;
        RECT 550.650 133.200 552.450 143.250 ;
        RECT 553.650 132.300 555.450 143.250 ;
        RECT 565.650 137.400 567.450 143.250 ;
        RECT 568.650 137.400 570.450 143.250 ;
        RECT 581.400 137.400 583.200 143.250 ;
        RECT 547.650 131.400 555.450 132.300 ;
        RECT 510.450 130.350 513.000 131.400 ;
        RECT 528.450 130.350 531.000 131.400 ;
        RECT 487.950 125.850 490.050 127.950 ;
        RECT 490.950 127.050 493.050 129.150 ;
        RECT 452.100 123.150 453.900 124.950 ;
        RECT 451.950 121.050 454.050 123.150 ;
        RECT 454.950 122.850 457.050 124.950 ;
        RECT 469.950 122.850 472.050 124.950 ;
        RECT 473.100 123.150 474.900 124.950 ;
        RECT 488.100 124.050 489.900 125.850 ;
        RECT 398.250 118.800 401.550 119.700 ;
        RECT 416.550 118.800 420.150 119.700 ;
        RECT 382.350 111.750 384.150 117.600 ;
        RECT 394.650 111.750 396.450 117.600 ;
        RECT 400.650 114.600 401.550 118.800 ;
        RECT 397.650 111.750 399.450 114.600 ;
        RECT 400.650 111.750 402.450 114.600 ;
        RECT 403.650 111.750 405.450 114.600 ;
        RECT 413.850 111.750 415.650 117.600 ;
        RECT 418.350 111.750 420.150 118.800 ;
        RECT 434.850 118.800 438.450 119.700 ;
        RECT 434.850 111.750 436.650 118.800 ;
        RECT 439.350 111.750 441.150 117.600 ;
        RECT 455.400 114.600 456.600 122.850 ;
        RECT 470.400 114.600 471.600 122.850 ;
        RECT 472.950 121.050 475.050 123.150 ;
        RECT 491.250 119.700 492.450 127.050 ;
        RECT 493.950 125.850 496.050 127.950 ;
        RECT 509.100 126.150 510.900 127.950 ;
        RECT 494.100 124.050 495.900 125.850 ;
        RECT 508.950 124.050 511.050 126.150 ;
        RECT 488.850 118.800 492.450 119.700 ;
        RECT 511.950 123.150 513.000 130.350 ;
        RECT 515.100 126.150 516.900 127.950 ;
        RECT 527.100 126.150 528.900 127.950 ;
        RECT 514.950 124.050 517.050 126.150 ;
        RECT 526.950 124.050 529.050 126.150 ;
        RECT 529.950 123.150 531.000 130.350 ;
        RECT 533.100 126.150 534.900 127.950 ;
        RECT 545.100 126.150 546.300 131.400 ;
        RECT 532.950 124.050 535.050 126.150 ;
        RECT 544.950 124.050 547.050 126.150 ;
        RECT 566.400 124.950 567.600 137.400 ;
        RECT 584.700 131.400 586.500 143.250 ;
        RECT 588.900 131.400 590.700 143.250 ;
        RECT 599.550 137.400 601.350 143.250 ;
        RECT 602.550 137.400 604.350 143.250 ;
        RECT 605.550 137.400 607.350 143.250 ;
        RECT 620.400 137.400 622.200 143.250 ;
        RECT 581.250 129.150 583.050 130.950 ;
        RECT 580.950 127.050 583.050 129.150 ;
        RECT 584.850 126.150 586.050 131.400 ;
        RECT 602.550 129.150 603.750 137.400 ;
        RECT 623.700 131.400 625.500 143.250 ;
        RECT 627.900 131.400 629.700 143.250 ;
        RECT 641.400 137.400 643.200 143.250 ;
        RECT 644.700 131.400 646.500 143.250 ;
        RECT 648.900 131.400 650.700 143.250 ;
        RECT 662.550 137.400 664.350 143.250 ;
        RECT 665.550 137.400 667.350 143.250 ;
        RECT 680.400 137.400 682.200 143.250 ;
        RECT 620.250 129.150 622.050 130.950 ;
        RECT 590.100 126.150 591.900 127.950 ;
        RECT 511.950 121.050 514.050 123.150 ;
        RECT 529.950 121.050 532.050 123.150 ;
        RECT 452.550 111.750 454.350 114.600 ;
        RECT 455.550 111.750 457.350 114.600 ;
        RECT 469.650 111.750 471.450 114.600 ;
        RECT 472.650 111.750 474.450 114.600 ;
        RECT 488.850 111.750 490.650 118.800 ;
        RECT 493.350 111.750 495.150 117.600 ;
        RECT 511.950 114.600 513.000 121.050 ;
        RECT 529.950 114.600 531.000 121.050 ;
        RECT 545.100 117.600 546.300 124.050 ;
        RECT 547.950 122.850 550.050 124.950 ;
        RECT 551.100 123.150 552.900 124.950 ;
        RECT 548.100 121.050 549.900 122.850 ;
        RECT 550.950 121.050 553.050 123.150 ;
        RECT 553.950 122.850 556.050 124.950 ;
        RECT 565.950 122.850 568.050 124.950 ;
        RECT 569.100 123.150 570.900 124.950 ;
        RECT 583.950 124.050 586.050 126.150 ;
        RECT 554.100 121.050 555.900 122.850 ;
        RECT 545.100 115.950 550.800 117.600 ;
        RECT 508.650 111.750 510.450 114.600 ;
        RECT 511.650 111.750 513.450 114.600 ;
        RECT 514.650 111.750 516.450 114.600 ;
        RECT 526.650 111.750 528.450 114.600 ;
        RECT 529.650 111.750 531.450 114.600 ;
        RECT 532.650 111.750 534.450 114.600 ;
        RECT 545.700 111.750 547.500 114.600 ;
        RECT 549.000 111.750 550.800 115.950 ;
        RECT 553.200 111.750 555.000 117.600 ;
        RECT 566.400 114.600 567.600 122.850 ;
        RECT 568.950 121.050 571.050 123.150 ;
        RECT 583.950 120.750 585.150 124.050 ;
        RECT 586.950 122.850 589.050 124.950 ;
        RECT 589.950 124.050 592.050 126.150 ;
        RECT 598.950 125.850 601.050 127.950 ;
        RECT 601.950 127.050 604.050 129.150 ;
        RECT 599.100 124.050 600.900 125.850 ;
        RECT 587.100 121.050 588.900 122.850 ;
        RECT 581.250 119.700 585.000 120.750 ;
        RECT 602.550 119.700 603.750 127.050 ;
        RECT 604.950 125.850 607.050 127.950 ;
        RECT 619.950 127.050 622.050 129.150 ;
        RECT 623.850 126.150 625.050 131.400 ;
        RECT 641.250 129.150 643.050 130.950 ;
        RECT 629.100 126.150 630.900 127.950 ;
        RECT 640.950 127.050 643.050 129.150 ;
        RECT 644.850 126.150 646.050 131.400 ;
        RECT 650.100 126.150 651.900 127.950 ;
        RECT 605.100 124.050 606.900 125.850 ;
        RECT 622.950 124.050 625.050 126.150 ;
        RECT 622.950 120.750 624.150 124.050 ;
        RECT 625.950 122.850 628.050 124.950 ;
        RECT 628.950 124.050 631.050 126.150 ;
        RECT 643.950 124.050 646.050 126.150 ;
        RECT 626.100 121.050 627.900 122.850 ;
        RECT 643.950 120.750 645.150 124.050 ;
        RECT 646.950 122.850 649.050 124.950 ;
        RECT 649.950 124.050 652.050 126.150 ;
        RECT 665.400 124.950 666.600 137.400 ;
        RECT 683.700 131.400 685.500 143.250 ;
        RECT 687.900 131.400 689.700 143.250 ;
        RECT 698.550 132.300 700.350 143.250 ;
        RECT 701.550 133.200 703.350 143.250 ;
        RECT 704.550 132.300 706.350 143.250 ;
        RECT 698.550 131.400 706.350 132.300 ;
        RECT 707.550 131.400 709.350 143.250 ;
        RECT 721.350 131.400 723.150 143.250 ;
        RECT 724.350 131.400 726.150 143.250 ;
        RECT 727.650 137.400 729.450 143.250 ;
        RECT 740.400 137.400 742.200 143.250 ;
        RECT 680.250 129.150 682.050 130.950 ;
        RECT 679.950 127.050 682.050 129.150 ;
        RECT 683.850 126.150 685.050 131.400 ;
        RECT 689.100 126.150 690.900 127.950 ;
        RECT 707.700 126.150 708.900 131.400 ;
        RECT 721.650 126.150 722.850 131.400 ;
        RECT 728.250 130.500 729.450 137.400 ;
        RECT 743.700 131.400 745.500 143.250 ;
        RECT 747.900 131.400 749.700 143.250 ;
        RECT 758.550 132.300 760.350 143.250 ;
        RECT 761.550 133.200 763.350 143.250 ;
        RECT 764.550 132.300 766.350 143.250 ;
        RECT 758.550 131.400 766.350 132.300 ;
        RECT 767.550 131.400 769.350 143.250 ;
        RECT 783.150 132.900 784.950 143.250 ;
        RECT 782.550 131.550 784.950 132.900 ;
        RECT 786.150 131.550 787.950 143.250 ;
        RECT 723.750 129.600 729.450 130.500 ;
        RECT 723.750 128.700 726.000 129.600 ;
        RECT 740.250 129.150 742.050 130.950 ;
        RECT 662.100 123.150 663.900 124.950 ;
        RECT 647.100 121.050 648.900 122.850 ;
        RECT 661.950 121.050 664.050 123.150 ;
        RECT 664.950 122.850 667.050 124.950 ;
        RECT 682.950 124.050 685.050 126.150 ;
        RECT 620.250 119.700 624.000 120.750 ;
        RECT 641.250 119.700 645.000 120.750 ;
        RECT 581.250 117.600 582.450 119.700 ;
        RECT 602.550 118.800 606.150 119.700 ;
        RECT 565.650 111.750 567.450 114.600 ;
        RECT 568.650 111.750 570.450 114.600 ;
        RECT 580.650 111.750 582.450 117.600 ;
        RECT 583.650 116.700 591.450 118.050 ;
        RECT 583.650 111.750 585.450 116.700 ;
        RECT 586.650 111.750 588.450 115.800 ;
        RECT 589.650 111.750 591.450 116.700 ;
        RECT 599.850 111.750 601.650 117.600 ;
        RECT 604.350 111.750 606.150 118.800 ;
        RECT 620.250 117.600 621.450 119.700 ;
        RECT 619.650 111.750 621.450 117.600 ;
        RECT 622.650 116.700 630.450 118.050 ;
        RECT 641.250 117.600 642.450 119.700 ;
        RECT 622.650 111.750 624.450 116.700 ;
        RECT 625.650 111.750 627.450 115.800 ;
        RECT 628.650 111.750 630.450 116.700 ;
        RECT 640.650 111.750 642.450 117.600 ;
        RECT 643.650 116.700 651.450 118.050 ;
        RECT 643.650 111.750 645.450 116.700 ;
        RECT 646.650 111.750 648.450 115.800 ;
        RECT 649.650 111.750 651.450 116.700 ;
        RECT 665.400 114.600 666.600 122.850 ;
        RECT 682.950 120.750 684.150 124.050 ;
        RECT 685.950 122.850 688.050 124.950 ;
        RECT 688.950 124.050 691.050 126.150 ;
        RECT 697.950 122.850 700.050 124.950 ;
        RECT 701.100 123.150 702.900 124.950 ;
        RECT 686.100 121.050 687.900 122.850 ;
        RECT 698.100 121.050 699.900 122.850 ;
        RECT 700.950 121.050 703.050 123.150 ;
        RECT 703.950 122.850 706.050 124.950 ;
        RECT 706.950 124.050 709.050 126.150 ;
        RECT 721.650 124.050 724.050 126.150 ;
        RECT 704.100 121.050 705.900 122.850 ;
        RECT 680.250 119.700 684.000 120.750 ;
        RECT 680.250 117.600 681.450 119.700 ;
        RECT 662.550 111.750 664.350 114.600 ;
        RECT 665.550 111.750 667.350 114.600 ;
        RECT 679.650 111.750 681.450 117.600 ;
        RECT 682.650 116.700 690.450 118.050 ;
        RECT 707.700 117.600 708.900 124.050 ;
        RECT 721.650 117.600 722.850 124.050 ;
        RECT 724.950 120.300 726.000 128.700 ;
        RECT 728.100 126.150 729.900 127.950 ;
        RECT 739.950 127.050 742.050 129.150 ;
        RECT 743.850 126.150 745.050 131.400 ;
        RECT 754.950 129.450 757.050 130.050 ;
        RECT 763.950 129.450 766.050 130.050 ;
        RECT 754.950 128.550 766.050 129.450 ;
        RECT 754.950 127.950 757.050 128.550 ;
        RECT 763.950 127.950 766.050 128.550 ;
        RECT 749.100 126.150 750.900 127.950 ;
        RECT 767.700 126.150 768.900 131.400 ;
        RECT 727.950 124.050 730.050 126.150 ;
        RECT 742.950 124.050 745.050 126.150 ;
        RECT 742.950 120.750 744.150 124.050 ;
        RECT 745.950 122.850 748.050 124.950 ;
        RECT 748.950 124.050 751.050 126.150 ;
        RECT 757.950 122.850 760.050 124.950 ;
        RECT 761.100 123.150 762.900 124.950 ;
        RECT 746.100 121.050 747.900 122.850 ;
        RECT 758.100 121.050 759.900 122.850 ;
        RECT 760.950 121.050 763.050 123.150 ;
        RECT 763.950 122.850 766.050 124.950 ;
        RECT 766.950 124.050 769.050 126.150 ;
        RECT 782.550 124.950 783.900 131.550 ;
        RECT 790.650 131.400 792.450 143.250 ;
        RECT 805.650 137.400 807.450 143.250 ;
        RECT 808.650 137.400 810.450 143.250 ;
        RECT 820.650 142.500 828.450 143.250 ;
        RECT 785.250 130.200 787.050 130.650 ;
        RECT 791.250 130.200 792.450 131.400 ;
        RECT 785.250 129.000 792.450 130.200 ;
        RECT 785.250 128.850 787.050 129.000 ;
        RECT 764.100 121.050 765.900 122.850 ;
        RECT 723.750 119.400 726.000 120.300 ;
        RECT 740.250 119.700 744.000 120.750 ;
        RECT 723.750 118.500 728.850 119.400 ;
        RECT 682.650 111.750 684.450 116.700 ;
        RECT 685.650 111.750 687.450 115.800 ;
        RECT 688.650 111.750 690.450 116.700 ;
        RECT 699.000 111.750 700.800 117.600 ;
        RECT 703.200 115.950 708.900 117.600 ;
        RECT 703.200 111.750 705.000 115.950 ;
        RECT 706.500 111.750 708.300 114.600 ;
        RECT 721.350 111.750 723.150 117.600 ;
        RECT 724.350 111.750 726.150 117.600 ;
        RECT 727.650 114.600 728.850 118.500 ;
        RECT 740.250 117.600 741.450 119.700 ;
        RECT 727.650 111.750 729.450 114.600 ;
        RECT 739.650 111.750 741.450 117.600 ;
        RECT 742.650 116.700 750.450 118.050 ;
        RECT 767.700 117.600 768.900 124.050 ;
        RECT 781.950 122.850 784.050 124.950 ;
        RECT 781.950 117.600 783.000 122.850 ;
        RECT 785.400 120.600 786.300 128.850 ;
        RECT 788.100 126.150 789.900 127.950 ;
        RECT 787.950 124.050 790.050 126.150 ;
        RECT 806.400 124.950 807.600 137.400 ;
        RECT 820.650 131.400 822.450 142.500 ;
        RECT 823.650 131.400 825.450 141.600 ;
        RECT 826.650 132.600 828.450 142.500 ;
        RECT 829.650 133.500 831.450 143.250 ;
        RECT 832.650 132.600 834.450 143.250 ;
        RECT 826.650 131.700 834.450 132.600 ;
        RECT 846.300 131.400 848.100 143.250 ;
        RECT 850.500 131.400 852.300 143.250 ;
        RECT 853.800 137.400 855.600 143.250 ;
        RECT 823.800 130.500 825.600 131.400 ;
        RECT 823.800 129.600 827.850 130.500 ;
        RECT 821.100 126.150 822.900 127.950 ;
        RECT 826.950 126.150 827.850 129.600 ;
        RECT 832.950 126.150 834.750 127.950 ;
        RECT 845.100 126.150 846.900 127.950 ;
        RECT 850.950 126.150 852.150 131.400 ;
        RECT 853.950 129.150 855.750 130.950 ;
        RECT 853.950 127.050 856.050 129.150 ;
        RECT 791.100 123.150 792.900 124.950 ;
        RECT 790.950 121.050 793.050 123.150 ;
        RECT 805.950 122.850 808.050 124.950 ;
        RECT 809.100 123.150 810.900 124.950 ;
        RECT 820.950 124.050 823.050 126.150 ;
        RECT 785.250 119.700 787.050 120.600 ;
        RECT 785.250 118.800 788.550 119.700 ;
        RECT 742.650 111.750 744.450 116.700 ;
        RECT 745.650 111.750 747.450 115.800 ;
        RECT 748.650 111.750 750.450 116.700 ;
        RECT 759.000 111.750 760.800 117.600 ;
        RECT 763.200 115.950 768.900 117.600 ;
        RECT 763.200 111.750 765.000 115.950 ;
        RECT 766.500 111.750 768.300 114.600 ;
        RECT 781.650 111.750 783.450 117.600 ;
        RECT 787.650 114.600 788.550 118.800 ;
        RECT 806.400 114.600 807.600 122.850 ;
        RECT 808.950 121.050 811.050 123.150 ;
        RECT 823.950 122.850 826.050 124.950 ;
        RECT 826.950 124.050 829.050 126.150 ;
        RECT 824.250 121.050 826.050 122.850 ;
        RECT 828.000 117.600 829.050 124.050 ;
        RECT 829.950 122.850 832.050 124.950 ;
        RECT 832.950 124.050 835.050 126.150 ;
        RECT 844.950 124.050 847.050 126.150 ;
        RECT 847.950 122.850 850.050 124.950 ;
        RECT 850.950 124.050 853.050 126.150 ;
        RECT 829.950 121.050 831.750 122.850 ;
        RECT 848.100 121.050 849.900 122.850 ;
        RECT 851.850 120.750 853.050 124.050 ;
        RECT 852.000 119.700 855.750 120.750 ;
        RECT 784.650 111.750 786.450 114.600 ;
        RECT 787.650 111.750 789.450 114.600 ;
        RECT 790.650 111.750 792.450 114.600 ;
        RECT 805.650 111.750 807.450 114.600 ;
        RECT 808.650 111.750 810.450 114.600 ;
        RECT 823.800 111.750 825.600 117.600 ;
        RECT 828.000 111.750 829.800 117.600 ;
        RECT 832.200 111.750 834.000 117.600 ;
        RECT 845.550 116.700 853.350 118.050 ;
        RECT 845.550 111.750 847.350 116.700 ;
        RECT 848.550 111.750 850.350 115.800 ;
        RECT 851.550 111.750 853.350 116.700 ;
        RECT 854.550 117.600 855.750 119.700 ;
        RECT 854.550 111.750 856.350 117.600 ;
        RECT 14.100 99.000 15.900 107.250 ;
        RECT 11.400 97.350 15.900 99.000 ;
        RECT 19.500 98.400 21.300 107.250 ;
        RECT 35.700 104.400 37.500 107.250 ;
        RECT 39.000 103.050 40.800 107.250 ;
        RECT 35.100 101.400 40.800 103.050 ;
        RECT 43.200 101.400 45.000 107.250 ;
        RECT 11.400 93.150 12.600 97.350 ;
        RECT 35.100 94.950 36.300 101.400 ;
        RECT 59.100 99.000 60.900 107.250 ;
        RECT 38.100 96.150 39.900 97.950 ;
        RECT 10.950 91.050 13.050 93.150 ;
        RECT 34.950 92.850 37.050 94.950 ;
        RECT 37.950 94.050 40.050 96.150 ;
        RECT 40.950 95.850 43.050 97.950 ;
        RECT 44.100 96.150 45.900 97.950 ;
        RECT 56.400 97.350 60.900 99.000 ;
        RECT 64.500 98.400 66.300 107.250 ;
        RECT 76.650 101.400 78.450 107.250 ;
        RECT 77.250 99.300 78.450 101.400 ;
        RECT 79.650 102.300 81.450 107.250 ;
        RECT 82.650 103.200 84.450 107.250 ;
        RECT 85.650 102.300 87.450 107.250 ;
        RECT 79.650 100.950 87.450 102.300 ;
        RECT 96.000 101.400 97.800 107.250 ;
        RECT 100.200 103.050 102.000 107.250 ;
        RECT 103.500 104.400 105.300 107.250 ;
        RECT 100.200 101.400 105.900 103.050 ;
        RECT 116.850 101.400 118.650 107.250 ;
        RECT 77.250 98.250 81.000 99.300 ;
        RECT 41.100 94.050 42.900 95.850 ;
        RECT 43.950 94.050 46.050 96.150 ;
        RECT 56.400 93.150 57.600 97.350 ;
        RECT 79.950 94.950 81.150 98.250 ;
        RECT 83.100 96.150 84.900 97.950 ;
        RECT 95.100 96.150 96.900 97.950 ;
        RECT 11.250 82.800 12.300 91.050 ;
        RECT 13.950 89.850 16.050 91.950 ;
        RECT 19.950 89.850 22.050 91.950 ;
        RECT 13.950 88.050 15.750 89.850 ;
        RECT 16.950 86.850 19.050 88.950 ;
        RECT 20.100 88.050 21.900 89.850 ;
        RECT 35.100 87.600 36.300 92.850 ;
        RECT 55.950 91.050 58.050 93.150 ;
        RECT 79.950 92.850 82.050 94.950 ;
        RECT 82.950 94.050 85.050 96.150 ;
        RECT 85.950 92.850 88.050 94.950 ;
        RECT 94.950 94.050 97.050 96.150 ;
        RECT 97.950 95.850 100.050 97.950 ;
        RECT 101.100 96.150 102.900 97.950 ;
        RECT 98.100 94.050 99.900 95.850 ;
        RECT 100.950 94.050 103.050 96.150 ;
        RECT 104.700 94.950 105.900 101.400 ;
        RECT 121.350 100.200 123.150 107.250 ;
        RECT 139.650 101.400 141.450 107.250 ;
        RECT 119.550 99.300 123.150 100.200 ;
        RECT 140.250 99.300 141.450 101.400 ;
        RECT 142.650 102.300 144.450 107.250 ;
        RECT 145.650 103.200 147.450 107.250 ;
        RECT 148.650 102.300 150.450 107.250 ;
        RECT 142.650 100.950 150.450 102.300 ;
        RECT 103.950 92.850 106.050 94.950 ;
        RECT 116.100 93.150 117.900 94.950 ;
        RECT 17.100 85.050 18.900 86.850 ;
        RECT 11.250 81.900 18.300 82.800 ;
        RECT 11.250 81.600 12.450 81.900 ;
        RECT 10.650 75.750 12.450 81.600 ;
        RECT 16.650 81.600 18.300 81.900 ;
        RECT 13.650 75.750 15.450 81.000 ;
        RECT 16.650 75.750 18.450 81.600 ;
        RECT 19.650 75.750 21.450 81.600 ;
        RECT 34.650 75.750 36.450 87.600 ;
        RECT 37.650 86.700 45.450 87.600 ;
        RECT 37.650 75.750 39.450 86.700 ;
        RECT 40.650 75.750 42.450 85.800 ;
        RECT 43.650 75.750 45.450 86.700 ;
        RECT 56.250 82.800 57.300 91.050 ;
        RECT 58.950 89.850 61.050 91.950 ;
        RECT 64.950 89.850 67.050 91.950 ;
        RECT 76.950 89.850 79.050 91.950 ;
        RECT 58.950 88.050 60.750 89.850 ;
        RECT 61.950 86.850 64.050 88.950 ;
        RECT 65.100 88.050 66.900 89.850 ;
        RECT 77.250 88.050 79.050 89.850 ;
        RECT 80.850 87.600 82.050 92.850 ;
        RECT 86.100 91.050 87.900 92.850 ;
        RECT 104.700 87.600 105.900 92.850 ;
        RECT 115.950 91.050 118.050 93.150 ;
        RECT 119.550 91.950 120.750 99.300 ;
        RECT 140.250 98.250 144.000 99.300 ;
        RECT 164.100 99.000 165.900 107.250 ;
        RECT 142.950 94.950 144.150 98.250 ;
        RECT 146.100 96.150 147.900 97.950 ;
        RECT 161.400 97.350 165.900 99.000 ;
        RECT 169.500 98.400 171.300 107.250 ;
        RECT 180.000 101.400 181.800 107.250 ;
        RECT 184.200 103.050 186.000 107.250 ;
        RECT 187.500 104.400 189.300 107.250 ;
        RECT 203.700 104.400 205.500 107.250 ;
        RECT 207.000 103.050 208.800 107.250 ;
        RECT 184.200 101.400 189.900 103.050 ;
        RECT 122.100 93.150 123.900 94.950 ;
        RECT 118.950 89.850 121.050 91.950 ;
        RECT 121.950 91.050 124.050 93.150 ;
        RECT 142.950 92.850 145.050 94.950 ;
        RECT 145.950 94.050 148.050 96.150 ;
        RECT 148.950 92.850 151.050 94.950 ;
        RECT 161.400 93.150 162.600 97.350 ;
        RECT 179.100 96.150 180.900 97.950 ;
        RECT 178.950 94.050 181.050 96.150 ;
        RECT 181.950 95.850 184.050 97.950 ;
        RECT 185.100 96.150 186.900 97.950 ;
        RECT 182.100 94.050 183.900 95.850 ;
        RECT 184.950 94.050 187.050 96.150 ;
        RECT 188.700 94.950 189.900 101.400 ;
        RECT 203.100 101.400 208.800 103.050 ;
        RECT 211.200 101.400 213.000 107.250 ;
        RECT 203.100 94.950 204.300 101.400 ;
        RECT 224.700 98.400 226.500 107.250 ;
        RECT 230.100 99.000 231.900 107.250 ;
        RECT 247.650 101.400 249.450 107.250 ;
        RECT 248.250 99.300 249.450 101.400 ;
        RECT 250.650 102.300 252.450 107.250 ;
        RECT 253.650 103.200 255.450 107.250 ;
        RECT 256.650 102.300 258.450 107.250 ;
        RECT 250.650 100.950 258.450 102.300 ;
        RECT 206.100 96.150 207.900 97.950 ;
        RECT 139.950 89.850 142.050 91.950 ;
        RECT 62.100 85.050 63.900 86.850 ;
        RECT 56.250 81.900 63.300 82.800 ;
        RECT 56.250 81.600 57.450 81.900 ;
        RECT 55.650 75.750 57.450 81.600 ;
        RECT 61.650 81.600 63.300 81.900 ;
        RECT 58.650 75.750 60.450 81.000 ;
        RECT 61.650 75.750 63.450 81.600 ;
        RECT 64.650 75.750 66.450 81.600 ;
        RECT 77.400 75.750 79.200 81.600 ;
        RECT 80.700 75.750 82.500 87.600 ;
        RECT 84.900 75.750 86.700 87.600 ;
        RECT 95.550 86.700 103.350 87.600 ;
        RECT 95.550 75.750 97.350 86.700 ;
        RECT 98.550 75.750 100.350 85.800 ;
        RECT 101.550 75.750 103.350 86.700 ;
        RECT 104.550 75.750 106.350 87.600 ;
        RECT 119.550 81.600 120.750 89.850 ;
        RECT 140.250 88.050 142.050 89.850 ;
        RECT 143.850 87.600 145.050 92.850 ;
        RECT 149.100 91.050 150.900 92.850 ;
        RECT 160.950 91.050 163.050 93.150 ;
        RECT 187.950 92.850 190.050 94.950 ;
        RECT 202.950 92.850 205.050 94.950 ;
        RECT 205.950 94.050 208.050 96.150 ;
        RECT 208.950 95.850 211.050 97.950 ;
        RECT 212.100 96.150 213.900 97.950 ;
        RECT 230.100 97.350 234.600 99.000 ;
        RECT 248.250 98.250 252.000 99.300 ;
        RECT 272.100 99.000 273.900 107.250 ;
        RECT 209.100 94.050 210.900 95.850 ;
        RECT 211.950 94.050 214.050 96.150 ;
        RECT 233.400 93.150 234.600 97.350 ;
        RECT 250.950 94.950 252.150 98.250 ;
        RECT 254.100 96.150 255.900 97.950 ;
        RECT 269.400 97.350 273.900 99.000 ;
        RECT 277.500 98.400 279.300 107.250 ;
        RECT 288.000 101.400 289.800 107.250 ;
        RECT 292.200 103.050 294.000 107.250 ;
        RECT 295.500 104.400 297.300 107.250 ;
        RECT 310.650 104.400 312.450 107.250 ;
        RECT 313.650 104.400 315.450 107.250 ;
        RECT 316.650 104.400 318.450 107.250 ;
        RECT 292.200 101.400 297.900 103.050 ;
        RECT 116.550 75.750 118.350 81.600 ;
        RECT 119.550 75.750 121.350 81.600 ;
        RECT 122.550 75.750 124.350 81.600 ;
        RECT 140.400 75.750 142.200 81.600 ;
        RECT 143.700 75.750 145.500 87.600 ;
        RECT 147.900 75.750 149.700 87.600 ;
        RECT 161.250 82.800 162.300 91.050 ;
        RECT 163.950 89.850 166.050 91.950 ;
        RECT 169.950 89.850 172.050 91.950 ;
        RECT 163.950 88.050 165.750 89.850 ;
        RECT 166.950 86.850 169.050 88.950 ;
        RECT 170.100 88.050 171.900 89.850 ;
        RECT 188.700 87.600 189.900 92.850 ;
        RECT 203.100 87.600 204.300 92.850 ;
        RECT 223.950 89.850 226.050 91.950 ;
        RECT 229.950 89.850 232.050 91.950 ;
        RECT 232.950 91.050 235.050 93.150 ;
        RECT 250.950 92.850 253.050 94.950 ;
        RECT 253.950 94.050 256.050 96.150 ;
        RECT 256.950 92.850 259.050 94.950 ;
        RECT 269.400 93.150 270.600 97.350 ;
        RECT 287.100 96.150 288.900 97.950 ;
        RECT 286.950 94.050 289.050 96.150 ;
        RECT 289.950 95.850 292.050 97.950 ;
        RECT 293.100 96.150 294.900 97.950 ;
        RECT 290.100 94.050 291.900 95.850 ;
        RECT 292.950 94.050 295.050 96.150 ;
        RECT 296.700 94.950 297.900 101.400 ;
        RECT 313.950 97.950 315.000 104.400 ;
        RECT 328.650 101.400 330.450 107.250 ;
        RECT 331.650 104.400 333.450 107.250 ;
        RECT 334.650 104.400 336.450 107.250 ;
        RECT 337.650 104.400 339.450 107.250 ;
        RECT 313.950 95.850 316.050 97.950 ;
        RECT 328.950 96.150 330.000 101.400 ;
        RECT 334.650 100.200 335.550 104.400 ;
        RECT 332.250 99.300 335.550 100.200 ;
        RECT 347.550 99.900 349.350 107.250 ;
        RECT 352.050 101.400 353.850 107.250 ;
        RECT 355.050 102.900 356.850 107.250 ;
        RECT 355.050 101.400 358.350 102.900 ;
        RECT 368.850 101.400 370.650 107.250 ;
        RECT 353.250 99.900 355.050 100.500 ;
        RECT 332.250 98.400 334.050 99.300 ;
        RECT 347.550 98.700 355.050 99.900 ;
        RECT 224.100 88.050 225.900 89.850 ;
        RECT 167.100 85.050 168.900 86.850 ;
        RECT 179.550 86.700 187.350 87.600 ;
        RECT 161.250 81.900 168.300 82.800 ;
        RECT 161.250 81.600 162.450 81.900 ;
        RECT 160.650 75.750 162.450 81.600 ;
        RECT 166.650 81.600 168.300 81.900 ;
        RECT 163.650 75.750 165.450 81.000 ;
        RECT 166.650 75.750 168.450 81.600 ;
        RECT 169.650 75.750 171.450 81.600 ;
        RECT 179.550 75.750 181.350 86.700 ;
        RECT 182.550 75.750 184.350 85.800 ;
        RECT 185.550 75.750 187.350 86.700 ;
        RECT 188.550 75.750 190.350 87.600 ;
        RECT 202.650 75.750 204.450 87.600 ;
        RECT 205.650 86.700 213.450 87.600 ;
        RECT 226.950 86.850 229.050 88.950 ;
        RECT 230.250 88.050 232.050 89.850 ;
        RECT 205.650 75.750 207.450 86.700 ;
        RECT 208.650 75.750 210.450 85.800 ;
        RECT 211.650 75.750 213.450 86.700 ;
        RECT 227.100 85.050 228.900 86.850 ;
        RECT 233.700 82.800 234.750 91.050 ;
        RECT 247.950 89.850 250.050 91.950 ;
        RECT 248.250 88.050 250.050 89.850 ;
        RECT 251.850 87.600 253.050 92.850 ;
        RECT 257.100 91.050 258.900 92.850 ;
        RECT 268.950 91.050 271.050 93.150 ;
        RECT 295.950 92.850 298.050 94.950 ;
        RECT 310.950 92.850 313.050 94.950 ;
        RECT 227.700 81.900 234.750 82.800 ;
        RECT 227.700 81.600 229.350 81.900 ;
        RECT 224.550 75.750 226.350 81.600 ;
        RECT 227.550 75.750 229.350 81.600 ;
        RECT 233.550 81.600 234.750 81.900 ;
        RECT 230.550 75.750 232.350 81.000 ;
        RECT 233.550 75.750 235.350 81.600 ;
        RECT 248.400 75.750 250.200 81.600 ;
        RECT 251.700 75.750 253.500 87.600 ;
        RECT 255.900 75.750 257.700 87.600 ;
        RECT 269.250 82.800 270.300 91.050 ;
        RECT 271.950 89.850 274.050 91.950 ;
        RECT 277.950 89.850 280.050 91.950 ;
        RECT 271.950 88.050 273.750 89.850 ;
        RECT 274.950 86.850 277.050 88.950 ;
        RECT 278.100 88.050 279.900 89.850 ;
        RECT 296.700 87.600 297.900 92.850 ;
        RECT 311.100 91.050 312.900 92.850 ;
        RECT 313.950 88.650 315.000 95.850 ;
        RECT 316.950 92.850 319.050 94.950 ;
        RECT 328.950 94.050 331.050 96.150 ;
        RECT 317.100 91.050 318.900 92.850 ;
        RECT 312.450 87.600 315.000 88.650 ;
        RECT 275.100 85.050 276.900 86.850 ;
        RECT 287.550 86.700 295.350 87.600 ;
        RECT 269.250 81.900 276.300 82.800 ;
        RECT 269.250 81.600 270.450 81.900 ;
        RECT 268.650 75.750 270.450 81.600 ;
        RECT 274.650 81.600 276.300 81.900 ;
        RECT 271.650 75.750 273.450 81.000 ;
        RECT 274.650 75.750 276.450 81.600 ;
        RECT 277.650 75.750 279.450 81.600 ;
        RECT 287.550 75.750 289.350 86.700 ;
        RECT 290.550 75.750 292.350 85.800 ;
        RECT 293.550 75.750 295.350 86.700 ;
        RECT 296.550 75.750 298.350 87.600 ;
        RECT 312.450 75.750 314.250 87.600 ;
        RECT 316.650 75.750 318.450 87.600 ;
        RECT 329.550 87.450 330.900 94.050 ;
        RECT 332.400 90.150 333.300 98.400 ;
        RECT 337.950 95.850 340.050 97.950 ;
        RECT 334.950 92.850 337.050 94.950 ;
        RECT 338.100 94.050 339.900 95.850 ;
        RECT 346.950 92.850 349.050 94.950 ;
        RECT 335.100 91.050 336.900 92.850 ;
        RECT 347.100 91.050 348.900 92.850 ;
        RECT 332.250 90.000 334.050 90.150 ;
        RECT 332.250 88.800 339.450 90.000 ;
        RECT 332.250 88.350 334.050 88.800 ;
        RECT 338.250 87.600 339.450 88.800 ;
        RECT 329.550 86.100 331.950 87.450 ;
        RECT 330.150 75.750 331.950 86.100 ;
        RECT 333.150 75.750 334.950 87.450 ;
        RECT 337.650 75.750 339.450 87.600 ;
        RECT 350.700 81.600 351.900 98.700 ;
        RECT 357.150 94.950 358.350 101.400 ;
        RECT 373.350 100.200 375.150 107.250 ;
        RECT 371.550 99.300 375.150 100.200 ;
        RECT 389.850 100.200 391.650 107.250 ;
        RECT 394.350 101.400 396.150 107.250 ;
        RECT 406.650 104.400 408.450 107.250 ;
        RECT 409.650 104.400 411.450 107.250 ;
        RECT 412.650 104.400 414.450 107.250 ;
        RECT 389.850 99.300 393.450 100.200 ;
        RECT 353.100 93.150 354.900 94.950 ;
        RECT 352.950 91.050 355.050 93.150 ;
        RECT 355.950 92.850 358.350 94.950 ;
        RECT 368.100 93.150 369.900 94.950 ;
        RECT 357.150 87.600 358.350 92.850 ;
        RECT 367.950 91.050 370.050 93.150 ;
        RECT 371.550 91.950 372.750 99.300 ;
        RECT 374.100 93.150 375.900 94.950 ;
        RECT 389.100 93.150 390.900 94.950 ;
        RECT 370.950 89.850 373.050 91.950 ;
        RECT 373.950 91.050 376.050 93.150 ;
        RECT 388.950 91.050 391.050 93.150 ;
        RECT 392.250 91.950 393.450 99.300 ;
        RECT 409.950 97.950 411.000 104.400 ;
        RECT 422.550 102.300 424.350 107.250 ;
        RECT 425.550 103.200 427.350 107.250 ;
        RECT 428.550 102.300 430.350 107.250 ;
        RECT 422.550 100.950 430.350 102.300 ;
        RECT 431.550 101.400 433.350 107.250 ;
        RECT 431.550 99.300 432.750 101.400 ;
        RECT 446.850 100.200 448.650 107.250 ;
        RECT 451.350 101.400 453.150 107.250 ;
        RECT 462.000 101.400 463.800 107.250 ;
        RECT 466.200 103.050 468.000 107.250 ;
        RECT 469.500 104.400 471.300 107.250 ;
        RECT 466.200 101.400 471.900 103.050 ;
        RECT 446.850 99.300 450.450 100.200 ;
        RECT 429.000 98.250 432.750 99.300 ;
        RECT 409.950 95.850 412.050 97.950 ;
        RECT 425.100 96.150 426.900 97.950 ;
        RECT 395.100 93.150 396.900 94.950 ;
        RECT 391.950 89.850 394.050 91.950 ;
        RECT 394.950 91.050 397.050 93.150 ;
        RECT 406.950 92.850 409.050 94.950 ;
        RECT 407.100 91.050 408.900 92.850 ;
        RECT 347.550 75.750 349.350 81.600 ;
        RECT 350.550 75.750 352.350 81.600 ;
        RECT 354.150 75.750 355.950 87.600 ;
        RECT 357.150 75.750 358.950 87.600 ;
        RECT 371.550 81.600 372.750 89.850 ;
        RECT 392.250 81.600 393.450 89.850 ;
        RECT 409.950 88.650 411.000 95.850 ;
        RECT 412.950 92.850 415.050 94.950 ;
        RECT 421.950 92.850 424.050 94.950 ;
        RECT 424.950 94.050 427.050 96.150 ;
        RECT 428.850 94.950 430.050 98.250 ;
        RECT 427.950 92.850 430.050 94.950 ;
        RECT 446.100 93.150 447.900 94.950 ;
        RECT 413.100 91.050 414.900 92.850 ;
        RECT 422.100 91.050 423.900 92.850 ;
        RECT 408.450 87.600 411.000 88.650 ;
        RECT 427.950 87.600 429.150 92.850 ;
        RECT 430.950 89.850 433.050 91.950 ;
        RECT 445.950 91.050 448.050 93.150 ;
        RECT 449.250 91.950 450.450 99.300 ;
        RECT 461.100 96.150 462.900 97.950 ;
        RECT 452.100 93.150 453.900 94.950 ;
        RECT 460.950 94.050 463.050 96.150 ;
        RECT 463.950 95.850 466.050 97.950 ;
        RECT 467.100 96.150 468.900 97.950 ;
        RECT 464.100 94.050 465.900 95.850 ;
        RECT 466.950 94.050 469.050 96.150 ;
        RECT 470.700 94.950 471.900 101.400 ;
        RECT 488.100 99.000 489.900 107.250 ;
        RECT 485.400 97.350 489.900 99.000 ;
        RECT 493.500 98.400 495.300 107.250 ;
        RECT 503.850 101.400 505.650 107.250 ;
        RECT 508.350 100.200 510.150 107.250 ;
        RECT 523.650 101.400 525.450 107.250 ;
        RECT 506.550 99.300 510.150 100.200 ;
        RECT 524.250 99.300 525.450 101.400 ;
        RECT 526.650 102.300 528.450 107.250 ;
        RECT 529.650 103.200 531.450 107.250 ;
        RECT 532.650 102.300 534.450 107.250 ;
        RECT 526.650 100.950 534.450 102.300 ;
        RECT 542.850 101.400 544.650 107.250 ;
        RECT 547.350 100.200 549.150 107.250 ;
        RECT 562.650 101.400 564.450 107.250 ;
        RECT 545.550 99.300 549.150 100.200 ;
        RECT 563.250 99.300 564.450 101.400 ;
        RECT 565.650 102.300 567.450 107.250 ;
        RECT 568.650 103.200 570.450 107.250 ;
        RECT 571.650 102.300 573.450 107.250 ;
        RECT 565.650 100.950 573.450 102.300 ;
        RECT 581.550 102.300 583.350 107.250 ;
        RECT 584.550 103.200 586.350 107.250 ;
        RECT 587.550 102.300 589.350 107.250 ;
        RECT 581.550 100.950 589.350 102.300 ;
        RECT 590.550 101.400 592.350 107.250 ;
        RECT 603.000 101.400 604.800 107.250 ;
        RECT 607.200 103.050 609.000 107.250 ;
        RECT 610.500 104.400 612.300 107.250 ;
        RECT 607.200 101.400 612.900 103.050 ;
        RECT 590.550 99.300 591.750 101.400 ;
        RECT 448.950 89.850 451.050 91.950 ;
        RECT 451.950 91.050 454.050 93.150 ;
        RECT 469.950 92.850 472.050 94.950 ;
        RECT 485.400 93.150 486.600 97.350 ;
        RECT 490.950 96.450 493.050 97.050 ;
        RECT 496.950 96.450 499.050 97.050 ;
        RECT 490.950 95.550 499.050 96.450 ;
        RECT 490.950 94.950 493.050 95.550 ;
        RECT 496.950 94.950 499.050 95.550 ;
        RECT 503.100 93.150 504.900 94.950 ;
        RECT 430.950 88.050 432.750 89.850 ;
        RECT 368.550 75.750 370.350 81.600 ;
        RECT 371.550 75.750 373.350 81.600 ;
        RECT 374.550 75.750 376.350 81.600 ;
        RECT 388.650 75.750 390.450 81.600 ;
        RECT 391.650 75.750 393.450 81.600 ;
        RECT 394.650 75.750 396.450 81.600 ;
        RECT 408.450 75.750 410.250 87.600 ;
        RECT 412.650 75.750 414.450 87.600 ;
        RECT 423.300 75.750 425.100 87.600 ;
        RECT 427.500 75.750 429.300 87.600 ;
        RECT 449.250 81.600 450.450 89.850 ;
        RECT 470.700 87.600 471.900 92.850 ;
        RECT 484.950 91.050 487.050 93.150 ;
        RECT 461.550 86.700 469.350 87.600 ;
        RECT 430.800 75.750 432.600 81.600 ;
        RECT 445.650 75.750 447.450 81.600 ;
        RECT 448.650 75.750 450.450 81.600 ;
        RECT 451.650 75.750 453.450 81.600 ;
        RECT 461.550 75.750 463.350 86.700 ;
        RECT 464.550 75.750 466.350 85.800 ;
        RECT 467.550 75.750 469.350 86.700 ;
        RECT 470.550 75.750 472.350 87.600 ;
        RECT 485.250 82.800 486.300 91.050 ;
        RECT 487.950 89.850 490.050 91.950 ;
        RECT 493.950 89.850 496.050 91.950 ;
        RECT 502.950 91.050 505.050 93.150 ;
        RECT 506.550 91.950 507.750 99.300 ;
        RECT 524.250 98.250 528.000 99.300 ;
        RECT 526.950 94.950 528.150 98.250 ;
        RECT 530.100 96.150 531.900 97.950 ;
        RECT 509.100 93.150 510.900 94.950 ;
        RECT 505.950 89.850 508.050 91.950 ;
        RECT 508.950 91.050 511.050 93.150 ;
        RECT 526.950 92.850 529.050 94.950 ;
        RECT 529.950 94.050 532.050 96.150 ;
        RECT 532.950 92.850 535.050 94.950 ;
        RECT 542.100 93.150 543.900 94.950 ;
        RECT 523.950 89.850 526.050 91.950 ;
        RECT 487.950 88.050 489.750 89.850 ;
        RECT 490.950 86.850 493.050 88.950 ;
        RECT 494.100 88.050 495.900 89.850 ;
        RECT 491.100 85.050 492.900 86.850 ;
        RECT 485.250 81.900 492.300 82.800 ;
        RECT 485.250 81.600 486.450 81.900 ;
        RECT 484.650 75.750 486.450 81.600 ;
        RECT 490.650 81.600 492.300 81.900 ;
        RECT 506.550 81.600 507.750 89.850 ;
        RECT 524.250 88.050 526.050 89.850 ;
        RECT 527.850 87.600 529.050 92.850 ;
        RECT 533.100 91.050 534.900 92.850 ;
        RECT 541.950 91.050 544.050 93.150 ;
        RECT 545.550 91.950 546.750 99.300 ;
        RECT 563.250 98.250 567.000 99.300 ;
        RECT 588.000 98.250 591.750 99.300 ;
        RECT 553.950 96.450 556.050 97.050 ;
        RECT 559.950 96.450 562.050 97.050 ;
        RECT 553.950 95.550 562.050 96.450 ;
        RECT 553.950 94.950 556.050 95.550 ;
        RECT 559.950 94.950 562.050 95.550 ;
        RECT 565.950 94.950 567.150 98.250 ;
        RECT 569.100 96.150 570.900 97.950 ;
        RECT 584.100 96.150 585.900 97.950 ;
        RECT 548.100 93.150 549.900 94.950 ;
        RECT 544.950 89.850 547.050 91.950 ;
        RECT 547.950 91.050 550.050 93.150 ;
        RECT 565.950 92.850 568.050 94.950 ;
        RECT 568.950 94.050 571.050 96.150 ;
        RECT 571.950 92.850 574.050 94.950 ;
        RECT 580.950 92.850 583.050 94.950 ;
        RECT 583.950 94.050 586.050 96.150 ;
        RECT 587.850 94.950 589.050 98.250 ;
        RECT 602.100 96.150 603.900 97.950 ;
        RECT 586.950 92.850 589.050 94.950 ;
        RECT 601.950 94.050 604.050 96.150 ;
        RECT 604.950 95.850 607.050 97.950 ;
        RECT 608.100 96.150 609.900 97.950 ;
        RECT 605.100 94.050 606.900 95.850 ;
        RECT 607.950 94.050 610.050 96.150 ;
        RECT 611.700 94.950 612.900 101.400 ;
        RECT 626.550 102.300 628.350 107.250 ;
        RECT 629.550 103.200 631.350 107.250 ;
        RECT 632.550 102.300 634.350 107.250 ;
        RECT 626.550 100.950 634.350 102.300 ;
        RECT 635.550 101.400 637.350 107.250 ;
        RECT 649.650 104.400 651.450 107.250 ;
        RECT 652.650 104.400 654.450 107.250 ;
        RECT 665.700 104.400 667.500 107.250 ;
        RECT 635.550 99.300 636.750 101.400 ;
        RECT 633.000 98.250 636.750 99.300 ;
        RECT 629.100 96.150 630.900 97.950 ;
        RECT 610.950 92.850 613.050 94.950 ;
        RECT 625.950 92.850 628.050 94.950 ;
        RECT 628.950 94.050 631.050 96.150 ;
        RECT 632.850 94.950 634.050 98.250 ;
        RECT 650.400 96.150 651.600 104.400 ;
        RECT 669.000 103.050 670.800 107.250 ;
        RECT 665.100 101.400 670.800 103.050 ;
        RECT 673.200 101.400 675.000 107.250 ;
        RECT 685.650 101.400 687.450 107.250 ;
        RECT 631.950 92.850 634.050 94.950 ;
        RECT 649.950 94.050 652.050 96.150 ;
        RECT 652.950 95.850 655.050 97.950 ;
        RECT 653.100 94.050 654.900 95.850 ;
        RECT 665.100 94.950 666.300 101.400 ;
        RECT 686.250 99.300 687.450 101.400 ;
        RECT 688.650 102.300 690.450 107.250 ;
        RECT 691.650 103.200 693.450 107.250 ;
        RECT 694.650 102.300 696.450 107.250 ;
        RECT 688.650 100.950 696.450 102.300 ;
        RECT 706.650 101.400 708.450 107.250 ;
        RECT 707.250 99.300 708.450 101.400 ;
        RECT 709.650 102.300 711.450 107.250 ;
        RECT 712.650 103.200 714.450 107.250 ;
        RECT 715.650 102.300 717.450 107.250 ;
        RECT 709.650 100.950 717.450 102.300 ;
        RECT 728.550 102.300 730.350 107.250 ;
        RECT 731.550 103.200 733.350 107.250 ;
        RECT 734.550 102.300 736.350 107.250 ;
        RECT 728.550 100.950 736.350 102.300 ;
        RECT 737.550 101.400 739.350 107.250 ;
        RECT 749.550 104.400 751.350 107.250 ;
        RECT 752.550 104.400 754.350 107.250 ;
        RECT 767.550 104.400 769.350 107.250 ;
        RECT 737.550 99.300 738.750 101.400 ;
        RECT 686.250 98.250 690.000 99.300 ;
        RECT 707.250 98.250 711.000 99.300 ;
        RECT 735.000 98.250 738.750 99.300 ;
        RECT 668.100 96.150 669.900 97.950 ;
        RECT 562.950 89.850 565.050 91.950 ;
        RECT 487.650 75.750 489.450 81.000 ;
        RECT 490.650 75.750 492.450 81.600 ;
        RECT 493.650 75.750 495.450 81.600 ;
        RECT 503.550 75.750 505.350 81.600 ;
        RECT 506.550 75.750 508.350 81.600 ;
        RECT 509.550 75.750 511.350 81.600 ;
        RECT 524.400 75.750 526.200 81.600 ;
        RECT 527.700 75.750 529.500 87.600 ;
        RECT 531.900 75.750 533.700 87.600 ;
        RECT 545.550 81.600 546.750 89.850 ;
        RECT 563.250 88.050 565.050 89.850 ;
        RECT 566.850 87.600 568.050 92.850 ;
        RECT 572.100 91.050 573.900 92.850 ;
        RECT 581.100 91.050 582.900 92.850 ;
        RECT 586.950 87.600 588.150 92.850 ;
        RECT 589.950 89.850 592.050 91.950 ;
        RECT 589.950 88.050 591.750 89.850 ;
        RECT 611.700 87.600 612.900 92.850 ;
        RECT 626.100 91.050 627.900 92.850 ;
        RECT 631.950 87.600 633.150 92.850 ;
        RECT 634.950 89.850 637.050 91.950 ;
        RECT 634.950 88.050 636.750 89.850 ;
        RECT 542.550 75.750 544.350 81.600 ;
        RECT 545.550 75.750 547.350 81.600 ;
        RECT 548.550 75.750 550.350 81.600 ;
        RECT 563.400 75.750 565.200 81.600 ;
        RECT 566.700 75.750 568.500 87.600 ;
        RECT 570.900 75.750 572.700 87.600 ;
        RECT 582.300 75.750 584.100 87.600 ;
        RECT 586.500 75.750 588.300 87.600 ;
        RECT 602.550 86.700 610.350 87.600 ;
        RECT 589.800 75.750 591.600 81.600 ;
        RECT 602.550 75.750 604.350 86.700 ;
        RECT 605.550 75.750 607.350 85.800 ;
        RECT 608.550 75.750 610.350 86.700 ;
        RECT 611.550 75.750 613.350 87.600 ;
        RECT 627.300 75.750 629.100 87.600 ;
        RECT 631.500 75.750 633.300 87.600 ;
        RECT 650.400 81.600 651.600 94.050 ;
        RECT 664.950 92.850 667.050 94.950 ;
        RECT 667.950 94.050 670.050 96.150 ;
        RECT 670.950 95.850 673.050 97.950 ;
        RECT 674.100 96.150 675.900 97.950 ;
        RECT 671.100 94.050 672.900 95.850 ;
        RECT 673.950 94.050 676.050 96.150 ;
        RECT 688.950 94.950 690.150 98.250 ;
        RECT 692.100 96.150 693.900 97.950 ;
        RECT 688.950 92.850 691.050 94.950 ;
        RECT 691.950 94.050 694.050 96.150 ;
        RECT 709.950 94.950 711.150 98.250 ;
        RECT 713.100 96.150 714.900 97.950 ;
        RECT 731.100 96.150 732.900 97.950 ;
        RECT 694.950 92.850 697.050 94.950 ;
        RECT 709.950 92.850 712.050 94.950 ;
        RECT 712.950 94.050 715.050 96.150 ;
        RECT 715.950 92.850 718.050 94.950 ;
        RECT 727.950 92.850 730.050 94.950 ;
        RECT 730.950 94.050 733.050 96.150 ;
        RECT 734.850 94.950 736.050 98.250 ;
        RECT 748.950 95.850 751.050 97.950 ;
        RECT 752.400 96.150 753.600 104.400 ;
        RECT 768.150 100.500 769.350 104.400 ;
        RECT 770.850 101.400 772.650 107.250 ;
        RECT 773.850 101.400 775.650 107.250 ;
        RECT 787.650 101.400 789.450 107.250 ;
        RECT 768.150 99.600 773.250 100.500 ;
        RECT 771.000 98.700 773.250 99.600 ;
        RECT 733.950 92.850 736.050 94.950 ;
        RECT 749.100 94.050 750.900 95.850 ;
        RECT 751.950 94.050 754.050 96.150 ;
        RECT 665.100 87.600 666.300 92.850 ;
        RECT 685.950 89.850 688.050 91.950 ;
        RECT 686.250 88.050 688.050 89.850 ;
        RECT 689.850 87.600 691.050 92.850 ;
        RECT 695.100 91.050 696.900 92.850 ;
        RECT 706.950 89.850 709.050 91.950 ;
        RECT 707.250 88.050 709.050 89.850 ;
        RECT 710.850 87.600 712.050 92.850 ;
        RECT 716.100 91.050 717.900 92.850 ;
        RECT 728.100 91.050 729.900 92.850 ;
        RECT 733.950 87.600 735.150 92.850 ;
        RECT 736.950 89.850 739.050 91.950 ;
        RECT 736.950 88.050 738.750 89.850 ;
        RECT 634.800 75.750 636.600 81.600 ;
        RECT 649.650 75.750 651.450 81.600 ;
        RECT 652.650 75.750 654.450 81.600 ;
        RECT 664.650 75.750 666.450 87.600 ;
        RECT 667.650 86.700 675.450 87.600 ;
        RECT 667.650 75.750 669.450 86.700 ;
        RECT 670.650 75.750 672.450 85.800 ;
        RECT 673.650 75.750 675.450 86.700 ;
        RECT 686.400 75.750 688.200 81.600 ;
        RECT 689.700 75.750 691.500 87.600 ;
        RECT 693.900 75.750 695.700 87.600 ;
        RECT 707.400 75.750 709.200 81.600 ;
        RECT 710.700 75.750 712.500 87.600 ;
        RECT 714.900 75.750 716.700 87.600 ;
        RECT 729.300 75.750 731.100 87.600 ;
        RECT 733.500 75.750 735.300 87.600 ;
        RECT 752.400 81.600 753.600 94.050 ;
        RECT 766.950 92.850 769.050 94.950 ;
        RECT 767.100 91.050 768.900 92.850 ;
        RECT 771.000 90.300 772.050 98.700 ;
        RECT 774.150 94.950 775.350 101.400 ;
        RECT 788.250 99.300 789.450 101.400 ;
        RECT 790.650 102.300 792.450 107.250 ;
        RECT 793.650 103.200 795.450 107.250 ;
        RECT 796.650 102.300 798.450 107.250 ;
        RECT 790.650 100.950 798.450 102.300 ;
        RECT 806.550 102.300 808.350 107.250 ;
        RECT 809.550 103.200 811.350 107.250 ;
        RECT 812.550 102.300 814.350 107.250 ;
        RECT 806.550 100.950 814.350 102.300 ;
        RECT 815.550 101.400 817.350 107.250 ;
        RECT 829.650 101.400 831.450 107.250 ;
        RECT 815.550 99.300 816.750 101.400 ;
        RECT 788.250 98.250 792.000 99.300 ;
        RECT 813.000 98.250 816.750 99.300 ;
        RECT 830.250 99.300 831.450 101.400 ;
        RECT 832.650 102.300 834.450 107.250 ;
        RECT 835.650 103.200 837.450 107.250 ;
        RECT 838.650 102.300 840.450 107.250 ;
        RECT 848.550 104.400 850.350 107.250 ;
        RECT 851.550 104.400 853.350 107.250 ;
        RECT 854.550 104.400 856.350 107.250 ;
        RECT 832.650 100.950 840.450 102.300 ;
        RECT 830.250 98.250 834.000 99.300 ;
        RECT 772.950 92.850 775.350 94.950 ;
        RECT 790.950 94.950 792.150 98.250 ;
        RECT 794.100 96.150 795.900 97.950 ;
        RECT 809.100 96.150 810.900 97.950 ;
        RECT 790.950 92.850 793.050 94.950 ;
        RECT 793.950 94.050 796.050 96.150 ;
        RECT 796.950 92.850 799.050 94.950 ;
        RECT 805.950 92.850 808.050 94.950 ;
        RECT 808.950 94.050 811.050 96.150 ;
        RECT 812.850 94.950 814.050 98.250 ;
        RECT 811.950 92.850 814.050 94.950 ;
        RECT 832.950 94.950 834.150 98.250 ;
        RECT 852.000 97.950 853.050 104.400 ;
        RECT 836.100 96.150 837.900 97.950 ;
        RECT 832.950 92.850 835.050 94.950 ;
        RECT 835.950 94.050 838.050 96.150 ;
        RECT 850.950 95.850 853.050 97.950 ;
        RECT 838.950 92.850 841.050 94.950 ;
        RECT 847.950 92.850 850.050 94.950 ;
        RECT 771.000 89.400 773.250 90.300 ;
        RECT 767.550 88.500 773.250 89.400 ;
        RECT 767.550 81.600 768.750 88.500 ;
        RECT 774.150 87.600 775.350 92.850 ;
        RECT 787.950 89.850 790.050 91.950 ;
        RECT 788.250 88.050 790.050 89.850 ;
        RECT 791.850 87.600 793.050 92.850 ;
        RECT 797.100 91.050 798.900 92.850 ;
        RECT 806.100 91.050 807.900 92.850 ;
        RECT 811.950 87.600 813.150 92.850 ;
        RECT 814.950 89.850 817.050 91.950 ;
        RECT 829.950 89.850 832.050 91.950 ;
        RECT 814.950 88.050 816.750 89.850 ;
        RECT 830.250 88.050 832.050 89.850 ;
        RECT 833.850 87.600 835.050 92.850 ;
        RECT 839.100 91.050 840.900 92.850 ;
        RECT 848.100 91.050 849.900 92.850 ;
        RECT 852.000 88.650 853.050 95.850 ;
        RECT 853.950 92.850 856.050 94.950 ;
        RECT 854.100 91.050 855.900 92.850 ;
        RECT 852.000 87.600 854.550 88.650 ;
        RECT 736.800 75.750 738.600 81.600 ;
        RECT 749.550 75.750 751.350 81.600 ;
        RECT 752.550 75.750 754.350 81.600 ;
        RECT 767.550 75.750 769.350 81.600 ;
        RECT 770.850 75.750 772.650 87.600 ;
        RECT 773.850 75.750 775.650 87.600 ;
        RECT 788.400 75.750 790.200 81.600 ;
        RECT 791.700 75.750 793.500 87.600 ;
        RECT 795.900 75.750 797.700 87.600 ;
        RECT 807.300 75.750 809.100 87.600 ;
        RECT 811.500 75.750 813.300 87.600 ;
        RECT 814.800 75.750 816.600 81.600 ;
        RECT 830.400 75.750 832.200 81.600 ;
        RECT 833.700 75.750 835.500 87.600 ;
        RECT 837.900 75.750 839.700 87.600 ;
        RECT 848.550 75.750 850.350 87.600 ;
        RECT 852.750 75.750 854.550 87.600 ;
        RECT 10.650 65.400 12.450 71.250 ;
        RECT 13.650 66.000 15.450 71.250 ;
        RECT 11.250 65.100 12.450 65.400 ;
        RECT 16.650 65.400 18.450 71.250 ;
        RECT 19.650 65.400 21.450 71.250 ;
        RECT 32.400 65.400 34.200 71.250 ;
        RECT 16.650 65.100 18.300 65.400 ;
        RECT 11.250 64.200 18.300 65.100 ;
        RECT 11.250 55.950 12.300 64.200 ;
        RECT 17.100 60.150 18.900 61.950 ;
        RECT 13.950 57.150 15.750 58.950 ;
        RECT 16.950 58.050 19.050 60.150 ;
        RECT 35.700 59.400 37.500 71.250 ;
        RECT 39.900 59.400 41.700 71.250 ;
        RECT 56.400 65.400 58.200 71.250 ;
        RECT 59.700 59.400 61.500 71.250 ;
        RECT 63.900 59.400 65.700 71.250 ;
        RECT 76.650 65.400 78.450 71.250 ;
        RECT 79.650 66.000 81.450 71.250 ;
        RECT 77.250 65.100 78.450 65.400 ;
        RECT 82.650 65.400 84.450 71.250 ;
        RECT 85.650 65.400 87.450 71.250 ;
        RECT 82.650 65.100 84.300 65.400 ;
        RECT 77.250 64.200 84.300 65.100 ;
        RECT 20.100 57.150 21.900 58.950 ;
        RECT 32.250 57.150 34.050 58.950 ;
        RECT 10.950 53.850 13.050 55.950 ;
        RECT 13.950 55.050 16.050 57.150 ;
        RECT 19.950 55.050 22.050 57.150 ;
        RECT 31.950 55.050 34.050 57.150 ;
        RECT 35.850 54.150 37.050 59.400 ;
        RECT 56.250 57.150 58.050 58.950 ;
        RECT 41.100 54.150 42.900 55.950 ;
        RECT 55.950 55.050 58.050 57.150 ;
        RECT 59.850 54.150 61.050 59.400 ;
        RECT 77.250 55.950 78.300 64.200 ;
        RECT 83.100 60.150 84.900 61.950 ;
        RECT 79.950 57.150 81.750 58.950 ;
        RECT 82.950 58.050 85.050 60.150 ;
        RECT 97.050 59.400 98.850 71.250 ;
        RECT 100.050 59.400 101.850 71.250 ;
        RECT 103.650 65.400 105.450 71.250 ;
        RECT 106.650 65.400 108.450 71.250 ;
        RECT 118.650 65.400 120.450 71.250 ;
        RECT 121.650 66.000 123.450 71.250 ;
        RECT 86.100 57.150 87.900 58.950 ;
        RECT 65.100 54.150 66.900 55.950 ;
        RECT 11.400 49.650 12.600 53.850 ;
        RECT 34.950 52.050 37.050 54.150 ;
        RECT 11.400 48.000 15.900 49.650 ;
        RECT 34.950 48.750 36.150 52.050 ;
        RECT 37.950 50.850 40.050 52.950 ;
        RECT 40.950 52.050 43.050 54.150 ;
        RECT 58.950 52.050 61.050 54.150 ;
        RECT 38.100 49.050 39.900 50.850 ;
        RECT 58.950 48.750 60.150 52.050 ;
        RECT 61.950 50.850 64.050 52.950 ;
        RECT 64.950 52.050 67.050 54.150 ;
        RECT 76.950 53.850 79.050 55.950 ;
        RECT 79.950 55.050 82.050 57.150 ;
        RECT 85.950 55.050 88.050 57.150 ;
        RECT 97.650 54.150 98.850 59.400 ;
        RECT 62.100 49.050 63.900 50.850 ;
        RECT 77.400 49.650 78.600 53.850 ;
        RECT 97.650 52.050 100.050 54.150 ;
        RECT 100.950 53.850 103.050 55.950 ;
        RECT 101.100 52.050 102.900 53.850 ;
        RECT 14.100 39.750 15.900 48.000 ;
        RECT 19.500 39.750 21.300 48.600 ;
        RECT 32.250 47.700 36.000 48.750 ;
        RECT 56.250 47.700 60.000 48.750 ;
        RECT 77.400 48.000 81.900 49.650 ;
        RECT 32.250 45.600 33.450 47.700 ;
        RECT 31.650 39.750 33.450 45.600 ;
        RECT 34.650 44.700 42.450 46.050 ;
        RECT 56.250 45.600 57.450 47.700 ;
        RECT 34.650 39.750 36.450 44.700 ;
        RECT 37.650 39.750 39.450 43.800 ;
        RECT 40.650 39.750 42.450 44.700 ;
        RECT 55.650 39.750 57.450 45.600 ;
        RECT 58.650 44.700 66.450 46.050 ;
        RECT 58.650 39.750 60.450 44.700 ;
        RECT 61.650 39.750 63.450 43.800 ;
        RECT 64.650 39.750 66.450 44.700 ;
        RECT 80.100 39.750 81.900 48.000 ;
        RECT 85.500 39.750 87.300 48.600 ;
        RECT 97.650 45.600 98.850 52.050 ;
        RECT 104.100 48.300 105.300 65.400 ;
        RECT 119.250 65.100 120.450 65.400 ;
        RECT 124.650 65.400 126.450 71.250 ;
        RECT 127.650 65.400 129.450 71.250 ;
        RECT 124.650 65.100 126.300 65.400 ;
        RECT 119.250 64.200 126.300 65.100 ;
        RECT 119.250 55.950 120.300 64.200 ;
        RECT 125.100 60.150 126.900 61.950 ;
        RECT 121.950 57.150 123.750 58.950 ;
        RECT 124.950 58.050 127.050 60.150 ;
        RECT 139.650 59.400 141.450 71.250 ;
        RECT 142.650 60.300 144.450 71.250 ;
        RECT 145.650 61.200 147.450 71.250 ;
        RECT 148.650 60.300 150.450 71.250 ;
        RECT 158.550 65.400 160.350 71.250 ;
        RECT 161.550 65.400 163.350 71.250 ;
        RECT 164.550 66.000 166.350 71.250 ;
        RECT 161.700 65.100 163.350 65.400 ;
        RECT 167.550 65.400 169.350 71.250 ;
        RECT 167.550 65.100 168.750 65.400 ;
        RECT 161.700 64.200 168.750 65.100 ;
        RECT 142.650 59.400 150.450 60.300 ;
        RECT 161.100 60.150 162.900 61.950 ;
        RECT 128.100 57.150 129.900 58.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 106.950 52.050 109.050 54.150 ;
        RECT 118.950 53.850 121.050 55.950 ;
        RECT 121.950 55.050 124.050 57.150 ;
        RECT 127.950 55.050 130.050 57.150 ;
        RECT 140.100 54.150 141.300 59.400 ;
        RECT 158.100 57.150 159.900 58.950 ;
        RECT 160.950 58.050 163.050 60.150 ;
        RECT 164.250 57.150 166.050 58.950 ;
        RECT 157.950 55.050 160.050 57.150 ;
        RECT 163.950 55.050 166.050 57.150 ;
        RECT 167.700 55.950 168.750 64.200 ;
        RECT 183.150 60.900 184.950 71.250 ;
        RECT 182.550 59.550 184.950 60.900 ;
        RECT 186.150 59.550 187.950 71.250 ;
        RECT 119.400 49.650 120.600 53.850 ;
        RECT 139.950 52.050 142.050 54.150 ;
        RECT 166.950 53.850 169.050 55.950 ;
        RECT 100.950 47.100 108.450 48.300 ;
        RECT 119.400 48.000 123.900 49.650 ;
        RECT 100.950 46.500 102.750 47.100 ;
        RECT 97.650 44.100 100.950 45.600 ;
        RECT 99.150 39.750 100.950 44.100 ;
        RECT 102.150 39.750 103.950 45.600 ;
        RECT 106.650 39.750 108.450 47.100 ;
        RECT 122.100 39.750 123.900 48.000 ;
        RECT 127.500 39.750 129.300 48.600 ;
        RECT 140.100 45.600 141.300 52.050 ;
        RECT 142.950 50.850 145.050 52.950 ;
        RECT 146.100 51.150 147.900 52.950 ;
        RECT 143.100 49.050 144.900 50.850 ;
        RECT 145.950 49.050 148.050 51.150 ;
        RECT 148.950 50.850 151.050 52.950 ;
        RECT 149.100 49.050 150.900 50.850 ;
        RECT 167.400 49.650 168.600 53.850 ;
        RECT 182.550 52.950 183.900 59.550 ;
        RECT 190.650 59.400 192.450 71.250 ;
        RECT 202.650 65.400 204.450 71.250 ;
        RECT 205.650 66.000 207.450 71.250 ;
        RECT 185.250 58.200 187.050 58.650 ;
        RECT 191.250 58.200 192.450 59.400 ;
        RECT 185.250 57.000 192.450 58.200 ;
        RECT 203.250 65.100 204.450 65.400 ;
        RECT 208.650 65.400 210.450 71.250 ;
        RECT 211.650 65.400 213.450 71.250 ;
        RECT 226.650 65.400 228.450 71.250 ;
        RECT 229.650 65.400 231.450 71.250 ;
        RECT 242.400 65.400 244.200 71.250 ;
        RECT 208.650 65.100 210.300 65.400 ;
        RECT 203.250 64.200 210.300 65.100 ;
        RECT 185.250 56.850 187.050 57.000 ;
        RECT 140.100 43.950 145.800 45.600 ;
        RECT 140.700 39.750 142.500 42.600 ;
        RECT 144.000 39.750 145.800 43.950 ;
        RECT 148.200 39.750 150.000 45.600 ;
        RECT 158.700 39.750 160.500 48.600 ;
        RECT 164.100 48.000 168.600 49.650 ;
        RECT 181.950 50.850 184.050 52.950 ;
        RECT 164.100 39.750 165.900 48.000 ;
        RECT 181.950 45.600 183.000 50.850 ;
        RECT 185.400 48.600 186.300 56.850 ;
        RECT 203.250 55.950 204.300 64.200 ;
        RECT 209.100 60.150 210.900 61.950 ;
        RECT 205.950 57.150 207.750 58.950 ;
        RECT 208.950 58.050 211.050 60.150 ;
        RECT 212.100 57.150 213.900 58.950 ;
        RECT 188.100 54.150 189.900 55.950 ;
        RECT 187.950 52.050 190.050 54.150 ;
        RECT 202.950 53.850 205.050 55.950 ;
        RECT 205.950 55.050 208.050 57.150 ;
        RECT 211.950 55.050 214.050 57.150 ;
        RECT 191.100 51.150 192.900 52.950 ;
        RECT 190.950 49.050 193.050 51.150 ;
        RECT 203.400 49.650 204.600 53.850 ;
        RECT 227.400 52.950 228.600 65.400 ;
        RECT 245.700 59.400 247.500 71.250 ;
        RECT 249.900 59.400 251.700 71.250 ;
        RECT 262.050 59.400 263.850 71.250 ;
        RECT 265.050 59.400 266.850 71.250 ;
        RECT 268.650 65.400 270.450 71.250 ;
        RECT 271.650 65.400 273.450 71.250 ;
        RECT 242.250 57.150 244.050 58.950 ;
        RECT 241.950 55.050 244.050 57.150 ;
        RECT 245.850 54.150 247.050 59.400 ;
        RECT 251.100 54.150 252.900 55.950 ;
        RECT 262.650 54.150 263.850 59.400 ;
        RECT 211.950 51.450 214.050 52.050 ;
        RECT 220.950 51.450 223.050 52.050 ;
        RECT 211.950 50.550 223.050 51.450 ;
        RECT 226.950 50.850 229.050 52.950 ;
        RECT 230.100 51.150 231.900 52.950 ;
        RECT 244.950 52.050 247.050 54.150 ;
        RECT 211.950 49.950 214.050 50.550 ;
        RECT 220.950 49.950 223.050 50.550 ;
        RECT 185.250 47.700 187.050 48.600 ;
        RECT 203.400 48.000 207.900 49.650 ;
        RECT 185.250 46.800 188.550 47.700 ;
        RECT 181.650 39.750 183.450 45.600 ;
        RECT 187.650 42.600 188.550 46.800 ;
        RECT 184.650 39.750 186.450 42.600 ;
        RECT 187.650 39.750 189.450 42.600 ;
        RECT 190.650 39.750 192.450 42.600 ;
        RECT 206.100 39.750 207.900 48.000 ;
        RECT 211.500 39.750 213.300 48.600 ;
        RECT 227.400 42.600 228.600 50.850 ;
        RECT 229.950 49.050 232.050 51.150 ;
        RECT 244.950 48.750 246.150 52.050 ;
        RECT 247.950 50.850 250.050 52.950 ;
        RECT 250.950 52.050 253.050 54.150 ;
        RECT 262.650 52.050 265.050 54.150 ;
        RECT 265.950 53.850 268.050 55.950 ;
        RECT 266.100 52.050 267.900 53.850 ;
        RECT 248.100 49.050 249.900 50.850 ;
        RECT 242.250 47.700 246.000 48.750 ;
        RECT 242.250 45.600 243.450 47.700 ;
        RECT 226.650 39.750 228.450 42.600 ;
        RECT 229.650 39.750 231.450 42.600 ;
        RECT 241.650 39.750 243.450 45.600 ;
        RECT 244.650 44.700 252.450 46.050 ;
        RECT 244.650 39.750 246.450 44.700 ;
        RECT 247.650 39.750 249.450 43.800 ;
        RECT 250.650 39.750 252.450 44.700 ;
        RECT 262.650 45.600 263.850 52.050 ;
        RECT 269.100 48.300 270.300 65.400 ;
        RECT 281.550 59.400 283.350 71.250 ;
        RECT 285.750 59.400 287.550 71.250 ;
        RECT 302.550 65.400 304.350 71.250 ;
        RECT 305.550 65.400 307.350 71.250 ;
        RECT 320.400 65.400 322.200 71.250 ;
        RECT 285.000 58.350 287.550 59.400 ;
        RECT 272.100 54.150 273.900 55.950 ;
        RECT 281.100 54.150 282.900 55.950 ;
        RECT 271.950 52.050 274.050 54.150 ;
        RECT 280.950 52.050 283.050 54.150 ;
        RECT 285.000 51.150 286.050 58.350 ;
        RECT 287.100 54.150 288.900 55.950 ;
        RECT 286.950 52.050 289.050 54.150 ;
        RECT 305.400 52.950 306.600 65.400 ;
        RECT 323.700 59.400 325.500 71.250 ;
        RECT 327.900 59.400 329.700 71.250 ;
        RECT 340.650 59.400 342.450 71.250 ;
        RECT 343.650 60.300 345.450 71.250 ;
        RECT 346.650 61.200 348.450 71.250 ;
        RECT 349.650 60.300 351.450 71.250 ;
        RECT 361.650 65.400 363.450 71.250 ;
        RECT 364.650 65.400 366.450 71.250 ;
        RECT 376.650 65.400 378.450 71.250 ;
        RECT 379.650 66.000 381.450 71.250 ;
        RECT 343.650 59.400 351.450 60.300 ;
        RECT 320.250 57.150 322.050 58.950 ;
        RECT 319.950 55.050 322.050 57.150 ;
        RECT 323.850 54.150 325.050 59.400 ;
        RECT 329.100 54.150 330.900 55.950 ;
        RECT 341.100 54.150 342.300 59.400 ;
        RECT 302.100 51.150 303.900 52.950 ;
        RECT 283.950 49.050 286.050 51.150 ;
        RECT 301.950 49.050 304.050 51.150 ;
        RECT 304.950 50.850 307.050 52.950 ;
        RECT 322.950 52.050 325.050 54.150 ;
        RECT 265.950 47.100 273.450 48.300 ;
        RECT 265.950 46.500 267.750 47.100 ;
        RECT 262.650 44.100 265.950 45.600 ;
        RECT 264.150 39.750 265.950 44.100 ;
        RECT 267.150 39.750 268.950 45.600 ;
        RECT 271.650 39.750 273.450 47.100 ;
        RECT 285.000 42.600 286.050 49.050 ;
        RECT 305.400 42.600 306.600 50.850 ;
        RECT 322.950 48.750 324.150 52.050 ;
        RECT 325.950 50.850 328.050 52.950 ;
        RECT 328.950 52.050 331.050 54.150 ;
        RECT 340.950 52.050 343.050 54.150 ;
        RECT 362.400 52.950 363.600 65.400 ;
        RECT 377.250 65.100 378.450 65.400 ;
        RECT 382.650 65.400 384.450 71.250 ;
        RECT 385.650 65.400 387.450 71.250 ;
        RECT 382.650 65.100 384.300 65.400 ;
        RECT 377.250 64.200 384.300 65.100 ;
        RECT 377.250 55.950 378.300 64.200 ;
        RECT 383.100 60.150 384.900 61.950 ;
        RECT 379.950 57.150 381.750 58.950 ;
        RECT 382.950 58.050 385.050 60.150 ;
        RECT 396.300 59.400 398.100 71.250 ;
        RECT 400.500 59.400 402.300 71.250 ;
        RECT 403.800 65.400 405.600 71.250 ;
        RECT 418.650 65.400 420.450 71.250 ;
        RECT 421.650 65.400 423.450 71.250 ;
        RECT 386.100 57.150 387.900 58.950 ;
        RECT 376.950 53.850 379.050 55.950 ;
        RECT 379.950 55.050 382.050 57.150 ;
        RECT 385.950 55.050 388.050 57.150 ;
        RECT 395.100 54.150 396.900 55.950 ;
        RECT 400.950 54.150 402.150 59.400 ;
        RECT 403.950 57.150 405.750 58.950 ;
        RECT 403.950 55.050 406.050 57.150 ;
        RECT 326.100 49.050 327.900 50.850 ;
        RECT 320.250 47.700 324.000 48.750 ;
        RECT 320.250 45.600 321.450 47.700 ;
        RECT 281.550 39.750 283.350 42.600 ;
        RECT 284.550 39.750 286.350 42.600 ;
        RECT 287.550 39.750 289.350 42.600 ;
        RECT 302.550 39.750 304.350 42.600 ;
        RECT 305.550 39.750 307.350 42.600 ;
        RECT 319.650 39.750 321.450 45.600 ;
        RECT 322.650 44.700 330.450 46.050 ;
        RECT 322.650 39.750 324.450 44.700 ;
        RECT 325.650 39.750 327.450 43.800 ;
        RECT 328.650 39.750 330.450 44.700 ;
        RECT 341.100 45.600 342.300 52.050 ;
        RECT 343.950 50.850 346.050 52.950 ;
        RECT 347.100 51.150 348.900 52.950 ;
        RECT 344.100 49.050 345.900 50.850 ;
        RECT 346.950 49.050 349.050 51.150 ;
        RECT 349.950 50.850 352.050 52.950 ;
        RECT 361.950 50.850 364.050 52.950 ;
        RECT 365.100 51.150 366.900 52.950 ;
        RECT 350.100 49.050 351.900 50.850 ;
        RECT 341.100 43.950 346.800 45.600 ;
        RECT 341.700 39.750 343.500 42.600 ;
        RECT 345.000 39.750 346.800 43.950 ;
        RECT 349.200 39.750 351.000 45.600 ;
        RECT 362.400 42.600 363.600 50.850 ;
        RECT 364.950 49.050 367.050 51.150 ;
        RECT 377.400 49.650 378.600 53.850 ;
        RECT 394.950 52.050 397.050 54.150 ;
        RECT 397.950 50.850 400.050 52.950 ;
        RECT 400.950 52.050 403.050 54.150 ;
        RECT 419.400 52.950 420.600 65.400 ;
        RECT 435.450 59.400 437.250 71.250 ;
        RECT 439.650 59.400 441.450 71.250 ;
        RECT 449.550 65.400 451.350 71.250 ;
        RECT 452.550 65.400 454.350 71.250 ;
        RECT 435.450 58.350 438.000 59.400 ;
        RECT 434.100 54.150 435.900 55.950 ;
        RECT 377.400 48.000 381.900 49.650 ;
        RECT 398.100 49.050 399.900 50.850 ;
        RECT 401.850 48.750 403.050 52.050 ;
        RECT 418.950 50.850 421.050 52.950 ;
        RECT 422.100 51.150 423.900 52.950 ;
        RECT 433.950 52.050 436.050 54.150 ;
        RECT 436.950 51.150 438.000 58.350 ;
        RECT 440.100 54.150 441.900 55.950 ;
        RECT 439.950 52.050 442.050 54.150 ;
        RECT 452.400 52.950 453.600 65.400 ;
        RECT 466.650 59.400 468.450 71.250 ;
        RECT 469.650 60.300 471.450 71.250 ;
        RECT 472.650 61.200 474.450 71.250 ;
        RECT 475.650 60.300 477.450 71.250 ;
        RECT 469.650 59.400 477.450 60.300 ;
        RECT 488.550 60.300 490.350 71.250 ;
        RECT 491.550 61.200 493.350 71.250 ;
        RECT 494.550 60.300 496.350 71.250 ;
        RECT 488.550 59.400 496.350 60.300 ;
        RECT 497.550 59.400 499.350 71.250 ;
        RECT 511.650 65.400 513.450 71.250 ;
        RECT 514.650 65.400 516.450 71.250 ;
        RECT 467.100 54.150 468.300 59.400 ;
        RECT 472.950 57.450 475.050 58.050 ;
        RECT 493.950 57.450 496.050 58.050 ;
        RECT 472.950 56.550 496.050 57.450 ;
        RECT 472.950 55.950 475.050 56.550 ;
        RECT 493.950 55.950 496.050 56.550 ;
        RECT 497.700 54.150 498.900 59.400 ;
        RECT 449.100 51.150 450.900 52.950 ;
        RECT 361.650 39.750 363.450 42.600 ;
        RECT 364.650 39.750 366.450 42.600 ;
        RECT 380.100 39.750 381.900 48.000 ;
        RECT 385.500 39.750 387.300 48.600 ;
        RECT 402.000 47.700 405.750 48.750 ;
        RECT 395.550 44.700 403.350 46.050 ;
        RECT 395.550 39.750 397.350 44.700 ;
        RECT 398.550 39.750 400.350 43.800 ;
        RECT 401.550 39.750 403.350 44.700 ;
        RECT 404.550 45.600 405.750 47.700 ;
        RECT 404.550 39.750 406.350 45.600 ;
        RECT 419.400 42.600 420.600 50.850 ;
        RECT 421.950 49.050 424.050 51.150 ;
        RECT 436.950 49.050 439.050 51.150 ;
        RECT 448.950 49.050 451.050 51.150 ;
        RECT 451.950 50.850 454.050 52.950 ;
        RECT 466.950 52.050 469.050 54.150 ;
        RECT 436.950 42.600 438.000 49.050 ;
        RECT 452.400 42.600 453.600 50.850 ;
        RECT 467.100 45.600 468.300 52.050 ;
        RECT 469.950 50.850 472.050 52.950 ;
        RECT 473.100 51.150 474.900 52.950 ;
        RECT 470.100 49.050 471.900 50.850 ;
        RECT 472.950 49.050 475.050 51.150 ;
        RECT 475.950 50.850 478.050 52.950 ;
        RECT 487.950 50.850 490.050 52.950 ;
        RECT 491.100 51.150 492.900 52.950 ;
        RECT 476.100 49.050 477.900 50.850 ;
        RECT 488.100 49.050 489.900 50.850 ;
        RECT 490.950 49.050 493.050 51.150 ;
        RECT 493.950 50.850 496.050 52.950 ;
        RECT 496.950 52.050 499.050 54.150 ;
        RECT 512.400 52.950 513.600 65.400 ;
        RECT 528.300 59.400 530.100 71.250 ;
        RECT 532.500 59.400 534.300 71.250 ;
        RECT 535.800 65.400 537.600 71.250 ;
        RECT 548.550 60.300 550.350 71.250 ;
        RECT 551.550 61.200 553.350 71.250 ;
        RECT 554.550 60.300 556.350 71.250 ;
        RECT 548.550 59.400 556.350 60.300 ;
        RECT 557.550 59.400 559.350 71.250 ;
        RECT 571.650 65.400 573.450 71.250 ;
        RECT 574.650 66.000 576.450 71.250 ;
        RECT 572.250 65.100 573.450 65.400 ;
        RECT 577.650 65.400 579.450 71.250 ;
        RECT 580.650 65.400 582.450 71.250 ;
        RECT 590.550 65.400 592.350 71.250 ;
        RECT 593.550 65.400 595.350 71.250 ;
        RECT 596.550 65.400 598.350 71.250 ;
        RECT 613.650 65.400 615.450 71.250 ;
        RECT 616.650 66.000 618.450 71.250 ;
        RECT 577.650 65.100 579.300 65.400 ;
        RECT 572.250 64.200 579.300 65.100 ;
        RECT 527.100 54.150 528.900 55.950 ;
        RECT 532.950 54.150 534.150 59.400 ;
        RECT 535.950 57.150 537.750 58.950 ;
        RECT 535.950 55.050 538.050 57.150 ;
        RECT 557.700 54.150 558.900 59.400 ;
        RECT 572.250 55.950 573.300 64.200 ;
        RECT 578.100 60.150 579.900 61.950 ;
        RECT 574.950 57.150 576.750 58.950 ;
        RECT 577.950 58.050 580.050 60.150 ;
        RECT 581.100 57.150 582.900 58.950 ;
        RECT 593.550 57.150 594.750 65.400 ;
        RECT 614.250 65.100 615.450 65.400 ;
        RECT 619.650 65.400 621.450 71.250 ;
        RECT 622.650 65.400 624.450 71.250 ;
        RECT 635.400 65.400 637.200 71.250 ;
        RECT 619.650 65.100 621.300 65.400 ;
        RECT 614.250 64.200 621.300 65.100 ;
        RECT 494.100 49.050 495.900 50.850 ;
        RECT 497.700 45.600 498.900 52.050 ;
        RECT 511.950 50.850 514.050 52.950 ;
        RECT 515.100 51.150 516.900 52.950 ;
        RECT 526.950 52.050 529.050 54.150 ;
        RECT 467.100 43.950 472.800 45.600 ;
        RECT 418.650 39.750 420.450 42.600 ;
        RECT 421.650 39.750 423.450 42.600 ;
        RECT 433.650 39.750 435.450 42.600 ;
        RECT 436.650 39.750 438.450 42.600 ;
        RECT 439.650 39.750 441.450 42.600 ;
        RECT 449.550 39.750 451.350 42.600 ;
        RECT 452.550 39.750 454.350 42.600 ;
        RECT 467.700 39.750 469.500 42.600 ;
        RECT 471.000 39.750 472.800 43.950 ;
        RECT 475.200 39.750 477.000 45.600 ;
        RECT 489.000 39.750 490.800 45.600 ;
        RECT 493.200 43.950 498.900 45.600 ;
        RECT 493.200 39.750 495.000 43.950 ;
        RECT 512.400 42.600 513.600 50.850 ;
        RECT 514.950 49.050 517.050 51.150 ;
        RECT 529.950 50.850 532.050 52.950 ;
        RECT 532.950 52.050 535.050 54.150 ;
        RECT 530.100 49.050 531.900 50.850 ;
        RECT 533.850 48.750 535.050 52.050 ;
        RECT 547.950 50.850 550.050 52.950 ;
        RECT 551.100 51.150 552.900 52.950 ;
        RECT 548.100 49.050 549.900 50.850 ;
        RECT 550.950 49.050 553.050 51.150 ;
        RECT 553.950 50.850 556.050 52.950 ;
        RECT 556.950 52.050 559.050 54.150 ;
        RECT 571.950 53.850 574.050 55.950 ;
        RECT 574.950 55.050 577.050 57.150 ;
        RECT 580.950 55.050 583.050 57.150 ;
        RECT 589.950 53.850 592.050 55.950 ;
        RECT 592.950 55.050 595.050 57.150 ;
        RECT 614.250 55.950 615.300 64.200 ;
        RECT 620.100 60.150 621.900 61.950 ;
        RECT 616.950 57.150 618.750 58.950 ;
        RECT 619.950 58.050 622.050 60.150 ;
        RECT 638.700 59.400 640.500 71.250 ;
        RECT 642.900 59.400 644.700 71.250 ;
        RECT 655.650 65.400 657.450 71.250 ;
        RECT 658.650 65.400 660.450 71.250 ;
        RECT 670.650 65.400 672.450 71.250 ;
        RECT 673.650 65.400 675.450 71.250 ;
        RECT 676.650 65.400 678.450 71.250 ;
        RECT 689.400 65.400 691.200 71.250 ;
        RECT 623.100 57.150 624.900 58.950 ;
        RECT 635.250 57.150 637.050 58.950 ;
        RECT 554.100 49.050 555.900 50.850 ;
        RECT 534.000 47.700 537.750 48.750 ;
        RECT 527.550 44.700 535.350 46.050 ;
        RECT 496.500 39.750 498.300 42.600 ;
        RECT 511.650 39.750 513.450 42.600 ;
        RECT 514.650 39.750 516.450 42.600 ;
        RECT 527.550 39.750 529.350 44.700 ;
        RECT 530.550 39.750 532.350 43.800 ;
        RECT 533.550 39.750 535.350 44.700 ;
        RECT 536.550 45.600 537.750 47.700 ;
        RECT 557.700 45.600 558.900 52.050 ;
        RECT 572.400 49.650 573.600 53.850 ;
        RECT 590.100 52.050 591.900 53.850 ;
        RECT 572.400 48.000 576.900 49.650 ;
        RECT 536.550 39.750 538.350 45.600 ;
        RECT 549.000 39.750 550.800 45.600 ;
        RECT 553.200 43.950 558.900 45.600 ;
        RECT 553.200 39.750 555.000 43.950 ;
        RECT 556.500 39.750 558.300 42.600 ;
        RECT 575.100 39.750 576.900 48.000 ;
        RECT 580.500 39.750 582.300 48.600 ;
        RECT 593.550 47.700 594.750 55.050 ;
        RECT 595.950 53.850 598.050 55.950 ;
        RECT 613.950 53.850 616.050 55.950 ;
        RECT 616.950 55.050 619.050 57.150 ;
        RECT 622.950 55.050 625.050 57.150 ;
        RECT 634.950 55.050 637.050 57.150 ;
        RECT 638.850 54.150 640.050 59.400 ;
        RECT 644.100 54.150 645.900 55.950 ;
        RECT 596.100 52.050 597.900 53.850 ;
        RECT 614.400 49.650 615.600 53.850 ;
        RECT 637.950 52.050 640.050 54.150 ;
        RECT 614.400 48.000 618.900 49.650 ;
        RECT 637.950 48.750 639.150 52.050 ;
        RECT 640.950 50.850 643.050 52.950 ;
        RECT 643.950 52.050 646.050 54.150 ;
        RECT 656.400 52.950 657.600 65.400 ;
        RECT 674.250 57.150 675.450 65.400 ;
        RECT 692.700 59.400 694.500 71.250 ;
        RECT 696.900 59.400 698.700 71.250 ;
        RECT 709.650 65.400 711.450 71.250 ;
        RECT 712.650 65.400 714.450 71.250 ;
        RECT 725.400 65.400 727.200 71.250 ;
        RECT 689.250 57.150 691.050 58.950 ;
        RECT 670.950 53.850 673.050 55.950 ;
        RECT 673.950 55.050 676.050 57.150 ;
        RECT 655.950 50.850 658.050 52.950 ;
        RECT 659.100 51.150 660.900 52.950 ;
        RECT 671.100 52.050 672.900 53.850 ;
        RECT 641.100 49.050 642.900 50.850 ;
        RECT 593.550 46.800 597.150 47.700 ;
        RECT 590.850 39.750 592.650 45.600 ;
        RECT 595.350 39.750 597.150 46.800 ;
        RECT 617.100 39.750 618.900 48.000 ;
        RECT 622.500 39.750 624.300 48.600 ;
        RECT 635.250 47.700 639.000 48.750 ;
        RECT 635.250 45.600 636.450 47.700 ;
        RECT 634.650 39.750 636.450 45.600 ;
        RECT 637.650 44.700 645.450 46.050 ;
        RECT 637.650 39.750 639.450 44.700 ;
        RECT 640.650 39.750 642.450 43.800 ;
        RECT 643.650 39.750 645.450 44.700 ;
        RECT 656.400 42.600 657.600 50.850 ;
        RECT 658.950 49.050 661.050 51.150 ;
        RECT 674.250 47.700 675.450 55.050 ;
        RECT 676.950 53.850 679.050 55.950 ;
        RECT 688.950 55.050 691.050 57.150 ;
        RECT 692.850 54.150 694.050 59.400 ;
        RECT 698.100 54.150 699.900 55.950 ;
        RECT 677.100 52.050 678.900 53.850 ;
        RECT 691.950 52.050 694.050 54.150 ;
        RECT 691.950 48.750 693.150 52.050 ;
        RECT 694.950 50.850 697.050 52.950 ;
        RECT 697.950 52.050 700.050 54.150 ;
        RECT 710.400 52.950 711.600 65.400 ;
        RECT 728.700 59.400 730.500 71.250 ;
        RECT 732.900 59.400 734.700 71.250 ;
        RECT 743.550 64.200 745.350 70.200 ;
        RECT 746.550 64.200 748.350 71.250 ;
        RECT 725.250 57.150 727.050 58.950 ;
        RECT 724.950 55.050 727.050 57.150 ;
        RECT 728.850 54.150 730.050 59.400 ;
        RECT 744.450 59.100 745.350 64.200 ;
        RECT 751.050 60.900 752.850 70.200 ;
        RECT 751.050 60.000 753.150 60.900 ;
        RECT 744.450 58.200 750.600 59.100 ;
        RECT 734.100 54.150 735.900 55.950 ;
        RECT 746.250 54.150 748.050 55.950 ;
        RECT 709.950 50.850 712.050 52.950 ;
        RECT 713.100 51.150 714.900 52.950 ;
        RECT 727.950 52.050 730.050 54.150 ;
        RECT 695.100 49.050 696.900 50.850 ;
        RECT 671.850 46.800 675.450 47.700 ;
        RECT 689.250 47.700 693.000 48.750 ;
        RECT 655.650 39.750 657.450 42.600 ;
        RECT 658.650 39.750 660.450 42.600 ;
        RECT 671.850 39.750 673.650 46.800 ;
        RECT 689.250 45.600 690.450 47.700 ;
        RECT 676.350 39.750 678.150 45.600 ;
        RECT 688.650 39.750 690.450 45.600 ;
        RECT 691.650 44.700 699.450 46.050 ;
        RECT 691.650 39.750 693.450 44.700 ;
        RECT 694.650 39.750 696.450 43.800 ;
        RECT 697.650 39.750 699.450 44.700 ;
        RECT 710.400 42.600 711.600 50.850 ;
        RECT 712.950 49.050 715.050 51.150 ;
        RECT 727.950 48.750 729.150 52.050 ;
        RECT 730.950 50.850 733.050 52.950 ;
        RECT 733.950 52.050 736.050 54.150 ;
        RECT 742.950 50.850 745.050 52.950 ;
        RECT 745.950 52.050 748.050 54.150 ;
        RECT 749.250 55.500 750.600 58.200 ;
        RECT 749.250 53.700 751.050 55.500 ;
        RECT 731.100 49.050 732.900 50.850 ;
        RECT 743.250 49.050 745.050 50.850 ;
        RECT 725.250 47.700 729.000 48.750 ;
        RECT 749.250 48.000 750.600 53.700 ;
        RECT 752.250 52.950 753.150 60.000 ;
        RECT 755.550 59.400 757.350 71.250 ;
        RECT 770.400 65.400 772.200 71.250 ;
        RECT 773.700 59.400 775.500 71.250 ;
        RECT 777.900 59.400 779.700 71.250 ;
        RECT 792.300 59.400 794.100 71.250 ;
        RECT 796.500 59.400 798.300 71.250 ;
        RECT 799.800 65.400 801.600 71.250 ;
        RECT 817.650 59.400 819.450 71.250 ;
        RECT 820.650 60.300 822.450 71.250 ;
        RECT 823.650 61.200 825.450 71.250 ;
        RECT 826.650 60.300 828.450 71.250 ;
        RECT 820.650 59.400 828.450 60.300 ;
        RECT 837.300 59.400 839.100 71.250 ;
        RECT 841.500 59.400 843.300 71.250 ;
        RECT 844.800 65.400 846.600 71.250 ;
        RECT 857.550 65.400 859.350 71.250 ;
        RECT 860.550 65.400 862.350 71.250 ;
        RECT 863.550 65.400 865.350 71.250 ;
        RECT 770.250 57.150 772.050 58.950 ;
        RECT 755.100 54.150 756.900 55.950 ;
        RECT 769.950 55.050 772.050 57.150 ;
        RECT 773.850 54.150 775.050 59.400 ;
        RECT 779.100 54.150 780.900 55.950 ;
        RECT 791.100 54.150 792.900 55.950 ;
        RECT 796.950 54.150 798.150 59.400 ;
        RECT 799.950 57.150 801.750 58.950 ;
        RECT 799.950 55.050 802.050 57.150 ;
        RECT 818.100 54.150 819.300 59.400 ;
        RECT 836.100 54.150 837.900 55.950 ;
        RECT 841.950 54.150 843.150 59.400 ;
        RECT 844.950 57.150 846.750 58.950 ;
        RECT 860.550 57.150 861.750 65.400 ;
        RECT 844.950 55.050 847.050 57.150 ;
        RECT 751.950 50.850 754.050 52.950 ;
        RECT 754.950 52.050 757.050 54.150 ;
        RECT 772.950 52.050 775.050 54.150 ;
        RECT 725.250 45.600 726.450 47.700 ;
        RECT 744.300 47.100 750.600 48.000 ;
        RECT 709.650 39.750 711.450 42.600 ;
        RECT 712.650 39.750 714.450 42.600 ;
        RECT 724.650 39.750 726.450 45.600 ;
        RECT 727.650 44.700 735.450 46.050 ;
        RECT 727.650 39.750 729.450 44.700 ;
        RECT 730.650 39.750 732.450 43.800 ;
        RECT 733.650 39.750 735.450 44.700 ;
        RECT 744.300 43.800 745.350 47.100 ;
        RECT 752.250 46.200 753.150 50.850 ;
        RECT 772.950 48.750 774.150 52.050 ;
        RECT 775.950 50.850 778.050 52.950 ;
        RECT 778.950 52.050 781.050 54.150 ;
        RECT 790.950 52.050 793.050 54.150 ;
        RECT 793.950 50.850 796.050 52.950 ;
        RECT 796.950 52.050 799.050 54.150 ;
        RECT 817.950 52.050 820.050 54.150 ;
        RECT 776.100 49.050 777.900 50.850 ;
        RECT 794.100 49.050 795.900 50.850 ;
        RECT 797.850 48.750 799.050 52.050 ;
        RECT 770.250 47.700 774.000 48.750 ;
        RECT 798.000 47.700 801.750 48.750 ;
        RECT 751.050 45.300 753.150 46.200 ;
        RECT 743.550 40.800 745.350 43.800 ;
        RECT 746.550 39.750 748.350 43.800 ;
        RECT 751.050 40.800 752.850 45.300 ;
        RECT 755.550 39.750 757.350 46.800 ;
        RECT 770.250 45.600 771.450 47.700 ;
        RECT 769.650 39.750 771.450 45.600 ;
        RECT 772.650 44.700 780.450 46.050 ;
        RECT 772.650 39.750 774.450 44.700 ;
        RECT 775.650 39.750 777.450 43.800 ;
        RECT 778.650 39.750 780.450 44.700 ;
        RECT 791.550 44.700 799.350 46.050 ;
        RECT 791.550 39.750 793.350 44.700 ;
        RECT 794.550 39.750 796.350 43.800 ;
        RECT 797.550 39.750 799.350 44.700 ;
        RECT 800.550 45.600 801.750 47.700 ;
        RECT 818.100 45.600 819.300 52.050 ;
        RECT 820.950 50.850 823.050 52.950 ;
        RECT 824.100 51.150 825.900 52.950 ;
        RECT 821.100 49.050 822.900 50.850 ;
        RECT 823.950 49.050 826.050 51.150 ;
        RECT 826.950 50.850 829.050 52.950 ;
        RECT 835.950 52.050 838.050 54.150 ;
        RECT 838.950 50.850 841.050 52.950 ;
        RECT 841.950 52.050 844.050 54.150 ;
        RECT 856.950 53.850 859.050 55.950 ;
        RECT 859.950 55.050 862.050 57.150 ;
        RECT 857.100 52.050 858.900 53.850 ;
        RECT 827.100 49.050 828.900 50.850 ;
        RECT 839.100 49.050 840.900 50.850 ;
        RECT 842.850 48.750 844.050 52.050 ;
        RECT 843.000 47.700 846.750 48.750 ;
        RECT 800.550 39.750 802.350 45.600 ;
        RECT 818.100 43.950 823.800 45.600 ;
        RECT 818.700 39.750 820.500 42.600 ;
        RECT 822.000 39.750 823.800 43.950 ;
        RECT 826.200 39.750 828.000 45.600 ;
        RECT 836.550 44.700 844.350 46.050 ;
        RECT 836.550 39.750 838.350 44.700 ;
        RECT 839.550 39.750 841.350 43.800 ;
        RECT 842.550 39.750 844.350 44.700 ;
        RECT 845.550 45.600 846.750 47.700 ;
        RECT 860.550 47.700 861.750 55.050 ;
        RECT 862.950 53.850 865.050 55.950 ;
        RECT 863.100 52.050 864.900 53.850 ;
        RECT 860.550 46.800 864.150 47.700 ;
        RECT 845.550 39.750 847.350 45.600 ;
        RECT 857.850 39.750 859.650 45.600 ;
        RECT 862.350 39.750 864.150 46.800 ;
        RECT 14.100 27.000 15.900 35.250 ;
        RECT 11.400 25.350 15.900 27.000 ;
        RECT 19.500 26.400 21.300 35.250 ;
        RECT 30.000 29.400 31.800 35.250 ;
        RECT 34.200 31.050 36.000 35.250 ;
        RECT 37.500 32.400 39.300 35.250 ;
        RECT 56.700 32.400 58.500 35.250 ;
        RECT 60.000 31.050 61.800 35.250 ;
        RECT 34.200 29.400 39.900 31.050 ;
        RECT 11.400 21.150 12.600 25.350 ;
        RECT 29.100 24.150 30.900 25.950 ;
        RECT 28.950 22.050 31.050 24.150 ;
        RECT 31.950 23.850 34.050 25.950 ;
        RECT 35.100 24.150 36.900 25.950 ;
        RECT 32.100 22.050 33.900 23.850 ;
        RECT 34.950 22.050 37.050 24.150 ;
        RECT 38.700 22.950 39.900 29.400 ;
        RECT 56.100 29.400 61.800 31.050 ;
        RECT 64.200 29.400 66.000 35.250 ;
        RECT 76.650 29.400 78.450 35.250 ;
        RECT 56.100 22.950 57.300 29.400 ;
        RECT 77.250 27.300 78.450 29.400 ;
        RECT 79.650 30.300 81.450 35.250 ;
        RECT 82.650 31.200 84.450 35.250 ;
        RECT 85.650 30.300 87.450 35.250 ;
        RECT 79.650 28.950 87.450 30.300 ;
        RECT 95.550 30.300 97.350 35.250 ;
        RECT 98.550 31.200 100.350 35.250 ;
        RECT 101.550 30.300 103.350 35.250 ;
        RECT 95.550 28.950 103.350 30.300 ;
        RECT 104.550 29.400 106.350 35.250 ;
        RECT 104.550 27.300 105.750 29.400 ;
        RECT 77.250 26.250 81.000 27.300 ;
        RECT 102.000 26.250 105.750 27.300 ;
        RECT 122.100 27.000 123.900 35.250 ;
        RECT 59.100 24.150 60.900 25.950 ;
        RECT 10.950 19.050 13.050 21.150 ;
        RECT 37.950 20.850 40.050 22.950 ;
        RECT 55.950 20.850 58.050 22.950 ;
        RECT 58.950 22.050 61.050 24.150 ;
        RECT 61.950 23.850 64.050 25.950 ;
        RECT 65.100 24.150 66.900 25.950 ;
        RECT 62.100 22.050 63.900 23.850 ;
        RECT 64.950 22.050 67.050 24.150 ;
        RECT 79.950 22.950 81.150 26.250 ;
        RECT 83.100 24.150 84.900 25.950 ;
        RECT 98.100 24.150 99.900 25.950 ;
        RECT 79.950 20.850 82.050 22.950 ;
        RECT 82.950 22.050 85.050 24.150 ;
        RECT 85.950 20.850 88.050 22.950 ;
        RECT 94.950 20.850 97.050 22.950 ;
        RECT 97.950 22.050 100.050 24.150 ;
        RECT 101.850 22.950 103.050 26.250 ;
        RECT 100.950 20.850 103.050 22.950 ;
        RECT 119.400 25.350 123.900 27.000 ;
        RECT 127.500 26.400 129.300 35.250 ;
        RECT 137.550 32.400 139.350 35.250 ;
        RECT 140.550 32.400 142.350 35.250 ;
        RECT 119.400 21.150 120.600 25.350 ;
        RECT 136.950 23.850 139.050 25.950 ;
        RECT 140.400 24.150 141.600 32.400 ;
        RECT 152.550 30.300 154.350 35.250 ;
        RECT 155.550 31.200 157.350 35.250 ;
        RECT 158.550 30.300 160.350 35.250 ;
        RECT 152.550 28.950 160.350 30.300 ;
        RECT 161.550 29.400 163.350 35.250 ;
        RECT 174.000 29.400 175.800 35.250 ;
        RECT 178.200 31.050 180.000 35.250 ;
        RECT 181.500 32.400 183.300 35.250 ;
        RECT 194.550 32.400 196.350 35.250 ;
        RECT 197.550 32.400 199.350 35.250 ;
        RECT 200.550 32.400 202.350 35.250 ;
        RECT 178.200 29.400 183.900 31.050 ;
        RECT 161.550 27.300 162.750 29.400 ;
        RECT 159.000 26.250 162.750 27.300 ;
        RECT 155.100 24.150 156.900 25.950 ;
        RECT 137.100 22.050 138.900 23.850 ;
        RECT 139.950 22.050 142.050 24.150 ;
        RECT 11.250 10.800 12.300 19.050 ;
        RECT 13.950 17.850 16.050 19.950 ;
        RECT 19.950 17.850 22.050 19.950 ;
        RECT 13.950 16.050 15.750 17.850 ;
        RECT 16.950 14.850 19.050 16.950 ;
        RECT 20.100 16.050 21.900 17.850 ;
        RECT 38.700 15.600 39.900 20.850 ;
        RECT 56.100 15.600 57.300 20.850 ;
        RECT 76.950 17.850 79.050 19.950 ;
        RECT 77.250 16.050 79.050 17.850 ;
        RECT 80.850 15.600 82.050 20.850 ;
        RECT 86.100 19.050 87.900 20.850 ;
        RECT 95.100 19.050 96.900 20.850 ;
        RECT 100.950 15.600 102.150 20.850 ;
        RECT 103.950 17.850 106.050 19.950 ;
        RECT 118.950 19.050 121.050 21.150 ;
        RECT 103.950 16.050 105.750 17.850 ;
        RECT 17.100 13.050 18.900 14.850 ;
        RECT 29.550 14.700 37.350 15.600 ;
        RECT 11.250 9.900 18.300 10.800 ;
        RECT 11.250 9.600 12.450 9.900 ;
        RECT 10.650 3.750 12.450 9.600 ;
        RECT 16.650 9.600 18.300 9.900 ;
        RECT 13.650 3.750 15.450 9.000 ;
        RECT 16.650 3.750 18.450 9.600 ;
        RECT 19.650 3.750 21.450 9.600 ;
        RECT 29.550 3.750 31.350 14.700 ;
        RECT 32.550 3.750 34.350 13.800 ;
        RECT 35.550 3.750 37.350 14.700 ;
        RECT 38.550 3.750 40.350 15.600 ;
        RECT 55.650 3.750 57.450 15.600 ;
        RECT 58.650 14.700 66.450 15.600 ;
        RECT 58.650 3.750 60.450 14.700 ;
        RECT 61.650 3.750 63.450 13.800 ;
        RECT 64.650 3.750 66.450 14.700 ;
        RECT 77.400 3.750 79.200 9.600 ;
        RECT 80.700 3.750 82.500 15.600 ;
        RECT 84.900 3.750 86.700 15.600 ;
        RECT 96.300 3.750 98.100 15.600 ;
        RECT 100.500 3.750 102.300 15.600 ;
        RECT 119.250 10.800 120.300 19.050 ;
        RECT 121.950 17.850 124.050 19.950 ;
        RECT 127.950 17.850 130.050 19.950 ;
        RECT 121.950 16.050 123.750 17.850 ;
        RECT 124.950 14.850 127.050 16.950 ;
        RECT 128.100 16.050 129.900 17.850 ;
        RECT 125.100 13.050 126.900 14.850 ;
        RECT 119.250 9.900 126.300 10.800 ;
        RECT 119.250 9.600 120.450 9.900 ;
        RECT 103.800 3.750 105.600 9.600 ;
        RECT 118.650 3.750 120.450 9.600 ;
        RECT 124.650 9.600 126.300 9.900 ;
        RECT 140.400 9.600 141.600 22.050 ;
        RECT 151.950 20.850 154.050 22.950 ;
        RECT 154.950 22.050 157.050 24.150 ;
        RECT 158.850 22.950 160.050 26.250 ;
        RECT 173.100 24.150 174.900 25.950 ;
        RECT 157.950 20.850 160.050 22.950 ;
        RECT 172.950 22.050 175.050 24.150 ;
        RECT 175.950 23.850 178.050 25.950 ;
        RECT 179.100 24.150 180.900 25.950 ;
        RECT 176.100 22.050 177.900 23.850 ;
        RECT 178.950 22.050 181.050 24.150 ;
        RECT 182.700 22.950 183.900 29.400 ;
        RECT 198.000 25.950 199.050 32.400 ;
        RECT 212.550 27.900 214.350 35.250 ;
        RECT 217.050 29.400 218.850 35.250 ;
        RECT 220.050 30.900 221.850 35.250 ;
        RECT 235.650 32.400 237.450 35.250 ;
        RECT 238.650 32.400 240.450 35.250 ;
        RECT 220.050 29.400 223.350 30.900 ;
        RECT 218.250 27.900 220.050 28.500 ;
        RECT 212.550 26.700 220.050 27.900 ;
        RECT 196.950 23.850 199.050 25.950 ;
        RECT 181.950 20.850 184.050 22.950 ;
        RECT 193.950 20.850 196.050 22.950 ;
        RECT 152.100 19.050 153.900 20.850 ;
        RECT 157.950 15.600 159.150 20.850 ;
        RECT 160.950 17.850 163.050 19.950 ;
        RECT 160.950 16.050 162.750 17.850 ;
        RECT 182.700 15.600 183.900 20.850 ;
        RECT 194.100 19.050 195.900 20.850 ;
        RECT 198.000 16.650 199.050 23.850 ;
        RECT 199.950 20.850 202.050 22.950 ;
        RECT 211.950 20.850 214.050 22.950 ;
        RECT 200.100 19.050 201.900 20.850 ;
        RECT 212.100 19.050 213.900 20.850 ;
        RECT 198.000 15.600 200.550 16.650 ;
        RECT 121.650 3.750 123.450 9.000 ;
        RECT 124.650 3.750 126.450 9.600 ;
        RECT 127.650 3.750 129.450 9.600 ;
        RECT 137.550 3.750 139.350 9.600 ;
        RECT 140.550 3.750 142.350 9.600 ;
        RECT 153.300 3.750 155.100 15.600 ;
        RECT 157.500 3.750 159.300 15.600 ;
        RECT 173.550 14.700 181.350 15.600 ;
        RECT 160.800 3.750 162.600 9.600 ;
        RECT 173.550 3.750 175.350 14.700 ;
        RECT 176.550 3.750 178.350 13.800 ;
        RECT 179.550 3.750 181.350 14.700 ;
        RECT 182.550 3.750 184.350 15.600 ;
        RECT 194.550 3.750 196.350 15.600 ;
        RECT 198.750 3.750 200.550 15.600 ;
        RECT 215.700 9.600 216.900 26.700 ;
        RECT 222.150 22.950 223.350 29.400 ;
        RECT 236.400 24.150 237.600 32.400 ;
        RECT 250.650 29.400 252.450 35.250 ;
        RECT 251.250 27.300 252.450 29.400 ;
        RECT 253.650 30.300 255.450 35.250 ;
        RECT 256.650 31.200 258.450 35.250 ;
        RECT 259.650 30.300 261.450 35.250 ;
        RECT 253.650 28.950 261.450 30.300 ;
        RECT 272.850 28.200 274.650 35.250 ;
        RECT 277.350 29.400 279.150 35.250 ;
        RECT 272.850 27.300 276.450 28.200 ;
        RECT 251.250 26.250 255.000 27.300 ;
        RECT 218.100 21.150 219.900 22.950 ;
        RECT 217.950 19.050 220.050 21.150 ;
        RECT 220.950 20.850 223.350 22.950 ;
        RECT 235.950 22.050 238.050 24.150 ;
        RECT 238.950 23.850 241.050 25.950 ;
        RECT 239.100 22.050 240.900 23.850 ;
        RECT 253.950 22.950 255.150 26.250 ;
        RECT 257.100 24.150 258.900 25.950 ;
        RECT 222.150 15.600 223.350 20.850 ;
        RECT 212.550 3.750 214.350 9.600 ;
        RECT 215.550 3.750 217.350 9.600 ;
        RECT 219.150 3.750 220.950 15.600 ;
        RECT 222.150 3.750 223.950 15.600 ;
        RECT 236.400 9.600 237.600 22.050 ;
        RECT 253.950 20.850 256.050 22.950 ;
        RECT 256.950 22.050 259.050 24.150 ;
        RECT 259.950 20.850 262.050 22.950 ;
        RECT 272.100 21.150 273.900 22.950 ;
        RECT 250.950 17.850 253.050 19.950 ;
        RECT 251.250 16.050 253.050 17.850 ;
        RECT 254.850 15.600 256.050 20.850 ;
        RECT 260.100 19.050 261.900 20.850 ;
        RECT 271.950 19.050 274.050 21.150 ;
        RECT 275.250 19.950 276.450 27.300 ;
        RECT 287.700 26.400 289.500 35.250 ;
        RECT 293.100 27.000 294.900 35.250 ;
        RECT 317.100 27.000 318.900 35.250 ;
        RECT 293.100 25.350 297.600 27.000 ;
        RECT 278.100 21.150 279.900 22.950 ;
        RECT 296.400 21.150 297.600 25.350 ;
        RECT 314.400 25.350 318.900 27.000 ;
        RECT 322.500 26.400 324.300 35.250 ;
        RECT 332.550 32.400 334.350 35.250 ;
        RECT 333.150 28.500 334.350 32.400 ;
        RECT 335.850 29.400 337.650 35.250 ;
        RECT 338.850 29.400 340.650 35.250 ;
        RECT 333.150 27.600 338.250 28.500 ;
        RECT 336.000 26.700 338.250 27.600 ;
        RECT 314.400 21.150 315.600 25.350 ;
        RECT 274.950 17.850 277.050 19.950 ;
        RECT 277.950 19.050 280.050 21.150 ;
        RECT 286.950 17.850 289.050 19.950 ;
        RECT 292.950 17.850 295.050 19.950 ;
        RECT 295.950 19.050 298.050 21.150 ;
        RECT 313.950 19.050 316.050 21.150 ;
        RECT 331.950 20.850 334.050 22.950 ;
        RECT 235.650 3.750 237.450 9.600 ;
        RECT 238.650 3.750 240.450 9.600 ;
        RECT 251.400 3.750 253.200 9.600 ;
        RECT 254.700 3.750 256.500 15.600 ;
        RECT 258.900 3.750 260.700 15.600 ;
        RECT 275.250 9.600 276.450 17.850 ;
        RECT 287.100 16.050 288.900 17.850 ;
        RECT 289.950 14.850 292.050 16.950 ;
        RECT 293.250 16.050 295.050 17.850 ;
        RECT 290.100 13.050 291.900 14.850 ;
        RECT 296.700 10.800 297.750 19.050 ;
        RECT 290.700 9.900 297.750 10.800 ;
        RECT 290.700 9.600 292.350 9.900 ;
        RECT 271.650 3.750 273.450 9.600 ;
        RECT 274.650 3.750 276.450 9.600 ;
        RECT 277.650 3.750 279.450 9.600 ;
        RECT 287.550 3.750 289.350 9.600 ;
        RECT 290.550 3.750 292.350 9.600 ;
        RECT 296.550 9.600 297.750 9.900 ;
        RECT 314.250 10.800 315.300 19.050 ;
        RECT 316.950 17.850 319.050 19.950 ;
        RECT 322.950 17.850 325.050 19.950 ;
        RECT 332.100 19.050 333.900 20.850 ;
        RECT 336.000 18.300 337.050 26.700 ;
        RECT 339.150 22.950 340.350 29.400 ;
        RECT 353.850 28.200 355.650 35.250 ;
        RECT 358.350 29.400 360.150 35.250 ;
        RECT 353.850 27.300 357.450 28.200 ;
        RECT 337.950 20.850 340.350 22.950 ;
        RECT 353.100 21.150 354.900 22.950 ;
        RECT 316.950 16.050 318.750 17.850 ;
        RECT 319.950 14.850 322.050 16.950 ;
        RECT 323.100 16.050 324.900 17.850 ;
        RECT 336.000 17.400 338.250 18.300 ;
        RECT 332.550 16.500 338.250 17.400 ;
        RECT 320.100 13.050 321.900 14.850 ;
        RECT 314.250 9.900 321.300 10.800 ;
        RECT 314.250 9.600 315.450 9.900 ;
        RECT 293.550 3.750 295.350 9.000 ;
        RECT 296.550 3.750 298.350 9.600 ;
        RECT 313.650 3.750 315.450 9.600 ;
        RECT 319.650 9.600 321.300 9.900 ;
        RECT 332.550 9.600 333.750 16.500 ;
        RECT 339.150 15.600 340.350 20.850 ;
        RECT 352.950 19.050 355.050 21.150 ;
        RECT 356.250 19.950 357.450 27.300 ;
        RECT 368.550 27.900 370.350 35.250 ;
        RECT 373.050 29.400 374.850 35.250 ;
        RECT 376.050 30.900 377.850 35.250 ;
        RECT 392.700 32.400 394.500 35.250 ;
        RECT 396.000 31.050 397.800 35.250 ;
        RECT 376.050 29.400 379.350 30.900 ;
        RECT 374.250 27.900 376.050 28.500 ;
        RECT 368.550 26.700 376.050 27.900 ;
        RECT 359.100 21.150 360.900 22.950 ;
        RECT 355.950 17.850 358.050 19.950 ;
        RECT 358.950 19.050 361.050 21.150 ;
        RECT 367.950 20.850 370.050 22.950 ;
        RECT 368.100 19.050 369.900 20.850 ;
        RECT 316.650 3.750 318.450 9.000 ;
        RECT 319.650 3.750 321.450 9.600 ;
        RECT 322.650 3.750 324.450 9.600 ;
        RECT 332.550 3.750 334.350 9.600 ;
        RECT 335.850 3.750 337.650 15.600 ;
        RECT 338.850 3.750 340.650 15.600 ;
        RECT 356.250 9.600 357.450 17.850 ;
        RECT 371.700 9.600 372.900 26.700 ;
        RECT 378.150 22.950 379.350 29.400 ;
        RECT 392.100 29.400 397.800 31.050 ;
        RECT 400.200 29.400 402.000 35.250 ;
        RECT 414.150 30.900 415.950 35.250 ;
        RECT 412.650 29.400 415.950 30.900 ;
        RECT 417.150 29.400 418.950 35.250 ;
        RECT 392.100 22.950 393.300 29.400 ;
        RECT 395.100 24.150 396.900 25.950 ;
        RECT 374.100 21.150 375.900 22.950 ;
        RECT 373.950 19.050 376.050 21.150 ;
        RECT 376.950 20.850 379.350 22.950 ;
        RECT 391.950 20.850 394.050 22.950 ;
        RECT 394.950 22.050 397.050 24.150 ;
        RECT 397.950 23.850 400.050 25.950 ;
        RECT 401.100 24.150 402.900 25.950 ;
        RECT 398.100 22.050 399.900 23.850 ;
        RECT 400.950 22.050 403.050 24.150 ;
        RECT 412.650 22.950 413.850 29.400 ;
        RECT 415.950 27.900 417.750 28.500 ;
        RECT 421.650 27.900 423.450 35.250 ;
        RECT 434.850 29.400 436.650 35.250 ;
        RECT 439.350 28.200 441.150 35.250 ;
        RECT 415.950 26.700 423.450 27.900 ;
        RECT 437.550 27.300 441.150 28.200 ;
        RECT 455.850 28.200 457.650 35.250 ;
        RECT 460.350 29.400 462.150 35.250 ;
        RECT 455.850 27.300 459.450 28.200 ;
        RECT 412.650 20.850 415.050 22.950 ;
        RECT 416.100 21.150 417.900 22.950 ;
        RECT 378.150 15.600 379.350 20.850 ;
        RECT 392.100 15.600 393.300 20.850 ;
        RECT 412.650 15.600 413.850 20.850 ;
        RECT 415.950 19.050 418.050 21.150 ;
        RECT 352.650 3.750 354.450 9.600 ;
        RECT 355.650 3.750 357.450 9.600 ;
        RECT 358.650 3.750 360.450 9.600 ;
        RECT 368.550 3.750 370.350 9.600 ;
        RECT 371.550 3.750 373.350 9.600 ;
        RECT 375.150 3.750 376.950 15.600 ;
        RECT 378.150 3.750 379.950 15.600 ;
        RECT 391.650 3.750 393.450 15.600 ;
        RECT 394.650 14.700 402.450 15.600 ;
        RECT 394.650 3.750 396.450 14.700 ;
        RECT 397.650 3.750 399.450 13.800 ;
        RECT 400.650 3.750 402.450 14.700 ;
        RECT 412.050 3.750 413.850 15.600 ;
        RECT 415.050 3.750 416.850 15.600 ;
        RECT 419.100 9.600 420.300 26.700 ;
        RECT 421.950 20.850 424.050 22.950 ;
        RECT 434.100 21.150 435.900 22.950 ;
        RECT 422.100 19.050 423.900 20.850 ;
        RECT 433.950 19.050 436.050 21.150 ;
        RECT 437.550 19.950 438.750 27.300 ;
        RECT 440.100 21.150 441.900 22.950 ;
        RECT 455.100 21.150 456.900 22.950 ;
        RECT 436.950 17.850 439.050 19.950 ;
        RECT 439.950 19.050 442.050 21.150 ;
        RECT 454.950 19.050 457.050 21.150 ;
        RECT 458.250 19.950 459.450 27.300 ;
        RECT 476.100 27.000 477.900 35.250 ;
        RECT 473.400 25.350 477.900 27.000 ;
        RECT 481.500 26.400 483.300 35.250 ;
        RECT 493.650 32.400 495.450 35.250 ;
        RECT 496.650 32.400 498.450 35.250 ;
        RECT 461.100 21.150 462.900 22.950 ;
        RECT 473.400 21.150 474.600 25.350 ;
        RECT 494.400 24.150 495.600 32.400 ;
        RECT 506.550 30.300 508.350 35.250 ;
        RECT 509.550 31.200 511.350 35.250 ;
        RECT 512.550 30.300 514.350 35.250 ;
        RECT 506.550 28.950 514.350 30.300 ;
        RECT 515.550 29.400 517.350 35.250 ;
        RECT 529.650 32.400 531.450 35.250 ;
        RECT 532.650 32.400 534.450 35.250 ;
        RECT 515.550 27.300 516.750 29.400 ;
        RECT 513.000 26.250 516.750 27.300 ;
        RECT 493.950 22.050 496.050 24.150 ;
        RECT 496.950 23.850 499.050 25.950 ;
        RECT 509.100 24.150 510.900 25.950 ;
        RECT 497.100 22.050 498.900 23.850 ;
        RECT 457.950 17.850 460.050 19.950 ;
        RECT 460.950 19.050 463.050 21.150 ;
        RECT 472.950 19.050 475.050 21.150 ;
        RECT 437.550 9.600 438.750 17.850 ;
        RECT 445.950 15.450 448.050 16.050 ;
        RECT 454.950 15.450 457.050 16.050 ;
        RECT 445.950 14.550 457.050 15.450 ;
        RECT 445.950 13.950 448.050 14.550 ;
        RECT 454.950 13.950 457.050 14.550 ;
        RECT 458.250 9.600 459.450 17.850 ;
        RECT 473.250 10.800 474.300 19.050 ;
        RECT 475.950 17.850 478.050 19.950 ;
        RECT 481.950 17.850 484.050 19.950 ;
        RECT 475.950 16.050 477.750 17.850 ;
        RECT 478.950 14.850 481.050 16.950 ;
        RECT 482.100 16.050 483.900 17.850 ;
        RECT 479.100 13.050 480.900 14.850 ;
        RECT 473.250 9.900 480.300 10.800 ;
        RECT 473.250 9.600 474.450 9.900 ;
        RECT 418.650 3.750 420.450 9.600 ;
        RECT 421.650 3.750 423.450 9.600 ;
        RECT 434.550 3.750 436.350 9.600 ;
        RECT 437.550 3.750 439.350 9.600 ;
        RECT 440.550 3.750 442.350 9.600 ;
        RECT 454.650 3.750 456.450 9.600 ;
        RECT 457.650 3.750 459.450 9.600 ;
        RECT 460.650 3.750 462.450 9.600 ;
        RECT 472.650 3.750 474.450 9.600 ;
        RECT 478.650 9.600 480.300 9.900 ;
        RECT 494.400 9.600 495.600 22.050 ;
        RECT 505.950 20.850 508.050 22.950 ;
        RECT 508.950 22.050 511.050 24.150 ;
        RECT 512.850 22.950 514.050 26.250 ;
        RECT 530.400 24.150 531.600 32.400 ;
        RECT 545.850 28.200 547.650 35.250 ;
        RECT 550.350 29.400 552.150 35.250 ;
        RECT 562.350 29.400 564.150 35.250 ;
        RECT 565.350 29.400 567.150 35.250 ;
        RECT 568.650 32.400 570.450 35.250 ;
        RECT 578.550 32.400 580.350 35.250 ;
        RECT 545.850 27.300 549.450 28.200 ;
        RECT 511.950 20.850 514.050 22.950 ;
        RECT 529.950 22.050 532.050 24.150 ;
        RECT 532.950 23.850 535.050 25.950 ;
        RECT 533.100 22.050 534.900 23.850 ;
        RECT 506.100 19.050 507.900 20.850 ;
        RECT 511.950 15.600 513.150 20.850 ;
        RECT 514.950 17.850 517.050 19.950 ;
        RECT 514.950 16.050 516.750 17.850 ;
        RECT 475.650 3.750 477.450 9.000 ;
        RECT 478.650 3.750 480.450 9.600 ;
        RECT 481.650 3.750 483.450 9.600 ;
        RECT 493.650 3.750 495.450 9.600 ;
        RECT 496.650 3.750 498.450 9.600 ;
        RECT 507.300 3.750 509.100 15.600 ;
        RECT 511.500 3.750 513.300 15.600 ;
        RECT 530.400 9.600 531.600 22.050 ;
        RECT 545.100 21.150 546.900 22.950 ;
        RECT 544.950 19.050 547.050 21.150 ;
        RECT 548.250 19.950 549.450 27.300 ;
        RECT 562.650 22.950 563.850 29.400 ;
        RECT 568.650 28.500 569.850 32.400 ;
        RECT 564.750 27.600 569.850 28.500 ;
        RECT 579.150 28.500 580.350 32.400 ;
        RECT 581.850 29.400 583.650 35.250 ;
        RECT 584.850 29.400 586.650 35.250 ;
        RECT 579.150 27.600 584.250 28.500 ;
        RECT 564.750 26.700 567.000 27.600 ;
        RECT 551.100 21.150 552.900 22.950 ;
        RECT 547.950 17.850 550.050 19.950 ;
        RECT 550.950 19.050 553.050 21.150 ;
        RECT 562.650 20.850 565.050 22.950 ;
        RECT 548.250 9.600 549.450 17.850 ;
        RECT 562.650 15.600 563.850 20.850 ;
        RECT 565.950 18.300 567.000 26.700 ;
        RECT 582.000 26.700 584.250 27.600 ;
        RECT 568.950 20.850 571.050 22.950 ;
        RECT 577.950 20.850 580.050 22.950 ;
        RECT 569.100 19.050 570.900 20.850 ;
        RECT 578.100 19.050 579.900 20.850 ;
        RECT 564.750 17.400 567.000 18.300 ;
        RECT 582.000 18.300 583.050 26.700 ;
        RECT 585.150 22.950 586.350 29.400 ;
        RECT 599.850 28.200 601.650 35.250 ;
        RECT 604.350 29.400 606.150 35.250 ;
        RECT 599.850 27.300 603.450 28.200 ;
        RECT 583.950 20.850 586.350 22.950 ;
        RECT 599.100 21.150 600.900 22.950 ;
        RECT 582.000 17.400 584.250 18.300 ;
        RECT 564.750 16.500 570.450 17.400 ;
        RECT 514.800 3.750 516.600 9.600 ;
        RECT 529.650 3.750 531.450 9.600 ;
        RECT 532.650 3.750 534.450 9.600 ;
        RECT 544.650 3.750 546.450 9.600 ;
        RECT 547.650 3.750 549.450 9.600 ;
        RECT 550.650 3.750 552.450 9.600 ;
        RECT 562.350 3.750 564.150 15.600 ;
        RECT 565.350 3.750 567.150 15.600 ;
        RECT 569.250 9.600 570.450 16.500 ;
        RECT 568.650 3.750 570.450 9.600 ;
        RECT 578.550 16.500 584.250 17.400 ;
        RECT 578.550 9.600 579.750 16.500 ;
        RECT 585.150 15.600 586.350 20.850 ;
        RECT 598.950 19.050 601.050 21.150 ;
        RECT 602.250 19.950 603.450 27.300 ;
        RECT 617.550 27.900 619.350 35.250 ;
        RECT 622.050 29.400 623.850 35.250 ;
        RECT 625.050 30.900 626.850 35.250 ;
        RECT 643.650 32.400 645.450 35.250 ;
        RECT 646.650 32.400 648.450 35.250 ;
        RECT 649.650 32.400 651.450 35.250 ;
        RECT 625.050 29.400 628.350 30.900 ;
        RECT 623.250 27.900 625.050 28.500 ;
        RECT 617.550 26.700 625.050 27.900 ;
        RECT 605.100 21.150 606.900 22.950 ;
        RECT 601.950 17.850 604.050 19.950 ;
        RECT 604.950 19.050 607.050 21.150 ;
        RECT 616.950 20.850 619.050 22.950 ;
        RECT 617.100 19.050 618.900 20.850 ;
        RECT 578.550 3.750 580.350 9.600 ;
        RECT 581.850 3.750 583.650 15.600 ;
        RECT 584.850 3.750 586.650 15.600 ;
        RECT 602.250 9.600 603.450 17.850 ;
        RECT 620.700 9.600 621.900 26.700 ;
        RECT 627.150 22.950 628.350 29.400 ;
        RECT 646.950 25.950 648.000 32.400 ;
        RECT 659.850 29.400 661.650 35.250 ;
        RECT 664.350 28.200 666.150 35.250 ;
        RECT 662.550 27.300 666.150 28.200 ;
        RECT 646.950 23.850 649.050 25.950 ;
        RECT 623.100 21.150 624.900 22.950 ;
        RECT 622.950 19.050 625.050 21.150 ;
        RECT 625.950 20.850 628.350 22.950 ;
        RECT 643.950 20.850 646.050 22.950 ;
        RECT 627.150 15.600 628.350 20.850 ;
        RECT 644.100 19.050 645.900 20.850 ;
        RECT 646.950 16.650 648.000 23.850 ;
        RECT 649.950 20.850 652.050 22.950 ;
        RECT 659.100 21.150 660.900 22.950 ;
        RECT 650.100 19.050 651.900 20.850 ;
        RECT 658.950 19.050 661.050 21.150 ;
        RECT 662.550 19.950 663.750 27.300 ;
        RECT 683.100 27.000 684.900 35.250 ;
        RECT 680.400 25.350 684.900 27.000 ;
        RECT 688.500 26.400 690.300 35.250 ;
        RECT 703.650 29.400 705.450 35.250 ;
        RECT 704.250 27.300 705.450 29.400 ;
        RECT 706.650 30.300 708.450 35.250 ;
        RECT 709.650 31.200 711.450 35.250 ;
        RECT 712.650 30.300 714.450 35.250 ;
        RECT 706.650 28.950 714.450 30.300 ;
        RECT 722.850 29.400 724.650 35.250 ;
        RECT 727.350 28.200 729.150 35.250 ;
        RECT 742.650 29.400 744.450 35.250 ;
        RECT 725.550 27.300 729.150 28.200 ;
        RECT 743.250 27.300 744.450 29.400 ;
        RECT 745.650 30.300 747.450 35.250 ;
        RECT 748.650 31.200 750.450 35.250 ;
        RECT 751.650 30.300 753.450 35.250 ;
        RECT 761.550 32.400 763.350 35.250 ;
        RECT 764.550 32.400 766.350 35.250 ;
        RECT 767.550 32.400 769.350 35.250 ;
        RECT 745.650 28.950 753.450 30.300 ;
        RECT 704.250 26.250 708.000 27.300 ;
        RECT 665.100 21.150 666.900 22.950 ;
        RECT 680.400 21.150 681.600 25.350 ;
        RECT 685.950 24.450 688.050 25.050 ;
        RECT 691.950 24.450 694.050 25.050 ;
        RECT 685.950 23.550 694.050 24.450 ;
        RECT 685.950 22.950 688.050 23.550 ;
        RECT 691.950 22.950 694.050 23.550 ;
        RECT 706.950 22.950 708.150 26.250 ;
        RECT 710.100 24.150 711.900 25.950 ;
        RECT 661.950 17.850 664.050 19.950 ;
        RECT 664.950 19.050 667.050 21.150 ;
        RECT 679.950 19.050 682.050 21.150 ;
        RECT 706.950 20.850 709.050 22.950 ;
        RECT 709.950 22.050 712.050 24.150 ;
        RECT 712.950 20.850 715.050 22.950 ;
        RECT 722.100 21.150 723.900 22.950 ;
        RECT 645.450 15.600 648.000 16.650 ;
        RECT 598.650 3.750 600.450 9.600 ;
        RECT 601.650 3.750 603.450 9.600 ;
        RECT 604.650 3.750 606.450 9.600 ;
        RECT 617.550 3.750 619.350 9.600 ;
        RECT 620.550 3.750 622.350 9.600 ;
        RECT 624.150 3.750 625.950 15.600 ;
        RECT 627.150 3.750 628.950 15.600 ;
        RECT 645.450 3.750 647.250 15.600 ;
        RECT 649.650 3.750 651.450 15.600 ;
        RECT 662.550 9.600 663.750 17.850 ;
        RECT 680.250 10.800 681.300 19.050 ;
        RECT 682.950 17.850 685.050 19.950 ;
        RECT 688.950 17.850 691.050 19.950 ;
        RECT 703.950 17.850 706.050 19.950 ;
        RECT 682.950 16.050 684.750 17.850 ;
        RECT 685.950 14.850 688.050 16.950 ;
        RECT 689.100 16.050 690.900 17.850 ;
        RECT 704.250 16.050 706.050 17.850 ;
        RECT 707.850 15.600 709.050 20.850 ;
        RECT 713.100 19.050 714.900 20.850 ;
        RECT 721.950 19.050 724.050 21.150 ;
        RECT 725.550 19.950 726.750 27.300 ;
        RECT 743.250 26.250 747.000 27.300 ;
        RECT 745.950 22.950 747.150 26.250 ;
        RECT 765.000 25.950 766.050 32.400 ;
        RECT 782.850 28.200 784.650 35.250 ;
        RECT 787.350 29.400 789.150 35.250 ;
        RECT 797.550 31.200 799.350 34.200 ;
        RECT 800.550 31.200 802.350 35.250 ;
        RECT 782.850 27.300 786.450 28.200 ;
        RECT 749.100 24.150 750.900 25.950 ;
        RECT 728.100 21.150 729.900 22.950 ;
        RECT 724.950 17.850 727.050 19.950 ;
        RECT 727.950 19.050 730.050 21.150 ;
        RECT 745.950 20.850 748.050 22.950 ;
        RECT 748.950 22.050 751.050 24.150 ;
        RECT 763.950 23.850 766.050 25.950 ;
        RECT 751.950 20.850 754.050 22.950 ;
        RECT 760.950 20.850 763.050 22.950 ;
        RECT 742.950 17.850 745.050 19.950 ;
        RECT 686.100 13.050 687.900 14.850 ;
        RECT 680.250 9.900 687.300 10.800 ;
        RECT 680.250 9.600 681.450 9.900 ;
        RECT 659.550 3.750 661.350 9.600 ;
        RECT 662.550 3.750 664.350 9.600 ;
        RECT 665.550 3.750 667.350 9.600 ;
        RECT 679.650 3.750 681.450 9.600 ;
        RECT 685.650 9.600 687.300 9.900 ;
        RECT 682.650 3.750 684.450 9.000 ;
        RECT 685.650 3.750 687.450 9.600 ;
        RECT 688.650 3.750 690.450 9.600 ;
        RECT 704.400 3.750 706.200 9.600 ;
        RECT 707.700 3.750 709.500 15.600 ;
        RECT 711.900 3.750 713.700 15.600 ;
        RECT 725.550 9.600 726.750 17.850 ;
        RECT 743.250 16.050 745.050 17.850 ;
        RECT 746.850 15.600 748.050 20.850 ;
        RECT 752.100 19.050 753.900 20.850 ;
        RECT 761.100 19.050 762.900 20.850 ;
        RECT 765.000 16.650 766.050 23.850 ;
        RECT 766.950 20.850 769.050 22.950 ;
        RECT 782.100 21.150 783.900 22.950 ;
        RECT 767.100 19.050 768.900 20.850 ;
        RECT 781.950 19.050 784.050 21.150 ;
        RECT 785.250 19.950 786.450 27.300 ;
        RECT 798.300 27.900 799.350 31.200 ;
        RECT 805.050 29.700 806.850 34.200 ;
        RECT 805.050 28.800 807.150 29.700 ;
        RECT 798.300 27.000 804.600 27.900 ;
        RECT 797.250 24.150 799.050 25.950 ;
        RECT 788.100 21.150 789.900 22.950 ;
        RECT 796.950 22.050 799.050 24.150 ;
        RECT 784.950 17.850 787.050 19.950 ;
        RECT 787.950 19.050 790.050 21.150 ;
        RECT 799.950 20.850 802.050 22.950 ;
        RECT 800.250 19.050 802.050 20.850 ;
        RECT 803.250 21.300 804.600 27.000 ;
        RECT 806.250 24.150 807.150 28.800 ;
        RECT 809.550 28.200 811.350 35.250 ;
        RECT 821.550 32.400 823.350 35.250 ;
        RECT 824.550 32.400 826.350 35.250 ;
        RECT 838.650 32.400 840.450 35.250 ;
        RECT 841.650 32.400 843.450 35.250 ;
        RECT 805.950 22.050 808.050 24.150 ;
        RECT 820.950 23.850 823.050 25.950 ;
        RECT 824.400 24.150 825.600 32.400 ;
        RECT 839.400 24.150 840.600 32.400 ;
        RECT 851.850 29.400 853.650 35.250 ;
        RECT 856.350 28.200 858.150 35.250 ;
        RECT 854.550 27.300 858.150 28.200 ;
        RECT 803.250 19.500 805.050 21.300 ;
        RECT 765.000 15.600 767.550 16.650 ;
        RECT 722.550 3.750 724.350 9.600 ;
        RECT 725.550 3.750 727.350 9.600 ;
        RECT 728.550 3.750 730.350 9.600 ;
        RECT 743.400 3.750 745.200 9.600 ;
        RECT 746.700 3.750 748.500 15.600 ;
        RECT 750.900 3.750 752.700 15.600 ;
        RECT 761.550 3.750 763.350 15.600 ;
        RECT 765.750 3.750 767.550 15.600 ;
        RECT 785.250 9.600 786.450 17.850 ;
        RECT 803.250 16.800 804.600 19.500 ;
        RECT 798.450 15.900 804.600 16.800 ;
        RECT 798.450 10.800 799.350 15.900 ;
        RECT 806.250 15.000 807.150 22.050 ;
        RECT 808.950 20.850 811.050 22.950 ;
        RECT 821.100 22.050 822.900 23.850 ;
        RECT 823.950 22.050 826.050 24.150 ;
        RECT 838.950 22.050 841.050 24.150 ;
        RECT 841.950 23.850 844.050 25.950 ;
        RECT 842.100 22.050 843.900 23.850 ;
        RECT 809.100 19.050 810.900 20.850 ;
        RECT 805.050 14.100 807.150 15.000 ;
        RECT 781.650 3.750 783.450 9.600 ;
        RECT 784.650 3.750 786.450 9.600 ;
        RECT 787.650 3.750 789.450 9.600 ;
        RECT 797.550 4.800 799.350 10.800 ;
        RECT 800.550 3.750 802.350 10.800 ;
        RECT 805.050 4.800 806.850 14.100 ;
        RECT 809.550 3.750 811.350 15.600 ;
        RECT 824.400 9.600 825.600 22.050 ;
        RECT 839.400 9.600 840.600 22.050 ;
        RECT 851.100 21.150 852.900 22.950 ;
        RECT 850.950 19.050 853.050 21.150 ;
        RECT 854.550 19.950 855.750 27.300 ;
        RECT 857.100 21.150 858.900 22.950 ;
        RECT 853.950 17.850 856.050 19.950 ;
        RECT 856.950 19.050 859.050 21.150 ;
        RECT 854.550 9.600 855.750 17.850 ;
        RECT 821.550 3.750 823.350 9.600 ;
        RECT 824.550 3.750 826.350 9.600 ;
        RECT 838.650 3.750 840.450 9.600 ;
        RECT 841.650 3.750 843.450 9.600 ;
        RECT 851.550 3.750 853.350 9.600 ;
        RECT 854.550 3.750 856.350 9.600 ;
        RECT 857.550 3.750 859.350 9.600 ;
      LAYER metal2 ;
        RECT 625.950 855.300 628.050 857.400 ;
        RECT 76.950 851.250 79.050 852.150 ;
        RECT 229.950 851.250 232.050 852.150 ;
        RECT 274.950 851.250 277.050 852.150 ;
        RECT 391.950 851.250 394.050 852.150 ;
        RECT 412.950 851.250 415.050 852.150 ;
        RECT 529.950 851.250 532.050 852.150 ;
        RECT 626.550 851.700 627.750 855.300 ;
        RECT 646.950 854.400 649.050 856.500 ;
        RECT 10.950 848.250 13.050 849.150 ;
        RECT 37.950 848.250 40.050 849.150 ;
        RECT 67.950 847.950 70.050 850.050 ;
        RECT 73.950 848.250 75.750 849.150 ;
        RECT 76.950 847.950 79.050 850.050 ;
        RECT 82.950 849.450 85.050 850.050 ;
        RECT 118.950 849.450 121.050 850.050 ;
        RECT 80.250 848.250 81.750 849.150 ;
        RECT 82.950 848.400 87.450 849.450 ;
        RECT 82.950 847.950 85.050 848.400 ;
        RECT 10.950 844.950 13.050 847.050 ;
        RECT 14.250 845.250 15.750 846.150 ;
        RECT 16.950 844.950 19.050 847.050 ;
        RECT 20.250 845.250 22.050 846.150 ;
        RECT 28.950 845.250 30.750 846.150 ;
        RECT 31.950 844.950 34.050 847.050 ;
        RECT 35.250 845.250 36.750 846.150 ;
        RECT 37.950 844.950 40.050 847.050 ;
        RECT 55.950 845.250 57.750 846.150 ;
        RECT 58.950 844.950 61.050 847.050 ;
        RECT 64.950 846.450 67.050 847.050 ;
        RECT 68.400 846.450 69.450 847.950 ;
        RECT 64.950 845.400 69.450 846.450 ;
        RECT 64.950 844.950 67.050 845.400 ;
        RECT 11.400 820.050 12.450 844.950 ;
        RECT 13.950 841.950 16.050 844.050 ;
        RECT 17.250 842.850 18.750 843.750 ;
        RECT 19.950 841.950 22.050 844.050 ;
        RECT 28.950 841.950 31.050 844.050 ;
        RECT 32.250 842.850 33.750 843.750 ;
        RECT 34.950 841.950 37.050 844.050 ;
        RECT 14.400 823.050 15.450 841.950 ;
        RECT 13.950 820.950 16.050 823.050 ;
        RECT 10.950 817.950 13.050 820.050 ;
        RECT 19.950 817.950 22.050 820.050 ;
        RECT 20.400 817.050 21.450 817.950 ;
        RECT 13.950 814.950 16.050 817.050 ;
        RECT 17.250 815.250 18.750 816.150 ;
        RECT 19.950 814.950 22.050 817.050 ;
        RECT 29.400 814.050 30.450 841.950 ;
        RECT 35.400 816.450 36.450 841.950 ;
        RECT 38.400 832.050 39.450 844.950 ;
        RECT 55.950 841.950 58.050 844.050 ;
        RECT 59.250 842.850 61.050 843.750 ;
        RECT 61.950 842.250 64.050 843.150 ;
        RECT 64.950 842.850 67.050 843.750 ;
        RECT 61.950 838.950 64.050 841.050 ;
        RECT 37.950 829.950 40.050 832.050 ;
        RECT 58.950 820.950 61.050 823.050 ;
        RECT 35.400 815.400 39.450 816.450 ;
        RECT 38.400 814.050 39.450 815.400 ;
        RECT 40.950 814.950 43.050 817.050 ;
        RECT 10.950 813.450 13.050 814.050 ;
        RECT 8.400 812.400 13.050 813.450 ;
        RECT 14.250 812.850 15.750 813.750 ;
        RECT 8.400 808.050 9.450 812.400 ;
        RECT 10.950 811.950 13.050 812.400 ;
        RECT 16.950 811.950 19.050 814.050 ;
        RECT 20.250 812.850 22.050 813.750 ;
        RECT 28.950 811.950 31.050 814.050 ;
        RECT 34.950 812.250 36.750 813.150 ;
        RECT 37.950 811.950 40.050 814.050 ;
        RECT 10.950 809.850 13.050 810.750 ;
        RECT 13.950 808.950 16.050 811.050 ;
        RECT 7.950 805.950 10.050 808.050 ;
        RECT 10.950 805.950 13.050 808.050 ;
        RECT 7.950 796.950 10.050 799.050 ;
        RECT 4.950 751.950 7.050 754.050 ;
        RECT 5.400 718.050 6.450 751.950 ;
        RECT 4.950 715.950 7.050 718.050 ;
        RECT 4.950 700.950 7.050 703.050 ;
        RECT 5.400 628.050 6.450 700.950 ;
        RECT 8.400 676.050 9.450 796.950 ;
        RECT 11.400 778.050 12.450 805.950 ;
        RECT 14.400 799.050 15.450 808.950 ;
        RECT 13.950 796.950 16.050 799.050 ;
        RECT 25.950 784.950 28.050 787.050 ;
        RECT 22.950 781.950 25.050 784.050 ;
        RECT 16.950 779.250 19.050 780.150 ;
        RECT 23.400 778.050 24.450 781.950 ;
        RECT 10.950 775.950 13.050 778.050 ;
        RECT 14.250 776.250 15.750 777.150 ;
        RECT 16.950 775.950 19.050 778.050 ;
        RECT 20.250 776.250 22.050 777.150 ;
        RECT 22.950 775.950 25.050 778.050 ;
        RECT 17.400 775.050 18.450 775.950 ;
        RECT 10.950 773.850 12.750 774.750 ;
        RECT 13.950 772.950 16.050 775.050 ;
        RECT 16.950 772.950 19.050 775.050 ;
        RECT 19.950 772.950 22.050 775.050 ;
        RECT 10.950 745.950 13.050 748.050 ;
        RECT 17.400 747.450 18.450 772.950 ;
        RECT 20.400 769.050 21.450 772.950 ;
        RECT 19.950 766.950 22.050 769.050 ;
        RECT 14.400 746.400 18.450 747.450 ;
        RECT 11.400 742.050 12.450 745.950 ;
        RECT 14.400 745.050 15.450 746.400 ;
        RECT 13.950 742.950 16.050 745.050 ;
        RECT 19.950 744.450 22.050 745.050 ;
        RECT 17.250 743.250 18.750 744.150 ;
        RECT 19.950 743.400 24.450 744.450 ;
        RECT 19.950 742.950 22.050 743.400 ;
        RECT 10.950 739.950 13.050 742.050 ;
        RECT 14.250 740.850 15.750 741.750 ;
        RECT 16.950 739.950 19.050 742.050 ;
        RECT 20.250 740.850 22.050 741.750 ;
        RECT 10.950 737.850 13.050 738.750 ;
        RECT 17.400 733.050 18.450 739.950 ;
        RECT 16.950 730.950 19.050 733.050 ;
        RECT 19.950 724.950 22.050 727.050 ;
        RECT 16.950 715.950 19.050 718.050 ;
        RECT 13.950 712.950 16.050 715.050 ;
        RECT 14.400 703.050 15.450 712.950 ;
        RECT 17.400 706.050 18.450 715.950 ;
        RECT 16.950 703.950 19.050 706.050 ;
        RECT 20.400 703.050 21.450 724.950 ;
        RECT 23.400 715.050 24.450 743.400 ;
        RECT 26.400 720.450 27.450 784.950 ;
        RECT 29.400 778.050 30.450 811.950 ;
        RECT 41.400 811.050 42.450 814.950 ;
        RECT 59.400 814.050 60.450 820.950 ;
        RECT 43.950 813.450 46.050 814.050 ;
        RECT 43.950 812.400 48.450 813.450 ;
        RECT 43.950 811.950 46.050 812.400 ;
        RECT 34.950 808.950 37.050 811.050 ;
        RECT 38.250 809.850 39.750 810.750 ;
        RECT 40.950 808.950 43.050 811.050 ;
        RECT 44.250 809.850 46.050 810.750 ;
        RECT 35.400 787.050 36.450 808.950 ;
        RECT 40.950 806.850 43.050 807.750 ;
        RECT 34.950 784.950 37.050 787.050 ;
        RECT 34.950 781.950 37.050 784.050 ;
        RECT 28.950 775.950 31.050 778.050 ;
        RECT 35.400 775.050 36.450 781.950 ;
        RECT 47.400 778.050 48.450 812.400 ;
        RECT 55.950 812.250 57.750 813.150 ;
        RECT 58.950 811.950 61.050 814.050 ;
        RECT 64.950 811.950 67.050 814.050 ;
        RECT 52.950 808.950 55.050 811.050 ;
        RECT 55.950 808.950 58.050 811.050 ;
        RECT 59.250 809.850 60.750 810.750 ;
        RECT 61.950 808.950 64.050 811.050 ;
        RECT 65.250 809.850 67.050 810.750 ;
        RECT 40.950 775.950 43.050 778.050 ;
        RECT 46.950 775.950 49.050 778.050 ;
        RECT 28.950 772.950 31.050 775.050 ;
        RECT 34.950 772.950 37.050 775.050 ;
        RECT 38.250 773.250 40.050 774.150 ;
        RECT 28.950 770.850 31.050 771.750 ;
        RECT 31.950 770.250 34.050 771.150 ;
        RECT 34.950 770.850 36.750 771.750 ;
        RECT 37.950 771.450 40.050 772.050 ;
        RECT 41.400 771.450 42.450 775.950 ;
        RECT 37.950 770.400 42.450 771.450 ;
        RECT 37.950 769.950 40.050 770.400 ;
        RECT 31.950 766.950 34.050 769.050 ;
        RECT 47.400 768.450 48.450 775.950 ;
        RECT 53.400 775.050 54.450 808.950 ;
        RECT 52.950 772.950 55.050 775.050 ;
        RECT 49.950 770.250 52.050 771.150 ;
        RECT 52.950 770.850 55.050 771.750 ;
        RECT 49.950 768.450 52.050 769.050 ;
        RECT 47.400 767.400 52.050 768.450 ;
        RECT 49.950 766.950 52.050 767.400 ;
        RECT 32.400 745.050 33.450 766.950 ;
        RECT 56.400 754.050 57.450 808.950 ;
        RECT 61.950 806.850 64.050 807.750 ;
        RECT 68.400 805.050 69.450 845.400 ;
        RECT 73.950 844.950 76.050 847.050 ;
        RECT 79.950 844.950 82.050 847.050 ;
        RECT 83.250 845.850 85.050 846.750 ;
        RECT 74.400 841.050 75.450 844.950 ;
        RECT 80.400 841.050 81.450 844.950 ;
        RECT 73.950 838.950 76.050 841.050 ;
        RECT 79.950 838.950 82.050 841.050 ;
        RECT 74.400 816.450 75.450 838.950 ;
        RECT 86.400 823.050 87.450 848.400 ;
        RECT 97.950 848.250 100.050 849.150 ;
        RECT 116.400 848.400 121.050 849.450 ;
        RECT 97.950 844.950 100.050 847.050 ;
        RECT 101.250 845.250 102.750 846.150 ;
        RECT 103.950 844.950 106.050 847.050 ;
        RECT 107.250 845.250 109.050 846.150 ;
        RECT 109.950 844.950 112.050 847.050 ;
        RECT 98.400 835.050 99.450 844.950 ;
        RECT 100.950 841.950 103.050 844.050 ;
        RECT 104.250 842.850 105.750 843.750 ;
        RECT 106.950 841.950 109.050 844.050 ;
        RECT 97.950 832.950 100.050 835.050 ;
        RECT 97.950 829.950 100.050 832.050 ;
        RECT 79.950 820.950 82.050 823.050 ;
        RECT 85.950 820.950 88.050 823.050 ;
        RECT 71.400 815.400 75.450 816.450 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 67.950 802.950 70.050 805.050 ;
        RECT 58.950 799.950 61.050 802.050 ;
        RECT 55.950 751.950 58.050 754.050 ;
        RECT 55.950 745.950 58.050 748.050 ;
        RECT 31.950 742.950 34.050 745.050 ;
        RECT 56.400 742.050 57.450 745.950 ;
        RECT 59.400 745.050 60.450 799.950 ;
        RECT 62.400 772.050 63.450 802.950 ;
        RECT 71.400 802.050 72.450 815.400 ;
        RECT 80.400 814.050 81.450 820.950 ;
        RECT 85.950 817.950 88.050 820.050 ;
        RECT 86.400 814.050 87.450 817.950 ;
        RECT 91.950 814.950 94.050 817.050 ;
        RECT 73.950 811.950 76.050 814.050 ;
        RECT 76.950 812.250 78.750 813.150 ;
        RECT 79.950 811.950 82.050 814.050 ;
        RECT 85.950 811.950 88.050 814.050 ;
        RECT 88.950 811.950 91.050 814.050 ;
        RECT 74.400 805.050 75.450 811.950 ;
        RECT 76.950 808.950 79.050 811.050 ;
        RECT 80.250 809.850 81.750 810.750 ;
        RECT 82.950 808.950 85.050 811.050 ;
        RECT 86.250 809.850 88.050 810.750 ;
        RECT 82.950 806.850 85.050 807.750 ;
        RECT 73.950 802.950 76.050 805.050 ;
        RECT 70.950 799.950 73.050 802.050 ;
        RECT 73.950 779.250 76.050 780.150 ;
        RECT 79.950 778.950 82.050 781.050 ;
        RECT 67.950 775.950 70.050 778.050 ;
        RECT 71.250 776.250 72.750 777.150 ;
        RECT 73.950 775.950 76.050 778.050 ;
        RECT 77.250 776.250 79.050 777.150 ;
        RECT 64.950 772.950 67.050 775.050 ;
        RECT 67.950 773.850 69.750 774.750 ;
        RECT 70.950 772.950 73.050 775.050 ;
        RECT 61.950 769.950 64.050 772.050 ;
        RECT 61.950 745.950 64.050 748.050 ;
        RECT 58.950 742.950 61.050 745.050 ;
        RECT 28.950 739.950 31.050 742.050 ;
        RECT 31.950 740.250 33.750 741.150 ;
        RECT 34.950 739.950 37.050 742.050 ;
        RECT 40.950 741.450 43.050 742.050 ;
        RECT 43.950 741.450 46.050 742.050 ;
        RECT 40.950 740.400 46.050 741.450 ;
        RECT 40.950 739.950 43.050 740.400 ;
        RECT 43.950 739.950 46.050 740.400 ;
        RECT 49.950 739.950 52.050 742.050 ;
        RECT 55.950 739.950 58.050 742.050 ;
        RECT 59.250 740.250 61.050 741.150 ;
        RECT 29.400 727.050 30.450 739.950 ;
        RECT 31.950 736.950 34.050 739.050 ;
        RECT 35.250 737.850 36.750 738.750 ;
        RECT 37.950 736.950 40.050 739.050 ;
        RECT 41.250 737.850 43.050 738.750 ;
        RECT 44.400 736.050 45.450 739.950 ;
        RECT 46.950 736.950 49.050 739.050 ;
        RECT 49.950 737.850 51.750 738.750 ;
        RECT 52.950 736.950 55.050 739.050 ;
        RECT 56.250 737.850 57.750 738.750 ;
        RECT 58.950 736.950 61.050 739.050 ;
        RECT 31.950 733.950 34.050 736.050 ;
        RECT 37.950 734.850 40.050 735.750 ;
        RECT 43.950 733.950 46.050 736.050 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 26.400 719.400 30.450 720.450 ;
        RECT 25.950 715.950 28.050 718.050 ;
        RECT 22.950 712.950 25.050 715.050 ;
        RECT 22.950 706.950 25.050 709.050 ;
        RECT 10.950 701.250 12.750 702.150 ;
        RECT 13.950 700.950 16.050 703.050 ;
        RECT 19.950 700.950 22.050 703.050 ;
        RECT 10.950 697.950 13.050 700.050 ;
        RECT 14.250 698.850 16.050 699.750 ;
        RECT 16.950 698.250 19.050 699.150 ;
        RECT 19.950 698.850 22.050 699.750 ;
        RECT 7.950 673.950 10.050 676.050 ;
        RECT 11.400 672.450 12.450 697.950 ;
        RECT 16.950 694.950 19.050 697.050 ;
        RECT 19.950 685.950 22.050 688.050 ;
        RECT 13.950 673.950 16.050 676.050 ;
        RECT 14.400 673.050 15.450 673.950 ;
        RECT 20.400 673.050 21.450 685.950 ;
        RECT 23.400 679.050 24.450 706.950 ;
        RECT 22.950 676.950 25.050 679.050 ;
        RECT 22.950 673.950 25.050 676.050 ;
        RECT 8.400 671.400 12.450 672.450 ;
        RECT 4.950 625.950 7.050 628.050 ;
        RECT 8.400 619.050 9.450 671.400 ;
        RECT 13.950 670.950 16.050 673.050 ;
        RECT 17.250 671.250 18.750 672.150 ;
        RECT 19.950 670.950 22.050 673.050 ;
        RECT 10.950 667.950 13.050 670.050 ;
        RECT 14.250 668.850 15.750 669.750 ;
        RECT 16.950 667.950 19.050 670.050 ;
        RECT 20.250 668.850 22.050 669.750 ;
        RECT 10.950 665.850 13.050 666.750 ;
        RECT 10.950 661.950 13.050 664.050 ;
        RECT 23.400 663.450 24.450 673.950 ;
        RECT 26.400 667.050 27.450 715.950 ;
        RECT 29.400 709.050 30.450 719.400 ;
        RECT 28.950 706.950 31.050 709.050 ;
        RECT 32.400 706.050 33.450 733.950 ;
        RECT 43.950 730.950 46.050 733.050 ;
        RECT 37.950 707.250 40.050 708.150 ;
        RECT 31.950 705.450 34.050 706.050 ;
        RECT 29.400 704.400 34.050 705.450 ;
        RECT 29.400 697.050 30.450 704.400 ;
        RECT 31.950 703.950 34.050 704.400 ;
        RECT 35.250 704.250 36.750 705.150 ;
        RECT 37.950 703.950 40.050 706.050 ;
        RECT 41.250 704.250 43.050 705.150 ;
        RECT 31.950 701.850 33.750 702.750 ;
        RECT 34.950 700.950 37.050 703.050 ;
        RECT 35.400 697.050 36.450 700.950 ;
        RECT 28.950 694.950 31.050 697.050 ;
        RECT 34.950 694.950 37.050 697.050 ;
        RECT 38.400 694.050 39.450 703.950 ;
        RECT 40.950 700.950 43.050 703.050 ;
        RECT 40.950 697.950 43.050 700.050 ;
        RECT 37.950 691.950 40.050 694.050 ;
        RECT 34.950 682.950 37.050 685.050 ;
        RECT 28.950 676.950 31.050 679.050 ;
        RECT 25.950 664.950 28.050 667.050 ;
        RECT 23.400 662.400 27.450 663.450 ;
        RECT 7.950 616.950 10.050 619.050 ;
        RECT 7.950 613.950 10.050 616.050 ;
        RECT 8.400 597.450 9.450 613.950 ;
        RECT 11.400 604.050 12.450 661.950 ;
        RECT 13.950 632.250 16.050 633.150 ;
        RECT 13.950 628.950 16.050 631.050 ;
        RECT 17.250 629.250 18.750 630.150 ;
        RECT 19.950 628.950 22.050 631.050 ;
        RECT 23.250 629.250 25.050 630.150 ;
        RECT 14.400 616.050 15.450 628.950 ;
        RECT 26.400 628.050 27.450 662.400 ;
        RECT 16.950 625.950 19.050 628.050 ;
        RECT 20.250 626.850 21.750 627.750 ;
        RECT 22.950 625.950 25.050 628.050 ;
        RECT 25.950 625.950 28.050 628.050 ;
        RECT 19.950 622.950 22.050 625.050 ;
        RECT 16.950 616.950 19.050 619.050 ;
        RECT 13.950 613.950 16.050 616.050 ;
        RECT 10.950 601.950 13.050 604.050 ;
        RECT 13.950 601.950 16.050 604.050 ;
        RECT 10.950 599.250 13.050 600.150 ;
        RECT 13.950 599.850 16.050 600.750 ;
        RECT 10.950 597.450 13.050 598.050 ;
        RECT 8.400 596.400 13.050 597.450 ;
        RECT 10.950 595.950 13.050 596.400 ;
        RECT 13.950 595.950 16.050 598.050 ;
        RECT 14.400 592.050 15.450 595.950 ;
        RECT 13.950 589.950 16.050 592.050 ;
        RECT 13.950 586.950 16.050 589.050 ;
        RECT 7.950 565.950 10.050 568.050 ;
        RECT 4.950 235.950 7.050 238.050 ;
        RECT 5.400 172.050 6.450 235.950 ;
        RECT 4.950 169.950 7.050 172.050 ;
        RECT 5.400 91.050 6.450 169.950 ;
        RECT 8.400 94.050 9.450 565.950 ;
        RECT 14.400 564.450 15.450 586.950 ;
        RECT 17.400 568.050 18.450 616.950 ;
        RECT 20.400 595.050 21.450 622.950 ;
        RECT 23.400 613.050 24.450 625.950 ;
        RECT 25.950 622.950 28.050 625.050 ;
        RECT 22.950 610.950 25.050 613.050 ;
        RECT 22.950 604.950 25.050 607.050 ;
        RECT 23.400 604.050 24.450 604.950 ;
        RECT 26.400 604.050 27.450 622.950 ;
        RECT 29.400 607.050 30.450 676.950 ;
        RECT 35.400 670.050 36.450 682.950 ;
        RECT 37.950 673.950 40.050 676.050 ;
        RECT 31.950 668.250 33.750 669.150 ;
        RECT 34.950 667.950 37.050 670.050 ;
        RECT 38.400 667.050 39.450 673.950 ;
        RECT 41.400 673.050 42.450 697.950 ;
        RECT 44.400 673.050 45.450 730.950 ;
        RECT 47.400 718.050 48.450 736.950 ;
        RECT 52.950 734.850 55.050 735.750 ;
        RECT 46.950 715.950 49.050 718.050 ;
        RECT 62.400 717.450 63.450 745.950 ;
        RECT 59.400 716.400 63.450 717.450 ;
        RECT 55.950 706.950 58.050 709.050 ;
        RECT 56.400 703.050 57.450 706.950 ;
        RECT 59.400 706.050 60.450 716.400 ;
        RECT 61.950 712.950 64.050 715.050 ;
        RECT 58.950 703.950 61.050 706.050 ;
        RECT 49.950 702.450 52.050 703.050 ;
        RECT 47.400 701.400 52.050 702.450 ;
        RECT 47.400 697.050 48.450 701.400 ;
        RECT 49.950 700.950 52.050 701.400 ;
        RECT 55.950 700.950 58.050 703.050 ;
        RECT 59.250 701.250 61.050 702.150 ;
        RECT 49.950 698.850 52.050 699.750 ;
        RECT 52.950 698.250 55.050 699.150 ;
        RECT 55.950 698.850 57.750 699.750 ;
        RECT 58.950 699.450 61.050 700.050 ;
        RECT 62.400 699.450 63.450 712.950 ;
        RECT 58.950 698.400 63.450 699.450 ;
        RECT 58.950 697.950 61.050 698.400 ;
        RECT 46.950 694.950 49.050 697.050 ;
        RECT 52.950 694.950 55.050 697.050 ;
        RECT 53.400 694.050 54.450 694.950 ;
        RECT 52.950 691.950 55.050 694.050 ;
        RECT 61.950 682.950 64.050 685.050 ;
        RECT 52.950 673.950 55.050 676.050 ;
        RECT 40.950 670.950 43.050 673.050 ;
        RECT 43.950 670.950 46.050 673.050 ;
        RECT 46.950 670.950 49.050 673.050 ;
        RECT 49.950 671.250 52.050 672.150 ;
        RECT 52.950 671.850 55.050 672.750 ;
        RECT 55.950 671.250 57.750 672.150 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 40.950 667.950 43.050 670.050 ;
        RECT 31.950 664.950 34.050 667.050 ;
        RECT 35.250 665.850 36.750 666.750 ;
        RECT 37.950 664.950 40.050 667.050 ;
        RECT 41.250 665.850 43.050 666.750 ;
        RECT 37.950 662.850 40.050 663.750 ;
        RECT 34.950 632.250 37.050 633.150 ;
        RECT 31.950 628.950 34.050 631.050 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 38.250 629.250 39.750 630.150 ;
        RECT 40.950 628.950 43.050 631.050 ;
        RECT 44.250 629.250 46.050 630.150 ;
        RECT 32.400 622.050 33.450 628.950 ;
        RECT 35.400 625.050 36.450 628.950 ;
        RECT 37.950 625.950 40.050 628.050 ;
        RECT 41.250 626.850 42.750 627.750 ;
        RECT 43.950 625.950 46.050 628.050 ;
        RECT 34.950 622.950 37.050 625.050 ;
        RECT 31.950 619.950 34.050 622.050 ;
        RECT 37.950 619.950 40.050 622.050 ;
        RECT 34.950 616.950 37.050 619.050 ;
        RECT 28.950 604.950 31.050 607.050 ;
        RECT 22.950 601.950 25.050 604.050 ;
        RECT 25.950 601.950 28.050 604.050 ;
        RECT 26.400 601.050 27.450 601.950 ;
        RECT 22.950 598.950 25.050 601.050 ;
        RECT 25.950 598.950 28.050 601.050 ;
        RECT 29.250 599.250 30.750 600.150 ;
        RECT 31.950 598.950 34.050 601.050 ;
        RECT 19.950 592.950 22.050 595.050 ;
        RECT 19.950 589.950 22.050 592.050 ;
        RECT 16.950 565.950 19.050 568.050 ;
        RECT 11.400 563.400 15.450 564.450 ;
        RECT 11.400 562.050 12.450 563.400 ;
        RECT 16.950 562.950 19.050 565.050 ;
        RECT 17.400 562.050 18.450 562.950 ;
        RECT 10.950 559.950 13.050 562.050 ;
        RECT 14.250 560.250 15.750 561.150 ;
        RECT 16.950 559.950 19.050 562.050 ;
        RECT 10.950 557.850 12.750 558.750 ;
        RECT 13.950 556.950 16.050 559.050 ;
        RECT 17.250 557.850 19.050 558.750 ;
        RECT 10.950 553.950 13.050 556.050 ;
        RECT 11.400 529.050 12.450 553.950 ;
        RECT 14.400 541.050 15.450 556.950 ;
        RECT 20.400 556.050 21.450 589.950 ;
        RECT 19.950 553.950 22.050 556.050 ;
        RECT 13.950 538.950 16.050 541.050 ;
        RECT 13.950 535.950 16.050 538.050 ;
        RECT 14.400 529.050 15.450 535.950 ;
        RECT 19.950 532.950 22.050 535.050 ;
        RECT 20.400 529.050 21.450 532.950 ;
        RECT 10.950 526.950 13.050 529.050 ;
        RECT 13.950 526.950 16.050 529.050 ;
        RECT 17.250 527.250 18.750 528.150 ;
        RECT 19.950 526.950 22.050 529.050 ;
        RECT 14.250 524.850 15.750 525.750 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 20.250 524.850 22.050 525.750 ;
        RECT 10.950 521.850 13.050 522.750 ;
        RECT 19.950 517.950 22.050 520.050 ;
        RECT 10.950 516.450 13.050 517.050 ;
        RECT 13.950 516.450 16.050 517.050 ;
        RECT 10.950 515.400 16.050 516.450 ;
        RECT 10.950 514.950 13.050 515.400 ;
        RECT 13.950 514.950 16.050 515.400 ;
        RECT 16.950 514.950 19.050 517.050 ;
        RECT 10.950 487.950 13.050 490.050 ;
        RECT 13.950 487.950 16.050 490.050 ;
        RECT 11.400 487.050 12.450 487.950 ;
        RECT 14.400 487.050 15.450 487.950 ;
        RECT 10.950 484.950 13.050 487.050 ;
        RECT 13.950 484.950 16.050 487.050 ;
        RECT 10.950 482.850 13.050 483.750 ;
        RECT 13.950 482.250 16.050 483.150 ;
        RECT 13.950 478.950 16.050 481.050 ;
        RECT 17.400 478.050 18.450 514.950 ;
        RECT 20.400 484.050 21.450 517.950 ;
        RECT 19.950 481.950 22.050 484.050 ;
        RECT 10.950 475.950 13.050 478.050 ;
        RECT 13.950 475.950 16.050 478.050 ;
        RECT 16.950 475.950 19.050 478.050 ;
        RECT 11.400 448.050 12.450 475.950 ;
        RECT 14.400 457.050 15.450 475.950 ;
        RECT 23.400 459.450 24.450 598.950 ;
        RECT 35.400 598.050 36.450 616.950 ;
        RECT 38.400 598.050 39.450 619.950 ;
        RECT 44.400 613.050 45.450 625.950 ;
        RECT 43.950 610.950 46.050 613.050 ;
        RECT 44.400 607.050 45.450 610.950 ;
        RECT 43.950 604.950 46.050 607.050 ;
        RECT 25.950 596.850 27.750 597.750 ;
        RECT 28.950 595.950 31.050 598.050 ;
        RECT 32.250 596.850 33.750 597.750 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 37.950 595.950 40.050 598.050 ;
        RECT 25.950 592.950 28.050 595.050 ;
        RECT 34.950 593.850 37.050 594.750 ;
        RECT 26.400 520.050 27.450 592.950 ;
        RECT 34.950 563.250 37.050 564.150 ;
        RECT 47.400 562.050 48.450 670.950 ;
        RECT 62.400 670.050 63.450 682.950 ;
        RECT 49.950 667.950 52.050 670.050 ;
        RECT 55.950 667.950 58.050 670.050 ;
        RECT 59.250 668.850 61.050 669.750 ;
        RECT 61.950 667.950 64.050 670.050 ;
        RECT 50.400 667.050 51.450 667.950 ;
        RECT 49.950 664.950 52.050 667.050 ;
        RECT 58.950 664.950 61.050 667.050 ;
        RECT 49.950 661.950 52.050 664.050 ;
        RECT 50.400 628.050 51.450 661.950 ;
        RECT 55.950 637.950 58.050 640.050 ;
        RECT 49.950 625.950 52.050 628.050 ;
        RECT 52.950 607.950 55.050 610.050 ;
        RECT 53.400 604.050 54.450 607.950 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 49.950 599.250 52.050 600.150 ;
        RECT 52.950 599.850 55.050 600.750 ;
        RECT 49.950 595.950 52.050 598.050 ;
        RECT 28.950 559.950 31.050 562.050 ;
        RECT 32.250 560.250 33.750 561.150 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 38.250 560.250 40.050 561.150 ;
        RECT 46.950 559.950 49.050 562.050 ;
        RECT 28.950 557.850 30.750 558.750 ;
        RECT 31.950 556.950 34.050 559.050 ;
        RECT 37.950 556.950 40.050 559.050 ;
        RECT 43.950 556.950 46.050 559.050 ;
        RECT 32.400 556.050 33.450 556.950 ;
        RECT 38.400 556.050 39.450 556.950 ;
        RECT 31.950 553.950 34.050 556.050 ;
        RECT 37.950 553.950 40.050 556.050 ;
        RECT 31.950 538.950 34.050 541.050 ;
        RECT 32.400 532.050 33.450 538.950 ;
        RECT 44.400 538.050 45.450 556.950 ;
        RECT 40.950 535.950 43.050 538.050 ;
        RECT 43.950 535.950 46.050 538.050 ;
        RECT 31.950 529.950 34.050 532.050 ;
        RECT 28.950 527.250 31.050 528.150 ;
        RECT 31.950 527.850 34.050 528.750 ;
        RECT 34.950 527.250 36.750 528.150 ;
        RECT 37.950 526.950 40.050 529.050 ;
        RECT 41.400 526.050 42.450 535.950 ;
        RECT 43.950 526.950 46.050 529.050 ;
        RECT 28.950 523.950 31.050 526.050 ;
        RECT 34.950 523.950 37.050 526.050 ;
        RECT 38.250 524.850 40.050 525.750 ;
        RECT 40.950 523.950 43.050 526.050 ;
        RECT 25.950 517.950 28.050 520.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 25.950 488.250 28.050 489.150 ;
        RECT 25.950 484.950 28.050 487.050 ;
        RECT 29.250 485.250 30.750 486.150 ;
        RECT 31.950 484.950 34.050 487.050 ;
        RECT 35.250 485.250 37.050 486.150 ;
        RECT 25.950 481.950 28.050 484.050 ;
        RECT 28.950 481.950 31.050 484.050 ;
        RECT 32.250 482.850 33.750 483.750 ;
        RECT 34.950 481.950 37.050 484.050 ;
        RECT 20.400 458.400 24.450 459.450 ;
        RECT 13.950 454.950 16.050 457.050 ;
        RECT 13.950 452.850 16.050 453.750 ;
        RECT 16.950 452.250 19.050 453.150 ;
        RECT 16.950 448.950 19.050 451.050 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 10.950 418.950 13.050 421.050 ;
        RECT 11.400 418.050 12.450 418.950 ;
        RECT 17.400 418.050 18.450 445.950 ;
        RECT 10.950 415.950 13.050 418.050 ;
        RECT 14.250 416.250 15.750 417.150 ;
        RECT 16.950 415.950 19.050 418.050 ;
        RECT 10.950 413.850 12.750 414.750 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 17.250 413.850 19.050 414.750 ;
        RECT 13.950 409.950 16.050 412.050 ;
        RECT 16.950 409.950 19.050 412.050 ;
        RECT 14.400 388.050 15.450 409.950 ;
        RECT 13.950 385.950 16.050 388.050 ;
        RECT 10.950 383.250 13.050 384.150 ;
        RECT 13.950 383.850 16.050 384.750 ;
        RECT 10.950 379.950 13.050 382.050 ;
        RECT 11.400 346.050 12.450 379.950 ;
        RECT 17.400 379.050 18.450 409.950 ;
        RECT 16.950 376.950 19.050 379.050 ;
        RECT 10.950 343.950 13.050 346.050 ;
        RECT 10.950 341.250 13.050 342.150 ;
        RECT 16.950 341.250 19.050 342.150 ;
        RECT 16.950 337.950 19.050 340.050 ;
        RECT 17.400 325.050 18.450 337.950 ;
        RECT 16.950 322.950 19.050 325.050 ;
        RECT 10.950 316.950 13.050 319.050 ;
        RECT 11.400 274.050 12.450 316.950 ;
        RECT 20.400 315.450 21.450 458.400 ;
        RECT 22.950 454.950 25.050 457.050 ;
        RECT 22.950 452.850 25.050 453.750 ;
        RECT 26.400 450.450 27.450 481.950 ;
        RECT 23.400 449.400 27.450 450.450 ;
        RECT 23.400 412.050 24.450 449.400 ;
        RECT 29.400 415.050 30.450 481.950 ;
        RECT 38.400 481.050 39.450 490.950 ;
        RECT 40.950 487.950 43.050 490.050 ;
        RECT 41.400 484.050 42.450 487.950 ;
        RECT 40.950 481.950 43.050 484.050 ;
        RECT 37.950 478.950 40.050 481.050 ;
        RECT 37.950 454.950 40.050 457.050 ;
        RECT 34.950 453.450 37.050 454.050 ;
        RECT 32.400 452.400 37.050 453.450 ;
        RECT 32.400 451.050 33.450 452.400 ;
        RECT 34.950 451.950 37.050 452.400 ;
        RECT 38.400 451.050 39.450 454.950 ;
        RECT 41.400 454.050 42.450 481.950 ;
        RECT 44.400 457.050 45.450 526.950 ;
        RECT 47.400 493.050 48.450 559.950 ;
        RECT 52.950 558.450 55.050 559.050 ;
        RECT 50.400 557.400 55.050 558.450 ;
        RECT 50.400 556.050 51.450 557.400 ;
        RECT 52.950 556.950 55.050 557.400 ;
        RECT 49.950 553.950 52.050 556.050 ;
        RECT 52.950 554.850 55.050 555.750 ;
        RECT 56.400 555.450 57.450 637.950 ;
        RECT 59.400 634.050 60.450 664.950 ;
        RECT 65.400 640.050 66.450 772.950 ;
        RECT 74.400 766.050 75.450 775.950 ;
        RECT 76.950 774.450 79.050 775.050 ;
        RECT 80.400 774.450 81.450 778.950 ;
        RECT 76.950 773.400 81.450 774.450 ;
        RECT 76.950 772.950 79.050 773.400 ;
        RECT 76.950 769.950 79.050 772.050 ;
        RECT 73.950 763.950 76.050 766.050 ;
        RECT 77.400 745.050 78.450 769.950 ;
        RECT 80.400 769.050 81.450 773.400 ;
        RECT 85.950 774.450 88.050 775.050 ;
        RECT 89.400 774.450 90.450 811.950 ;
        RECT 92.400 784.050 93.450 814.950 ;
        RECT 98.400 814.050 99.450 829.950 ;
        RECT 101.400 814.050 102.450 841.950 ;
        RECT 107.400 838.050 108.450 841.950 ;
        RECT 106.950 835.950 109.050 838.050 ;
        RECT 103.950 820.950 106.050 823.050 ;
        RECT 104.400 814.050 105.450 820.950 ;
        RECT 110.400 814.050 111.450 844.950 ;
        RECT 116.400 844.050 117.450 848.400 ;
        RECT 118.950 847.950 121.050 848.400 ;
        RECT 122.250 848.250 123.750 849.150 ;
        RECT 124.950 847.950 127.050 850.050 ;
        RECT 199.950 847.950 202.050 850.050 ;
        RECT 205.950 849.450 208.050 850.050 ;
        RECT 205.950 848.400 210.450 849.450 ;
        RECT 205.950 847.950 208.050 848.400 ;
        RECT 118.950 845.850 120.750 846.750 ;
        RECT 121.950 844.950 124.050 847.050 ;
        RECT 125.250 845.850 127.050 846.750 ;
        RECT 133.950 844.950 136.050 847.050 ;
        RECT 136.950 845.250 138.750 846.150 ;
        RECT 139.950 844.950 142.050 847.050 ;
        RECT 145.950 846.450 148.050 847.050 ;
        RECT 145.950 845.400 150.450 846.450 ;
        RECT 145.950 844.950 148.050 845.400 ;
        RECT 115.950 841.950 118.050 844.050 ;
        RECT 116.400 820.050 117.450 841.950 ;
        RECT 122.400 835.050 123.450 844.950 ;
        RECT 134.400 838.050 135.450 844.950 ;
        RECT 136.950 841.950 139.050 844.050 ;
        RECT 140.250 842.850 142.050 843.750 ;
        RECT 142.950 842.250 145.050 843.150 ;
        RECT 145.950 842.850 148.050 843.750 ;
        RECT 137.400 841.050 138.450 841.950 ;
        RECT 149.400 841.050 150.450 845.400 ;
        RECT 157.950 845.250 160.050 846.150 ;
        RECT 163.950 845.250 166.050 846.150 ;
        RECT 181.950 844.950 184.050 847.050 ;
        RECT 187.950 845.250 190.050 846.150 ;
        RECT 157.950 841.950 160.050 844.050 ;
        RECT 161.250 842.250 162.750 843.150 ;
        RECT 163.950 841.950 166.050 844.050 ;
        RECT 181.950 842.850 184.050 843.750 ;
        RECT 187.950 841.950 190.050 844.050 ;
        RECT 191.250 842.250 193.050 843.150 ;
        RECT 136.950 838.950 139.050 841.050 ;
        RECT 142.950 838.950 145.050 841.050 ;
        RECT 148.950 838.950 151.050 841.050 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 118.950 832.950 121.050 835.050 ;
        RECT 121.950 832.950 124.050 835.050 ;
        RECT 115.950 817.950 118.050 820.050 ;
        RECT 119.400 817.050 120.450 832.950 ;
        RECT 143.400 817.050 144.450 838.950 ;
        RECT 158.400 832.050 159.450 841.950 ;
        RECT 160.950 838.950 163.050 841.050 ;
        RECT 164.400 840.450 165.450 841.950 ;
        RECT 164.400 839.400 168.450 840.450 ;
        RECT 157.950 829.950 160.050 832.050 ;
        RECT 118.950 814.950 121.050 817.050 ;
        RECT 122.250 815.250 123.750 816.150 ;
        RECT 124.950 814.950 127.050 817.050 ;
        RECT 142.950 814.950 145.050 817.050 ;
        RECT 97.950 811.950 100.050 814.050 ;
        RECT 100.950 811.950 103.050 814.050 ;
        RECT 103.950 811.950 106.050 814.050 ;
        RECT 107.250 812.250 109.050 813.150 ;
        RECT 109.950 811.950 112.050 814.050 ;
        RECT 118.950 812.850 120.750 813.750 ;
        RECT 121.950 811.950 124.050 814.050 ;
        RECT 125.250 812.850 126.750 813.750 ;
        RECT 127.950 811.950 130.050 814.050 ;
        RECT 136.950 811.950 139.050 814.050 ;
        RECT 139.950 811.950 142.050 814.050 ;
        RECT 97.950 809.850 99.750 810.750 ;
        RECT 100.950 808.950 103.050 811.050 ;
        RECT 104.250 809.850 105.750 810.750 ;
        RECT 106.950 808.950 109.050 811.050 ;
        RECT 100.950 806.850 103.050 807.750 ;
        RECT 107.400 805.050 108.450 808.950 ;
        RECT 106.950 802.950 109.050 805.050 ;
        RECT 91.950 781.950 94.050 784.050 ;
        RECT 91.950 775.950 94.050 778.050 ;
        RECT 118.950 775.950 121.050 778.050 ;
        RECT 92.400 775.050 93.450 775.950 ;
        RECT 119.400 775.050 120.450 775.950 ;
        RECT 85.950 773.400 90.450 774.450 ;
        RECT 85.950 772.950 88.050 773.400 ;
        RECT 91.950 772.950 94.050 775.050 ;
        RECT 95.250 773.250 97.050 774.150 ;
        RECT 109.950 773.250 111.750 774.150 ;
        RECT 112.950 772.950 115.050 775.050 ;
        RECT 118.950 772.950 121.050 775.050 ;
        RECT 122.400 772.050 123.450 811.950 ;
        RECT 127.950 809.850 130.050 810.750 ;
        RECT 130.950 779.250 133.050 780.150 ;
        RECT 137.400 778.050 138.450 811.950 ;
        RECT 143.400 811.050 144.450 814.950 ;
        RECT 161.400 814.050 162.450 838.950 ;
        RECT 167.400 838.050 168.450 839.400 ;
        RECT 190.950 838.950 193.050 841.050 ;
        RECT 163.950 835.950 166.050 838.050 ;
        RECT 166.950 835.950 169.050 838.050 ;
        RECT 164.400 817.050 165.450 835.950 ;
        RECT 169.950 817.950 172.050 820.050 ;
        RECT 175.950 817.950 178.050 820.050 ;
        RECT 163.950 814.950 166.050 817.050 ;
        RECT 167.250 815.250 169.050 816.150 ;
        RECT 169.950 815.850 172.050 816.750 ;
        RECT 172.950 815.250 175.050 816.150 ;
        RECT 145.950 811.950 148.050 814.050 ;
        RECT 149.250 812.250 151.050 813.150 ;
        RECT 160.950 811.950 163.050 814.050 ;
        RECT 163.950 812.850 165.750 813.750 ;
        RECT 166.950 811.950 169.050 814.050 ;
        RECT 172.950 811.950 175.050 814.050 ;
        RECT 167.400 811.050 168.450 811.950 ;
        RECT 139.950 809.850 141.750 810.750 ;
        RECT 142.950 808.950 145.050 811.050 ;
        RECT 146.250 809.850 147.750 810.750 ;
        RECT 148.950 808.950 151.050 811.050 ;
        RECT 166.950 808.950 169.050 811.050 ;
        RECT 142.950 806.850 145.050 807.750 ;
        RECT 149.400 781.050 150.450 808.950 ;
        RECT 148.950 778.950 151.050 781.050 ;
        RECT 157.950 779.250 160.050 780.150 ;
        RECT 127.950 776.250 129.750 777.150 ;
        RECT 130.950 775.950 133.050 778.050 ;
        RECT 134.250 776.250 135.750 777.150 ;
        RECT 136.950 775.950 139.050 778.050 ;
        RECT 151.950 775.950 154.050 778.050 ;
        RECT 155.250 776.250 156.750 777.150 ;
        RECT 157.950 775.950 160.050 778.050 ;
        RECT 161.250 776.250 163.050 777.150 ;
        RECT 131.400 775.050 132.450 775.950 ;
        RECT 127.950 772.950 130.050 775.050 ;
        RECT 130.950 772.950 133.050 775.050 ;
        RECT 133.950 772.950 136.050 775.050 ;
        RECT 137.250 773.850 139.050 774.750 ;
        RECT 151.950 773.850 153.750 774.750 ;
        RECT 154.950 772.950 157.050 775.050 ;
        RECT 128.400 772.050 129.450 772.950 ;
        RECT 85.950 770.850 88.050 771.750 ;
        RECT 88.950 770.250 91.050 771.150 ;
        RECT 91.950 770.850 93.750 771.750 ;
        RECT 94.950 769.950 97.050 772.050 ;
        RECT 109.950 769.950 112.050 772.050 ;
        RECT 113.250 770.850 115.050 771.750 ;
        RECT 115.950 770.250 118.050 771.150 ;
        RECT 118.950 770.850 121.050 771.750 ;
        RECT 121.950 769.950 124.050 772.050 ;
        RECT 127.950 769.950 130.050 772.050 ;
        RECT 79.950 766.950 82.050 769.050 ;
        RECT 88.950 766.950 91.050 769.050 ;
        RECT 95.400 745.050 96.450 769.950 ;
        RECT 128.400 769.050 129.450 769.950 ;
        RECT 115.950 766.950 118.050 769.050 ;
        RECT 127.950 766.950 130.050 769.050 ;
        RECT 109.950 763.950 112.050 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 70.950 744.450 73.050 745.050 ;
        RECT 68.400 743.400 73.050 744.450 ;
        RECT 68.400 715.050 69.450 743.400 ;
        RECT 70.950 742.950 73.050 743.400 ;
        RECT 74.250 743.250 75.750 744.150 ;
        RECT 76.950 742.950 79.050 745.050 ;
        RECT 85.950 742.950 88.050 745.050 ;
        RECT 94.950 742.950 97.050 745.050 ;
        RECT 103.950 742.950 106.050 745.050 ;
        RECT 70.950 740.850 72.750 741.750 ;
        RECT 73.950 739.950 76.050 742.050 ;
        RECT 77.250 740.850 78.750 741.750 ;
        RECT 79.950 741.450 82.050 742.050 ;
        RECT 82.950 741.450 85.050 742.050 ;
        RECT 79.950 740.400 85.050 741.450 ;
        RECT 79.950 739.950 82.050 740.400 ;
        RECT 82.950 739.950 85.050 740.400 ;
        RECT 74.400 733.050 75.450 739.950 ;
        RECT 79.950 737.850 82.050 738.750 ;
        RECT 73.950 730.950 76.050 733.050 ;
        RECT 83.400 727.050 84.450 739.950 ;
        RECT 82.950 724.950 85.050 727.050 ;
        RECT 67.950 712.950 70.050 715.050 ;
        RECT 70.950 705.450 73.050 706.050 ;
        RECT 68.400 704.400 73.050 705.450 ;
        RECT 68.400 700.050 69.450 704.400 ;
        RECT 70.950 703.950 73.050 704.400 ;
        RECT 74.250 704.250 75.750 705.150 ;
        RECT 76.950 703.950 79.050 706.050 ;
        RECT 70.950 701.850 72.750 702.750 ;
        RECT 73.950 700.950 76.050 703.050 ;
        RECT 77.250 701.850 79.050 702.750 ;
        RECT 67.950 697.950 70.050 700.050 ;
        RECT 67.950 694.950 70.050 697.050 ;
        RECT 68.400 667.050 69.450 694.950 ;
        RECT 74.400 688.050 75.450 700.950 ;
        RECT 79.950 697.950 82.050 700.050 ;
        RECT 76.950 688.950 79.050 691.050 ;
        RECT 73.950 685.950 76.050 688.050 ;
        RECT 73.950 679.950 76.050 682.050 ;
        RECT 67.950 664.950 70.050 667.050 ;
        RECT 64.950 637.950 67.050 640.050 ;
        RECT 64.950 635.250 67.050 636.150 ;
        RECT 58.950 631.950 61.050 634.050 ;
        RECT 62.250 632.250 63.750 633.150 ;
        RECT 64.950 631.950 67.050 634.050 ;
        RECT 68.250 632.250 70.050 633.150 ;
        RECT 58.950 629.850 60.750 630.750 ;
        RECT 61.950 628.950 64.050 631.050 ;
        RECT 62.400 619.050 63.450 628.950 ;
        RECT 61.950 616.950 64.050 619.050 ;
        RECT 65.400 616.050 66.450 631.950 ;
        RECT 67.950 628.950 70.050 631.050 ;
        RECT 74.400 622.050 75.450 679.950 ;
        RECT 77.400 670.050 78.450 688.950 ;
        RECT 80.400 673.050 81.450 697.950 ;
        RECT 86.400 682.050 87.450 742.950 ;
        RECT 94.950 740.250 96.750 741.150 ;
        RECT 97.950 739.950 100.050 742.050 ;
        RECT 101.250 740.250 103.050 741.150 ;
        RECT 94.950 736.950 97.050 739.050 ;
        RECT 98.250 737.850 99.750 738.750 ;
        RECT 100.950 736.950 103.050 739.050 ;
        RECT 95.400 736.050 96.450 736.950 ;
        RECT 88.950 733.950 91.050 736.050 ;
        RECT 94.950 733.950 97.050 736.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 85.950 676.950 88.050 679.050 ;
        RECT 86.400 673.050 87.450 676.950 ;
        RECT 89.400 673.050 90.450 733.950 ;
        RECT 97.950 707.250 100.050 708.150 ;
        RECT 91.950 703.950 94.050 706.050 ;
        RECT 95.250 704.250 96.750 705.150 ;
        RECT 97.950 703.950 100.050 706.050 ;
        RECT 101.250 704.250 103.050 705.150 ;
        RECT 98.400 703.050 99.450 703.950 ;
        RECT 91.950 701.850 93.750 702.750 ;
        RECT 94.950 700.950 97.050 703.050 ;
        RECT 97.950 700.950 100.050 703.050 ;
        RECT 100.950 700.950 103.050 703.050 ;
        RECT 95.400 682.050 96.450 700.950 ;
        RECT 94.950 679.950 97.050 682.050 ;
        RECT 97.950 679.950 100.050 682.050 ;
        RECT 79.950 670.950 82.050 673.050 ;
        RECT 83.250 671.250 84.750 672.150 ;
        RECT 85.950 670.950 88.050 673.050 ;
        RECT 88.950 670.950 91.050 673.050 ;
        RECT 98.400 670.050 99.450 679.950 ;
        RECT 101.400 676.050 102.450 700.950 ;
        RECT 104.400 685.050 105.450 742.950 ;
        RECT 103.950 682.950 106.050 685.050 ;
        RECT 106.950 676.950 109.050 679.050 ;
        RECT 100.950 673.950 103.050 676.050 ;
        RECT 107.400 673.050 108.450 676.950 ;
        RECT 100.950 670.950 103.050 673.050 ;
        RECT 104.250 671.250 105.750 672.150 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 76.950 667.950 79.050 670.050 ;
        RECT 80.250 668.850 81.750 669.750 ;
        RECT 82.950 667.950 85.050 670.050 ;
        RECT 86.250 668.850 88.050 669.750 ;
        RECT 97.950 667.950 100.050 670.050 ;
        RECT 101.250 668.850 102.750 669.750 ;
        RECT 103.950 667.950 106.050 670.050 ;
        RECT 107.250 668.850 109.050 669.750 ;
        RECT 76.950 665.850 79.050 666.750 ;
        RECT 79.950 664.950 82.050 667.050 ;
        RECT 97.950 665.850 100.050 666.750 ;
        RECT 80.400 634.050 81.450 664.950 ;
        RECT 85.950 635.250 88.050 636.150 ;
        RECT 79.950 631.950 82.050 634.050 ;
        RECT 83.250 632.250 84.750 633.150 ;
        RECT 85.950 631.950 88.050 634.050 ;
        RECT 89.250 632.250 91.050 633.150 ;
        RECT 79.950 629.850 81.750 630.750 ;
        RECT 82.950 628.950 85.050 631.050 ;
        RECT 73.950 619.950 76.050 622.050 ;
        RECT 79.950 619.950 82.050 622.050 ;
        RECT 64.950 613.950 67.050 616.050 ;
        RECT 67.950 613.950 70.050 616.050 ;
        RECT 61.950 607.950 64.050 610.050 ;
        RECT 62.400 597.450 63.450 607.950 ;
        RECT 68.400 604.050 69.450 613.950 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 64.950 599.250 67.050 600.150 ;
        RECT 67.950 599.850 70.050 600.750 ;
        RECT 73.950 600.450 76.050 601.050 ;
        RECT 70.950 599.250 72.750 600.150 ;
        RECT 73.950 599.400 78.450 600.450 ;
        RECT 73.950 598.950 76.050 599.400 ;
        RECT 64.950 597.450 67.050 598.050 ;
        RECT 62.400 596.400 67.050 597.450 ;
        RECT 64.950 595.950 67.050 596.400 ;
        RECT 70.950 595.950 73.050 598.050 ;
        RECT 74.250 596.850 76.050 597.750 ;
        RECT 58.950 557.250 60.750 558.150 ;
        RECT 61.950 556.950 64.050 559.050 ;
        RECT 67.950 557.250 70.050 558.150 ;
        RECT 73.950 556.950 76.050 559.050 ;
        RECT 58.950 555.450 61.050 556.050 ;
        RECT 56.400 554.400 61.050 555.450 ;
        RECT 62.250 554.850 64.050 555.750 ;
        RECT 58.950 553.950 61.050 554.400 ;
        RECT 64.950 553.950 67.050 556.050 ;
        RECT 67.950 553.950 70.050 556.050 ;
        RECT 50.400 532.050 51.450 553.950 ;
        RECT 55.950 532.950 58.050 535.050 ;
        RECT 56.400 532.050 57.450 532.950 ;
        RECT 49.950 529.950 52.050 532.050 ;
        RECT 55.950 529.950 58.050 532.050 ;
        RECT 49.950 527.850 52.050 528.750 ;
        RECT 52.950 527.250 55.050 528.150 ;
        RECT 52.950 525.450 55.050 526.050 ;
        RECT 56.400 525.450 57.450 529.950 ;
        RECT 59.400 526.050 60.450 553.950 ;
        RECT 61.950 535.950 64.050 538.050 ;
        RECT 52.950 524.400 57.450 525.450 ;
        RECT 52.950 523.950 55.050 524.400 ;
        RECT 58.950 523.950 61.050 526.050 ;
        RECT 62.400 496.050 63.450 535.950 ;
        RECT 65.400 529.050 66.450 553.950 ;
        RECT 74.400 535.050 75.450 556.950 ;
        RECT 73.950 532.950 76.050 535.050 ;
        RECT 64.950 526.950 67.050 529.050 ;
        RECT 68.250 527.250 69.750 528.150 ;
        RECT 70.950 526.950 73.050 529.050 ;
        RECT 74.400 526.050 75.450 532.950 ;
        RECT 64.950 524.850 66.750 525.750 ;
        RECT 67.950 523.950 70.050 526.050 ;
        RECT 71.250 524.850 72.750 525.750 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 73.950 521.850 76.050 522.750 ;
        RECT 77.400 519.450 78.450 599.400 ;
        RECT 80.400 556.050 81.450 619.950 ;
        RECT 83.400 619.050 84.450 628.950 ;
        RECT 86.400 625.050 87.450 631.950 ;
        RECT 110.400 631.050 111.450 763.950 ;
        RECT 113.400 742.050 114.450 763.950 ;
        RECT 115.950 742.950 118.050 745.050 ;
        RECT 119.250 743.250 120.750 744.150 ;
        RECT 121.950 742.950 124.050 745.050 ;
        RECT 112.950 739.950 115.050 742.050 ;
        RECT 116.250 740.850 117.750 741.750 ;
        RECT 118.950 739.950 121.050 742.050 ;
        RECT 122.250 740.850 124.050 741.750 ;
        RECT 112.950 737.850 115.050 738.750 ;
        RECT 115.950 736.950 118.050 739.050 ;
        RECT 116.400 706.050 117.450 736.950 ;
        RECT 121.950 707.250 124.050 708.150 ;
        RECT 115.950 703.950 118.050 706.050 ;
        RECT 119.250 704.250 120.750 705.150 ;
        RECT 121.950 703.950 124.050 706.050 ;
        RECT 125.250 704.250 127.050 705.150 ;
        RECT 115.950 701.850 117.750 702.750 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 122.400 676.050 123.450 703.950 ;
        RECT 124.950 700.950 127.050 703.050 ;
        RECT 125.400 691.050 126.450 700.950 ;
        RECT 131.400 700.050 132.450 772.950 ;
        RECT 136.950 769.950 139.050 772.050 ;
        RECT 133.950 766.950 136.050 769.050 ;
        RECT 134.400 745.050 135.450 766.950 ;
        RECT 137.400 745.050 138.450 769.950 ;
        RECT 155.400 766.050 156.450 772.950 ;
        RECT 154.950 763.950 157.050 766.050 ;
        RECT 142.950 745.950 145.050 748.050 ;
        RECT 148.950 745.950 151.050 748.050 ;
        RECT 158.400 747.450 159.450 775.950 ;
        RECT 160.950 772.950 163.050 775.050 ;
        RECT 167.400 763.050 168.450 808.950 ;
        RECT 173.400 808.050 174.450 811.950 ;
        RECT 176.400 811.050 177.450 817.950 ;
        RECT 193.950 814.950 196.050 817.050 ;
        RECT 181.950 813.450 184.050 814.050 ;
        RECT 179.400 812.400 184.050 813.450 ;
        RECT 179.400 811.050 180.450 812.400 ;
        RECT 181.950 811.950 184.050 812.400 ;
        RECT 187.950 811.950 190.050 814.050 ;
        RECT 191.250 812.250 193.050 813.150 ;
        RECT 175.950 808.950 178.050 811.050 ;
        RECT 178.950 808.950 181.050 811.050 ;
        RECT 181.950 809.850 183.750 810.750 ;
        RECT 184.950 808.950 187.050 811.050 ;
        RECT 188.250 809.850 189.750 810.750 ;
        RECT 190.950 810.450 193.050 811.050 ;
        RECT 194.400 810.450 195.450 814.950 ;
        RECT 190.950 809.400 195.450 810.450 ;
        RECT 190.950 808.950 193.050 809.400 ;
        RECT 172.950 805.950 175.050 808.050 ;
        RECT 176.400 807.450 177.450 808.950 ;
        RECT 176.400 806.400 180.450 807.450 ;
        RECT 184.950 806.850 187.050 807.750 ;
        RECT 172.950 774.450 175.050 775.050 ;
        RECT 172.950 773.400 177.450 774.450 ;
        RECT 172.950 772.950 175.050 773.400 ;
        RECT 169.950 770.250 172.050 771.150 ;
        RECT 172.950 770.850 175.050 771.750 ;
        RECT 169.950 766.950 172.050 769.050 ;
        RECT 169.950 763.950 172.050 766.050 ;
        RECT 166.950 760.950 169.050 763.050 ;
        RECT 160.950 747.450 163.050 748.050 ;
        RECT 158.400 746.400 163.050 747.450 ;
        RECT 160.950 745.950 163.050 746.400 ;
        RECT 143.400 745.050 144.450 745.950 ;
        RECT 133.950 742.950 136.050 745.050 ;
        RECT 136.950 742.950 139.050 745.050 ;
        RECT 140.250 743.250 141.750 744.150 ;
        RECT 142.950 742.950 145.050 745.050 ;
        RECT 134.400 742.050 135.450 742.950 ;
        RECT 149.400 742.050 150.450 745.950 ;
        RECT 154.950 744.450 157.050 745.050 ;
        RECT 152.400 743.400 157.050 744.450 ;
        RECT 133.950 739.950 136.050 742.050 ;
        RECT 137.250 740.850 138.750 741.750 ;
        RECT 139.950 739.950 142.050 742.050 ;
        RECT 143.250 740.850 145.050 741.750 ;
        RECT 148.950 739.950 151.050 742.050 ;
        RECT 133.950 737.850 136.050 738.750 ;
        RECT 152.400 709.050 153.450 743.400 ;
        RECT 154.950 742.950 157.050 743.400 ;
        RECT 158.250 743.250 160.050 744.150 ;
        RECT 160.950 743.850 163.050 744.750 ;
        RECT 163.950 743.250 166.050 744.150 ;
        RECT 166.950 742.950 169.050 745.050 ;
        RECT 154.950 740.850 156.750 741.750 ;
        RECT 157.950 739.950 160.050 742.050 ;
        RECT 163.950 741.450 166.050 742.050 ;
        RECT 167.400 741.450 168.450 742.950 ;
        RECT 163.950 740.400 168.450 741.450 ;
        RECT 163.950 739.950 166.050 740.400 ;
        RECT 151.950 706.950 154.050 709.050 ;
        RECT 136.950 702.450 139.050 703.050 ;
        RECT 136.950 701.400 141.450 702.450 ;
        RECT 136.950 700.950 139.050 701.400 ;
        RECT 130.950 697.950 133.050 700.050 ;
        RECT 133.950 698.250 136.050 699.150 ;
        RECT 136.950 698.850 139.050 699.750 ;
        RECT 133.950 694.950 136.050 697.050 ;
        RECT 134.400 691.050 135.450 694.950 ;
        RECT 124.950 688.950 127.050 691.050 ;
        RECT 133.950 688.950 136.050 691.050 ;
        RECT 140.400 682.050 141.450 701.400 ;
        RECT 151.950 700.950 154.050 703.050 ;
        RECT 148.950 698.250 151.050 699.150 ;
        RECT 151.950 698.850 154.050 699.750 ;
        RECT 158.400 697.050 159.450 739.950 ;
        RECT 163.950 730.950 166.050 733.050 ;
        RECT 148.950 694.950 151.050 697.050 ;
        RECT 157.950 694.950 160.050 697.050 ;
        RECT 149.400 685.050 150.450 694.950 ;
        RECT 148.950 682.950 151.050 685.050 ;
        RECT 127.950 679.950 130.050 682.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 115.950 673.950 118.050 676.050 ;
        RECT 121.950 673.950 124.050 676.050 ;
        RECT 115.950 671.850 118.050 672.750 ;
        RECT 118.950 671.250 121.050 672.150 ;
        RECT 118.950 667.950 121.050 670.050 ;
        RECT 128.400 669.450 129.450 679.950 ;
        RECT 133.950 676.950 136.050 679.050 ;
        RECT 134.400 676.050 135.450 676.950 ;
        RECT 133.950 673.950 136.050 676.050 ;
        RECT 130.950 671.250 133.050 672.150 ;
        RECT 133.950 671.850 136.050 672.750 ;
        RECT 136.950 671.250 138.750 672.150 ;
        RECT 139.950 670.950 142.050 673.050 ;
        RECT 149.400 670.050 150.450 682.950 ;
        RECT 157.950 675.450 160.050 676.050 ;
        RECT 157.950 674.400 162.450 675.450 ;
        RECT 157.950 673.950 160.050 674.400 ;
        RECT 151.950 670.950 154.050 673.050 ;
        RECT 154.950 671.250 157.050 672.150 ;
        RECT 157.950 671.850 160.050 672.750 ;
        RECT 130.950 669.450 133.050 670.050 ;
        RECT 128.400 668.400 133.050 669.450 ;
        RECT 130.950 667.950 133.050 668.400 ;
        RECT 136.950 667.950 139.050 670.050 ;
        RECT 140.250 668.850 142.050 669.750 ;
        RECT 148.950 667.950 151.050 670.050 ;
        RECT 133.950 643.950 136.050 646.050 ;
        RECT 121.950 632.250 124.050 633.150 ;
        RECT 88.950 628.950 91.050 631.050 ;
        RECT 100.950 630.450 103.050 631.050 ;
        RECT 98.400 629.400 103.050 630.450 ;
        RECT 85.950 622.950 88.050 625.050 ;
        RECT 86.400 622.050 87.450 622.950 ;
        RECT 85.950 619.950 88.050 622.050 ;
        RECT 82.950 616.950 85.050 619.050 ;
        RECT 89.400 610.050 90.450 628.950 ;
        RECT 98.400 619.050 99.450 629.400 ;
        RECT 100.950 628.950 103.050 629.400 ;
        RECT 106.950 629.250 109.050 630.150 ;
        RECT 109.950 628.950 112.050 631.050 ;
        RECT 112.950 628.950 115.050 631.050 ;
        RECT 121.950 628.950 124.050 631.050 ;
        RECT 125.250 629.250 126.750 630.150 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 131.250 629.250 133.050 630.150 ;
        RECT 100.950 626.850 103.050 627.750 ;
        RECT 106.950 625.950 109.050 628.050 ;
        RECT 110.250 626.250 112.050 627.150 ;
        RECT 97.950 616.950 100.050 619.050 ;
        RECT 94.950 613.950 97.050 616.050 ;
        RECT 88.950 607.950 91.050 610.050 ;
        RECT 82.950 604.950 85.050 607.050 ;
        RECT 91.950 604.950 94.050 607.050 ;
        RECT 83.400 598.050 84.450 604.950 ;
        RECT 92.400 604.050 93.450 604.950 ;
        RECT 91.950 601.950 94.050 604.050 ;
        RECT 95.400 601.050 96.450 613.950 ;
        RECT 107.400 601.050 108.450 625.950 ;
        RECT 109.950 622.950 112.050 625.050 ;
        RECT 110.400 616.050 111.450 622.950 ;
        RECT 109.950 613.950 112.050 616.050 ;
        RECT 113.400 604.050 114.450 628.950 ;
        RECT 124.950 625.950 127.050 628.050 ;
        RECT 128.250 626.850 129.750 627.750 ;
        RECT 130.950 625.950 133.050 628.050 ;
        RECT 121.950 622.950 124.050 625.050 ;
        RECT 112.950 601.950 115.050 604.050 ;
        RECT 122.400 601.050 123.450 622.950 ;
        RECT 131.400 607.050 132.450 625.950 ;
        RECT 130.950 604.950 133.050 607.050 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 92.250 599.850 93.750 600.750 ;
        RECT 94.950 598.950 97.050 601.050 ;
        RECT 106.950 598.950 109.050 601.050 ;
        RECT 109.950 599.250 112.050 600.150 ;
        RECT 112.950 599.850 115.050 600.750 ;
        RECT 121.950 598.950 124.050 601.050 ;
        RECT 125.250 599.250 126.750 600.150 ;
        RECT 127.950 598.950 130.050 601.050 ;
        RECT 82.950 595.950 85.050 598.050 ;
        RECT 88.950 596.850 91.050 597.750 ;
        RECT 94.950 596.850 97.050 597.750 ;
        RECT 107.400 595.050 108.450 598.950 ;
        RECT 131.400 598.050 132.450 604.950 ;
        RECT 109.950 595.950 112.050 598.050 ;
        RECT 121.950 596.850 123.750 597.750 ;
        RECT 124.950 595.950 127.050 598.050 ;
        RECT 128.250 596.850 129.750 597.750 ;
        RECT 130.950 595.950 133.050 598.050 ;
        RECT 106.950 592.950 109.050 595.050 ;
        RECT 130.950 593.850 133.050 594.750 ;
        RECT 82.950 560.250 85.050 561.150 ;
        RECT 97.950 559.950 100.050 562.050 ;
        RECT 103.950 561.450 106.050 562.050 ;
        RECT 101.400 560.400 106.050 561.450 ;
        RECT 82.950 556.950 85.050 559.050 ;
        RECT 86.250 557.250 87.750 558.150 ;
        RECT 88.950 556.950 91.050 559.050 ;
        RECT 92.250 557.250 94.050 558.150 ;
        RECT 83.400 556.050 84.450 556.950 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 82.950 553.950 85.050 556.050 ;
        RECT 85.950 553.950 88.050 556.050 ;
        RECT 89.250 554.850 90.750 555.750 ;
        RECT 91.950 553.950 94.050 556.050 ;
        RECT 86.400 550.050 87.450 553.950 ;
        RECT 92.400 553.050 93.450 553.950 ;
        RECT 91.950 550.950 94.050 553.050 ;
        RECT 85.950 547.950 88.050 550.050 ;
        RECT 91.950 529.950 94.050 532.050 ;
        RECT 88.950 526.950 91.050 529.050 ;
        RECT 89.400 523.050 90.450 526.950 ;
        RECT 92.400 526.050 93.450 529.950 ;
        RECT 91.950 523.950 94.050 526.050 ;
        RECT 95.250 524.250 97.050 525.150 ;
        RECT 85.950 521.850 87.750 522.750 ;
        RECT 88.950 520.950 91.050 523.050 ;
        RECT 92.250 521.850 93.750 522.750 ;
        RECT 94.950 520.950 97.050 523.050 ;
        RECT 74.400 518.400 78.450 519.450 ;
        RECT 88.950 518.850 91.050 519.750 ;
        RECT 52.950 493.950 55.050 496.050 ;
        RECT 61.950 493.950 64.050 496.050 ;
        RECT 46.950 490.950 49.050 493.050 ;
        RECT 46.950 487.950 49.050 490.050 ;
        RECT 47.400 487.050 48.450 487.950 ;
        RECT 46.950 484.950 49.050 487.050 ;
        RECT 46.950 482.850 49.050 483.750 ;
        RECT 49.950 482.250 52.050 483.150 ;
        RECT 49.950 480.450 52.050 481.050 ;
        RECT 53.400 480.450 54.450 493.950 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 59.400 490.050 60.450 490.950 ;
        RECT 58.950 487.950 61.050 490.050 ;
        RECT 64.950 489.450 67.050 490.050 ;
        RECT 62.250 488.250 63.750 489.150 ;
        RECT 64.950 488.400 69.450 489.450 ;
        RECT 64.950 487.950 67.050 488.400 ;
        RECT 58.950 485.850 60.750 486.750 ;
        RECT 61.950 484.950 64.050 487.050 ;
        RECT 65.250 485.850 67.050 486.750 ;
        RECT 68.400 484.050 69.450 488.400 ;
        RECT 58.950 481.950 61.050 484.050 ;
        RECT 67.950 481.950 70.050 484.050 ;
        RECT 49.950 479.400 54.450 480.450 ;
        RECT 49.950 478.950 52.050 479.400 ;
        RECT 53.400 460.050 54.450 479.400 ;
        RECT 59.400 463.050 60.450 481.950 ;
        RECT 58.950 460.950 61.050 463.050 ;
        RECT 52.950 457.950 55.050 460.050 ;
        RECT 43.950 454.950 46.050 457.050 ;
        RECT 59.400 454.050 60.450 460.950 ;
        RECT 70.950 454.950 73.050 457.050 ;
        RECT 40.950 451.950 43.050 454.050 ;
        RECT 44.250 452.250 46.050 453.150 ;
        RECT 46.950 451.950 49.050 454.050 ;
        RECT 55.950 452.250 57.750 453.150 ;
        RECT 58.950 451.950 61.050 454.050 ;
        RECT 62.250 452.250 64.050 453.150 ;
        RECT 31.950 448.950 34.050 451.050 ;
        RECT 34.950 449.850 36.750 450.750 ;
        RECT 37.950 448.950 40.050 451.050 ;
        RECT 41.250 449.850 42.750 450.750 ;
        RECT 43.950 450.450 46.050 451.050 ;
        RECT 47.400 450.450 48.450 451.950 ;
        RECT 43.950 449.400 48.450 450.450 ;
        RECT 43.950 448.950 46.050 449.400 ;
        RECT 55.950 448.950 58.050 451.050 ;
        RECT 59.250 449.850 60.750 450.750 ;
        RECT 61.950 448.950 64.050 451.050 ;
        RECT 32.400 448.050 33.450 448.950 ;
        RECT 56.400 448.050 57.450 448.950 ;
        RECT 31.950 445.950 34.050 448.050 ;
        RECT 37.950 446.850 40.050 447.750 ;
        RECT 55.950 445.950 58.050 448.050 ;
        RECT 37.950 418.950 40.050 421.050 ;
        RECT 34.950 416.250 37.050 417.150 ;
        RECT 25.950 413.250 27.750 414.150 ;
        RECT 28.950 412.950 31.050 415.050 ;
        RECT 32.250 413.250 33.750 414.150 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 22.950 409.950 25.050 412.050 ;
        RECT 25.950 409.950 28.050 412.050 ;
        RECT 29.250 410.850 30.750 411.750 ;
        RECT 31.950 409.950 34.050 412.050 ;
        RECT 26.400 400.050 27.450 409.950 ;
        RECT 28.950 406.950 31.050 409.050 ;
        RECT 25.950 397.950 28.050 400.050 ;
        RECT 22.950 388.950 25.050 391.050 ;
        RECT 23.400 388.050 24.450 388.950 ;
        RECT 22.950 385.950 25.050 388.050 ;
        RECT 22.950 383.850 25.050 384.750 ;
        RECT 25.950 383.250 28.050 384.150 ;
        RECT 25.950 379.950 28.050 382.050 ;
        RECT 25.950 376.950 28.050 379.050 ;
        RECT 22.950 364.950 25.050 367.050 ;
        RECT 23.400 340.050 24.450 364.950 ;
        RECT 22.950 337.950 25.050 340.050 ;
        RECT 20.400 314.400 24.450 315.450 ;
        RECT 19.950 312.450 22.050 313.050 ;
        RECT 17.400 311.400 22.050 312.450 ;
        RECT 13.950 308.850 16.050 309.750 ;
        RECT 17.400 301.050 18.450 311.400 ;
        RECT 19.950 310.950 22.050 311.400 ;
        RECT 19.950 308.850 22.050 309.750 ;
        RECT 16.950 298.950 19.050 301.050 ;
        RECT 16.950 275.250 19.050 276.150 ;
        RECT 10.950 271.950 13.050 274.050 ;
        RECT 14.250 272.250 15.750 273.150 ;
        RECT 16.950 271.950 19.050 274.050 ;
        RECT 20.250 272.250 22.050 273.150 ;
        RECT 10.950 269.850 12.750 270.750 ;
        RECT 13.950 268.950 16.050 271.050 ;
        RECT 17.400 265.050 18.450 271.950 ;
        RECT 19.950 268.950 22.050 271.050 ;
        RECT 20.400 268.050 21.450 268.950 ;
        RECT 19.950 265.950 22.050 268.050 ;
        RECT 16.950 262.950 19.050 265.050 ;
        RECT 20.400 256.050 21.450 265.950 ;
        RECT 19.950 253.950 22.050 256.050 ;
        RECT 10.950 244.950 13.050 247.050 ;
        RECT 11.400 238.050 12.450 244.950 ;
        RECT 10.950 235.950 13.050 238.050 ;
        RECT 16.950 235.950 19.050 238.050 ;
        RECT 20.250 236.250 22.050 237.150 ;
        RECT 10.950 233.850 12.750 234.750 ;
        RECT 13.950 232.950 16.050 235.050 ;
        RECT 17.250 233.850 18.750 234.750 ;
        RECT 19.950 232.950 22.050 235.050 ;
        RECT 13.950 230.850 16.050 231.750 ;
        RECT 16.950 229.950 19.050 232.050 ;
        RECT 10.950 226.950 13.050 229.050 ;
        RECT 11.400 202.050 12.450 226.950 ;
        RECT 17.400 214.050 18.450 229.950 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 16.950 203.250 19.050 204.150 ;
        RECT 10.950 199.950 13.050 202.050 ;
        RECT 14.250 200.250 15.750 201.150 ;
        RECT 16.950 199.950 19.050 202.050 ;
        RECT 20.250 200.250 22.050 201.150 ;
        RECT 10.950 197.850 12.750 198.750 ;
        RECT 13.950 196.950 16.050 199.050 ;
        RECT 17.400 187.050 18.450 199.950 ;
        RECT 19.950 196.950 22.050 199.050 ;
        RECT 16.950 184.950 19.050 187.050 ;
        RECT 20.400 184.050 21.450 196.950 ;
        RECT 19.950 181.950 22.050 184.050 ;
        RECT 13.950 175.950 16.050 178.050 ;
        RECT 14.400 172.050 15.450 175.950 ;
        RECT 13.950 169.950 16.050 172.050 ;
        RECT 23.400 171.450 24.450 314.400 ;
        RECT 26.400 190.050 27.450 376.950 ;
        RECT 29.400 346.050 30.450 406.950 ;
        RECT 35.400 388.050 36.450 412.950 ;
        RECT 34.950 385.950 37.050 388.050 ;
        RECT 38.400 367.050 39.450 418.950 ;
        RECT 56.400 418.050 57.450 445.950 ;
        RECT 62.400 429.450 63.450 448.950 ;
        RECT 71.400 436.050 72.450 454.950 ;
        RECT 70.950 433.950 73.050 436.050 ;
        RECT 74.400 432.450 75.450 518.400 ;
        RECT 82.950 487.950 85.050 490.050 ;
        RECT 83.400 487.050 84.450 487.950 ;
        RECT 76.950 484.950 79.050 487.050 ;
        RECT 82.950 484.950 85.050 487.050 ;
        RECT 86.250 485.250 88.050 486.150 ;
        RECT 76.950 482.850 79.050 483.750 ;
        RECT 79.950 482.250 82.050 483.150 ;
        RECT 82.950 482.850 84.750 483.750 ;
        RECT 85.950 481.950 88.050 484.050 ;
        RECT 79.950 480.450 82.050 481.050 ;
        RECT 77.400 479.400 82.050 480.450 ;
        RECT 77.400 454.050 78.450 479.400 ;
        RECT 79.950 478.950 82.050 479.400 ;
        RECT 86.400 469.050 87.450 481.950 ;
        RECT 95.400 478.050 96.450 520.950 ;
        RECT 98.400 496.050 99.450 559.950 ;
        RECT 101.400 538.050 102.450 560.400 ;
        RECT 103.950 559.950 106.050 560.400 ;
        RECT 107.250 560.250 108.750 561.150 ;
        RECT 109.950 559.950 112.050 562.050 ;
        RECT 127.950 560.250 130.050 561.150 ;
        RECT 103.950 557.850 105.750 558.750 ;
        RECT 106.950 556.950 109.050 559.050 ;
        RECT 110.250 557.850 112.050 558.750 ;
        RECT 118.950 557.250 120.750 558.150 ;
        RECT 121.950 556.950 124.050 559.050 ;
        RECT 125.250 557.250 126.750 558.150 ;
        RECT 127.950 556.950 130.050 559.050 ;
        RECT 107.400 556.050 108.450 556.950 ;
        RECT 134.400 556.050 135.450 643.950 ;
        RECT 136.950 628.950 139.050 631.050 ;
        RECT 142.950 630.450 145.050 631.050 ;
        RECT 142.950 629.400 147.450 630.450 ;
        RECT 142.950 628.950 145.050 629.400 ;
        RECT 137.400 625.050 138.450 628.950 ;
        RECT 139.950 626.250 142.050 627.150 ;
        RECT 142.950 626.850 145.050 627.750 ;
        RECT 136.950 622.950 139.050 625.050 ;
        RECT 139.950 622.950 142.050 625.050 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 143.400 604.050 144.450 604.950 ;
        RECT 146.400 604.050 147.450 629.400 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 145.950 601.950 148.050 604.050 ;
        RECT 136.950 598.950 139.050 601.050 ;
        RECT 142.950 599.850 145.050 600.750 ;
        RECT 145.950 599.250 148.050 600.150 ;
        RECT 106.950 553.950 109.050 556.050 ;
        RECT 109.950 553.950 112.050 556.050 ;
        RECT 118.950 555.450 121.050 556.050 ;
        RECT 116.400 554.400 121.050 555.450 ;
        RECT 122.250 554.850 123.750 555.750 ;
        RECT 107.400 547.050 108.450 553.950 ;
        RECT 106.950 544.950 109.050 547.050 ;
        RECT 100.950 535.950 103.050 538.050 ;
        RECT 97.950 493.950 100.050 496.050 ;
        RECT 100.950 493.950 103.050 496.050 ;
        RECT 97.950 485.250 100.050 486.150 ;
        RECT 97.950 483.450 100.050 484.050 ;
        RECT 101.400 483.450 102.450 493.950 ;
        RECT 103.950 487.950 106.050 490.050 ;
        RECT 103.950 485.850 106.050 486.750 ;
        RECT 106.950 485.250 109.050 486.150 ;
        RECT 97.950 482.400 102.450 483.450 ;
        RECT 97.950 481.950 100.050 482.400 ;
        RECT 106.950 481.950 109.050 484.050 ;
        RECT 94.950 475.950 97.050 478.050 ;
        RECT 85.950 466.950 88.050 469.050 ;
        RECT 85.950 457.950 88.050 460.050 ;
        RECT 94.950 457.950 97.050 460.050 ;
        RECT 100.950 457.950 103.050 460.050 ;
        RECT 86.400 457.050 87.450 457.950 ;
        RECT 95.400 457.050 96.450 457.950 ;
        RECT 101.400 457.050 102.450 457.950 ;
        RECT 79.950 454.950 82.050 457.050 ;
        RECT 83.250 455.250 84.750 456.150 ;
        RECT 85.950 454.950 88.050 457.050 ;
        RECT 91.950 454.950 94.050 457.050 ;
        RECT 94.950 454.950 97.050 457.050 ;
        RECT 98.250 455.250 99.750 456.150 ;
        RECT 100.950 454.950 103.050 457.050 ;
        RECT 76.950 451.950 79.050 454.050 ;
        RECT 80.250 452.850 81.750 453.750 ;
        RECT 82.950 451.950 85.050 454.050 ;
        RECT 86.250 452.850 88.050 453.750 ;
        RECT 76.950 449.850 79.050 450.750 ;
        RECT 74.400 431.400 78.450 432.450 ;
        RECT 59.400 428.400 63.450 429.450 ;
        RECT 55.950 415.950 58.050 418.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 49.950 410.850 52.050 411.750 ;
        RECT 52.950 410.250 55.050 411.150 ;
        RECT 52.950 406.950 55.050 409.050 ;
        RECT 53.400 400.050 54.450 406.950 ;
        RECT 40.950 397.950 43.050 400.050 ;
        RECT 52.950 397.950 55.050 400.050 ;
        RECT 41.400 385.050 42.450 397.950 ;
        RECT 56.400 391.050 57.450 415.950 ;
        RECT 59.400 409.050 60.450 428.400 ;
        RECT 73.950 421.950 76.050 424.050 ;
        RECT 61.950 412.950 64.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 71.250 413.250 73.050 414.150 ;
        RECT 74.400 412.050 75.450 421.950 ;
        RECT 61.950 410.850 64.050 411.750 ;
        RECT 64.950 410.250 67.050 411.150 ;
        RECT 67.950 410.850 69.750 411.750 ;
        RECT 70.950 409.950 73.050 412.050 ;
        RECT 73.950 409.950 76.050 412.050 ;
        RECT 71.400 409.050 72.450 409.950 ;
        RECT 58.950 406.950 61.050 409.050 ;
        RECT 64.950 406.950 67.050 409.050 ;
        RECT 70.950 406.950 73.050 409.050 ;
        RECT 65.400 406.050 66.450 406.950 ;
        RECT 64.950 403.950 67.050 406.050 ;
        RECT 55.950 388.950 58.050 391.050 ;
        RECT 46.950 387.450 49.050 388.050 ;
        RECT 46.950 386.400 54.450 387.450 ;
        RECT 46.950 385.950 49.050 386.400 ;
        RECT 40.950 382.950 43.050 385.050 ;
        RECT 44.250 383.250 46.050 384.150 ;
        RECT 46.950 383.850 49.050 384.750 ;
        RECT 49.950 383.250 52.050 384.150 ;
        RECT 40.950 380.850 42.750 381.750 ;
        RECT 43.950 379.950 46.050 382.050 ;
        RECT 49.950 379.950 52.050 382.050 ;
        RECT 53.400 379.050 54.450 386.400 ;
        RECT 70.950 385.950 73.050 388.050 ;
        RECT 58.950 382.950 61.050 385.050 ;
        RECT 59.400 382.050 60.450 382.950 ;
        RECT 55.950 379.950 58.050 382.050 ;
        RECT 58.950 379.950 61.050 382.050 ;
        RECT 64.950 379.950 67.050 382.050 ;
        RECT 68.250 380.250 70.050 381.150 ;
        RECT 40.950 376.950 43.050 379.050 ;
        RECT 52.950 376.950 55.050 379.050 ;
        RECT 37.950 364.950 40.050 367.050 ;
        RECT 34.950 347.250 37.050 348.150 ;
        RECT 28.950 343.950 31.050 346.050 ;
        RECT 32.250 344.250 33.750 345.150 ;
        RECT 34.950 343.950 37.050 346.050 ;
        RECT 38.250 344.250 40.050 345.150 ;
        RECT 28.950 341.850 30.750 342.750 ;
        RECT 31.950 340.950 34.050 343.050 ;
        RECT 35.400 339.450 36.450 343.950 ;
        RECT 37.950 340.950 40.050 343.050 ;
        RECT 38.400 340.050 39.450 340.950 ;
        RECT 32.400 338.400 36.450 339.450 ;
        RECT 28.950 313.950 31.050 316.050 ;
        RECT 29.400 307.050 30.450 313.950 ;
        RECT 28.950 304.950 31.050 307.050 ;
        RECT 32.400 303.450 33.450 338.400 ;
        RECT 37.950 337.950 40.050 340.050 ;
        RECT 41.400 316.050 42.450 376.950 ;
        RECT 43.950 346.950 46.050 349.050 ;
        RECT 52.950 346.950 55.050 349.050 ;
        RECT 44.400 340.050 45.450 346.950 ;
        RECT 53.400 346.050 54.450 346.950 ;
        RECT 46.950 343.950 49.050 346.050 ;
        RECT 50.250 344.250 51.750 345.150 ;
        RECT 52.950 343.950 55.050 346.050 ;
        RECT 46.950 341.850 48.750 342.750 ;
        RECT 49.950 340.950 52.050 343.050 ;
        RECT 53.250 341.850 55.050 342.750 ;
        RECT 43.950 337.950 46.050 340.050 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 40.950 313.950 43.050 316.050 ;
        RECT 43.950 313.950 46.050 316.050 ;
        RECT 40.950 310.950 43.050 313.050 ;
        RECT 34.950 308.250 36.750 309.150 ;
        RECT 37.950 307.950 40.050 310.050 ;
        RECT 41.400 307.050 42.450 310.950 ;
        RECT 44.400 310.050 45.450 313.950 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 34.950 304.950 37.050 307.050 ;
        RECT 38.250 305.850 39.750 306.750 ;
        RECT 40.950 304.950 43.050 307.050 ;
        RECT 44.250 305.850 46.050 306.750 ;
        RECT 32.400 302.400 36.450 303.450 ;
        RECT 40.950 302.850 43.050 303.750 ;
        RECT 31.950 277.950 34.050 280.050 ;
        RECT 28.950 274.950 31.050 277.050 ;
        RECT 29.400 271.050 30.450 274.950 ;
        RECT 32.400 274.050 33.450 277.950 ;
        RECT 35.400 274.050 36.450 302.400 ;
        RECT 43.950 301.950 46.050 304.050 ;
        RECT 40.950 292.950 43.050 295.050 ;
        RECT 31.950 271.950 34.050 274.050 ;
        RECT 34.950 271.950 37.050 274.050 ;
        RECT 28.950 268.950 31.050 271.050 ;
        RECT 34.950 268.950 37.050 271.050 ;
        RECT 38.250 269.250 40.050 270.150 ;
        RECT 28.950 266.850 31.050 267.750 ;
        RECT 31.950 266.250 34.050 267.150 ;
        RECT 34.950 266.850 36.750 267.750 ;
        RECT 37.950 265.950 40.050 268.050 ;
        RECT 31.950 262.950 34.050 265.050 ;
        RECT 31.950 259.950 34.050 262.050 ;
        RECT 28.950 250.950 31.050 253.050 ;
        RECT 29.400 232.050 30.450 250.950 ;
        RECT 32.400 235.050 33.450 259.950 ;
        RECT 38.400 259.050 39.450 265.950 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 41.400 241.050 42.450 292.950 ;
        RECT 44.400 253.050 45.450 301.950 ;
        RECT 47.400 267.450 48.450 337.950 ;
        RECT 56.400 337.050 57.450 379.950 ;
        RECT 58.950 377.850 60.750 378.750 ;
        RECT 61.950 376.950 64.050 379.050 ;
        RECT 65.250 377.850 66.750 378.750 ;
        RECT 67.950 378.450 70.050 379.050 ;
        RECT 71.400 378.450 72.450 385.950 ;
        RECT 67.950 377.400 72.450 378.450 ;
        RECT 67.950 376.950 70.050 377.400 ;
        RECT 61.950 374.850 64.050 375.750 ;
        RECT 73.950 344.250 76.050 345.150 ;
        RECT 61.950 340.950 64.050 343.050 ;
        RECT 64.950 341.250 66.750 342.150 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 71.250 341.250 72.750 342.150 ;
        RECT 73.950 340.950 76.050 343.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 49.950 328.950 52.050 331.050 ;
        RECT 50.400 313.050 51.450 328.950 ;
        RECT 62.400 328.050 63.450 340.950 ;
        RECT 64.950 337.950 67.050 340.050 ;
        RECT 68.250 338.850 69.750 339.750 ;
        RECT 70.950 337.950 73.050 340.050 ;
        RECT 61.950 325.950 64.050 328.050 ;
        RECT 55.950 313.950 58.050 316.050 ;
        RECT 49.950 310.950 52.050 313.050 ;
        RECT 52.950 311.250 55.050 312.150 ;
        RECT 55.950 311.850 58.050 312.750 ;
        RECT 58.950 311.250 60.750 312.150 ;
        RECT 61.950 310.950 64.050 313.050 ;
        RECT 50.400 295.050 51.450 310.950 ;
        RECT 52.950 307.950 55.050 310.050 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 62.250 308.850 64.050 309.750 ;
        RECT 53.400 304.050 54.450 307.950 ;
        RECT 52.950 301.950 55.050 304.050 ;
        RECT 61.950 301.950 64.050 304.050 ;
        RECT 49.950 292.950 52.050 295.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 49.950 274.950 52.050 277.050 ;
        RECT 50.400 270.450 51.450 274.950 ;
        RECT 56.400 274.050 57.450 289.950 ;
        RECT 58.950 280.950 61.050 283.050 ;
        RECT 52.950 272.250 55.050 273.150 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 59.400 271.050 60.450 280.950 ;
        RECT 62.400 274.050 63.450 301.950 ;
        RECT 61.950 271.950 64.050 274.050 ;
        RECT 52.950 270.450 55.050 271.050 ;
        RECT 50.400 269.400 55.050 270.450 ;
        RECT 52.950 268.950 55.050 269.400 ;
        RECT 56.250 269.250 57.750 270.150 ;
        RECT 58.950 268.950 61.050 271.050 ;
        RECT 62.250 269.250 64.050 270.150 ;
        RECT 47.400 266.400 51.450 267.450 ;
        RECT 43.950 250.950 46.050 253.050 ;
        RECT 46.950 241.950 49.050 244.050 ;
        RECT 40.950 238.950 43.050 241.050 ;
        RECT 34.950 236.250 36.750 237.150 ;
        RECT 37.950 235.950 40.050 238.050 ;
        RECT 40.950 235.950 43.050 238.050 ;
        RECT 43.950 237.450 46.050 238.050 ;
        RECT 47.400 237.450 48.450 241.950 ;
        RECT 43.950 236.400 48.450 237.450 ;
        RECT 43.950 235.950 46.050 236.400 ;
        RECT 41.400 235.050 42.450 235.950 ;
        RECT 31.950 232.950 34.050 235.050 ;
        RECT 34.950 232.950 37.050 235.050 ;
        RECT 38.250 233.850 39.750 234.750 ;
        RECT 40.950 232.950 43.050 235.050 ;
        RECT 44.250 233.850 46.050 234.750 ;
        RECT 35.400 232.050 36.450 232.950 ;
        RECT 28.950 229.950 31.050 232.050 ;
        RECT 34.950 229.950 37.050 232.050 ;
        RECT 40.950 230.850 43.050 231.750 ;
        RECT 43.950 220.950 46.050 223.050 ;
        RECT 28.950 199.950 31.050 202.050 ;
        RECT 29.400 199.050 30.450 199.950 ;
        RECT 28.950 196.950 31.050 199.050 ;
        RECT 34.950 196.950 37.050 199.050 ;
        RECT 38.250 197.250 40.050 198.150 ;
        RECT 40.950 196.950 43.050 199.050 ;
        RECT 28.950 194.850 31.050 195.750 ;
        RECT 31.950 194.250 34.050 195.150 ;
        RECT 34.950 194.850 36.750 195.750 ;
        RECT 37.950 193.950 40.050 196.050 ;
        RECT 31.950 190.950 34.050 193.050 ;
        RECT 25.950 187.950 28.050 190.050 ;
        RECT 32.400 184.050 33.450 190.950 ;
        RECT 34.950 187.950 37.050 190.050 ;
        RECT 31.950 181.950 34.050 184.050 ;
        RECT 31.950 172.950 34.050 175.050 ;
        RECT 20.400 170.400 24.450 171.450 ;
        RECT 10.950 167.250 13.050 168.150 ;
        RECT 13.950 167.850 16.050 168.750 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 10.950 160.950 13.050 163.050 ;
        RECT 11.400 130.050 12.450 160.950 ;
        RECT 20.400 133.050 21.450 170.400 ;
        RECT 25.950 169.950 28.050 172.050 ;
        RECT 32.400 169.050 33.450 172.950 ;
        RECT 22.950 167.250 25.050 168.150 ;
        RECT 25.950 167.850 28.050 168.750 ;
        RECT 28.950 167.250 30.750 168.150 ;
        RECT 31.950 166.950 34.050 169.050 ;
        RECT 22.950 163.950 25.050 166.050 ;
        RECT 28.950 163.950 31.050 166.050 ;
        RECT 32.250 164.850 34.050 165.750 ;
        RECT 16.950 131.250 19.050 132.150 ;
        RECT 19.950 130.950 22.050 133.050 ;
        RECT 25.950 130.950 28.050 133.050 ;
        RECT 10.950 127.950 13.050 130.050 ;
        RECT 14.250 128.250 15.750 129.150 ;
        RECT 16.950 127.950 19.050 130.050 ;
        RECT 20.250 128.250 22.050 129.150 ;
        RECT 10.950 125.850 12.750 126.750 ;
        RECT 13.950 124.950 16.050 127.050 ;
        RECT 17.400 121.050 18.450 127.950 ;
        RECT 19.950 124.950 22.050 127.050 ;
        RECT 16.950 118.950 19.050 121.050 ;
        RECT 20.400 109.050 21.450 124.950 ;
        RECT 19.950 106.950 22.050 109.050 ;
        RECT 22.950 97.950 25.050 100.050 ;
        RECT 16.950 94.950 19.050 97.050 ;
        RECT 7.950 91.950 10.050 94.050 ;
        RECT 10.950 92.250 12.750 93.150 ;
        RECT 13.950 91.950 16.050 94.050 ;
        RECT 17.400 91.050 18.450 94.950 ;
        RECT 19.950 93.450 22.050 94.050 ;
        RECT 23.400 93.450 24.450 97.950 ;
        RECT 19.950 92.400 24.450 93.450 ;
        RECT 19.950 91.950 22.050 92.400 ;
        RECT 4.950 88.950 7.050 91.050 ;
        RECT 10.950 88.950 13.050 91.050 ;
        RECT 14.250 89.850 15.750 90.750 ;
        RECT 16.950 88.950 19.050 91.050 ;
        RECT 20.250 89.850 22.050 90.750 ;
        RECT 23.400 88.050 24.450 92.400 ;
        RECT 10.950 85.950 13.050 88.050 ;
        RECT 16.950 86.850 19.050 87.750 ;
        RECT 22.950 85.950 25.050 88.050 ;
        RECT 11.400 58.050 12.450 85.950 ;
        RECT 22.950 79.950 25.050 82.050 ;
        RECT 16.950 59.250 19.050 60.150 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 14.250 56.250 15.750 57.150 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 20.250 56.250 22.050 57.150 ;
        RECT 10.950 53.850 12.750 54.750 ;
        RECT 13.950 52.950 16.050 55.050 ;
        RECT 17.400 52.050 18.450 55.950 ;
        RECT 19.950 54.450 22.050 55.050 ;
        RECT 23.400 54.450 24.450 79.950 ;
        RECT 19.950 53.400 24.450 54.450 ;
        RECT 19.950 52.950 22.050 53.400 ;
        RECT 16.950 49.950 19.050 52.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 14.400 22.050 15.450 22.950 ;
        RECT 17.400 22.050 18.450 49.950 ;
        RECT 22.950 25.950 25.050 28.050 ;
        RECT 10.950 20.250 12.750 21.150 ;
        RECT 13.950 19.950 16.050 22.050 ;
        RECT 16.950 19.950 19.050 22.050 ;
        RECT 19.950 19.950 22.050 22.050 ;
        RECT 23.400 19.050 24.450 25.950 ;
        RECT 26.400 25.050 27.450 130.950 ;
        RECT 35.400 130.050 36.450 187.950 ;
        RECT 41.400 187.050 42.450 196.950 ;
        RECT 40.950 184.950 43.050 187.050 ;
        RECT 44.400 175.050 45.450 220.950 ;
        RECT 47.400 220.050 48.450 236.400 ;
        RECT 46.950 217.950 49.050 220.050 ;
        RECT 46.950 211.950 49.050 214.050 ;
        RECT 47.400 190.050 48.450 211.950 ;
        RECT 46.950 187.950 49.050 190.050 ;
        RECT 43.950 172.950 46.050 175.050 ;
        RECT 50.400 169.050 51.450 266.400 ;
        RECT 52.950 265.950 55.050 268.050 ;
        RECT 55.950 265.950 58.050 268.050 ;
        RECT 59.250 266.850 60.750 267.750 ;
        RECT 61.950 265.950 64.050 268.050 ;
        RECT 53.400 259.050 54.450 265.950 ;
        RECT 62.400 265.050 63.450 265.950 ;
        RECT 61.950 262.950 64.050 265.050 ;
        RECT 61.950 259.950 64.050 262.050 ;
        RECT 52.950 256.950 55.050 259.050 ;
        RECT 55.950 241.950 58.050 244.050 ;
        RECT 62.400 241.050 63.450 259.950 ;
        RECT 52.950 239.250 55.050 240.150 ;
        RECT 55.950 239.850 58.050 240.750 ;
        RECT 58.950 239.250 60.750 240.150 ;
        RECT 61.950 238.950 64.050 241.050 ;
        RECT 52.950 235.950 55.050 238.050 ;
        RECT 55.950 235.950 58.050 238.050 ;
        RECT 58.950 235.950 61.050 238.050 ;
        RECT 62.250 236.850 64.050 237.750 ;
        RECT 53.400 232.050 54.450 235.950 ;
        RECT 52.950 229.950 55.050 232.050 ;
        RECT 56.400 229.050 57.450 235.950 ;
        RECT 59.400 235.050 60.450 235.950 ;
        RECT 58.950 232.950 61.050 235.050 ;
        RECT 55.950 226.950 58.050 229.050 ;
        RECT 59.400 223.050 60.450 232.950 ;
        RECT 58.950 220.950 61.050 223.050 ;
        RECT 52.950 217.950 55.050 220.050 ;
        RECT 53.400 202.050 54.450 217.950 ;
        RECT 58.950 203.250 61.050 204.150 ;
        RECT 52.950 199.950 55.050 202.050 ;
        RECT 56.250 200.250 57.750 201.150 ;
        RECT 58.950 199.950 61.050 202.050 ;
        RECT 62.250 200.250 64.050 201.150 ;
        RECT 59.400 199.050 60.450 199.950 ;
        RECT 52.950 197.850 54.750 198.750 ;
        RECT 55.950 196.950 58.050 199.050 ;
        RECT 58.950 196.950 61.050 199.050 ;
        RECT 61.950 196.950 64.050 199.050 ;
        RECT 56.400 193.050 57.450 196.950 ;
        RECT 55.950 190.950 58.050 193.050 ;
        RECT 55.950 187.950 58.050 190.050 ;
        RECT 43.950 168.450 46.050 169.050 ;
        RECT 41.400 167.400 46.050 168.450 ;
        RECT 41.400 166.050 42.450 167.400 ;
        RECT 43.950 166.950 46.050 167.400 ;
        RECT 47.250 167.250 48.750 168.150 ;
        RECT 49.950 166.950 52.050 169.050 ;
        RECT 52.950 166.950 55.050 169.050 ;
        RECT 53.400 166.050 54.450 166.950 ;
        RECT 56.400 166.050 57.450 187.950 ;
        RECT 59.400 169.050 60.450 196.950 ;
        RECT 58.950 166.950 61.050 169.050 ;
        RECT 40.950 163.950 43.050 166.050 ;
        RECT 43.950 164.850 45.750 165.750 ;
        RECT 46.950 163.950 49.050 166.050 ;
        RECT 50.250 164.850 51.750 165.750 ;
        RECT 52.950 163.950 55.050 166.050 ;
        RECT 55.950 163.950 58.050 166.050 ;
        RECT 34.950 127.950 37.050 130.050 ;
        RECT 35.400 127.050 36.450 127.950 ;
        RECT 28.950 124.950 31.050 127.050 ;
        RECT 34.950 124.950 37.050 127.050 ;
        RECT 38.250 125.250 40.050 126.150 ;
        RECT 28.950 122.850 31.050 123.750 ;
        RECT 31.950 122.250 34.050 123.150 ;
        RECT 34.950 122.850 36.750 123.750 ;
        RECT 37.950 121.950 40.050 124.050 ;
        RECT 41.400 121.050 42.450 163.950 ;
        RECT 47.400 163.050 48.450 163.950 ;
        RECT 46.950 160.950 49.050 163.050 ;
        RECT 52.950 161.850 55.050 162.750 ;
        RECT 47.400 124.050 48.450 160.950 ;
        RECT 59.400 154.050 60.450 166.950 ;
        RECT 62.400 154.050 63.450 196.950 ;
        RECT 65.400 196.050 66.450 337.950 ;
        RECT 71.400 337.050 72.450 337.950 ;
        RECT 74.400 337.050 75.450 340.950 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 77.400 334.050 78.450 431.400 ;
        RECT 92.400 420.450 93.450 454.950 ;
        RECT 110.400 454.050 111.450 553.950 ;
        RECT 116.400 553.050 117.450 554.400 ;
        RECT 118.950 553.950 121.050 554.400 ;
        RECT 124.950 553.950 127.050 556.050 ;
        RECT 133.950 553.950 136.050 556.050 ;
        RECT 115.950 550.950 118.050 553.050 ;
        RECT 116.400 526.050 117.450 550.950 ;
        RECT 133.950 535.950 136.050 538.050 ;
        RECT 134.400 526.050 135.450 535.950 ;
        RECT 137.400 529.050 138.450 598.950 ;
        RECT 145.950 595.950 148.050 598.050 ;
        RECT 146.400 595.050 147.450 595.950 ;
        RECT 145.950 592.950 148.050 595.050 ;
        RECT 152.400 565.050 153.450 670.950 ;
        RECT 154.950 667.950 157.050 670.050 ;
        RECT 161.400 667.050 162.450 674.400 ;
        RECT 160.950 664.950 163.050 667.050 ;
        RECT 164.400 664.050 165.450 730.950 ;
        RECT 166.950 702.450 169.050 703.050 ;
        RECT 170.400 702.450 171.450 763.950 ;
        RECT 172.950 760.950 175.050 763.050 ;
        RECT 173.400 735.450 174.450 760.950 ;
        RECT 176.400 745.050 177.450 773.400 ;
        RECT 179.400 745.050 180.450 806.400 ;
        RECT 187.950 805.950 190.050 808.050 ;
        RECT 188.400 778.050 189.450 805.950 ;
        RECT 193.950 779.250 196.050 780.150 ;
        RECT 187.950 775.950 190.050 778.050 ;
        RECT 191.250 776.250 192.750 777.150 ;
        RECT 193.950 775.950 196.050 778.050 ;
        RECT 197.250 776.250 199.050 777.150 ;
        RECT 187.950 773.850 189.750 774.750 ;
        RECT 190.950 772.950 193.050 775.050 ;
        RECT 191.400 766.050 192.450 772.950 ;
        RECT 190.950 763.950 193.050 766.050 ;
        RECT 194.400 748.050 195.450 775.950 ;
        RECT 196.950 772.950 199.050 775.050 ;
        RECT 197.400 769.050 198.450 772.950 ;
        RECT 200.400 772.050 201.450 847.950 ;
        RECT 202.950 845.250 205.050 846.150 ;
        RECT 205.950 845.850 208.050 846.750 ;
        RECT 209.400 844.050 210.450 848.400 ;
        RECT 223.950 847.950 226.050 850.050 ;
        RECT 227.250 848.250 228.750 849.150 ;
        RECT 229.950 847.950 232.050 850.050 ;
        RECT 233.250 848.250 235.050 849.150 ;
        RECT 244.950 847.950 247.050 850.050 ;
        RECT 268.950 849.450 271.050 850.050 ;
        RECT 266.400 848.400 271.050 849.450 ;
        RECT 211.950 845.250 214.050 846.150 ;
        RECT 223.950 845.850 225.750 846.750 ;
        RECT 226.950 844.950 229.050 847.050 ;
        RECT 202.950 841.950 205.050 844.050 ;
        RECT 205.950 841.950 208.050 844.050 ;
        RECT 208.950 841.950 211.050 844.050 ;
        RECT 211.950 841.950 214.050 844.050 ;
        RECT 203.400 838.050 204.450 841.950 ;
        RECT 202.950 835.950 205.050 838.050 ;
        RECT 206.400 826.050 207.450 841.950 ;
        RECT 212.400 841.050 213.450 841.950 ;
        RECT 230.400 841.050 231.450 847.950 ;
        RECT 232.950 844.950 235.050 847.050 ;
        RECT 233.400 844.050 234.450 844.950 ;
        RECT 232.950 841.950 235.050 844.050 ;
        RECT 211.950 838.950 214.050 841.050 ;
        RECT 229.950 838.950 232.050 841.050 ;
        RECT 208.950 829.950 211.050 832.050 ;
        RECT 205.950 823.950 208.050 826.050 ;
        RECT 206.400 817.050 207.450 823.950 ;
        RECT 209.400 820.050 210.450 829.950 ;
        RECT 208.950 817.950 211.050 820.050 ;
        RECT 212.400 817.050 213.450 838.950 ;
        RECT 245.400 823.050 246.450 847.950 ;
        RECT 247.950 845.250 249.750 846.150 ;
        RECT 250.950 844.950 253.050 847.050 ;
        RECT 256.950 846.450 259.050 847.050 ;
        RECT 256.950 845.400 261.450 846.450 ;
        RECT 256.950 844.950 259.050 845.400 ;
        RECT 260.400 844.050 261.450 845.400 ;
        RECT 262.950 844.950 265.050 847.050 ;
        RECT 247.950 841.950 250.050 844.050 ;
        RECT 251.250 842.850 253.050 843.750 ;
        RECT 253.950 842.250 256.050 843.150 ;
        RECT 256.950 842.850 259.050 843.750 ;
        RECT 259.950 841.950 262.050 844.050 ;
        RECT 241.950 820.950 244.050 823.050 ;
        RECT 244.950 820.950 247.050 823.050 ;
        RECT 202.950 814.950 205.050 817.050 ;
        RECT 205.950 814.950 208.050 817.050 ;
        RECT 209.250 815.850 210.750 816.750 ;
        RECT 211.950 814.950 214.050 817.050 ;
        RECT 232.950 814.950 235.050 817.050 ;
        RECT 238.950 814.950 241.050 817.050 ;
        RECT 203.400 775.050 204.450 814.950 ;
        RECT 205.950 812.850 208.050 813.750 ;
        RECT 211.950 812.850 214.050 813.750 ;
        RECT 226.950 812.250 228.750 813.150 ;
        RECT 229.950 811.950 232.050 814.050 ;
        RECT 233.400 811.050 234.450 814.950 ;
        RECT 235.950 813.450 238.050 814.050 ;
        RECT 239.400 813.450 240.450 814.950 ;
        RECT 235.950 812.400 240.450 813.450 ;
        RECT 235.950 811.950 238.050 812.400 ;
        RECT 226.950 808.950 229.050 811.050 ;
        RECT 230.250 809.850 231.750 810.750 ;
        RECT 232.950 808.950 235.050 811.050 ;
        RECT 236.250 809.850 238.050 810.750 ;
        RECT 227.400 777.450 228.450 808.950 ;
        RECT 229.950 805.950 232.050 808.050 ;
        RECT 232.950 806.850 235.050 807.750 ;
        RECT 211.950 776.250 214.050 777.150 ;
        RECT 224.400 776.400 228.450 777.450 ;
        RECT 202.950 772.950 205.050 775.050 ;
        RECT 211.950 772.950 214.050 775.050 ;
        RECT 215.250 773.250 216.750 774.150 ;
        RECT 217.950 772.950 220.050 775.050 ;
        RECT 221.250 773.250 223.050 774.150 ;
        RECT 199.950 769.950 202.050 772.050 ;
        RECT 196.950 766.950 199.050 769.050 ;
        RECT 202.950 766.950 205.050 769.050 ;
        RECT 184.950 745.950 187.050 748.050 ;
        RECT 193.950 745.950 196.050 748.050 ;
        RECT 199.950 745.950 202.050 748.050 ;
        RECT 185.400 745.050 186.450 745.950 ;
        RECT 175.950 742.950 178.050 745.050 ;
        RECT 178.950 742.950 181.050 745.050 ;
        RECT 182.250 743.250 183.750 744.150 ;
        RECT 184.950 742.950 187.050 745.050 ;
        RECT 176.400 742.050 177.450 742.950 ;
        RECT 175.950 739.950 178.050 742.050 ;
        RECT 179.250 740.850 180.750 741.750 ;
        RECT 181.950 739.950 184.050 742.050 ;
        RECT 185.250 740.850 187.050 741.750 ;
        RECT 175.950 737.850 178.050 738.750 ;
        RECT 173.400 734.400 177.450 735.450 ;
        RECT 166.950 701.400 171.450 702.450 ;
        RECT 166.950 700.950 169.050 701.400 ;
        RECT 172.950 700.950 175.050 703.050 ;
        RECT 166.950 698.850 169.050 699.750 ;
        RECT 169.950 698.250 172.050 699.150 ;
        RECT 169.950 694.950 172.050 697.050 ;
        RECT 173.400 670.050 174.450 700.950 ;
        RECT 176.400 676.050 177.450 734.400 ;
        RECT 194.400 718.050 195.450 745.950 ;
        RECT 196.950 743.250 199.050 744.150 ;
        RECT 199.950 743.850 202.050 744.750 ;
        RECT 196.950 739.950 199.050 742.050 ;
        RECT 193.950 715.950 196.050 718.050 ;
        RECT 203.400 712.050 204.450 766.950 ;
        RECT 212.400 754.050 213.450 772.950 ;
        RECT 214.950 769.950 217.050 772.050 ;
        RECT 218.250 770.850 219.750 771.750 ;
        RECT 220.950 769.950 223.050 772.050 ;
        RECT 211.950 751.950 214.050 754.050 ;
        RECT 208.950 739.950 211.050 742.050 ;
        RECT 211.950 740.250 213.750 741.150 ;
        RECT 214.950 739.950 217.050 742.050 ;
        RECT 218.250 740.250 220.050 741.150 ;
        RECT 202.950 709.950 205.050 712.050 ;
        RECT 209.400 708.450 210.450 739.950 ;
        RECT 211.950 736.950 214.050 739.050 ;
        RECT 215.250 737.850 216.750 738.750 ;
        RECT 217.950 736.950 220.050 739.050 ;
        RECT 212.400 736.050 213.450 736.950 ;
        RECT 211.950 733.950 214.050 736.050 ;
        RECT 221.400 733.050 222.450 769.950 ;
        RECT 224.400 739.050 225.450 776.400 ;
        RECT 226.950 772.950 229.050 775.050 ;
        RECT 223.950 736.950 226.050 739.050 ;
        RECT 220.950 730.950 223.050 733.050 ;
        RECT 209.400 707.400 213.450 708.450 ;
        RECT 181.950 704.250 184.050 705.150 ;
        RECT 208.950 704.250 211.050 705.150 ;
        RECT 181.950 700.950 184.050 703.050 ;
        RECT 185.250 701.250 186.750 702.150 ;
        RECT 187.950 700.950 190.050 703.050 ;
        RECT 191.250 701.250 193.050 702.150 ;
        RECT 199.950 701.250 201.750 702.150 ;
        RECT 202.950 700.950 205.050 703.050 ;
        RECT 206.250 701.250 207.750 702.150 ;
        RECT 208.950 700.950 211.050 703.050 ;
        RECT 184.950 697.950 187.050 700.050 ;
        RECT 188.250 698.850 189.750 699.750 ;
        RECT 190.950 697.950 193.050 700.050 ;
        RECT 199.950 697.950 202.050 700.050 ;
        RECT 203.250 698.850 204.750 699.750 ;
        RECT 205.950 697.950 208.050 700.050 ;
        RECT 181.950 694.950 184.050 697.050 ;
        RECT 187.950 694.950 190.050 697.050 ;
        RECT 175.950 673.950 178.050 676.050 ;
        RECT 175.950 670.950 178.050 673.050 ;
        RECT 169.950 668.250 171.750 669.150 ;
        RECT 172.950 667.950 175.050 670.050 ;
        RECT 176.400 667.050 177.450 670.950 ;
        RECT 178.950 667.950 181.050 670.050 ;
        RECT 169.950 664.950 172.050 667.050 ;
        RECT 173.250 665.850 174.750 666.750 ;
        RECT 175.950 664.950 178.050 667.050 ;
        RECT 179.250 665.850 181.050 666.750 ;
        RECT 163.950 661.950 166.050 664.050 ;
        RECT 154.950 631.950 157.050 634.050 ;
        RECT 155.400 597.450 156.450 631.950 ;
        RECT 170.400 631.050 171.450 664.950 ;
        RECT 172.950 661.950 175.050 664.050 ;
        RECT 175.950 662.850 178.050 663.750 ;
        RECT 157.950 629.250 159.750 630.150 ;
        RECT 160.950 628.950 163.050 631.050 ;
        RECT 166.950 630.450 169.050 631.050 ;
        RECT 169.950 630.450 172.050 631.050 ;
        RECT 166.950 629.400 172.050 630.450 ;
        RECT 166.950 628.950 169.050 629.400 ;
        RECT 169.950 628.950 172.050 629.400 ;
        RECT 157.950 625.950 160.050 628.050 ;
        RECT 161.250 626.850 163.050 627.750 ;
        RECT 163.950 626.250 166.050 627.150 ;
        RECT 166.950 626.850 169.050 627.750 ;
        RECT 158.400 625.050 159.450 625.950 ;
        RECT 157.950 622.950 160.050 625.050 ;
        RECT 163.950 622.950 166.050 625.050 ;
        RECT 164.400 619.050 165.450 622.950 ;
        RECT 163.950 616.950 166.050 619.050 ;
        RECT 163.950 601.950 166.050 604.050 ;
        RECT 164.400 598.050 165.450 601.950 ;
        RECT 157.950 597.450 160.050 598.050 ;
        RECT 155.400 596.400 160.050 597.450 ;
        RECT 157.950 595.950 160.050 596.400 ;
        RECT 163.950 595.950 166.050 598.050 ;
        RECT 167.250 596.250 169.050 597.150 ;
        RECT 157.950 593.850 159.750 594.750 ;
        RECT 160.950 592.950 163.050 595.050 ;
        RECT 164.250 593.850 165.750 594.750 ;
        RECT 166.950 592.950 169.050 595.050 ;
        RECT 160.950 590.850 163.050 591.750 ;
        RECT 163.950 577.950 166.050 580.050 ;
        RECT 160.950 571.950 163.050 574.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 142.950 562.950 145.050 565.050 ;
        RECT 151.950 562.950 154.050 565.050 ;
        RECT 143.400 532.050 144.450 562.950 ;
        RECT 148.950 559.950 151.050 562.050 ;
        RECT 149.400 559.050 150.450 559.950 ;
        RECT 155.400 559.050 156.450 568.950 ;
        RECT 145.950 557.250 147.750 558.150 ;
        RECT 148.950 556.950 151.050 559.050 ;
        RECT 152.250 557.250 153.750 558.150 ;
        RECT 154.950 556.950 157.050 559.050 ;
        RECT 158.250 557.250 160.050 558.150 ;
        RECT 145.950 553.950 148.050 556.050 ;
        RECT 149.250 554.850 150.750 555.750 ;
        RECT 151.950 553.950 154.050 556.050 ;
        RECT 155.250 554.850 156.750 555.750 ;
        RECT 157.950 555.450 160.050 556.050 ;
        RECT 161.400 555.450 162.450 571.950 ;
        RECT 157.950 554.400 162.450 555.450 ;
        RECT 157.950 553.950 160.050 554.400 ;
        RECT 146.400 538.050 147.450 553.950 ;
        RECT 164.400 553.050 165.450 577.950 ;
        RECT 167.400 565.050 168.450 592.950 ;
        RECT 173.400 592.050 174.450 661.950 ;
        RECT 175.950 634.950 178.050 637.050 ;
        RECT 182.400 636.450 183.450 694.950 ;
        RECT 188.400 640.050 189.450 694.950 ;
        RECT 191.400 682.050 192.450 697.950 ;
        RECT 200.400 696.450 201.450 697.950 ;
        RECT 206.400 697.050 207.450 697.950 ;
        RECT 200.400 695.400 204.450 696.450 ;
        RECT 196.950 691.950 199.050 694.050 ;
        RECT 190.950 679.950 193.050 682.050 ;
        RECT 197.400 676.050 198.450 691.950 ;
        RECT 190.950 673.950 193.050 676.050 ;
        RECT 196.950 673.950 199.050 676.050 ;
        RECT 191.400 673.050 192.450 673.950 ;
        RECT 190.950 670.950 193.050 673.050 ;
        RECT 194.250 671.250 196.050 672.150 ;
        RECT 196.950 671.850 199.050 672.750 ;
        RECT 199.950 671.250 202.050 672.150 ;
        RECT 190.950 668.850 192.750 669.750 ;
        RECT 193.950 667.950 196.050 670.050 ;
        RECT 199.950 667.950 202.050 670.050 ;
        RECT 194.400 667.050 195.450 667.950 ;
        RECT 203.400 667.050 204.450 695.400 ;
        RECT 205.950 694.950 208.050 697.050 ;
        RECT 205.950 685.950 208.050 688.050 ;
        RECT 193.950 664.950 196.050 667.050 ;
        RECT 202.950 664.950 205.050 667.050 ;
        RECT 203.400 655.050 204.450 664.950 ;
        RECT 202.950 652.950 205.050 655.050 ;
        RECT 187.950 637.950 190.050 640.050 ;
        RECT 193.950 637.950 196.050 640.050 ;
        RECT 196.950 637.950 199.050 640.050 ;
        RECT 179.400 635.400 183.450 636.450 ;
        RECT 176.400 600.450 177.450 634.950 ;
        RECT 179.400 625.050 180.450 635.400 ;
        RECT 187.950 635.250 190.050 636.150 ;
        RECT 194.400 634.050 195.450 637.950 ;
        RECT 181.950 631.950 184.050 634.050 ;
        RECT 185.250 632.250 186.750 633.150 ;
        RECT 187.950 631.950 190.050 634.050 ;
        RECT 191.250 632.250 193.050 633.150 ;
        RECT 193.950 631.950 196.050 634.050 ;
        RECT 181.950 629.850 183.750 630.750 ;
        RECT 184.950 628.950 187.050 631.050 ;
        RECT 178.950 622.950 181.050 625.050 ;
        RECT 188.400 619.050 189.450 631.950 ;
        RECT 190.950 630.450 193.050 631.050 ;
        RECT 190.950 629.400 195.450 630.450 ;
        RECT 190.950 628.950 193.050 629.400 ;
        RECT 191.400 628.050 192.450 628.950 ;
        RECT 190.950 625.950 193.050 628.050 ;
        RECT 187.950 616.950 190.050 619.050 ;
        RECT 184.950 610.950 187.050 613.050 ;
        RECT 185.400 601.050 186.450 610.950 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 191.400 601.050 192.450 601.950 ;
        RECT 178.950 600.450 181.050 601.050 ;
        RECT 176.400 599.400 181.050 600.450 ;
        RECT 172.950 589.950 175.050 592.050 ;
        RECT 176.400 574.050 177.450 599.400 ;
        RECT 178.950 598.950 181.050 599.400 ;
        RECT 182.250 599.250 183.750 600.150 ;
        RECT 184.950 598.950 187.050 601.050 ;
        RECT 188.250 599.250 189.750 600.150 ;
        RECT 190.950 598.950 193.050 601.050 ;
        RECT 178.950 596.850 180.750 597.750 ;
        RECT 181.950 595.950 184.050 598.050 ;
        RECT 185.250 596.850 186.750 597.750 ;
        RECT 187.950 595.950 190.050 598.050 ;
        RECT 191.250 596.850 193.050 597.750 ;
        RECT 182.400 595.050 183.450 595.950 ;
        RECT 181.950 592.950 184.050 595.050 ;
        RECT 175.950 571.950 178.050 574.050 ;
        RECT 182.400 571.050 183.450 592.950 ;
        RECT 188.400 580.050 189.450 595.950 ;
        RECT 194.400 586.050 195.450 629.400 ;
        RECT 197.400 595.050 198.450 637.950 ;
        RECT 206.400 637.050 207.450 685.950 ;
        RECT 209.400 682.050 210.450 700.950 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 212.400 675.450 213.450 707.400 ;
        RECT 214.950 706.950 217.050 709.050 ;
        RECT 215.400 688.050 216.450 706.950 ;
        RECT 223.950 700.950 226.050 703.050 ;
        RECT 220.950 698.250 223.050 699.150 ;
        RECT 223.950 698.850 226.050 699.750 ;
        RECT 227.400 697.050 228.450 772.950 ;
        RECT 230.400 772.050 231.450 805.950 ;
        RECT 239.400 793.050 240.450 812.400 ;
        RECT 232.950 790.950 235.050 793.050 ;
        RECT 238.950 790.950 241.050 793.050 ;
        RECT 233.400 775.050 234.450 790.950 ;
        RECT 232.950 772.950 235.050 775.050 ;
        RECT 242.400 774.450 243.450 820.950 ;
        RECT 248.400 820.050 249.450 841.950 ;
        RECT 253.950 838.950 256.050 841.050 ;
        RECT 253.950 820.950 256.050 823.050 ;
        RECT 247.950 817.950 250.050 820.050 ;
        RECT 244.950 814.950 247.050 817.050 ;
        RECT 248.250 815.250 249.750 816.150 ;
        RECT 250.950 814.950 253.050 817.050 ;
        RECT 254.400 814.050 255.450 820.950 ;
        RECT 260.400 820.050 261.450 841.950 ;
        RECT 259.950 817.950 262.050 820.050 ;
        RECT 244.950 812.850 246.750 813.750 ;
        RECT 247.950 811.950 250.050 814.050 ;
        RECT 251.250 812.850 252.750 813.750 ;
        RECT 253.950 811.950 256.050 814.050 ;
        RECT 253.950 809.850 256.050 810.750 ;
        RECT 247.950 776.250 250.050 777.150 ;
        RECT 253.950 775.950 256.050 778.050 ;
        RECT 254.400 775.050 255.450 775.950 ;
        RECT 263.400 775.050 264.450 844.950 ;
        RECT 266.400 841.050 267.450 848.400 ;
        RECT 268.950 847.950 271.050 848.400 ;
        RECT 272.250 848.250 273.750 849.150 ;
        RECT 274.950 847.950 277.050 850.050 ;
        RECT 278.250 848.250 280.050 849.150 ;
        RECT 289.950 847.950 292.050 850.050 ;
        RECT 304.950 848.250 307.050 849.150 ;
        RECT 310.950 847.950 313.050 850.050 ;
        RECT 316.950 847.950 319.050 850.050 ;
        RECT 331.950 848.250 334.050 849.150 ;
        RECT 355.950 847.950 358.050 850.050 ;
        RECT 367.950 847.950 370.050 850.050 ;
        RECT 373.950 849.450 376.050 850.050 ;
        RECT 385.950 849.450 388.050 850.050 ;
        RECT 371.250 848.250 372.750 849.150 ;
        RECT 373.950 848.400 378.450 849.450 ;
        RECT 373.950 847.950 376.050 848.400 ;
        RECT 268.950 845.850 270.750 846.750 ;
        RECT 271.950 844.950 274.050 847.050 ;
        RECT 265.950 838.950 268.050 841.050 ;
        RECT 272.400 835.050 273.450 844.950 ;
        RECT 275.400 843.450 276.450 847.950 ;
        RECT 290.400 847.050 291.450 847.950 ;
        RECT 311.400 847.050 312.450 847.950 ;
        RECT 277.950 846.450 280.050 847.050 ;
        RECT 277.950 845.400 282.450 846.450 ;
        RECT 277.950 844.950 280.050 845.400 ;
        RECT 281.400 844.050 282.450 845.400 ;
        RECT 289.950 844.950 292.050 847.050 ;
        RECT 304.950 844.950 307.050 847.050 ;
        RECT 308.250 845.250 309.750 846.150 ;
        RECT 310.950 844.950 313.050 847.050 ;
        RECT 314.250 845.250 316.050 846.150 ;
        RECT 275.400 842.400 279.450 843.450 ;
        RECT 278.400 841.050 279.450 842.400 ;
        RECT 280.950 841.950 283.050 844.050 ;
        RECT 286.950 842.250 289.050 843.150 ;
        RECT 289.950 842.850 292.050 843.750 ;
        RECT 307.950 841.950 310.050 844.050 ;
        RECT 311.250 842.850 312.750 843.750 ;
        RECT 313.950 841.950 316.050 844.050 ;
        RECT 274.950 838.950 277.050 841.050 ;
        RECT 277.950 838.950 280.050 841.050 ;
        RECT 286.950 838.950 289.050 841.050 ;
        RECT 271.950 832.950 274.050 835.050 ;
        RECT 265.950 811.950 268.050 814.050 ;
        RECT 268.950 812.250 270.750 813.150 ;
        RECT 271.950 811.950 274.050 814.050 ;
        RECT 239.400 773.400 243.450 774.450 ;
        RECT 229.950 769.950 232.050 772.050 ;
        RECT 232.950 770.850 235.050 771.750 ;
        RECT 235.950 770.250 238.050 771.150 ;
        RECT 235.950 766.950 238.050 769.050 ;
        RECT 236.400 766.050 237.450 766.950 ;
        RECT 235.950 763.950 238.050 766.050 ;
        RECT 235.950 745.950 238.050 748.050 ;
        RECT 236.400 742.050 237.450 745.950 ;
        RECT 232.950 740.250 234.750 741.150 ;
        RECT 235.950 739.950 238.050 742.050 ;
        RECT 239.400 739.050 240.450 773.400 ;
        RECT 247.950 772.950 250.050 775.050 ;
        RECT 251.250 773.250 252.750 774.150 ;
        RECT 253.950 772.950 256.050 775.050 ;
        RECT 257.250 773.250 259.050 774.150 ;
        RECT 262.950 772.950 265.050 775.050 ;
        RECT 241.950 763.950 244.050 766.050 ;
        RECT 242.400 742.050 243.450 763.950 ;
        RECT 241.950 741.450 244.050 742.050 ;
        RECT 241.950 740.400 246.450 741.450 ;
        RECT 241.950 739.950 244.050 740.400 ;
        RECT 245.400 739.050 246.450 740.400 ;
        RECT 229.950 736.950 232.050 739.050 ;
        RECT 232.950 736.950 235.050 739.050 ;
        RECT 236.250 737.850 237.750 738.750 ;
        RECT 238.950 736.950 241.050 739.050 ;
        RECT 242.250 737.850 244.050 738.750 ;
        RECT 244.950 736.950 247.050 739.050 ;
        RECT 230.400 703.050 231.450 736.950 ;
        RECT 233.400 736.050 234.450 736.950 ;
        RECT 232.950 733.950 235.050 736.050 ;
        RECT 238.950 734.850 241.050 735.750 ;
        RECT 233.400 706.050 234.450 733.950 ;
        RECT 238.950 707.250 241.050 708.150 ;
        RECT 232.950 703.950 235.050 706.050 ;
        RECT 235.950 704.250 237.750 705.150 ;
        RECT 238.950 703.950 241.050 706.050 ;
        RECT 242.250 704.250 243.750 705.150 ;
        RECT 244.950 703.950 247.050 706.050 ;
        RECT 229.950 700.950 232.050 703.050 ;
        RECT 235.950 700.950 238.050 703.050 ;
        RECT 241.950 702.450 244.050 703.050 ;
        RECT 239.400 701.400 244.050 702.450 ;
        RECT 245.250 701.850 247.050 702.750 ;
        RECT 239.400 699.450 240.450 701.400 ;
        RECT 241.950 700.950 244.050 701.400 ;
        RECT 236.400 698.400 240.450 699.450 ;
        RECT 220.950 694.950 223.050 697.050 ;
        RECT 226.950 694.950 229.050 697.050 ;
        RECT 221.400 694.050 222.450 694.950 ;
        RECT 220.950 691.950 223.050 694.050 ;
        RECT 214.950 685.950 217.050 688.050 ;
        RECT 214.950 679.950 217.050 682.050 ;
        RECT 215.400 676.050 216.450 679.950 ;
        RECT 209.400 674.400 213.450 675.450 ;
        RECT 209.400 639.450 210.450 674.400 ;
        RECT 214.950 673.950 217.050 676.050 ;
        RECT 211.950 671.250 214.050 672.150 ;
        RECT 214.950 671.850 217.050 672.750 ;
        RECT 217.950 670.950 220.050 673.050 ;
        RECT 211.950 667.950 214.050 670.050 ;
        RECT 214.950 667.950 217.050 670.050 ;
        RECT 209.400 638.400 213.450 639.450 ;
        RECT 205.950 636.450 208.050 637.050 ;
        RECT 205.950 635.400 210.450 636.450 ;
        RECT 205.950 634.950 208.050 635.400 ;
        RECT 209.400 634.050 210.450 635.400 ;
        RECT 202.950 631.950 205.050 634.050 ;
        RECT 206.250 632.250 207.750 633.150 ;
        RECT 208.950 631.950 211.050 634.050 ;
        RECT 202.950 629.850 204.750 630.750 ;
        RECT 205.950 628.950 208.050 631.050 ;
        RECT 209.250 629.850 211.050 630.750 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 199.950 601.950 202.050 604.050 ;
        RECT 196.950 592.950 199.050 595.050 ;
        RECT 196.950 589.950 199.050 592.050 ;
        RECT 193.950 583.950 196.050 586.050 ;
        RECT 187.950 577.950 190.050 580.050 ;
        RECT 193.950 574.950 196.050 577.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 166.950 562.950 169.050 565.050 ;
        RECT 175.950 562.950 178.050 565.050 ;
        RECT 187.950 563.250 190.050 564.150 ;
        RECT 166.950 559.950 169.050 562.050 ;
        RECT 170.250 560.250 171.750 561.150 ;
        RECT 172.950 559.950 175.050 562.050 ;
        RECT 166.950 557.850 168.750 558.750 ;
        RECT 169.950 556.950 172.050 559.050 ;
        RECT 173.250 557.850 175.050 558.750 ;
        RECT 170.400 556.050 171.450 556.950 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 151.950 550.950 154.050 553.050 ;
        RECT 163.950 550.950 166.050 553.050 ;
        RECT 145.950 535.950 148.050 538.050 ;
        RECT 142.950 529.950 145.050 532.050 ;
        RECT 152.400 529.050 153.450 550.950 ;
        RECT 166.950 532.950 169.050 535.050 ;
        RECT 157.950 529.950 160.050 532.050 ;
        RECT 136.950 526.950 139.050 529.050 ;
        RECT 145.950 528.450 148.050 529.050 ;
        RECT 143.400 527.400 148.050 528.450 ;
        RECT 112.950 524.250 114.750 525.150 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 119.250 524.250 121.050 525.150 ;
        RECT 130.950 524.250 132.750 525.150 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 137.250 524.250 139.050 525.150 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 116.250 521.850 117.750 522.750 ;
        RECT 118.950 520.950 121.050 523.050 ;
        RECT 130.950 520.950 133.050 523.050 ;
        RECT 134.250 521.850 135.750 522.750 ;
        RECT 136.950 520.950 139.050 523.050 ;
        RECT 113.400 484.050 114.450 520.950 ;
        RECT 119.400 520.050 120.450 520.950 ;
        RECT 118.950 517.950 121.050 520.050 ;
        RECT 131.400 517.050 132.450 520.950 ;
        RECT 133.950 517.950 136.050 520.050 ;
        RECT 121.950 514.950 124.050 517.050 ;
        RECT 130.950 514.950 133.050 517.050 ;
        RECT 112.950 481.950 115.050 484.050 ;
        RECT 122.400 483.450 123.450 514.950 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 125.400 490.050 126.450 493.950 ;
        RECT 124.950 487.950 127.050 490.050 ;
        RECT 128.250 488.250 129.750 489.150 ;
        RECT 130.950 487.950 133.050 490.050 ;
        RECT 124.950 485.850 126.750 486.750 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 131.250 485.850 133.050 486.750 ;
        RECT 122.400 482.400 126.450 483.450 ;
        RECT 115.950 454.950 118.050 457.050 ;
        RECT 119.250 455.250 120.750 456.150 ;
        RECT 121.950 454.950 124.050 457.050 ;
        RECT 125.400 454.050 126.450 482.400 ;
        RECT 128.400 475.050 129.450 484.950 ;
        RECT 130.950 478.950 133.050 481.050 ;
        RECT 127.950 472.950 130.050 475.050 ;
        RECT 127.950 463.950 130.050 466.050 ;
        RECT 94.950 452.850 96.750 453.750 ;
        RECT 97.950 451.950 100.050 454.050 ;
        RECT 101.250 452.850 102.750 453.750 ;
        RECT 109.950 451.950 112.050 454.050 ;
        RECT 112.950 451.950 115.050 454.050 ;
        RECT 115.950 452.850 117.750 453.750 ;
        RECT 118.950 451.950 121.050 454.050 ;
        RECT 122.250 452.850 123.750 453.750 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 97.950 448.950 100.050 451.050 ;
        RECT 103.950 449.850 106.050 450.750 ;
        RECT 98.400 445.050 99.450 448.950 ;
        RECT 113.400 448.050 114.450 451.950 ;
        RECT 118.950 448.950 121.050 451.050 ;
        RECT 124.950 449.850 127.050 450.750 ;
        RECT 112.950 445.950 115.050 448.050 ;
        RECT 97.950 442.950 100.050 445.050 ;
        RECT 92.400 419.400 96.450 420.450 ;
        RECT 85.950 417.450 88.050 418.050 ;
        RECT 83.400 416.400 88.050 417.450 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 80.400 403.050 81.450 412.950 ;
        RECT 83.400 412.050 84.450 416.400 ;
        RECT 85.950 415.950 88.050 416.400 ;
        RECT 89.250 416.250 90.750 417.150 ;
        RECT 91.950 415.950 94.050 418.050 ;
        RECT 85.950 413.850 87.750 414.750 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 92.250 413.850 94.050 414.750 ;
        RECT 82.950 409.950 85.050 412.050 ;
        RECT 85.950 409.950 88.050 412.050 ;
        RECT 79.950 400.950 82.050 403.050 ;
        RECT 79.950 385.950 82.050 388.050 ;
        RECT 79.950 383.850 82.050 384.750 ;
        RECT 82.950 383.250 85.050 384.150 ;
        RECT 82.950 379.950 85.050 382.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 67.950 331.950 70.050 334.050 ;
        RECT 76.950 331.950 79.050 334.050 ;
        RECT 64.950 193.950 67.050 196.050 ;
        RECT 68.400 190.050 69.450 331.950 ;
        RECT 70.950 325.950 73.050 328.050 ;
        RECT 71.400 310.050 72.450 325.950 ;
        RECT 80.400 316.050 81.450 334.950 ;
        RECT 86.400 334.050 87.450 409.950 ;
        RECT 95.400 406.050 96.450 419.400 ;
        RECT 98.400 415.050 99.450 442.950 ;
        RECT 106.950 415.950 109.050 418.050 ;
        RECT 97.950 412.950 100.050 415.050 ;
        RECT 100.950 413.250 103.050 414.150 ;
        RECT 106.950 413.850 109.050 414.750 ;
        RECT 109.950 413.250 112.050 414.150 ;
        RECT 100.950 409.950 103.050 412.050 ;
        RECT 109.950 409.950 112.050 412.050 ;
        RECT 113.400 409.050 114.450 445.950 ;
        RECT 115.950 418.950 118.050 421.050 ;
        RECT 116.400 412.050 117.450 418.950 ;
        RECT 119.400 418.050 120.450 448.950 ;
        RECT 128.400 424.050 129.450 463.950 ;
        RECT 127.950 421.950 130.050 424.050 ;
        RECT 121.950 418.950 124.050 421.050 ;
        RECT 122.400 418.050 123.450 418.950 ;
        RECT 128.400 418.050 129.450 421.950 ;
        RECT 118.950 415.950 121.050 418.050 ;
        RECT 121.950 415.950 124.050 418.050 ;
        RECT 125.250 416.250 126.750 417.150 ;
        RECT 127.950 415.950 130.050 418.050 ;
        RECT 121.950 413.850 123.750 414.750 ;
        RECT 124.950 412.950 127.050 415.050 ;
        RECT 128.250 413.850 130.050 414.750 ;
        RECT 115.950 409.950 118.050 412.050 ;
        RECT 112.950 406.950 115.050 409.050 ;
        RECT 94.950 403.950 97.050 406.050 ;
        RECT 109.950 403.950 112.050 406.050 ;
        RECT 100.950 400.950 103.050 403.050 ;
        RECT 106.950 400.950 109.050 403.050 ;
        RECT 94.950 397.950 97.050 400.050 ;
        RECT 95.400 385.050 96.450 397.950 ;
        RECT 97.950 385.950 100.050 388.050 ;
        RECT 101.400 385.050 102.450 400.950 ;
        RECT 94.950 382.950 97.050 385.050 ;
        RECT 98.250 383.850 99.750 384.750 ;
        RECT 100.950 382.950 103.050 385.050 ;
        RECT 94.950 380.850 97.050 381.750 ;
        RECT 100.950 380.850 103.050 381.750 ;
        RECT 88.950 344.250 91.050 345.150 ;
        RECT 100.950 343.950 103.050 346.050 ;
        RECT 88.950 340.950 91.050 343.050 ;
        RECT 92.250 341.250 93.750 342.150 ;
        RECT 94.950 340.950 97.050 343.050 ;
        RECT 98.250 341.250 100.050 342.150 ;
        RECT 85.950 331.950 88.050 334.050 ;
        RECT 89.400 331.050 90.450 340.950 ;
        RECT 91.950 337.950 94.050 340.050 ;
        RECT 95.250 338.850 96.750 339.750 ;
        RECT 97.950 339.450 100.050 340.050 ;
        RECT 101.400 339.450 102.450 343.950 ;
        RECT 97.950 338.400 102.450 339.450 ;
        RECT 97.950 337.950 100.050 338.400 ;
        RECT 92.400 331.050 93.450 337.950 ;
        RECT 98.400 337.050 99.450 337.950 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 94.950 331.950 97.050 334.050 ;
        RECT 88.950 328.950 91.050 331.050 ;
        RECT 91.950 328.950 94.050 331.050 ;
        RECT 85.950 319.950 88.050 322.050 ;
        RECT 79.950 313.950 82.050 316.050 ;
        RECT 76.950 311.250 79.050 312.150 ;
        RECT 79.950 311.850 82.050 312.750 ;
        RECT 70.950 307.950 73.050 310.050 ;
        RECT 76.950 307.950 79.050 310.050 ;
        RECT 71.400 262.050 72.450 307.950 ;
        RECT 77.400 307.050 78.450 307.950 ;
        RECT 76.950 304.950 79.050 307.050 ;
        RECT 76.950 280.950 79.050 283.050 ;
        RECT 77.400 277.050 78.450 280.950 ;
        RECT 73.950 274.950 76.050 277.050 ;
        RECT 76.950 274.950 79.050 277.050 ;
        RECT 79.950 275.250 82.050 276.150 ;
        RECT 74.400 274.050 75.450 274.950 ;
        RECT 73.950 271.950 76.050 274.050 ;
        RECT 77.250 272.250 78.750 273.150 ;
        RECT 79.950 271.950 82.050 274.050 ;
        RECT 83.250 272.250 85.050 273.150 ;
        RECT 73.950 269.850 75.750 270.750 ;
        RECT 76.950 268.950 79.050 271.050 ;
        RECT 77.400 262.050 78.450 268.950 ;
        RECT 70.950 259.950 73.050 262.050 ;
        RECT 76.950 261.450 79.050 262.050 ;
        RECT 74.400 260.400 79.050 261.450 ;
        RECT 74.400 238.050 75.450 260.400 ;
        RECT 76.950 259.950 79.050 260.400 ;
        RECT 76.950 256.950 79.050 259.050 ;
        RECT 77.400 241.050 78.450 256.950 ;
        RECT 80.400 243.450 81.450 271.950 ;
        RECT 82.950 268.950 85.050 271.050 ;
        RECT 82.950 265.950 85.050 268.050 ;
        RECT 83.400 259.050 84.450 265.950 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 86.400 247.050 87.450 319.950 ;
        RECT 95.400 313.050 96.450 331.950 ;
        RECT 91.950 310.950 94.050 313.050 ;
        RECT 94.950 310.950 97.050 313.050 ;
        RECT 98.250 311.250 99.750 312.150 ;
        RECT 100.950 310.950 103.050 313.050 ;
        RECT 92.400 310.050 93.450 310.950 ;
        RECT 91.950 307.950 94.050 310.050 ;
        RECT 95.250 308.850 96.750 309.750 ;
        RECT 97.950 307.950 100.050 310.050 ;
        RECT 101.250 308.850 103.050 309.750 ;
        RECT 91.950 305.850 94.050 306.750 ;
        RECT 98.400 292.050 99.450 307.950 ;
        RECT 107.400 304.050 108.450 400.950 ;
        RECT 110.400 382.050 111.450 403.950 ;
        RECT 131.400 403.050 132.450 478.950 ;
        RECT 134.400 421.050 135.450 517.950 ;
        RECT 137.400 490.050 138.450 520.950 ;
        RECT 136.950 487.950 139.050 490.050 ;
        RECT 136.950 481.950 139.050 484.050 ;
        RECT 137.400 457.050 138.450 481.950 ;
        RECT 140.400 475.050 141.450 523.950 ;
        RECT 143.400 517.050 144.450 527.400 ;
        RECT 145.950 526.950 148.050 527.400 ;
        RECT 149.250 527.250 150.750 528.150 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 145.950 524.850 147.750 525.750 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 152.250 524.850 153.750 525.750 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 154.950 521.850 157.050 522.750 ;
        RECT 142.950 514.950 145.050 517.050 ;
        RECT 148.950 491.250 151.050 492.150 ;
        RECT 142.950 487.950 145.050 490.050 ;
        RECT 146.250 488.250 147.750 489.150 ;
        RECT 148.950 487.950 151.050 490.050 ;
        RECT 152.250 488.250 154.050 489.150 ;
        RECT 142.950 485.850 144.750 486.750 ;
        RECT 145.950 484.950 148.050 487.050 ;
        RECT 151.950 484.950 154.050 487.050 ;
        RECT 146.400 481.050 147.450 484.950 ;
        RECT 145.950 478.950 148.050 481.050 ;
        RECT 145.950 475.950 148.050 478.050 ;
        RECT 139.950 472.950 142.050 475.050 ;
        RECT 146.400 457.050 147.450 475.950 ;
        RECT 148.950 472.950 151.050 475.050 ;
        RECT 136.950 454.950 139.050 457.050 ;
        RECT 140.250 455.250 141.750 456.150 ;
        RECT 142.950 454.950 145.050 457.050 ;
        RECT 145.950 454.950 148.050 457.050 ;
        RECT 136.950 452.850 138.750 453.750 ;
        RECT 139.950 451.950 142.050 454.050 ;
        RECT 143.250 452.850 144.750 453.750 ;
        RECT 145.950 449.850 148.050 450.750 ;
        RECT 149.400 432.450 150.450 472.950 ;
        RECT 152.400 463.050 153.450 484.950 ;
        RECT 151.950 460.950 154.050 463.050 ;
        RECT 151.950 454.950 154.050 457.050 ;
        RECT 146.400 431.400 150.450 432.450 ;
        RECT 133.950 418.950 136.050 421.050 ;
        RECT 133.950 415.950 136.050 418.050 ;
        RECT 139.950 415.950 142.050 418.050 ;
        RECT 134.400 409.050 135.450 415.950 ;
        RECT 140.400 415.050 141.450 415.950 ;
        RECT 146.400 415.050 147.450 431.400 ;
        RECT 139.950 412.950 142.050 415.050 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 149.250 413.250 151.050 414.150 ;
        RECT 139.950 410.850 142.050 411.750 ;
        RECT 142.950 410.250 145.050 411.150 ;
        RECT 145.950 410.850 147.750 411.750 ;
        RECT 148.950 409.950 151.050 412.050 ;
        RECT 133.950 406.950 136.050 409.050 ;
        RECT 142.950 406.950 145.050 409.050 ;
        RECT 130.950 400.950 133.050 403.050 ;
        RECT 118.950 388.950 121.050 391.050 ;
        RECT 112.950 385.950 115.050 388.050 ;
        RECT 113.400 385.050 114.450 385.950 ;
        RECT 119.400 385.050 120.450 388.950 ;
        RECT 130.950 385.950 133.050 388.050 ;
        RECT 112.950 382.950 115.050 385.050 ;
        RECT 116.250 383.250 117.750 384.150 ;
        RECT 118.950 382.950 121.050 385.050 ;
        RECT 121.950 382.950 124.050 385.050 ;
        RECT 122.400 382.050 123.450 382.950 ;
        RECT 131.400 382.050 132.450 385.950 ;
        RECT 109.950 379.950 112.050 382.050 ;
        RECT 112.950 380.850 114.750 381.750 ;
        RECT 115.950 379.950 118.050 382.050 ;
        RECT 119.250 380.850 120.750 381.750 ;
        RECT 121.950 379.950 124.050 382.050 ;
        RECT 130.950 379.950 133.050 382.050 ;
        RECT 121.950 377.850 124.050 378.750 ;
        RECT 134.400 367.050 135.450 406.950 ;
        RECT 139.950 403.950 142.050 406.050 ;
        RECT 140.400 388.050 141.450 403.950 ;
        RECT 148.950 388.950 151.050 391.050 ;
        RECT 139.950 385.950 142.050 388.050 ;
        RECT 136.950 383.250 139.050 384.150 ;
        RECT 139.950 383.850 142.050 384.750 ;
        RECT 142.950 383.250 144.750 384.150 ;
        RECT 145.950 382.950 148.050 385.050 ;
        RECT 136.950 379.950 139.050 382.050 ;
        RECT 139.950 379.950 142.050 382.050 ;
        RECT 142.950 379.950 145.050 382.050 ;
        RECT 146.250 380.850 148.050 381.750 ;
        RECT 112.950 364.950 115.050 367.050 ;
        RECT 133.950 364.950 136.050 367.050 ;
        RECT 113.400 346.050 114.450 364.950 ;
        RECT 118.950 347.250 121.050 348.150 ;
        RECT 140.400 346.050 141.450 379.950 ;
        RECT 112.950 343.950 115.050 346.050 ;
        RECT 116.250 344.250 117.750 345.150 ;
        RECT 118.950 343.950 121.050 346.050 ;
        RECT 122.250 344.250 124.050 345.150 ;
        RECT 133.950 343.950 136.050 346.050 ;
        RECT 137.250 344.250 138.750 345.150 ;
        RECT 139.950 343.950 142.050 346.050 ;
        RECT 112.950 341.850 114.750 342.750 ;
        RECT 115.950 340.950 118.050 343.050 ;
        RECT 116.400 331.050 117.450 340.950 ;
        RECT 115.950 328.950 118.050 331.050 ;
        RECT 119.400 319.050 120.450 343.950 ;
        RECT 121.950 340.950 124.050 343.050 ;
        RECT 127.950 340.950 130.050 343.050 ;
        RECT 133.950 341.850 135.750 342.750 ;
        RECT 136.950 340.950 139.050 343.050 ;
        RECT 140.250 341.850 142.050 342.750 ;
        RECT 118.950 316.950 121.050 319.050 ;
        RECT 118.950 313.950 121.050 316.050 ;
        RECT 128.400 313.050 129.450 340.950 ;
        RECT 137.400 322.050 138.450 340.950 ;
        RECT 143.400 340.050 144.450 379.950 ;
        RECT 145.950 376.950 148.050 379.050 ;
        RECT 142.950 337.950 145.050 340.050 ;
        RECT 136.950 319.950 139.050 322.050 ;
        RECT 136.950 316.950 139.050 319.050 ;
        RECT 133.950 313.950 136.050 316.050 ;
        RECT 112.950 310.950 115.050 313.050 ;
        RECT 116.250 311.250 118.050 312.150 ;
        RECT 118.950 311.850 121.050 312.750 ;
        RECT 121.950 311.250 124.050 312.150 ;
        RECT 124.950 310.950 127.050 313.050 ;
        RECT 127.950 310.950 130.050 313.050 ;
        RECT 112.950 308.850 114.750 309.750 ;
        RECT 115.950 307.950 118.050 310.050 ;
        RECT 121.950 307.950 124.050 310.050 ;
        RECT 116.400 307.050 117.450 307.950 ;
        RECT 115.950 304.950 118.050 307.050 ;
        RECT 121.950 304.950 124.050 307.050 ;
        RECT 122.400 304.050 123.450 304.950 ;
        RECT 106.950 301.950 109.050 304.050 ;
        RECT 121.950 301.950 124.050 304.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 106.950 277.950 109.050 280.050 ;
        RECT 107.400 277.050 108.450 277.950 ;
        RECT 106.950 274.950 109.050 277.050 ;
        RECT 88.950 268.950 91.050 271.050 ;
        RECT 97.950 269.250 100.050 270.150 ;
        RECT 103.950 269.250 106.050 270.150 ;
        RECT 85.950 244.950 88.050 247.050 ;
        RECT 82.950 243.450 85.050 244.050 ;
        RECT 80.400 242.400 85.050 243.450 ;
        RECT 82.950 241.950 85.050 242.400 ;
        RECT 76.950 238.950 79.050 241.050 ;
        RECT 80.250 239.250 82.050 240.150 ;
        RECT 82.950 239.850 85.050 240.750 ;
        RECT 85.950 239.250 88.050 240.150 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 76.950 236.850 78.750 237.750 ;
        RECT 79.950 235.950 82.050 238.050 ;
        RECT 85.950 237.450 88.050 238.050 ;
        RECT 89.400 237.450 90.450 268.950 ;
        RECT 97.950 265.950 100.050 268.050 ;
        RECT 101.250 266.250 102.750 267.150 ;
        RECT 103.950 265.950 106.050 268.050 ;
        RECT 91.950 244.950 94.050 247.050 ;
        RECT 85.950 236.400 90.450 237.450 ;
        RECT 85.950 235.950 88.050 236.400 ;
        RECT 80.400 202.050 81.450 235.950 ;
        RECT 89.400 235.050 90.450 236.400 ;
        RECT 88.950 232.950 91.050 235.050 ;
        RECT 70.950 199.950 73.050 202.050 ;
        RECT 73.950 200.250 76.050 201.150 ;
        RECT 79.950 199.950 82.050 202.050 ;
        RECT 71.400 195.450 72.450 199.950 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 77.250 197.250 78.750 198.150 ;
        RECT 79.950 196.950 82.050 199.050 ;
        RECT 83.250 197.250 85.050 198.150 ;
        RECT 85.950 196.950 88.050 199.050 ;
        RECT 71.400 194.400 75.450 195.450 ;
        RECT 74.400 192.450 75.450 194.400 ;
        RECT 76.950 193.950 79.050 196.050 ;
        RECT 80.250 194.850 81.750 195.750 ;
        RECT 82.950 193.950 85.050 196.050 ;
        RECT 83.400 193.050 84.450 193.950 ;
        RECT 74.400 191.400 81.450 192.450 ;
        RECT 80.400 190.050 81.450 191.400 ;
        RECT 82.950 190.950 85.050 193.050 ;
        RECT 67.950 187.950 70.050 190.050 ;
        RECT 76.950 187.950 79.050 190.050 ;
        RECT 79.950 187.950 82.050 190.050 ;
        RECT 70.950 184.950 73.050 187.050 ;
        RECT 64.950 175.950 67.050 178.050 ;
        RECT 65.400 172.050 66.450 175.950 ;
        RECT 64.950 169.950 67.050 172.050 ;
        RECT 65.400 169.050 66.450 169.950 ;
        RECT 71.400 169.050 72.450 184.950 ;
        RECT 64.950 166.950 67.050 169.050 ;
        RECT 68.250 167.250 69.750 168.150 ;
        RECT 70.950 166.950 73.050 169.050 ;
        RECT 64.950 164.850 66.750 165.750 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 71.250 164.850 72.750 165.750 ;
        RECT 73.950 163.950 76.050 166.050 ;
        RECT 68.400 163.050 69.450 163.950 ;
        RECT 67.950 160.950 70.050 163.050 ;
        RECT 73.950 161.850 76.050 162.750 ;
        RECT 52.950 151.950 55.050 154.050 ;
        RECT 58.950 151.950 61.050 154.050 ;
        RECT 61.950 151.950 64.050 154.050 ;
        RECT 53.400 130.050 54.450 151.950 ;
        RECT 77.400 145.050 78.450 187.950 ;
        RECT 79.950 181.950 82.050 184.050 ;
        RECT 80.400 163.050 81.450 181.950 ;
        RECT 79.950 160.950 82.050 163.050 ;
        RECT 70.950 142.950 73.050 145.050 ;
        RECT 76.950 142.950 79.050 145.050 ;
        RECT 58.950 131.250 61.050 132.150 ;
        RECT 52.950 127.950 55.050 130.050 ;
        RECT 56.250 128.250 57.750 129.150 ;
        RECT 58.950 127.950 61.050 130.050 ;
        RECT 62.250 128.250 64.050 129.150 ;
        RECT 64.950 127.950 67.050 130.050 ;
        RECT 52.950 125.850 54.750 126.750 ;
        RECT 55.950 124.950 58.050 127.050 ;
        RECT 46.950 121.950 49.050 124.050 ;
        RECT 56.400 121.050 57.450 124.950 ;
        RECT 59.400 121.050 60.450 127.950 ;
        RECT 61.950 126.450 64.050 127.050 ;
        RECT 65.400 126.450 66.450 127.950 ;
        RECT 61.950 125.400 66.450 126.450 ;
        RECT 61.950 124.950 64.050 125.400 ;
        RECT 31.950 118.950 34.050 121.050 ;
        RECT 34.950 118.950 37.050 121.050 ;
        RECT 40.950 118.950 43.050 121.050 ;
        RECT 49.950 118.950 52.050 121.050 ;
        RECT 55.950 118.950 58.050 121.050 ;
        RECT 58.950 118.950 61.050 121.050 ;
        RECT 32.400 69.450 33.450 118.950 ;
        RECT 35.400 97.050 36.450 118.950 ;
        RECT 40.950 97.950 43.050 100.050 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 38.250 95.250 40.050 96.150 ;
        RECT 40.950 95.850 43.050 96.750 ;
        RECT 43.950 95.250 46.050 96.150 ;
        RECT 34.950 92.850 36.750 93.750 ;
        RECT 37.950 91.950 40.050 94.050 ;
        RECT 43.950 91.950 46.050 94.050 ;
        RECT 46.950 91.950 49.050 94.050 ;
        RECT 29.400 68.400 33.450 69.450 ;
        RECT 29.400 51.450 30.450 68.400 ;
        RECT 43.950 61.950 46.050 64.050 ;
        RECT 31.950 56.250 34.050 57.150 ;
        RECT 44.400 55.050 45.450 61.950 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 35.250 53.250 36.750 54.150 ;
        RECT 37.950 52.950 40.050 55.050 ;
        RECT 41.250 53.250 43.050 54.150 ;
        RECT 43.950 52.950 46.050 55.050 ;
        RECT 34.950 51.450 37.050 52.050 ;
        RECT 29.400 50.400 37.050 51.450 ;
        RECT 38.250 50.850 39.750 51.750 ;
        RECT 34.950 49.950 37.050 50.400 ;
        RECT 40.950 49.950 43.050 52.050 ;
        RECT 37.950 46.950 40.050 49.050 ;
        RECT 31.950 25.950 34.050 28.050 ;
        RECT 38.400 25.050 39.450 46.950 ;
        RECT 41.400 40.050 42.450 49.950 ;
        RECT 44.400 49.050 45.450 52.950 ;
        RECT 47.400 52.050 48.450 91.950 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 43.950 46.950 46.050 49.050 ;
        RECT 50.400 46.050 51.450 118.950 ;
        RECT 52.950 106.950 55.050 109.050 ;
        RECT 53.400 90.450 54.450 106.950 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 55.950 92.250 57.750 93.150 ;
        RECT 58.950 91.950 61.050 94.050 ;
        RECT 64.950 93.450 67.050 94.050 ;
        RECT 68.400 93.450 69.450 97.950 ;
        RECT 64.950 92.400 69.450 93.450 ;
        RECT 64.950 91.950 67.050 92.400 ;
        RECT 55.950 90.450 58.050 91.050 ;
        RECT 53.400 89.400 58.050 90.450 ;
        RECT 59.250 89.850 60.750 90.750 ;
        RECT 55.950 88.950 58.050 89.400 ;
        RECT 61.950 88.950 64.050 91.050 ;
        RECT 65.250 89.850 67.050 90.750 ;
        RECT 61.950 86.850 64.050 87.750 ;
        RECT 68.400 82.050 69.450 92.400 ;
        RECT 67.950 79.950 70.050 82.050 ;
        RECT 55.950 56.250 58.050 57.150 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 62.400 55.050 63.450 55.950 ;
        RECT 55.950 52.950 58.050 55.050 ;
        RECT 59.250 53.250 60.750 54.150 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 65.250 53.250 67.050 54.150 ;
        RECT 67.950 52.950 70.050 55.050 ;
        RECT 56.400 52.050 57.450 52.950 ;
        RECT 55.950 49.950 58.050 52.050 ;
        RECT 58.950 49.950 61.050 52.050 ;
        RECT 62.250 50.850 63.750 51.750 ;
        RECT 64.950 49.950 67.050 52.050 ;
        RECT 59.400 46.050 60.450 49.950 ;
        RECT 65.400 49.050 66.450 49.950 ;
        RECT 64.950 46.950 67.050 49.050 ;
        RECT 49.950 43.950 52.050 46.050 ;
        RECT 58.950 43.950 61.050 46.050 ;
        RECT 40.950 37.950 43.050 40.050 ;
        RECT 55.950 37.950 58.050 40.050 ;
        RECT 56.400 25.050 57.450 37.950 ;
        RECT 61.950 28.950 64.050 31.050 ;
        RECT 62.400 28.050 63.450 28.950 ;
        RECT 61.950 25.950 64.050 28.050 ;
        RECT 25.950 22.950 28.050 25.050 ;
        RECT 28.950 23.250 31.050 24.150 ;
        RECT 31.950 23.850 34.050 24.750 ;
        RECT 34.950 23.250 36.750 24.150 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 59.250 23.250 61.050 24.150 ;
        RECT 61.950 23.850 64.050 24.750 ;
        RECT 64.950 23.250 67.050 24.150 ;
        RECT 26.400 19.050 27.450 22.950 ;
        RECT 28.950 19.950 31.050 22.050 ;
        RECT 34.950 19.950 37.050 22.050 ;
        RECT 38.250 20.850 40.050 21.750 ;
        RECT 55.950 20.850 57.750 21.750 ;
        RECT 58.950 19.950 61.050 22.050 ;
        RECT 64.950 21.450 67.050 22.050 ;
        RECT 68.400 21.450 69.450 52.950 ;
        RECT 71.400 37.050 72.450 142.950 ;
        RECT 86.400 136.050 87.450 196.950 ;
        RECT 92.400 172.050 93.450 244.950 ;
        RECT 98.400 238.050 99.450 265.950 ;
        RECT 107.400 265.050 108.450 274.950 ;
        RECT 118.950 271.950 121.050 274.050 ;
        RECT 119.400 271.050 120.450 271.950 ;
        RECT 125.400 271.050 126.450 310.950 ;
        RECT 130.950 309.450 133.050 310.050 ;
        RECT 128.400 308.400 133.050 309.450 ;
        RECT 128.400 307.050 129.450 308.400 ;
        RECT 130.950 307.950 133.050 308.400 ;
        RECT 134.400 307.050 135.450 313.950 ;
        RECT 137.400 310.050 138.450 316.950 ;
        RECT 136.950 307.950 139.050 310.050 ;
        RECT 140.250 308.250 142.050 309.150 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 130.950 305.850 132.750 306.750 ;
        RECT 133.950 304.950 136.050 307.050 ;
        RECT 137.250 305.850 138.750 306.750 ;
        RECT 139.950 304.950 142.050 307.050 ;
        RECT 112.950 270.450 115.050 271.050 ;
        RECT 110.400 269.400 115.050 270.450 ;
        RECT 100.950 264.450 103.050 265.050 ;
        RECT 103.950 264.450 106.050 265.050 ;
        RECT 100.950 263.400 106.050 264.450 ;
        RECT 100.950 262.950 103.050 263.400 ;
        RECT 103.950 262.950 106.050 263.400 ;
        RECT 106.950 262.950 109.050 265.050 ;
        RECT 110.400 256.050 111.450 269.400 ;
        RECT 112.950 268.950 115.050 269.400 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 122.250 269.250 124.050 270.150 ;
        RECT 124.950 268.950 127.050 271.050 ;
        RECT 112.950 266.850 115.050 267.750 ;
        RECT 115.950 266.250 118.050 267.150 ;
        RECT 118.950 266.850 120.750 267.750 ;
        RECT 121.950 265.950 124.050 268.050 ;
        RECT 115.950 262.950 118.050 265.050 ;
        RECT 128.400 262.050 129.450 304.950 ;
        RECT 140.400 304.050 141.450 304.950 ;
        RECT 133.950 302.850 136.050 303.750 ;
        RECT 139.950 301.950 142.050 304.050 ;
        RECT 142.950 301.950 145.050 304.050 ;
        RECT 143.400 274.050 144.450 301.950 ;
        RECT 142.950 271.950 145.050 274.050 ;
        RECT 139.950 268.950 142.050 271.050 ;
        RECT 146.400 268.050 147.450 376.950 ;
        RECT 149.400 364.050 150.450 388.950 ;
        RECT 148.950 361.950 151.050 364.050 ;
        RECT 152.400 348.450 153.450 454.950 ;
        RECT 154.950 436.950 157.050 439.050 ;
        RECT 155.400 379.050 156.450 436.950 ;
        RECT 158.400 381.450 159.450 529.950 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 164.400 520.050 165.450 526.950 ;
        RECT 167.400 522.450 168.450 532.950 ;
        RECT 172.950 526.950 175.050 529.050 ;
        RECT 173.400 526.050 174.450 526.950 ;
        RECT 169.950 524.250 171.750 525.150 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 176.400 523.050 177.450 562.950 ;
        RECT 194.400 562.050 195.450 574.950 ;
        RECT 178.950 559.950 181.050 562.050 ;
        RECT 184.950 560.250 186.750 561.150 ;
        RECT 187.950 559.950 190.050 562.050 ;
        RECT 191.250 560.250 192.750 561.150 ;
        RECT 193.950 559.950 196.050 562.050 ;
        RECT 179.400 544.050 180.450 559.950 ;
        RECT 184.950 556.950 187.050 559.050 ;
        RECT 190.950 556.950 193.050 559.050 ;
        RECT 194.250 557.850 196.050 558.750 ;
        RECT 178.950 541.950 181.050 544.050 ;
        RECT 181.950 541.950 184.050 544.050 ;
        RECT 182.400 529.050 183.450 541.950 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 178.950 525.450 181.050 526.050 ;
        RECT 178.950 524.400 183.450 525.450 ;
        RECT 178.950 523.950 181.050 524.400 ;
        RECT 169.950 522.450 172.050 523.050 ;
        RECT 167.400 521.400 172.050 522.450 ;
        RECT 173.250 521.850 174.750 522.750 ;
        RECT 169.950 520.950 172.050 521.400 ;
        RECT 175.950 520.950 178.050 523.050 ;
        RECT 179.250 521.850 181.050 522.750 ;
        RECT 163.950 517.950 166.050 520.050 ;
        RECT 175.950 518.850 178.050 519.750 ;
        RECT 182.400 519.450 183.450 524.400 ;
        RECT 179.400 518.400 183.450 519.450 ;
        RECT 160.950 496.950 163.050 499.050 ;
        RECT 161.400 466.050 162.450 496.950 ;
        RECT 169.950 491.250 172.050 492.150 ;
        RECT 175.950 490.950 178.050 493.050 ;
        RECT 163.950 487.950 166.050 490.050 ;
        RECT 167.250 488.250 168.750 489.150 ;
        RECT 169.950 487.950 172.050 490.050 ;
        RECT 173.250 488.250 175.050 489.150 ;
        RECT 163.950 485.850 165.750 486.750 ;
        RECT 166.950 484.950 169.050 487.050 ;
        RECT 170.400 478.050 171.450 487.950 ;
        RECT 172.950 486.450 175.050 487.050 ;
        RECT 176.400 486.450 177.450 490.950 ;
        RECT 172.950 485.400 177.450 486.450 ;
        RECT 172.950 484.950 175.050 485.400 ;
        RECT 175.950 481.950 178.050 484.050 ;
        RECT 169.950 475.950 172.050 478.050 ;
        RECT 176.400 472.050 177.450 481.950 ;
        RECT 175.950 469.950 178.050 472.050 ;
        RECT 169.950 466.950 172.050 469.050 ;
        RECT 160.950 463.950 163.050 466.050 ;
        RECT 160.950 452.250 162.750 453.150 ;
        RECT 163.950 451.950 166.050 454.050 ;
        RECT 167.250 452.250 169.050 453.150 ;
        RECT 160.950 448.950 163.050 451.050 ;
        RECT 164.250 449.850 165.750 450.750 ;
        RECT 166.950 448.950 169.050 451.050 ;
        RECT 161.400 448.050 162.450 448.950 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 164.400 420.450 165.450 445.950 ;
        RECT 167.400 445.050 168.450 448.950 ;
        RECT 166.950 442.950 169.050 445.050 ;
        RECT 164.400 419.400 168.450 420.450 ;
        RECT 167.400 418.050 168.450 419.400 ;
        RECT 160.950 415.950 163.050 418.050 ;
        RECT 164.250 416.250 165.750 417.150 ;
        RECT 166.950 415.950 169.050 418.050 ;
        RECT 160.950 413.850 162.750 414.750 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 167.250 413.850 169.050 414.750 ;
        RECT 164.400 388.050 165.450 412.950 ;
        RECT 163.950 385.950 166.050 388.050 ;
        RECT 170.400 385.050 171.450 466.950 ;
        RECT 172.950 460.950 175.050 463.050 ;
        RECT 173.400 451.050 174.450 460.950 ;
        RECT 175.950 457.950 178.050 460.050 ;
        RECT 172.950 448.950 175.050 451.050 ;
        RECT 176.400 391.050 177.450 457.950 ;
        RECT 179.400 403.050 180.450 518.400 ;
        RECT 185.400 499.050 186.450 556.950 ;
        RECT 191.400 544.050 192.450 556.950 ;
        RECT 197.400 547.050 198.450 589.950 ;
        RECT 200.400 565.050 201.450 601.950 ;
        RECT 199.950 562.950 202.050 565.050 ;
        RECT 203.400 562.050 204.450 625.950 ;
        RECT 208.950 598.950 211.050 601.050 ;
        RECT 212.400 600.450 213.450 638.400 ;
        RECT 215.400 631.050 216.450 667.950 ;
        RECT 214.950 628.950 217.050 631.050 ;
        RECT 218.400 627.450 219.450 670.950 ;
        RECT 221.400 652.050 222.450 691.950 ;
        RECT 229.950 676.950 232.050 679.050 ;
        RECT 230.400 673.050 231.450 676.950 ;
        RECT 223.950 670.950 226.050 673.050 ;
        RECT 227.250 671.250 228.750 672.150 ;
        RECT 229.950 670.950 232.050 673.050 ;
        RECT 232.950 670.950 235.050 673.050 ;
        RECT 233.400 670.050 234.450 670.950 ;
        RECT 223.950 668.850 225.750 669.750 ;
        RECT 226.950 667.950 229.050 670.050 ;
        RECT 230.250 668.850 231.750 669.750 ;
        RECT 232.950 667.950 235.050 670.050 ;
        RECT 227.400 664.050 228.450 667.950 ;
        RECT 232.950 665.850 235.050 666.750 ;
        RECT 226.950 661.950 229.050 664.050 ;
        RECT 232.950 661.950 235.050 664.050 ;
        RECT 220.950 649.950 223.050 652.050 ;
        RECT 226.950 634.950 229.050 637.050 ;
        RECT 227.400 634.050 228.450 634.950 ;
        RECT 220.950 631.950 223.050 634.050 ;
        RECT 224.250 632.250 225.750 633.150 ;
        RECT 226.950 631.950 229.050 634.050 ;
        RECT 220.950 629.850 222.750 630.750 ;
        RECT 223.950 628.950 226.050 631.050 ;
        RECT 227.250 629.850 229.050 630.750 ;
        RECT 229.950 628.950 232.050 631.050 ;
        RECT 218.400 626.400 222.450 627.450 ;
        RECT 212.400 599.400 216.450 600.450 ;
        RECT 209.400 598.050 210.450 598.950 ;
        RECT 205.950 596.250 207.750 597.150 ;
        RECT 208.950 595.950 211.050 598.050 ;
        RECT 212.250 596.250 214.050 597.150 ;
        RECT 205.950 592.950 208.050 595.050 ;
        RECT 209.250 593.850 210.750 594.750 ;
        RECT 211.950 592.950 214.050 595.050 ;
        RECT 206.400 592.050 207.450 592.950 ;
        RECT 205.950 589.950 208.050 592.050 ;
        RECT 208.950 562.950 211.050 565.050 ;
        RECT 199.950 559.950 202.050 562.050 ;
        RECT 202.950 559.950 205.050 562.050 ;
        RECT 196.950 544.950 199.050 547.050 ;
        RECT 190.950 541.950 193.050 544.050 ;
        RECT 200.400 529.050 201.450 559.950 ;
        RECT 199.950 526.950 202.050 529.050 ;
        RECT 187.950 524.250 189.750 525.150 ;
        RECT 190.950 523.950 193.050 526.050 ;
        RECT 194.250 524.250 196.050 525.150 ;
        RECT 199.950 523.950 202.050 526.050 ;
        RECT 187.950 520.950 190.050 523.050 ;
        RECT 191.250 521.850 192.750 522.750 ;
        RECT 193.950 520.950 196.050 523.050 ;
        RECT 194.400 520.050 195.450 520.950 ;
        RECT 187.950 517.950 190.050 520.050 ;
        RECT 193.950 517.950 196.050 520.050 ;
        RECT 184.950 496.950 187.050 499.050 ;
        RECT 188.400 495.450 189.450 517.950 ;
        RECT 193.950 514.950 196.050 517.050 ;
        RECT 185.400 494.400 189.450 495.450 ;
        RECT 181.950 487.950 184.050 490.050 ;
        RECT 182.400 487.050 183.450 487.950 ;
        RECT 185.400 487.050 186.450 494.400 ;
        RECT 187.950 490.950 190.050 493.050 ;
        RECT 188.400 487.050 189.450 490.950 ;
        RECT 181.950 484.950 184.050 487.050 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 187.950 484.950 190.050 487.050 ;
        RECT 191.250 485.250 193.050 486.150 ;
        RECT 181.950 482.850 184.050 483.750 ;
        RECT 184.950 482.250 187.050 483.150 ;
        RECT 187.950 482.850 189.750 483.750 ;
        RECT 190.950 481.950 193.050 484.050 ;
        RECT 184.950 478.950 187.050 481.050 ;
        RECT 185.400 478.050 186.450 478.950 ;
        RECT 184.950 475.950 187.050 478.050 ;
        RECT 181.950 472.950 184.050 475.050 ;
        RECT 182.400 457.050 183.450 472.950 ;
        RECT 184.950 469.950 187.050 472.050 ;
        RECT 185.400 460.050 186.450 469.950 ;
        RECT 191.400 460.050 192.450 481.950 ;
        RECT 194.400 469.050 195.450 514.950 ;
        RECT 200.400 472.050 201.450 523.950 ;
        RECT 203.400 523.050 204.450 559.950 ;
        RECT 209.400 559.050 210.450 562.950 ;
        RECT 212.400 562.050 213.450 592.950 ;
        RECT 215.400 562.050 216.450 599.400 ;
        RECT 217.950 598.950 220.050 601.050 ;
        RECT 211.950 559.950 214.050 562.050 ;
        RECT 214.950 559.950 217.050 562.050 ;
        RECT 218.400 559.050 219.450 598.950 ;
        RECT 205.950 556.950 208.050 559.050 ;
        RECT 208.950 556.950 211.050 559.050 ;
        RECT 211.950 556.950 214.050 559.050 ;
        RECT 215.250 557.250 217.050 558.150 ;
        RECT 217.950 556.950 220.050 559.050 ;
        RECT 205.950 554.850 208.050 555.750 ;
        RECT 208.950 554.250 211.050 555.150 ;
        RECT 211.950 554.850 213.750 555.750 ;
        RECT 214.950 553.950 217.050 556.050 ;
        RECT 208.950 550.950 211.050 553.050 ;
        RECT 209.400 550.050 210.450 550.950 ;
        RECT 208.950 547.950 211.050 550.050 ;
        RECT 205.950 544.950 208.050 547.050 ;
        RECT 206.400 541.050 207.450 544.950 ;
        RECT 205.950 538.950 208.050 541.050 ;
        RECT 202.950 520.950 205.050 523.050 ;
        RECT 206.400 517.050 207.450 538.950 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 212.400 526.050 213.450 526.950 ;
        RECT 208.950 524.250 210.750 525.150 ;
        RECT 211.950 523.950 214.050 526.050 ;
        RECT 217.950 523.950 220.050 526.050 ;
        RECT 208.950 520.950 211.050 523.050 ;
        RECT 212.250 521.850 213.750 522.750 ;
        RECT 214.950 520.950 217.050 523.050 ;
        RECT 218.250 521.850 220.050 522.750 ;
        RECT 211.950 517.950 214.050 520.050 ;
        RECT 214.950 518.850 217.050 519.750 ;
        RECT 205.950 514.950 208.050 517.050 ;
        RECT 202.950 493.950 205.050 496.050 ;
        RECT 199.950 469.950 202.050 472.050 ;
        RECT 193.950 466.950 196.050 469.050 ;
        RECT 184.950 457.950 187.050 460.050 ;
        RECT 190.950 457.950 193.050 460.050 ;
        RECT 196.950 457.950 199.050 460.050 ;
        RECT 197.400 457.050 198.450 457.950 ;
        RECT 203.400 457.050 204.450 493.950 ;
        RECT 205.950 484.950 208.050 487.050 ;
        RECT 205.950 482.850 208.050 483.750 ;
        RECT 208.950 482.250 211.050 483.150 ;
        RECT 208.950 478.950 211.050 481.050 ;
        RECT 209.400 469.050 210.450 478.950 ;
        RECT 208.950 466.950 211.050 469.050 ;
        RECT 181.950 454.950 184.050 457.050 ;
        RECT 185.250 455.850 186.750 456.750 ;
        RECT 187.950 456.450 190.050 457.050 ;
        RECT 187.950 455.400 192.450 456.450 ;
        RECT 187.950 454.950 190.050 455.400 ;
        RECT 181.950 452.850 184.050 453.750 ;
        RECT 187.950 452.850 190.050 453.750 ;
        RECT 191.400 445.050 192.450 455.400 ;
        RECT 193.950 454.950 196.050 457.050 ;
        RECT 196.950 454.950 199.050 457.050 ;
        RECT 200.250 455.250 201.750 456.150 ;
        RECT 202.950 454.950 205.050 457.050 ;
        RECT 190.950 442.950 193.050 445.050 ;
        RECT 194.400 424.050 195.450 454.950 ;
        RECT 196.950 452.850 198.750 453.750 ;
        RECT 199.950 451.950 202.050 454.050 ;
        RECT 203.250 452.850 204.750 453.750 ;
        RECT 205.950 453.450 208.050 454.050 ;
        RECT 205.950 452.400 210.450 453.450 ;
        RECT 205.950 451.950 208.050 452.400 ;
        RECT 205.950 449.850 208.050 450.750 ;
        RECT 209.400 439.050 210.450 452.400 ;
        RECT 212.400 451.050 213.450 517.950 ;
        RECT 221.400 511.050 222.450 626.400 ;
        RECT 224.400 607.050 225.450 628.950 ;
        RECT 230.400 607.050 231.450 628.950 ;
        RECT 233.400 619.050 234.450 661.950 ;
        RECT 236.400 624.450 237.450 698.400 ;
        RECT 241.950 697.950 244.050 700.050 ;
        RECT 238.950 694.950 241.050 697.050 ;
        RECT 239.400 694.050 240.450 694.950 ;
        RECT 238.950 691.950 241.050 694.050 ;
        RECT 239.400 664.050 240.450 691.950 ;
        RECT 238.950 661.950 241.050 664.050 ;
        RECT 242.400 631.050 243.450 697.950 ;
        RECT 248.400 679.050 249.450 772.950 ;
        RECT 250.950 769.950 253.050 772.050 ;
        RECT 254.250 770.850 255.750 771.750 ;
        RECT 256.950 769.950 259.050 772.050 ;
        RECT 262.950 769.950 265.050 772.050 ;
        RECT 253.950 766.950 256.050 769.050 ;
        RECT 254.400 742.050 255.450 766.950 ;
        RECT 256.950 745.950 259.050 748.050 ;
        RECT 257.400 745.050 258.450 745.950 ;
        RECT 263.400 745.050 264.450 769.950 ;
        RECT 266.400 769.050 267.450 811.950 ;
        RECT 275.400 811.050 276.450 838.950 ;
        RECT 287.400 838.050 288.450 838.950 ;
        RECT 286.950 835.950 289.050 838.050 ;
        RECT 277.950 817.950 280.050 820.050 ;
        RECT 278.400 814.050 279.450 817.950 ;
        RECT 277.950 811.950 280.050 814.050 ;
        RECT 268.950 808.950 271.050 811.050 ;
        RECT 272.250 809.850 273.750 810.750 ;
        RECT 274.950 808.950 277.050 811.050 ;
        RECT 278.250 809.850 280.050 810.750 ;
        RECT 274.950 806.850 277.050 807.750 ;
        RECT 287.400 778.050 288.450 835.950 ;
        RECT 295.950 820.950 298.050 823.050 ;
        RECT 292.950 814.950 295.050 817.050 ;
        RECT 293.400 814.050 294.450 814.950 ;
        RECT 289.950 812.250 291.750 813.150 ;
        RECT 292.950 811.950 295.050 814.050 ;
        RECT 296.400 811.050 297.450 820.950 ;
        RECT 308.400 820.050 309.450 841.950 ;
        RECT 314.400 820.050 315.450 841.950 ;
        RECT 317.400 841.050 318.450 847.950 ;
        RECT 319.950 844.950 322.050 847.050 ;
        RECT 322.950 845.250 324.750 846.150 ;
        RECT 325.950 844.950 328.050 847.050 ;
        RECT 329.250 845.250 330.750 846.150 ;
        RECT 331.950 844.950 334.050 847.050 ;
        RECT 343.950 846.450 346.050 847.050 ;
        RECT 341.400 845.400 346.050 846.450 ;
        RECT 316.950 838.950 319.050 841.050 ;
        RECT 307.950 817.950 310.050 820.050 ;
        RECT 313.950 817.950 316.050 820.050 ;
        RECT 298.950 813.450 301.050 814.050 ;
        RECT 298.950 812.400 303.450 813.450 ;
        RECT 298.950 811.950 301.050 812.400 ;
        RECT 289.950 808.950 292.050 811.050 ;
        RECT 293.250 809.850 294.750 810.750 ;
        RECT 295.950 808.950 298.050 811.050 ;
        RECT 299.250 809.850 301.050 810.750 ;
        RECT 283.950 775.950 286.050 778.050 ;
        RECT 286.950 775.950 289.050 778.050 ;
        RECT 290.400 777.450 291.450 808.950 ;
        RECT 302.400 808.050 303.450 812.400 ;
        RECT 304.950 811.950 307.050 814.050 ;
        RECT 307.950 812.250 309.750 813.150 ;
        RECT 310.950 811.950 313.050 814.050 ;
        RECT 314.250 812.250 316.050 813.150 ;
        RECT 295.950 806.850 298.050 807.750 ;
        RECT 301.950 805.950 304.050 808.050 ;
        RECT 301.950 781.950 304.050 784.050 ;
        RECT 298.950 778.950 301.050 781.050 ;
        RECT 290.400 776.400 294.450 777.450 ;
        RECT 284.400 775.050 285.450 775.950 ;
        RECT 268.950 772.950 271.050 775.050 ;
        RECT 274.950 772.950 277.050 775.050 ;
        RECT 283.950 774.450 286.050 775.050 ;
        RECT 280.950 773.250 282.750 774.150 ;
        RECT 283.950 773.400 288.450 774.450 ;
        RECT 283.950 772.950 286.050 773.400 ;
        RECT 265.950 766.950 268.050 769.050 ;
        RECT 265.950 754.950 268.050 757.050 ;
        RECT 256.950 742.950 259.050 745.050 ;
        RECT 260.250 743.250 261.750 744.150 ;
        RECT 262.950 742.950 265.050 745.050 ;
        RECT 266.400 742.050 267.450 754.950 ;
        RECT 269.400 742.050 270.450 772.950 ;
        RECT 274.950 770.850 277.050 771.750 ;
        RECT 280.950 769.950 283.050 772.050 ;
        RECT 284.250 770.850 286.050 771.750 ;
        RECT 281.400 769.050 282.450 769.950 ;
        RECT 280.950 766.950 283.050 769.050 ;
        RECT 287.400 757.050 288.450 773.400 ;
        RECT 289.950 773.250 292.050 774.150 ;
        RECT 289.950 769.950 292.050 772.050 ;
        RECT 286.950 754.950 289.050 757.050 ;
        RECT 274.950 745.950 277.050 748.050 ;
        RECT 271.950 743.250 274.050 744.150 ;
        RECT 274.950 743.850 277.050 744.750 ;
        RECT 277.950 743.250 279.750 744.150 ;
        RECT 280.950 742.950 283.050 745.050 ;
        RECT 286.950 742.950 289.050 745.050 ;
        RECT 293.400 744.450 294.450 776.400 ;
        RECT 299.400 747.450 300.450 778.950 ;
        RECT 302.400 771.450 303.450 781.950 ;
        RECT 305.400 781.050 306.450 811.950 ;
        RECT 307.950 808.950 310.050 811.050 ;
        RECT 311.250 809.850 312.750 810.750 ;
        RECT 313.950 808.950 316.050 811.050 ;
        RECT 314.400 808.050 315.450 808.950 ;
        RECT 313.950 805.950 316.050 808.050 ;
        RECT 304.950 778.950 307.050 781.050 ;
        RECT 313.950 778.950 316.050 781.050 ;
        RECT 307.950 775.950 310.050 778.050 ;
        RECT 308.400 775.050 309.450 775.950 ;
        RECT 314.400 775.050 315.450 778.950 ;
        RECT 320.400 775.050 321.450 844.950 ;
        RECT 332.400 844.050 333.450 844.950 ;
        RECT 322.950 841.950 325.050 844.050 ;
        RECT 326.250 842.850 327.750 843.750 ;
        RECT 328.950 841.950 331.050 844.050 ;
        RECT 331.950 841.950 334.050 844.050 ;
        RECT 323.400 841.050 324.450 841.950 ;
        RECT 329.400 841.050 330.450 841.950 ;
        RECT 322.950 838.950 325.050 841.050 ;
        RECT 328.950 838.950 331.050 841.050 ;
        RECT 332.400 834.450 333.450 841.950 ;
        RECT 341.400 835.050 342.450 845.400 ;
        RECT 343.950 844.950 346.050 845.400 ;
        RECT 349.950 844.950 352.050 847.050 ;
        RECT 353.250 845.250 355.050 846.150 ;
        RECT 343.950 842.850 346.050 843.750 ;
        RECT 346.950 842.250 349.050 843.150 ;
        RECT 349.950 842.850 351.750 843.750 ;
        RECT 352.950 843.450 355.050 844.050 ;
        RECT 356.400 843.450 357.450 847.950 ;
        RECT 361.950 844.950 364.050 847.050 ;
        RECT 367.950 845.850 369.750 846.750 ;
        RECT 370.950 844.950 373.050 847.050 ;
        RECT 374.250 845.850 376.050 846.750 ;
        RECT 352.950 842.400 357.450 843.450 ;
        RECT 352.950 841.950 355.050 842.400 ;
        RECT 346.950 838.950 349.050 841.050 ;
        RECT 347.400 838.050 348.450 838.950 ;
        RECT 346.950 835.950 349.050 838.050 ;
        RECT 329.400 833.400 333.450 834.450 ;
        RECT 329.400 813.450 330.450 833.400 ;
        RECT 340.950 832.950 343.050 835.050 ;
        RECT 346.950 832.950 349.050 835.050 ;
        RECT 334.950 817.950 337.050 820.050 ;
        RECT 347.400 817.050 348.450 832.950 ;
        RECT 356.400 832.050 357.450 842.400 ;
        RECT 355.950 829.950 358.050 832.050 ;
        RECT 362.400 820.050 363.450 844.950 ;
        RECT 377.400 820.050 378.450 848.400 ;
        RECT 383.400 848.400 388.050 849.450 ;
        RECT 383.400 823.050 384.450 848.400 ;
        RECT 385.950 847.950 388.050 848.400 ;
        RECT 389.250 848.250 390.750 849.150 ;
        RECT 391.950 847.950 394.050 850.050 ;
        RECT 395.250 848.250 397.050 849.150 ;
        RECT 406.950 847.950 409.050 850.050 ;
        RECT 410.250 848.250 411.750 849.150 ;
        RECT 412.950 847.950 415.050 850.050 ;
        RECT 416.250 848.250 418.050 849.150 ;
        RECT 418.950 847.950 421.050 850.050 ;
        RECT 424.950 849.450 427.050 850.050 ;
        RECT 422.400 848.400 427.050 849.450 ;
        RECT 385.950 845.850 387.750 846.750 ;
        RECT 388.950 844.950 391.050 847.050 ;
        RECT 394.950 844.950 397.050 847.050 ;
        RECT 403.950 844.950 406.050 847.050 ;
        RECT 406.950 845.850 408.750 846.750 ;
        RECT 409.950 844.950 412.050 847.050 ;
        RECT 415.950 844.950 418.050 847.050 ;
        RECT 382.950 820.950 385.050 823.050 ;
        RECT 361.950 817.950 364.050 820.050 ;
        RECT 373.950 817.950 376.050 820.050 ;
        RECT 376.950 817.950 379.050 820.050 ;
        RECT 331.950 815.250 334.050 816.150 ;
        RECT 334.950 815.850 337.050 816.750 ;
        RECT 346.950 814.950 349.050 817.050 ;
        RECT 355.950 816.450 358.050 817.050 ;
        RECT 362.400 816.450 363.450 817.950 ;
        RECT 364.950 816.450 367.050 817.050 ;
        RECT 355.950 815.400 360.450 816.450 ;
        RECT 355.950 814.950 358.050 815.400 ;
        RECT 331.950 813.450 334.050 814.050 ;
        RECT 329.400 812.400 334.050 813.450 ;
        RECT 346.950 812.850 349.050 813.750 ;
        RECT 325.950 793.950 328.050 796.050 ;
        RECT 326.400 778.050 327.450 793.950 ;
        RECT 329.400 784.050 330.450 812.400 ;
        RECT 331.950 811.950 334.050 812.400 ;
        RECT 349.950 812.250 352.050 813.150 ;
        RECT 355.950 812.850 358.050 813.750 ;
        RECT 349.950 808.950 352.050 811.050 ;
        RECT 350.400 796.050 351.450 808.950 ;
        RECT 349.950 793.950 352.050 796.050 ;
        RECT 328.950 781.950 331.050 784.050 ;
        RECT 359.400 781.050 360.450 815.400 ;
        RECT 362.400 815.400 367.050 816.450 ;
        RECT 331.950 778.950 334.050 781.050 ;
        RECT 352.950 779.250 355.050 780.150 ;
        RECT 358.950 778.950 361.050 781.050 ;
        RECT 332.400 778.050 333.450 778.950 ;
        RECT 325.950 777.450 328.050 778.050 ;
        RECT 323.400 776.400 328.050 777.450 ;
        RECT 304.950 773.250 306.750 774.150 ;
        RECT 307.950 772.950 310.050 775.050 ;
        RECT 311.250 773.250 312.750 774.150 ;
        RECT 313.950 772.950 316.050 775.050 ;
        RECT 317.250 773.250 319.050 774.150 ;
        RECT 319.950 772.950 322.050 775.050 ;
        RECT 304.950 771.450 307.050 772.050 ;
        RECT 302.400 770.400 307.050 771.450 ;
        RECT 308.250 770.850 309.750 771.750 ;
        RECT 304.950 769.950 307.050 770.400 ;
        RECT 310.950 769.950 313.050 772.050 ;
        RECT 314.250 770.850 315.750 771.750 ;
        RECT 316.950 769.950 319.050 772.050 ;
        RECT 317.400 766.050 318.450 769.950 ;
        RECT 323.400 766.050 324.450 776.400 ;
        RECT 325.950 775.950 328.050 776.400 ;
        RECT 329.250 776.250 330.750 777.150 ;
        RECT 331.950 775.950 334.050 778.050 ;
        RECT 346.950 775.950 349.050 778.050 ;
        RECT 350.250 776.250 351.750 777.150 ;
        RECT 352.950 775.950 355.050 778.050 ;
        RECT 356.250 776.250 358.050 777.150 ;
        RECT 325.950 773.850 327.750 774.750 ;
        RECT 328.950 772.950 331.050 775.050 ;
        RECT 332.250 773.850 334.050 774.750 ;
        RECT 340.950 772.950 343.050 775.050 ;
        RECT 346.950 773.850 348.750 774.750 ;
        RECT 349.950 772.950 352.050 775.050 ;
        RECT 316.950 763.950 319.050 766.050 ;
        RECT 322.950 763.950 325.050 766.050 ;
        RECT 313.950 754.950 316.050 757.050 ;
        RECT 299.400 746.400 303.450 747.450 ;
        RECT 290.400 743.400 294.450 744.450 ;
        RECT 253.950 741.450 256.050 742.050 ;
        RECT 251.400 740.400 256.050 741.450 ;
        RECT 257.250 740.850 258.750 741.750 ;
        RECT 251.400 736.050 252.450 740.400 ;
        RECT 253.950 739.950 256.050 740.400 ;
        RECT 259.950 739.950 262.050 742.050 ;
        RECT 263.250 740.850 265.050 741.750 ;
        RECT 265.950 739.950 268.050 742.050 ;
        RECT 268.950 739.950 271.050 742.050 ;
        RECT 271.950 739.950 274.050 742.050 ;
        RECT 277.950 739.950 280.050 742.050 ;
        RECT 281.250 740.850 283.050 741.750 ;
        RECT 283.950 739.950 286.050 742.050 ;
        RECT 272.400 739.050 273.450 739.950 ;
        RECT 253.950 737.850 256.050 738.750 ;
        RECT 271.950 736.950 274.050 739.050 ;
        RECT 250.950 733.950 253.050 736.050 ;
        RECT 272.400 721.050 273.450 736.950 ;
        RECT 277.950 733.950 280.050 736.050 ;
        RECT 271.950 718.950 274.050 721.050 ;
        RECT 256.950 703.950 259.050 706.050 ;
        RECT 259.950 704.250 262.050 705.150 ;
        RECT 257.400 702.450 258.450 703.950 ;
        RECT 259.950 702.450 262.050 703.050 ;
        RECT 257.400 701.400 262.050 702.450 ;
        RECT 257.400 700.050 258.450 701.400 ;
        RECT 259.950 700.950 262.050 701.400 ;
        RECT 263.250 701.250 264.750 702.150 ;
        RECT 265.950 700.950 268.050 703.050 ;
        RECT 269.250 701.250 271.050 702.150 ;
        RECT 256.950 697.950 259.050 700.050 ;
        RECT 262.950 697.950 265.050 700.050 ;
        RECT 266.250 698.850 267.750 699.750 ;
        RECT 268.950 697.950 271.050 700.050 ;
        RECT 256.950 694.950 259.050 697.050 ;
        RECT 250.950 688.950 253.050 691.050 ;
        RECT 247.950 676.950 250.050 679.050 ;
        RECT 251.400 670.050 252.450 688.950 ;
        RECT 257.400 670.050 258.450 694.950 ;
        RECT 263.400 684.450 264.450 697.950 ;
        RECT 274.950 685.950 277.050 688.050 ;
        RECT 260.400 683.400 264.450 684.450 ;
        RECT 247.950 668.250 249.750 669.150 ;
        RECT 250.950 667.950 253.050 670.050 ;
        RECT 254.250 668.250 256.050 669.150 ;
        RECT 256.950 667.950 259.050 670.050 ;
        RECT 247.950 664.950 250.050 667.050 ;
        RECT 251.250 665.850 252.750 666.750 ;
        RECT 253.950 664.950 256.050 667.050 ;
        RECT 248.400 634.050 249.450 664.950 ;
        RECT 254.400 661.050 255.450 664.950 ;
        RECT 253.950 658.950 256.050 661.050 ;
        RECT 250.950 640.950 253.050 643.050 ;
        RECT 247.950 631.950 250.050 634.050 ;
        RECT 238.950 629.250 241.050 630.150 ;
        RECT 241.950 628.950 244.050 631.050 ;
        RECT 244.950 629.250 247.050 630.150 ;
        RECT 238.950 625.950 241.050 628.050 ;
        RECT 242.250 626.250 243.750 627.150 ;
        RECT 244.950 625.950 247.050 628.050 ;
        RECT 236.400 623.400 240.450 624.450 ;
        RECT 232.950 616.950 235.050 619.050 ;
        RECT 223.950 604.950 226.050 607.050 ;
        RECT 229.950 604.950 232.050 607.050 ;
        RECT 232.950 604.950 235.050 607.050 ;
        RECT 230.400 604.050 231.450 604.950 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 226.950 599.250 229.050 600.150 ;
        RECT 229.950 599.850 232.050 600.750 ;
        RECT 226.950 595.950 229.050 598.050 ;
        RECT 227.400 562.050 228.450 595.950 ;
        RECT 233.400 592.050 234.450 604.950 ;
        RECT 232.950 589.950 235.050 592.050 ;
        RECT 229.950 562.950 232.050 565.050 ;
        RECT 226.950 559.950 229.050 562.050 ;
        RECT 230.400 559.050 231.450 562.950 ;
        RECT 235.950 560.250 238.050 561.150 ;
        RECT 223.950 556.950 226.050 559.050 ;
        RECT 226.950 557.250 228.750 558.150 ;
        RECT 229.950 556.950 232.050 559.050 ;
        RECT 233.250 557.250 234.750 558.150 ;
        RECT 235.950 556.950 238.050 559.050 ;
        RECT 224.400 553.050 225.450 556.950 ;
        RECT 226.950 553.950 229.050 556.050 ;
        RECT 230.250 554.850 231.750 555.750 ;
        RECT 232.950 553.950 235.050 556.050 ;
        RECT 223.950 550.950 226.050 553.050 ;
        RECT 239.400 547.050 240.450 623.400 ;
        RECT 241.950 622.950 244.050 625.050 ;
        RECT 245.400 619.050 246.450 625.950 ;
        RECT 248.400 624.450 249.450 631.950 ;
        RECT 251.400 628.050 252.450 640.950 ;
        RECT 260.400 640.050 261.450 683.400 ;
        RECT 262.950 679.950 265.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 263.400 666.450 264.450 679.950 ;
        RECT 268.950 673.950 271.050 676.050 ;
        RECT 269.400 670.050 270.450 673.950 ;
        RECT 265.950 668.250 267.750 669.150 ;
        RECT 268.950 667.950 271.050 670.050 ;
        RECT 272.400 667.050 273.450 679.950 ;
        RECT 275.400 670.050 276.450 685.950 ;
        RECT 274.950 667.950 277.050 670.050 ;
        RECT 265.950 666.450 268.050 667.050 ;
        RECT 263.400 665.400 268.050 666.450 ;
        RECT 269.250 665.850 270.750 666.750 ;
        RECT 265.950 664.950 268.050 665.400 ;
        RECT 271.950 664.950 274.050 667.050 ;
        RECT 275.250 665.850 277.050 666.750 ;
        RECT 268.950 661.950 271.050 664.050 ;
        RECT 271.950 662.850 274.050 663.750 ;
        RECT 259.950 637.950 262.050 640.050 ;
        RECT 262.950 635.250 265.050 636.150 ;
        RECT 269.400 634.050 270.450 661.950 ;
        RECT 278.400 658.050 279.450 733.950 ;
        RECT 280.950 708.450 283.050 709.050 ;
        RECT 284.400 708.450 285.450 739.950 ;
        RECT 287.400 739.050 288.450 742.950 ;
        RECT 286.950 736.950 289.050 739.050 ;
        RECT 280.950 707.400 285.450 708.450 ;
        RECT 280.950 706.950 283.050 707.400 ;
        RECT 281.400 706.050 282.450 706.950 ;
        RECT 280.950 703.950 283.050 706.050 ;
        RECT 286.950 705.450 289.050 706.050 ;
        RECT 290.400 705.450 291.450 743.400 ;
        RECT 292.950 740.250 294.750 741.150 ;
        RECT 295.950 739.950 298.050 742.050 ;
        RECT 299.250 740.250 301.050 741.150 ;
        RECT 292.950 736.950 295.050 739.050 ;
        RECT 296.250 737.850 297.750 738.750 ;
        RECT 298.950 738.450 301.050 739.050 ;
        RECT 302.400 738.450 303.450 746.400 ;
        RECT 314.400 745.050 315.450 754.950 ;
        RECT 319.950 745.950 322.050 748.050 ;
        RECT 313.950 742.950 316.050 745.050 ;
        RECT 317.250 743.250 319.050 744.150 ;
        RECT 319.950 743.850 322.050 744.750 ;
        RECT 322.950 743.250 325.050 744.150 ;
        RECT 329.400 742.050 330.450 772.950 ;
        RECT 341.400 748.050 342.450 772.950 ;
        RECT 353.400 760.050 354.450 775.950 ;
        RECT 355.950 772.950 358.050 775.050 ;
        RECT 356.400 769.050 357.450 772.950 ;
        RECT 362.400 772.050 363.450 815.400 ;
        RECT 364.950 814.950 367.050 815.400 ;
        RECT 368.250 815.250 369.750 816.150 ;
        RECT 370.950 814.950 373.050 817.050 ;
        RECT 374.400 814.050 375.450 817.950 ;
        RECT 382.950 814.950 385.050 817.050 ;
        RECT 388.950 814.950 391.050 817.050 ;
        RECT 400.950 814.950 403.050 817.050 ;
        RECT 364.950 812.850 366.750 813.750 ;
        RECT 367.950 811.950 370.050 814.050 ;
        RECT 371.250 812.850 372.750 813.750 ;
        RECT 373.950 811.950 376.050 814.050 ;
        RECT 368.400 810.450 369.450 811.950 ;
        RECT 365.400 809.400 369.450 810.450 ;
        RECT 373.950 809.850 376.050 810.750 ;
        RECT 361.950 769.950 364.050 772.050 ;
        RECT 355.950 766.950 358.050 769.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 340.950 745.950 343.050 748.050 ;
        RECT 337.950 743.250 340.050 744.150 ;
        RECT 340.950 743.850 343.050 744.750 ;
        RECT 353.400 742.050 354.450 757.950 ;
        RECT 365.400 757.050 366.450 809.400 ;
        RECT 383.400 808.050 384.450 814.950 ;
        RECT 382.950 805.950 385.050 808.050 ;
        RECT 382.950 778.950 385.050 781.050 ;
        RECT 370.950 775.950 373.050 778.050 ;
        RECT 371.400 775.050 372.450 775.950 ;
        RECT 367.950 773.250 369.750 774.150 ;
        RECT 370.950 772.950 373.050 775.050 ;
        RECT 376.950 774.450 379.050 775.050 ;
        RECT 376.950 773.400 381.450 774.450 ;
        RECT 376.950 772.950 379.050 773.400 ;
        RECT 367.950 769.950 370.050 772.050 ;
        RECT 371.250 770.850 373.050 771.750 ;
        RECT 373.950 770.250 376.050 771.150 ;
        RECT 376.950 770.850 379.050 771.750 ;
        RECT 373.950 766.950 376.050 769.050 ;
        RECT 364.950 754.950 367.050 757.050 ;
        RECT 364.950 751.950 367.050 754.050 ;
        RECT 355.950 745.950 358.050 748.050 ;
        RECT 356.400 745.050 357.450 745.950 ;
        RECT 355.950 742.950 358.050 745.050 ;
        RECT 359.250 743.250 360.750 744.150 ;
        RECT 361.950 742.950 364.050 745.050 ;
        RECT 313.950 740.850 315.750 741.750 ;
        RECT 316.950 739.950 319.050 742.050 ;
        RECT 322.950 739.950 325.050 742.050 ;
        RECT 328.950 739.950 331.050 742.050 ;
        RECT 337.950 739.950 340.050 742.050 ;
        RECT 352.950 739.950 355.050 742.050 ;
        RECT 356.250 740.850 357.750 741.750 ;
        RECT 358.950 739.950 361.050 742.050 ;
        RECT 362.250 740.850 364.050 741.750 ;
        RECT 323.400 739.050 324.450 739.950 ;
        RECT 298.950 737.400 303.450 738.450 ;
        RECT 298.950 736.950 301.050 737.400 ;
        RECT 322.950 736.950 325.050 739.050 ;
        RECT 352.950 737.850 355.050 738.750 ;
        RECT 284.250 704.250 285.750 705.150 ;
        RECT 286.950 704.400 291.450 705.450 ;
        RECT 286.950 703.950 289.050 704.400 ;
        RECT 280.950 701.850 282.750 702.750 ;
        RECT 283.950 700.950 286.050 703.050 ;
        RECT 287.250 701.850 289.050 702.750 ;
        RECT 271.950 655.950 274.050 658.050 ;
        RECT 277.950 655.950 280.050 658.050 ;
        RECT 256.950 633.450 259.050 634.050 ;
        RECT 254.400 632.400 259.050 633.450 ;
        RECT 250.950 625.950 253.050 628.050 ;
        RECT 248.400 623.400 252.450 624.450 ;
        RECT 241.950 616.950 244.050 619.050 ;
        RECT 244.950 616.950 247.050 619.050 ;
        RECT 242.400 615.450 243.450 616.950 ;
        RECT 242.400 614.400 249.450 615.450 ;
        RECT 248.400 607.050 249.450 614.400 ;
        RECT 247.950 604.950 250.050 607.050 ;
        RECT 244.950 601.950 247.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 248.400 601.050 249.450 601.950 ;
        RECT 241.950 598.950 244.050 601.050 ;
        RECT 245.250 599.850 246.750 600.750 ;
        RECT 247.950 598.950 250.050 601.050 ;
        RECT 241.950 596.850 244.050 597.750 ;
        RECT 244.950 595.950 247.050 598.050 ;
        RECT 247.950 596.850 250.050 597.750 ;
        RECT 232.950 544.950 235.050 547.050 ;
        RECT 238.950 544.950 241.050 547.050 ;
        RECT 233.400 529.050 234.450 544.950 ;
        RECT 238.950 541.950 241.050 544.050 ;
        RECT 226.950 528.450 229.050 529.050 ;
        RECT 224.400 527.400 229.050 528.450 ;
        RECT 220.950 508.950 223.050 511.050 ;
        RECT 224.400 493.050 225.450 527.400 ;
        RECT 226.950 526.950 229.050 527.400 ;
        RECT 230.250 527.250 231.750 528.150 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 226.950 524.850 228.750 525.750 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 233.250 524.850 234.750 525.750 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 235.950 521.850 238.050 522.750 ;
        RECT 223.950 490.950 226.050 493.050 ;
        RECT 226.950 491.250 229.050 492.150 ;
        RECT 232.950 490.950 235.050 493.050 ;
        RECT 220.950 487.950 223.050 490.050 ;
        RECT 224.250 488.250 225.750 489.150 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 230.250 488.250 232.050 489.150 ;
        RECT 214.950 484.950 217.050 487.050 ;
        RECT 220.950 485.850 222.750 486.750 ;
        RECT 223.950 484.950 226.050 487.050 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 208.950 436.950 211.050 439.050 ;
        RECT 193.950 421.950 196.050 424.050 ;
        RECT 184.950 416.250 187.050 417.150 ;
        RECT 196.950 415.950 199.050 418.050 ;
        RECT 211.950 416.250 214.050 417.150 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 188.250 413.250 189.750 414.150 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 194.250 413.250 196.050 414.150 ;
        RECT 178.950 400.950 181.050 403.050 ;
        RECT 185.400 400.050 186.450 412.950 ;
        RECT 197.400 412.050 198.450 415.950 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 413.250 204.750 414.150 ;
        RECT 205.950 412.950 208.050 415.050 ;
        RECT 209.250 413.250 210.750 414.150 ;
        RECT 211.950 412.950 214.050 415.050 ;
        RECT 187.950 409.950 190.050 412.050 ;
        RECT 191.250 410.850 192.750 411.750 ;
        RECT 193.950 409.950 196.050 412.050 ;
        RECT 196.950 409.950 199.050 412.050 ;
        RECT 184.950 397.950 187.050 400.050 ;
        RECT 175.950 388.950 178.050 391.050 ;
        RECT 175.950 385.950 178.050 388.050 ;
        RECT 163.950 382.950 166.050 385.050 ;
        RECT 167.250 383.250 168.750 384.150 ;
        RECT 169.950 382.950 172.050 385.050 ;
        RECT 160.950 381.450 163.050 382.050 ;
        RECT 158.400 380.400 163.050 381.450 ;
        RECT 164.250 380.850 165.750 381.750 ;
        RECT 154.950 376.950 157.050 379.050 ;
        RECT 149.400 347.400 153.450 348.450 ;
        RECT 149.400 312.450 150.450 347.400 ;
        RECT 151.950 343.950 154.050 346.050 ;
        RECT 158.400 345.450 159.450 380.400 ;
        RECT 160.950 379.950 163.050 380.400 ;
        RECT 166.950 379.950 169.050 382.050 ;
        RECT 170.250 380.850 172.050 381.750 ;
        RECT 160.950 377.850 163.050 378.750 ;
        RECT 163.950 358.950 166.050 361.050 ;
        RECT 155.400 344.400 159.450 345.450 ;
        RECT 152.400 343.050 153.450 343.950 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 151.950 338.850 154.050 339.750 ;
        RECT 155.400 337.050 156.450 344.400 ;
        RECT 157.950 341.250 160.050 342.150 ;
        RECT 157.950 337.950 160.050 340.050 ;
        RECT 161.250 338.250 163.050 339.150 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 158.400 334.050 159.450 337.950 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 164.400 334.050 165.450 358.950 ;
        RECT 166.950 343.950 169.050 346.050 ;
        RECT 157.950 331.950 160.050 334.050 ;
        RECT 163.950 331.950 166.050 334.050 ;
        RECT 167.400 313.050 168.450 343.950 ;
        RECT 173.250 341.250 175.050 342.150 ;
        RECT 169.950 338.850 171.750 339.750 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 149.400 311.400 153.450 312.450 ;
        RECT 148.950 307.950 151.050 310.050 ;
        RECT 139.950 266.850 142.050 267.750 ;
        RECT 142.950 266.250 145.050 267.150 ;
        RECT 145.950 265.950 148.050 268.050 ;
        RECT 149.400 265.050 150.450 307.950 ;
        RECT 152.400 283.050 153.450 311.400 ;
        RECT 166.950 310.950 169.050 313.050 ;
        RECT 169.950 310.950 172.050 313.050 ;
        RECT 167.400 310.050 168.450 310.950 ;
        RECT 157.950 308.250 159.750 309.150 ;
        RECT 160.950 307.950 163.050 310.050 ;
        RECT 166.950 307.950 169.050 310.050 ;
        RECT 157.950 304.950 160.050 307.050 ;
        RECT 161.250 305.850 162.750 306.750 ;
        RECT 163.950 304.950 166.050 307.050 ;
        RECT 167.250 305.850 169.050 306.750 ;
        RECT 163.950 302.850 166.050 303.750 ;
        RECT 151.950 280.950 154.050 283.050 ;
        RECT 170.400 277.050 171.450 310.950 ;
        RECT 169.950 274.950 172.050 277.050 ;
        RECT 157.950 272.250 160.050 273.150 ;
        RECT 154.950 268.950 157.050 271.050 ;
        RECT 157.950 268.950 160.050 271.050 ;
        RECT 161.250 269.250 162.750 270.150 ;
        RECT 163.950 268.950 166.050 271.050 ;
        RECT 167.250 269.250 169.050 270.150 ;
        RECT 155.400 265.050 156.450 268.950 ;
        RECT 142.950 262.950 145.050 265.050 ;
        RECT 148.950 262.950 151.050 265.050 ;
        RECT 154.950 262.950 157.050 265.050 ;
        RECT 143.400 262.050 144.450 262.950 ;
        RECT 127.950 259.950 130.050 262.050 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 109.950 253.950 112.050 256.050 ;
        RECT 110.400 244.050 111.450 253.950 ;
        RECT 103.950 241.950 106.050 244.050 ;
        RECT 109.950 241.950 112.050 244.050 ;
        RECT 112.950 241.950 115.050 244.050 ;
        RECT 94.950 236.250 96.750 237.150 ;
        RECT 97.950 235.950 100.050 238.050 ;
        RECT 101.250 236.250 103.050 237.150 ;
        RECT 94.950 232.950 97.050 235.050 ;
        RECT 98.250 233.850 99.750 234.750 ;
        RECT 100.950 234.450 103.050 235.050 ;
        RECT 104.400 234.450 105.450 241.950 ;
        RECT 112.950 239.850 115.050 240.750 ;
        RECT 115.950 239.250 118.050 240.150 ;
        RECT 128.400 238.050 129.450 259.950 ;
        RECT 139.950 247.950 142.050 250.050 ;
        RECT 133.950 241.950 136.050 244.050 ;
        RECT 134.400 241.050 135.450 241.950 ;
        RECT 140.400 241.050 141.450 247.950 ;
        RECT 130.950 238.950 133.050 241.050 ;
        RECT 133.950 238.950 136.050 241.050 ;
        RECT 137.250 239.250 138.750 240.150 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 131.400 238.050 132.450 238.950 ;
        RECT 115.950 235.950 118.050 238.050 ;
        RECT 127.950 235.950 130.050 238.050 ;
        RECT 130.950 235.950 133.050 238.050 ;
        RECT 134.250 236.850 135.750 237.750 ;
        RECT 136.950 235.950 139.050 238.050 ;
        RECT 140.250 236.850 142.050 237.750 ;
        RECT 100.950 233.400 105.450 234.450 ;
        RECT 130.950 233.850 133.050 234.750 ;
        RECT 100.950 232.950 103.050 233.400 ;
        RECT 112.950 229.950 115.050 232.050 ;
        RECT 94.950 200.250 97.050 201.150 ;
        RECT 94.950 196.950 97.050 199.050 ;
        RECT 98.250 197.250 99.750 198.150 ;
        RECT 100.950 196.950 103.050 199.050 ;
        RECT 104.250 197.250 106.050 198.150 ;
        RECT 95.400 196.050 96.450 196.950 ;
        RECT 94.950 193.950 97.050 196.050 ;
        RECT 97.950 193.950 100.050 196.050 ;
        RECT 101.250 194.850 102.750 195.750 ;
        RECT 103.950 193.950 106.050 196.050 ;
        RECT 98.400 190.050 99.450 193.950 ;
        RECT 97.950 187.950 100.050 190.050 ;
        RECT 97.950 172.950 100.050 175.050 ;
        RECT 91.950 169.950 94.050 172.050 ;
        RECT 91.950 166.950 94.050 169.050 ;
        RECT 92.400 166.050 93.450 166.950 ;
        RECT 98.400 166.050 99.450 172.950 ;
        RECT 100.950 169.950 103.050 172.050 ;
        RECT 88.950 164.250 90.750 165.150 ;
        RECT 91.950 163.950 94.050 166.050 ;
        RECT 97.950 163.950 100.050 166.050 ;
        RECT 101.400 163.050 102.450 169.950 ;
        RECT 104.400 168.450 105.450 193.950 ;
        RECT 113.400 169.050 114.450 229.950 ;
        RECT 143.400 229.050 144.450 259.950 ;
        RECT 145.950 241.950 148.050 244.050 ;
        RECT 146.400 238.050 147.450 241.950 ;
        RECT 145.950 235.950 148.050 238.050 ;
        RECT 142.950 226.950 145.050 229.050 ;
        RECT 121.950 202.950 124.050 205.050 ;
        RECT 136.950 202.950 139.050 205.050 ;
        RECT 122.400 202.050 123.450 202.950 ;
        RECT 137.400 202.050 138.450 202.950 ;
        RECT 121.950 199.950 124.050 202.050 ;
        RECT 130.950 199.950 133.050 202.050 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 140.250 200.250 141.750 201.150 ;
        RECT 142.950 199.950 145.050 202.050 ;
        RECT 118.950 197.250 121.050 198.150 ;
        RECT 121.950 197.850 124.050 198.750 ;
        RECT 127.950 197.250 130.050 198.150 ;
        RECT 118.950 193.950 121.050 196.050 ;
        RECT 127.950 195.450 130.050 196.050 ;
        RECT 131.400 195.450 132.450 199.950 ;
        RECT 136.950 197.850 138.750 198.750 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 143.250 197.850 145.050 198.750 ;
        RECT 127.950 194.400 132.450 195.450 ;
        RECT 127.950 193.950 130.050 194.400 ;
        RECT 140.400 175.050 141.450 196.950 ;
        RECT 115.950 172.950 118.050 175.050 ;
        RECT 139.950 172.950 142.050 175.050 ;
        RECT 106.950 168.450 109.050 169.050 ;
        RECT 104.400 167.400 109.050 168.450 ;
        RECT 104.400 163.050 105.450 167.400 ;
        RECT 106.950 166.950 109.050 167.400 ;
        RECT 110.250 167.250 111.750 168.150 ;
        RECT 112.950 166.950 115.050 169.050 ;
        RECT 116.400 166.050 117.450 172.950 ;
        RECT 149.400 172.050 150.450 262.950 ;
        RECT 158.400 262.050 159.450 268.950 ;
        RECT 160.950 265.950 163.050 268.050 ;
        RECT 164.250 266.850 165.750 267.750 ;
        RECT 166.950 265.950 169.050 268.050 ;
        RECT 157.950 259.950 160.050 262.050 ;
        RECT 154.950 238.950 157.050 241.050 ;
        RECT 161.400 240.450 162.450 265.950 ;
        RECT 169.950 262.950 172.050 265.050 ;
        RECT 170.400 253.050 171.450 262.950 ;
        RECT 169.950 250.950 172.050 253.050 ;
        RECT 163.950 247.950 166.050 250.050 ;
        RECT 158.400 239.400 162.450 240.450 ;
        RECT 155.400 238.050 156.450 238.950 ;
        RECT 151.950 236.250 153.750 237.150 ;
        RECT 154.950 235.950 157.050 238.050 ;
        RECT 158.400 235.050 159.450 239.400 ;
        RECT 160.950 237.450 163.050 238.050 ;
        RECT 164.400 237.450 165.450 247.950 ;
        RECT 160.950 236.400 165.450 237.450 ;
        RECT 160.950 235.950 163.050 236.400 ;
        RECT 151.950 232.950 154.050 235.050 ;
        RECT 155.250 233.850 156.750 234.750 ;
        RECT 157.950 232.950 160.050 235.050 ;
        RECT 161.250 233.850 163.050 234.750 ;
        RECT 152.400 205.050 153.450 232.950 ;
        RECT 157.950 230.850 160.050 231.750 ;
        RECT 151.950 202.950 154.050 205.050 ;
        RECT 157.950 196.950 160.050 199.050 ;
        RECT 157.950 194.850 160.050 195.750 ;
        RECT 160.950 194.250 163.050 195.150 ;
        RECT 160.950 192.450 163.050 193.050 ;
        RECT 164.400 192.450 165.450 236.400 ;
        RECT 170.400 234.450 171.450 250.950 ;
        RECT 173.400 241.050 174.450 337.950 ;
        RECT 176.400 334.050 177.450 385.950 ;
        RECT 188.400 384.450 189.450 409.950 ;
        RECT 194.400 406.050 195.450 409.950 ;
        RECT 200.400 409.050 201.450 412.950 ;
        RECT 202.950 409.950 205.050 412.050 ;
        RECT 206.250 410.850 207.750 411.750 ;
        RECT 208.950 409.950 211.050 412.050 ;
        RECT 199.950 406.950 202.050 409.050 ;
        RECT 193.950 403.950 196.050 406.050 ;
        RECT 203.400 400.050 204.450 409.950 ;
        RECT 202.950 397.950 205.050 400.050 ;
        RECT 196.950 384.450 199.050 385.050 ;
        RECT 205.950 384.450 208.050 385.050 ;
        RECT 188.400 383.400 192.450 384.450 ;
        RECT 178.950 379.950 181.050 382.050 ;
        RECT 181.950 380.250 183.750 381.150 ;
        RECT 184.950 379.950 187.050 382.050 ;
        RECT 188.250 380.250 190.050 381.150 ;
        RECT 179.400 367.050 180.450 379.950 ;
        RECT 191.400 379.050 192.450 383.400 ;
        RECT 196.950 383.400 201.450 384.450 ;
        RECT 196.950 382.950 199.050 383.400 ;
        RECT 196.950 380.850 199.050 381.750 ;
        RECT 181.950 376.950 184.050 379.050 ;
        RECT 185.250 377.850 186.750 378.750 ;
        RECT 187.950 378.450 190.050 379.050 ;
        RECT 190.950 378.450 193.050 379.050 ;
        RECT 187.950 377.400 193.050 378.450 ;
        RECT 187.950 376.950 190.050 377.400 ;
        RECT 190.950 376.950 193.050 377.400 ;
        RECT 182.400 376.050 183.450 376.950 ;
        RECT 200.400 376.050 201.450 383.400 ;
        RECT 205.950 383.400 210.450 384.450 ;
        RECT 205.950 382.950 208.050 383.400 ;
        RECT 202.950 380.250 205.050 381.150 ;
        RECT 205.950 380.850 208.050 381.750 ;
        RECT 202.950 376.950 205.050 379.050 ;
        RECT 181.950 373.950 184.050 376.050 ;
        RECT 199.950 373.950 202.050 376.050 ;
        RECT 178.950 364.950 181.050 367.050 ;
        RECT 175.950 331.950 178.050 334.050 ;
        RECT 179.400 330.450 180.450 364.950 ;
        RECT 209.400 352.050 210.450 383.400 ;
        RECT 211.950 382.950 214.050 385.050 ;
        RECT 212.400 382.050 213.450 382.950 ;
        RECT 211.950 379.950 214.050 382.050 ;
        RECT 208.950 349.950 211.050 352.050 ;
        RECT 193.950 347.250 196.050 348.150 ;
        RECT 212.400 346.050 213.450 379.950 ;
        RECT 215.400 346.050 216.450 484.950 ;
        RECT 224.400 481.050 225.450 484.950 ;
        RECT 227.400 484.050 228.450 487.950 ;
        RECT 229.950 486.450 232.050 487.050 ;
        RECT 233.400 486.450 234.450 490.950 ;
        RECT 235.950 487.950 238.050 490.050 ;
        RECT 229.950 485.400 234.450 486.450 ;
        RECT 229.950 484.950 232.050 485.400 ;
        RECT 226.950 481.950 229.050 484.050 ;
        RECT 223.950 478.950 226.050 481.050 ;
        RECT 232.950 478.950 235.050 481.050 ;
        RECT 229.950 466.950 232.050 469.050 ;
        RECT 223.950 460.950 226.050 463.050 ;
        RECT 224.400 454.050 225.450 460.950 ;
        RECT 226.950 457.950 229.050 460.050 ;
        RECT 220.950 452.250 222.750 453.150 ;
        RECT 223.950 451.950 226.050 454.050 ;
        RECT 227.400 451.050 228.450 457.950 ;
        RECT 230.400 454.050 231.450 466.950 ;
        RECT 229.950 451.950 232.050 454.050 ;
        RECT 220.950 448.950 223.050 451.050 ;
        RECT 224.250 449.850 225.750 450.750 ;
        RECT 226.950 448.950 229.050 451.050 ;
        RECT 230.250 449.850 232.050 450.750 ;
        RECT 233.400 448.050 234.450 478.950 ;
        RECT 236.400 460.050 237.450 487.950 ;
        RECT 239.400 487.050 240.450 541.950 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 242.400 523.050 243.450 523.950 ;
        RECT 241.950 520.950 244.050 523.050 ;
        RECT 242.400 490.050 243.450 520.950 ;
        RECT 245.400 520.050 246.450 595.950 ;
        RECT 251.400 580.050 252.450 623.400 ;
        RECT 254.400 622.050 255.450 632.400 ;
        RECT 256.950 631.950 259.050 632.400 ;
        RECT 260.250 632.250 261.750 633.150 ;
        RECT 262.950 631.950 265.050 634.050 ;
        RECT 266.250 632.250 268.050 633.150 ;
        RECT 268.950 631.950 271.050 634.050 ;
        RECT 256.950 629.850 258.750 630.750 ;
        RECT 259.950 628.950 262.050 631.050 ;
        RECT 265.950 628.950 268.050 631.050 ;
        RECT 260.400 628.050 261.450 628.950 ;
        RECT 259.950 625.950 262.050 628.050 ;
        RECT 272.400 625.050 273.450 655.950 ;
        RECT 277.950 640.950 280.050 643.050 ;
        RECT 274.950 637.950 277.050 640.050 ;
        RECT 256.950 622.950 259.050 625.050 ;
        RECT 271.950 622.950 274.050 625.050 ;
        RECT 253.950 619.950 256.050 622.050 ;
        RECT 253.950 604.950 256.050 607.050 ;
        RECT 254.400 598.050 255.450 604.950 ;
        RECT 253.950 595.950 256.050 598.050 ;
        RECT 250.950 577.950 253.050 580.050 ;
        RECT 250.950 559.950 253.050 562.050 ;
        RECT 251.400 559.050 252.450 559.950 ;
        RECT 250.950 556.950 253.050 559.050 ;
        RECT 247.950 554.250 250.050 555.150 ;
        RECT 250.950 554.850 253.050 555.750 ;
        RECT 247.950 550.950 250.050 553.050 ;
        RECT 257.400 535.050 258.450 622.950 ;
        RECT 271.950 604.950 274.050 607.050 ;
        RECT 262.950 601.950 265.050 604.050 ;
        RECT 259.950 599.250 262.050 600.150 ;
        RECT 262.950 599.850 265.050 600.750 ;
        RECT 272.400 598.050 273.450 604.950 ;
        RECT 275.400 604.050 276.450 637.950 ;
        RECT 278.400 634.050 279.450 640.950 ;
        RECT 284.400 640.050 285.450 700.950 ;
        RECT 293.400 700.050 294.450 736.950 ;
        RECT 299.400 703.050 300.450 736.950 ;
        RECT 316.950 715.950 319.050 718.050 ;
        RECT 304.950 704.250 307.050 705.150 ;
        RECT 295.950 701.250 297.750 702.150 ;
        RECT 298.950 700.950 301.050 703.050 ;
        RECT 302.250 701.250 303.750 702.150 ;
        RECT 304.950 700.950 307.050 703.050 ;
        RECT 310.950 700.950 313.050 703.050 ;
        RECT 292.950 699.450 295.050 700.050 ;
        RECT 295.950 699.450 298.050 700.050 ;
        RECT 292.950 698.400 298.050 699.450 ;
        RECT 299.250 698.850 300.750 699.750 ;
        RECT 292.950 697.950 295.050 698.400 ;
        RECT 295.950 697.950 298.050 698.400 ;
        RECT 301.950 697.950 304.050 700.050 ;
        RECT 289.950 682.950 292.050 685.050 ;
        RECT 290.400 676.050 291.450 682.950 ;
        RECT 302.400 679.050 303.450 697.950 ;
        RECT 305.400 697.050 306.450 700.950 ;
        RECT 304.950 694.950 307.050 697.050 ;
        RECT 295.950 676.950 298.050 679.050 ;
        RECT 301.950 676.950 304.050 679.050 ;
        RECT 289.950 673.950 292.050 676.050 ;
        RECT 292.950 673.950 295.050 676.050 ;
        RECT 293.400 673.050 294.450 673.950 ;
        RECT 286.950 670.950 289.050 673.050 ;
        RECT 290.250 671.850 291.750 672.750 ;
        RECT 292.950 670.950 295.050 673.050 ;
        RECT 286.950 668.850 289.050 669.750 ;
        RECT 289.950 667.950 292.050 670.050 ;
        RECT 292.950 668.850 295.050 669.750 ;
        RECT 290.400 640.050 291.450 667.950 ;
        RECT 296.400 654.450 297.450 676.950 ;
        RECT 301.950 675.450 304.050 676.050 ;
        RECT 301.950 674.400 306.450 675.450 ;
        RECT 301.950 673.950 304.050 674.400 ;
        RECT 305.400 673.050 306.450 674.400 ;
        RECT 301.950 670.950 304.050 673.050 ;
        RECT 304.950 670.950 307.050 673.050 ;
        RECT 302.400 666.450 303.450 670.950 ;
        RECT 304.950 668.250 306.750 669.150 ;
        RECT 307.950 667.950 310.050 670.050 ;
        RECT 311.400 667.050 312.450 700.950 ;
        RECT 313.950 697.950 316.050 700.050 ;
        RECT 314.400 688.050 315.450 697.950 ;
        RECT 313.950 685.950 316.050 688.050 ;
        RECT 314.400 670.050 315.450 685.950 ;
        RECT 313.950 667.950 316.050 670.050 ;
        RECT 304.950 666.450 307.050 667.050 ;
        RECT 302.400 665.400 307.050 666.450 ;
        RECT 308.250 665.850 309.750 666.750 ;
        RECT 304.950 664.950 307.050 665.400 ;
        RECT 310.950 664.950 313.050 667.050 ;
        RECT 314.250 665.850 316.050 666.750 ;
        RECT 307.950 661.950 310.050 664.050 ;
        RECT 310.950 662.850 313.050 663.750 ;
        RECT 293.400 653.400 297.450 654.450 ;
        RECT 283.950 637.950 286.050 640.050 ;
        RECT 289.950 637.950 292.050 640.050 ;
        RECT 283.950 635.250 286.050 636.150 ;
        RECT 277.950 631.950 280.050 634.050 ;
        RECT 281.250 632.250 282.750 633.150 ;
        RECT 283.950 631.950 286.050 634.050 ;
        RECT 287.250 632.250 289.050 633.150 ;
        RECT 277.950 629.850 279.750 630.750 ;
        RECT 280.950 628.950 283.050 631.050 ;
        RECT 281.400 628.050 282.450 628.950 ;
        RECT 280.950 625.950 283.050 628.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 259.950 595.950 262.050 598.050 ;
        RECT 271.950 595.950 274.050 598.050 ;
        RECT 260.400 559.050 261.450 595.950 ;
        RECT 275.400 595.050 276.450 601.950 ;
        RECT 281.400 601.050 282.450 625.950 ;
        RECT 284.400 625.050 285.450 631.950 ;
        RECT 290.400 631.050 291.450 637.950 ;
        RECT 286.950 630.450 289.050 631.050 ;
        RECT 289.950 630.450 292.050 631.050 ;
        RECT 286.950 629.400 292.050 630.450 ;
        RECT 286.950 628.950 289.050 629.400 ;
        RECT 289.950 628.950 292.050 629.400 ;
        RECT 283.950 622.950 286.050 625.050 ;
        RECT 280.950 598.950 283.050 601.050 ;
        RECT 277.950 595.950 280.050 598.050 ;
        RECT 281.250 596.250 283.050 597.150 ;
        RECT 283.950 595.950 286.050 598.050 ;
        RECT 271.950 593.850 273.750 594.750 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 278.250 593.850 279.750 594.750 ;
        RECT 280.950 592.950 283.050 595.050 ;
        RECT 274.950 590.850 277.050 591.750 ;
        RECT 281.400 565.050 282.450 592.950 ;
        RECT 284.400 565.050 285.450 595.950 ;
        RECT 271.950 562.950 274.050 565.050 ;
        RECT 280.950 562.950 283.050 565.050 ;
        RECT 283.950 562.950 286.050 565.050 ;
        RECT 272.400 562.050 273.450 562.950 ;
        RECT 265.950 561.450 268.050 562.050 ;
        RECT 263.400 560.400 268.050 561.450 ;
        RECT 259.950 556.950 262.050 559.050 ;
        RECT 263.400 556.050 264.450 560.400 ;
        RECT 265.950 559.950 268.050 560.400 ;
        RECT 269.250 560.250 270.750 561.150 ;
        RECT 271.950 559.950 274.050 562.050 ;
        RECT 280.950 559.950 283.050 562.050 ;
        RECT 286.950 561.450 289.050 562.050 ;
        RECT 284.250 560.250 285.750 561.150 ;
        RECT 286.950 560.400 291.450 561.450 ;
        RECT 286.950 559.950 289.050 560.400 ;
        RECT 265.950 557.850 267.750 558.750 ;
        RECT 268.950 556.950 271.050 559.050 ;
        RECT 272.250 557.850 274.050 558.750 ;
        RECT 280.950 557.850 282.750 558.750 ;
        RECT 283.950 556.950 286.050 559.050 ;
        RECT 287.250 557.850 289.050 558.750 ;
        RECT 262.950 553.950 265.050 556.050 ;
        RECT 262.950 535.950 265.050 538.050 ;
        RECT 256.950 532.950 259.050 535.050 ;
        RECT 247.950 529.950 250.050 532.050 ;
        RECT 256.950 529.950 259.050 532.050 ;
        RECT 248.400 523.050 249.450 529.950 ;
        RECT 250.950 526.950 253.050 529.050 ;
        RECT 254.250 527.250 256.050 528.150 ;
        RECT 256.950 527.850 259.050 528.750 ;
        RECT 259.950 527.250 262.050 528.150 ;
        RECT 250.950 524.850 252.750 525.750 ;
        RECT 253.950 525.450 256.050 526.050 ;
        RECT 259.950 525.450 262.050 526.050 ;
        RECT 263.400 525.450 264.450 535.950 ;
        RECT 253.950 524.400 258.450 525.450 ;
        RECT 253.950 523.950 256.050 524.400 ;
        RECT 247.950 520.950 250.050 523.050 ;
        RECT 253.950 520.950 256.050 523.050 ;
        RECT 244.950 517.950 247.050 520.050 ;
        RECT 247.950 491.250 250.050 492.150 ;
        RECT 241.950 487.950 244.050 490.050 ;
        RECT 245.250 488.250 246.750 489.150 ;
        RECT 247.950 487.950 250.050 490.050 ;
        RECT 251.250 488.250 253.050 489.150 ;
        RECT 238.950 484.950 241.050 487.050 ;
        RECT 241.950 485.850 243.750 486.750 ;
        RECT 244.950 484.950 247.050 487.050 ;
        RECT 250.950 486.450 253.050 487.050 ;
        RECT 254.400 486.450 255.450 520.950 ;
        RECT 257.400 487.050 258.450 524.400 ;
        RECT 259.950 524.400 264.450 525.450 ;
        RECT 259.950 523.950 262.050 524.400 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 260.400 493.050 261.450 523.950 ;
        RECT 262.950 517.950 265.050 520.050 ;
        RECT 259.950 490.950 262.050 493.050 ;
        RECT 263.400 489.450 264.450 517.950 ;
        RECT 266.400 496.050 267.450 523.950 ;
        RECT 265.950 493.950 268.050 496.050 ;
        RECT 260.400 488.400 264.450 489.450 ;
        RECT 250.950 485.400 255.450 486.450 ;
        RECT 250.950 484.950 253.050 485.400 ;
        RECT 256.950 484.950 259.050 487.050 ;
        RECT 251.400 484.050 252.450 484.950 ;
        RECT 250.950 481.950 253.050 484.050 ;
        RECT 241.950 469.950 244.050 472.050 ;
        RECT 238.950 463.950 241.050 466.050 ;
        RECT 235.950 457.950 238.050 460.050 ;
        RECT 226.950 446.850 229.050 447.750 ;
        RECT 232.950 445.950 235.050 448.050 ;
        RECT 223.950 442.950 226.050 445.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 221.400 384.450 222.450 412.950 ;
        RECT 224.400 412.050 225.450 442.950 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 232.950 413.250 235.050 414.150 ;
        RECT 223.950 409.950 226.050 412.050 ;
        RECT 226.950 410.850 229.050 411.750 ;
        RECT 232.950 409.950 235.050 412.050 ;
        RECT 236.250 410.250 238.050 411.150 ;
        RECT 235.950 406.950 238.050 409.050 ;
        RECT 236.400 397.050 237.450 406.950 ;
        RECT 239.400 406.050 240.450 463.950 ;
        RECT 242.400 433.050 243.450 469.950 ;
        RECT 250.950 457.950 253.050 460.050 ;
        RECT 244.950 454.950 247.050 457.050 ;
        RECT 248.250 455.250 250.050 456.150 ;
        RECT 250.950 455.850 253.050 456.750 ;
        RECT 253.950 455.250 256.050 456.150 ;
        RECT 257.400 454.050 258.450 484.950 ;
        RECT 260.400 468.450 261.450 488.400 ;
        RECT 266.400 487.050 267.450 493.950 ;
        RECT 269.400 487.050 270.450 556.950 ;
        RECT 290.400 550.050 291.450 560.400 ;
        RECT 293.400 556.050 294.450 653.400 ;
        RECT 308.400 637.050 309.450 661.950 ;
        RECT 317.400 640.050 318.450 715.950 ;
        RECT 319.950 709.950 322.050 712.050 ;
        RECT 361.950 709.950 364.050 712.050 ;
        RECT 320.400 706.050 321.450 709.950 ;
        RECT 325.950 707.250 328.050 708.150 ;
        RECT 334.950 706.950 337.050 709.050 ;
        RECT 319.950 703.950 322.050 706.050 ;
        RECT 323.250 704.250 324.750 705.150 ;
        RECT 325.950 703.950 328.050 706.050 ;
        RECT 329.250 704.250 331.050 705.150 ;
        RECT 319.950 701.850 321.750 702.750 ;
        RECT 322.950 700.950 325.050 703.050 ;
        RECT 323.400 670.050 324.450 700.950 ;
        RECT 326.400 697.050 327.450 703.950 ;
        RECT 328.950 700.950 331.050 703.050 ;
        RECT 329.400 700.050 330.450 700.950 ;
        RECT 328.950 697.950 331.050 700.050 ;
        RECT 325.950 694.950 328.050 697.050 ;
        RECT 326.400 682.050 327.450 694.950 ;
        RECT 325.950 679.950 328.050 682.050 ;
        RECT 331.950 673.950 334.050 676.050 ;
        RECT 332.400 673.050 333.450 673.950 ;
        RECT 325.950 670.950 328.050 673.050 ;
        RECT 331.950 670.950 334.050 673.050 ;
        RECT 322.950 667.950 325.050 670.050 ;
        RECT 323.400 643.050 324.450 667.950 ;
        RECT 326.400 666.450 327.450 670.950 ;
        RECT 332.400 670.050 333.450 670.950 ;
        RECT 328.950 668.250 330.750 669.150 ;
        RECT 331.950 667.950 334.050 670.050 ;
        RECT 335.400 667.050 336.450 706.950 ;
        RECT 362.400 706.050 363.450 709.950 ;
        RECT 355.950 705.450 358.050 706.050 ;
        RECT 353.400 704.400 358.050 705.450 ;
        RECT 353.400 703.050 354.450 704.400 ;
        RECT 355.950 703.950 358.050 704.400 ;
        RECT 359.250 704.250 360.750 705.150 ;
        RECT 361.950 703.950 364.050 706.050 ;
        RECT 365.400 703.050 366.450 751.950 ;
        RECT 367.950 742.950 370.050 745.050 ;
        RECT 340.950 701.250 343.050 702.150 ;
        RECT 346.950 701.250 349.050 702.150 ;
        RECT 352.950 700.950 355.050 703.050 ;
        RECT 355.950 701.850 357.750 702.750 ;
        RECT 358.950 700.950 361.050 703.050 ;
        RECT 362.250 701.850 364.050 702.750 ;
        RECT 364.950 700.950 367.050 703.050 ;
        RECT 337.950 697.950 340.050 700.050 ;
        RECT 340.950 697.950 343.050 700.050 ;
        RECT 346.950 697.950 349.050 700.050 ;
        RECT 358.950 697.950 361.050 700.050 ;
        RECT 338.400 670.050 339.450 697.950 ;
        RECT 347.400 694.050 348.450 697.950 ;
        RECT 346.950 691.950 349.050 694.050 ;
        RECT 340.950 682.950 343.050 685.050 ;
        RECT 337.950 667.950 340.050 670.050 ;
        RECT 328.950 666.450 331.050 667.050 ;
        RECT 326.400 665.400 331.050 666.450 ;
        RECT 332.250 665.850 333.750 666.750 ;
        RECT 328.950 664.950 331.050 665.400 ;
        RECT 334.950 664.950 337.050 667.050 ;
        RECT 338.250 665.850 340.050 666.750 ;
        RECT 334.950 662.850 337.050 663.750 ;
        RECT 331.950 646.950 334.050 649.050 ;
        RECT 322.950 640.950 325.050 643.050 ;
        RECT 328.950 640.950 331.050 643.050 ;
        RECT 313.950 637.950 316.050 640.050 ;
        RECT 316.950 637.950 319.050 640.050 ;
        RECT 298.950 635.250 301.050 636.150 ;
        RECT 307.950 634.950 310.050 637.050 ;
        RECT 295.950 632.250 297.750 633.150 ;
        RECT 298.950 631.950 301.050 634.050 ;
        RECT 302.250 632.250 303.750 633.150 ;
        RECT 304.950 631.950 307.050 634.050 ;
        RECT 295.950 628.950 298.050 631.050 ;
        RECT 299.400 625.050 300.450 631.950 ;
        RECT 301.950 628.950 304.050 631.050 ;
        RECT 305.250 629.850 307.050 630.750 ;
        RECT 308.400 628.050 309.450 634.950 ;
        RECT 310.950 631.950 313.050 634.050 ;
        RECT 307.950 625.950 310.050 628.050 ;
        RECT 298.950 622.950 301.050 625.050 ;
        RECT 295.950 613.950 298.050 616.050 ;
        RECT 307.950 613.950 310.050 616.050 ;
        RECT 296.400 598.050 297.450 613.950 ;
        RECT 298.950 607.950 301.050 610.050 ;
        RECT 304.950 607.950 307.050 610.050 ;
        RECT 299.400 601.050 300.450 607.950 ;
        RECT 305.400 601.050 306.450 607.950 ;
        RECT 298.950 598.950 301.050 601.050 ;
        RECT 302.250 599.250 303.750 600.150 ;
        RECT 304.950 598.950 307.050 601.050 ;
        RECT 295.950 595.950 298.050 598.050 ;
        RECT 299.250 596.850 300.750 597.750 ;
        RECT 301.950 595.950 304.050 598.050 ;
        RECT 305.250 596.850 307.050 597.750 ;
        RECT 295.950 593.850 298.050 594.750 ;
        RECT 302.400 592.050 303.450 595.950 ;
        RECT 295.950 589.950 298.050 592.050 ;
        RECT 301.950 589.950 304.050 592.050 ;
        RECT 292.950 553.950 295.050 556.050 ;
        RECT 296.400 553.050 297.450 589.950 ;
        RECT 308.400 571.050 309.450 613.950 ;
        RECT 311.400 598.050 312.450 631.950 ;
        RECT 314.400 630.450 315.450 637.950 ;
        RECT 319.950 635.250 322.050 636.150 ;
        RECT 325.950 634.950 328.050 637.050 ;
        RECT 326.400 634.050 327.450 634.950 ;
        RECT 316.950 632.250 318.750 633.150 ;
        RECT 319.950 631.950 322.050 634.050 ;
        RECT 323.250 632.250 324.750 633.150 ;
        RECT 325.950 631.950 328.050 634.050 ;
        RECT 316.950 630.450 319.050 631.050 ;
        RECT 314.400 629.400 319.050 630.450 ;
        RECT 316.950 628.950 319.050 629.400 ;
        RECT 313.950 625.950 316.050 628.050 ;
        RECT 316.950 625.950 319.050 628.050 ;
        RECT 310.950 595.950 313.050 598.050 ;
        RECT 307.950 568.950 310.050 571.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 298.950 562.950 301.050 565.050 ;
        RECT 299.400 559.050 300.450 562.950 ;
        RECT 304.950 559.950 307.050 562.050 ;
        RECT 307.950 559.950 310.050 562.050 ;
        RECT 298.950 556.950 301.050 559.050 ;
        RECT 301.950 557.250 304.050 558.150 ;
        RECT 301.950 555.450 304.050 556.050 ;
        RECT 305.400 555.450 306.450 559.950 ;
        RECT 308.400 559.050 309.450 559.950 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 298.950 554.250 300.750 555.150 ;
        RECT 301.950 554.400 306.450 555.450 ;
        RECT 307.950 554.850 310.050 555.750 ;
        RECT 301.950 553.950 304.050 554.400 ;
        RECT 295.950 550.950 298.050 553.050 ;
        RECT 298.950 550.950 301.050 553.050 ;
        RECT 304.950 550.950 307.050 553.050 ;
        RECT 299.400 550.050 300.450 550.950 ;
        RECT 289.950 547.950 292.050 550.050 ;
        RECT 298.950 547.950 301.050 550.050 ;
        RECT 283.950 544.950 286.050 547.050 ;
        RECT 274.950 526.950 277.050 529.050 ;
        RECT 275.400 526.050 276.450 526.950 ;
        RECT 271.950 524.250 273.750 525.150 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 278.400 523.050 279.450 523.950 ;
        RECT 271.950 520.950 274.050 523.050 ;
        RECT 275.250 521.850 276.750 522.750 ;
        RECT 277.950 520.950 280.050 523.050 ;
        RECT 281.250 521.850 283.050 522.750 ;
        RECT 277.950 518.850 280.050 519.750 ;
        RECT 284.400 496.050 285.450 544.950 ;
        RECT 298.950 532.950 301.050 535.050 ;
        RECT 286.950 529.950 289.050 532.050 ;
        RECT 292.950 529.950 295.050 532.050 ;
        RECT 287.400 526.050 288.450 529.950 ;
        RECT 299.400 529.050 300.450 532.950 ;
        RECT 289.950 527.250 292.050 528.150 ;
        RECT 292.950 527.850 295.050 528.750 ;
        RECT 295.950 527.250 297.750 528.150 ;
        RECT 298.950 526.950 301.050 529.050 ;
        RECT 301.950 526.950 304.050 529.050 ;
        RECT 302.400 526.050 303.450 526.950 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 289.950 523.950 292.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 299.250 524.850 301.050 525.750 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 277.950 493.950 280.050 496.050 ;
        RECT 283.950 493.950 286.050 496.050 ;
        RECT 271.950 490.950 274.050 493.050 ;
        RECT 272.400 487.050 273.450 490.950 ;
        RECT 262.950 485.250 264.750 486.150 ;
        RECT 265.950 484.950 268.050 487.050 ;
        RECT 268.950 484.950 271.050 487.050 ;
        RECT 271.950 484.950 274.050 487.050 ;
        RECT 262.950 481.950 265.050 484.050 ;
        RECT 266.250 482.850 268.050 483.750 ;
        RECT 268.950 482.250 271.050 483.150 ;
        RECT 271.950 482.850 274.050 483.750 ;
        RECT 263.400 475.050 264.450 481.950 ;
        RECT 268.950 478.950 271.050 481.050 ;
        RECT 268.950 475.950 271.050 478.050 ;
        RECT 262.950 472.950 265.050 475.050 ;
        RECT 260.400 467.400 264.450 468.450 ;
        RECT 259.950 460.950 262.050 463.050 ;
        RECT 244.950 452.850 246.750 453.750 ;
        RECT 247.950 451.950 250.050 454.050 ;
        RECT 253.950 451.950 256.050 454.050 ;
        RECT 256.950 451.950 259.050 454.050 ;
        RECT 248.400 445.050 249.450 451.950 ;
        RECT 254.400 451.050 255.450 451.950 ;
        RECT 253.950 448.950 256.050 451.050 ;
        RECT 253.950 445.950 256.050 448.050 ;
        RECT 257.400 447.450 258.450 451.950 ;
        RECT 260.400 451.050 261.450 460.950 ;
        RECT 259.950 448.950 262.050 451.050 ;
        RECT 257.400 446.400 261.450 447.450 ;
        RECT 247.950 442.950 250.050 445.050 ;
        RECT 241.950 430.950 244.050 433.050 ;
        RECT 244.950 413.250 247.050 414.150 ;
        RECT 250.950 413.250 253.050 414.150 ;
        RECT 244.950 409.950 247.050 412.050 ;
        RECT 248.250 410.250 249.750 411.150 ;
        RECT 250.950 409.950 253.050 412.050 ;
        RECT 251.400 409.050 252.450 409.950 ;
        RECT 247.950 406.950 250.050 409.050 ;
        RECT 250.950 406.950 253.050 409.050 ;
        RECT 248.400 406.050 249.450 406.950 ;
        RECT 238.950 403.950 241.050 406.050 ;
        RECT 244.950 403.950 247.050 406.050 ;
        RECT 247.950 403.950 250.050 406.050 ;
        RECT 238.950 397.950 241.050 400.050 ;
        RECT 235.950 394.950 238.050 397.050 ;
        RECT 235.950 391.950 238.050 394.050 ;
        RECT 221.400 383.400 225.450 384.450 ;
        RECT 224.400 382.050 225.450 383.400 ;
        RECT 220.950 380.250 222.750 381.150 ;
        RECT 223.950 379.950 226.050 382.050 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 220.950 376.950 223.050 379.050 ;
        RECT 224.250 377.850 225.750 378.750 ;
        RECT 226.950 376.950 229.050 379.050 ;
        RECT 230.250 377.850 232.050 378.750 ;
        RECT 232.950 376.950 235.050 379.050 ;
        RECT 221.400 376.050 222.450 376.950 ;
        RECT 220.950 373.950 223.050 376.050 ;
        RECT 226.950 374.850 229.050 375.750 ;
        RECT 229.950 373.950 232.050 376.050 ;
        RECT 223.950 367.950 226.050 370.050 ;
        RECT 217.950 355.950 220.050 358.050 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 191.250 344.250 192.750 345.150 ;
        RECT 193.950 343.950 196.050 346.050 ;
        RECT 197.250 344.250 199.050 345.150 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 211.950 343.950 214.050 346.050 ;
        RECT 214.950 343.950 217.050 346.050 ;
        RECT 187.950 341.850 189.750 342.750 ;
        RECT 190.950 340.950 193.050 343.050 ;
        RECT 194.400 337.050 195.450 343.950 ;
        RECT 196.950 342.450 199.050 343.050 ;
        RECT 200.400 342.450 201.450 343.950 ;
        RECT 212.400 343.050 213.450 343.950 ;
        RECT 218.400 343.050 219.450 355.950 ;
        RECT 220.950 343.950 223.050 346.050 ;
        RECT 196.950 341.400 201.450 342.450 ;
        RECT 196.950 340.950 199.050 341.400 ;
        RECT 208.950 341.250 210.750 342.150 ;
        RECT 211.950 340.950 214.050 343.050 ;
        RECT 217.950 340.950 220.050 343.050 ;
        RECT 208.950 337.950 211.050 340.050 ;
        RECT 212.250 338.850 214.050 339.750 ;
        RECT 214.950 338.250 217.050 339.150 ;
        RECT 217.950 338.850 220.050 339.750 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 193.950 331.950 196.050 334.050 ;
        RECT 176.400 329.400 180.450 330.450 ;
        RECT 176.400 271.050 177.450 329.400 ;
        RECT 190.950 313.950 193.050 316.050 ;
        RECT 181.950 310.950 184.050 313.050 ;
        RECT 185.250 311.250 186.750 312.150 ;
        RECT 187.950 310.950 190.050 313.050 ;
        RECT 191.400 310.050 192.450 313.950 ;
        RECT 178.950 307.950 181.050 310.050 ;
        RECT 182.250 308.850 183.750 309.750 ;
        RECT 184.950 307.950 187.050 310.050 ;
        RECT 188.250 308.850 190.050 309.750 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 178.950 305.850 181.050 306.750 ;
        RECT 184.950 274.950 187.050 277.050 ;
        RECT 178.950 272.250 181.050 273.150 ;
        RECT 185.400 271.050 186.450 274.950 ;
        RECT 175.950 268.950 178.050 271.050 ;
        RECT 178.950 268.950 181.050 271.050 ;
        RECT 182.250 269.250 183.750 270.150 ;
        RECT 184.950 268.950 187.050 271.050 ;
        RECT 188.250 269.250 190.050 270.150 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 179.400 265.050 180.450 268.950 ;
        RECT 181.950 265.950 184.050 268.050 ;
        RECT 185.250 266.850 186.750 267.750 ;
        RECT 187.950 265.950 190.050 268.050 ;
        RECT 178.950 262.950 181.050 265.050 ;
        RECT 172.950 238.950 175.050 241.050 ;
        RECT 172.950 236.250 174.750 237.150 ;
        RECT 175.950 235.950 178.050 238.050 ;
        RECT 179.250 236.250 181.050 237.150 ;
        RECT 172.950 234.450 175.050 235.050 ;
        RECT 170.400 233.400 175.050 234.450 ;
        RECT 176.250 233.850 177.750 234.750 ;
        RECT 172.950 232.950 175.050 233.400 ;
        RECT 178.950 232.950 181.050 235.050 ;
        RECT 172.950 203.250 175.050 204.150 ;
        RECT 169.950 200.250 171.750 201.150 ;
        RECT 172.950 199.950 175.050 202.050 ;
        RECT 176.250 200.250 177.750 201.150 ;
        RECT 178.950 199.950 181.050 202.050 ;
        RECT 169.950 196.950 172.050 199.050 ;
        RECT 173.400 196.050 174.450 199.950 ;
        RECT 182.400 199.050 183.450 265.950 ;
        RECT 191.400 241.050 192.450 268.950 ;
        RECT 194.400 247.050 195.450 331.950 ;
        RECT 202.950 316.950 205.050 319.050 ;
        RECT 203.400 313.050 204.450 316.950 ;
        RECT 209.400 316.050 210.450 337.950 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 211.950 331.950 214.050 334.050 ;
        RECT 208.950 313.950 211.050 316.050 ;
        RECT 202.950 310.950 205.050 313.050 ;
        RECT 206.250 311.250 207.750 312.150 ;
        RECT 208.950 310.950 211.050 313.050 ;
        RECT 199.950 309.450 202.050 310.050 ;
        RECT 197.400 308.400 202.050 309.450 ;
        RECT 203.250 308.850 204.750 309.750 ;
        RECT 197.400 259.050 198.450 308.400 ;
        RECT 199.950 307.950 202.050 308.400 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 209.250 308.850 211.050 309.750 ;
        RECT 199.950 305.850 202.050 306.750 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 199.950 268.950 202.050 271.050 ;
        RECT 209.400 268.050 210.450 289.950 ;
        RECT 199.950 266.850 202.050 267.750 ;
        RECT 202.950 266.250 205.050 267.150 ;
        RECT 208.950 265.950 211.050 268.050 ;
        RECT 202.950 264.450 205.050 265.050 ;
        RECT 202.950 263.400 207.450 264.450 ;
        RECT 202.950 262.950 205.050 263.400 ;
        RECT 202.950 259.950 205.050 262.050 ;
        RECT 196.950 256.950 199.050 259.050 ;
        RECT 196.950 250.950 199.050 253.050 ;
        RECT 193.950 244.950 196.050 247.050 ;
        RECT 193.950 241.950 196.050 244.050 ;
        RECT 197.400 241.050 198.450 250.950 ;
        RECT 199.950 241.950 202.050 244.050 ;
        RECT 190.950 240.450 193.050 241.050 ;
        RECT 188.400 239.400 193.050 240.450 ;
        RECT 194.250 239.850 195.750 240.750 ;
        RECT 188.400 235.050 189.450 239.400 ;
        RECT 190.950 238.950 193.050 239.400 ;
        RECT 196.950 238.950 199.050 241.050 ;
        RECT 190.950 236.850 193.050 237.750 ;
        RECT 196.950 236.850 199.050 237.750 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 196.950 232.950 199.050 235.050 ;
        RECT 187.950 226.950 190.050 229.050 ;
        RECT 188.400 201.450 189.450 226.950 ;
        RECT 197.400 202.050 198.450 232.950 ;
        RECT 190.950 201.450 193.050 202.050 ;
        RECT 188.400 200.400 193.050 201.450 ;
        RECT 175.950 196.950 178.050 199.050 ;
        RECT 179.250 197.850 181.050 198.750 ;
        RECT 181.950 196.950 184.050 199.050 ;
        RECT 172.950 193.950 175.050 196.050 ;
        RECT 188.400 193.050 189.450 200.400 ;
        RECT 190.950 199.950 193.050 200.400 ;
        RECT 194.250 200.250 195.750 201.150 ;
        RECT 196.950 199.950 199.050 202.050 ;
        RECT 190.950 197.850 192.750 198.750 ;
        RECT 193.950 196.950 196.050 199.050 ;
        RECT 197.250 197.850 199.050 198.750 ;
        RECT 194.400 196.050 195.450 196.950 ;
        RECT 193.950 193.950 196.050 196.050 ;
        RECT 160.950 191.400 165.450 192.450 ;
        RECT 160.950 190.950 163.050 191.400 ;
        RECT 187.950 190.950 190.050 193.050 ;
        RECT 196.950 190.950 199.050 193.050 ;
        RECT 169.950 172.950 172.050 175.050 ;
        RECT 133.950 169.950 136.050 172.050 ;
        RECT 139.950 169.950 142.050 172.050 ;
        RECT 148.950 169.950 151.050 172.050 ;
        RECT 140.400 169.050 141.450 169.950 ;
        RECT 124.950 166.950 127.050 169.050 ;
        RECT 130.950 167.250 133.050 168.150 ;
        RECT 133.950 167.850 136.050 168.750 ;
        RECT 136.950 167.250 138.750 168.150 ;
        RECT 139.950 166.950 142.050 169.050 ;
        RECT 157.950 166.950 160.050 169.050 ;
        RECT 163.950 168.450 166.050 169.050 ;
        RECT 161.250 167.250 162.750 168.150 ;
        RECT 163.950 167.400 168.450 168.450 ;
        RECT 163.950 166.950 166.050 167.400 ;
        RECT 106.950 164.850 108.750 165.750 ;
        RECT 109.950 163.950 112.050 166.050 ;
        RECT 113.250 164.850 114.750 165.750 ;
        RECT 115.950 163.950 118.050 166.050 ;
        RECT 88.950 160.950 91.050 163.050 ;
        RECT 92.250 161.850 93.750 162.750 ;
        RECT 94.950 160.950 97.050 163.050 ;
        RECT 98.250 161.850 100.050 162.750 ;
        RECT 100.950 160.950 103.050 163.050 ;
        RECT 103.950 160.950 106.050 163.050 ;
        RECT 94.950 158.850 97.050 159.750 ;
        RECT 101.400 154.050 102.450 160.950 ;
        RECT 94.950 151.950 97.050 154.050 ;
        RECT 100.950 151.950 103.050 154.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 82.950 127.950 85.050 130.050 ;
        RECT 83.400 127.050 84.450 127.950 ;
        RECT 73.950 125.250 75.750 126.150 ;
        RECT 76.950 124.950 79.050 127.050 ;
        RECT 82.950 124.950 85.050 127.050 ;
        RECT 92.400 124.050 93.450 133.950 ;
        RECT 95.400 130.050 96.450 151.950 ;
        RECT 110.400 136.050 111.450 163.950 ;
        RECT 115.950 161.850 118.050 162.750 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 100.950 131.250 103.050 132.150 ;
        RECT 94.950 127.950 97.050 130.050 ;
        RECT 98.250 128.250 99.750 129.150 ;
        RECT 100.950 127.950 103.050 130.050 ;
        RECT 104.250 128.250 106.050 129.150 ;
        RECT 106.950 127.950 109.050 130.050 ;
        RECT 118.950 127.950 121.050 130.050 ;
        RECT 94.950 125.850 96.750 126.750 ;
        RECT 97.950 124.950 100.050 127.050 ;
        RECT 103.950 126.450 106.050 127.050 ;
        RECT 101.400 125.400 106.050 126.450 ;
        RECT 73.950 121.950 76.050 124.050 ;
        RECT 77.250 122.850 79.050 123.750 ;
        RECT 79.950 122.250 82.050 123.150 ;
        RECT 82.950 122.850 85.050 123.750 ;
        RECT 91.950 121.950 94.050 124.050 ;
        RECT 79.950 118.950 82.050 121.050 ;
        RECT 98.400 118.050 99.450 124.950 ;
        RECT 97.950 115.950 100.050 118.050 ;
        RECT 101.400 115.050 102.450 125.400 ;
        RECT 103.950 124.950 106.050 125.400 ;
        RECT 107.400 123.450 108.450 127.950 ;
        RECT 119.400 127.050 120.450 127.950 ;
        RECT 112.950 126.450 115.050 127.050 ;
        RECT 104.400 122.400 108.450 123.450 ;
        RECT 110.400 125.400 115.050 126.450 ;
        RECT 100.950 112.950 103.050 115.050 ;
        RECT 97.950 97.950 100.050 100.050 ;
        RECT 104.400 97.050 105.450 122.400 ;
        RECT 110.400 118.050 111.450 125.400 ;
        RECT 112.950 124.950 115.050 125.400 ;
        RECT 118.950 124.950 121.050 127.050 ;
        RECT 122.250 125.250 124.050 126.150 ;
        RECT 112.950 122.850 115.050 123.750 ;
        RECT 115.950 122.250 118.050 123.150 ;
        RECT 118.950 122.850 120.750 123.750 ;
        RECT 121.950 121.950 124.050 124.050 ;
        RECT 115.950 118.950 118.050 121.050 ;
        RECT 109.950 115.950 112.050 118.050 ;
        RECT 116.400 115.050 117.450 118.950 ;
        RECT 115.950 112.950 118.050 115.050 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 85.950 96.450 88.050 97.050 ;
        RECT 83.250 95.250 84.750 96.150 ;
        RECT 85.950 95.400 90.450 96.450 ;
        RECT 85.950 94.950 88.050 95.400 ;
        RECT 89.400 94.050 90.450 95.400 ;
        RECT 94.950 95.250 97.050 96.150 ;
        RECT 97.950 95.850 100.050 96.750 ;
        RECT 100.950 95.250 102.750 96.150 ;
        RECT 103.950 94.950 106.050 97.050 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 80.250 92.850 81.750 93.750 ;
        RECT 82.950 91.950 85.050 94.050 ;
        RECT 86.250 92.850 88.050 93.750 ;
        RECT 88.950 91.950 91.050 94.050 ;
        RECT 94.950 91.950 97.050 94.050 ;
        RECT 100.950 91.950 103.050 94.050 ;
        RECT 104.250 92.850 106.050 93.750 ;
        RECT 115.950 92.250 117.750 93.150 ;
        RECT 118.950 91.950 121.050 94.050 ;
        RECT 122.250 92.250 124.050 93.150 ;
        RECT 76.950 89.850 79.050 90.750 ;
        RECT 76.950 79.950 79.050 82.050 ;
        RECT 77.400 58.050 78.450 79.950 ;
        RECT 83.400 64.050 84.450 91.950 ;
        RECT 82.950 61.950 85.050 64.050 ;
        RECT 82.950 59.250 85.050 60.150 ;
        RECT 76.950 55.950 79.050 58.050 ;
        RECT 80.250 56.250 81.750 57.150 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 86.250 56.250 88.050 57.150 ;
        RECT 76.950 53.850 78.750 54.750 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 70.950 34.950 73.050 37.050 ;
        RECT 71.400 22.050 72.450 34.950 ;
        RECT 76.950 31.950 79.050 34.050 ;
        RECT 77.400 22.050 78.450 31.950 ;
        RECT 83.400 31.050 84.450 55.950 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 86.400 37.050 87.450 52.950 ;
        RECT 89.400 40.050 90.450 91.950 ;
        RECT 95.400 91.050 96.450 91.950 ;
        RECT 94.950 88.950 97.050 91.050 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 119.250 89.850 120.750 90.750 ;
        RECT 121.950 90.450 124.050 91.050 ;
        RECT 125.400 90.450 126.450 166.950 ;
        RECT 167.400 166.050 168.450 167.400 ;
        RECT 130.950 163.950 133.050 166.050 ;
        RECT 136.950 165.450 139.050 166.050 ;
        RECT 134.400 164.400 139.050 165.450 ;
        RECT 140.250 164.850 142.050 165.750 ;
        RECT 134.400 163.050 135.450 164.400 ;
        RECT 136.950 163.950 139.050 164.400 ;
        RECT 154.950 163.950 157.050 166.050 ;
        RECT 158.250 164.850 159.750 165.750 ;
        RECT 160.950 163.950 163.050 166.050 ;
        RECT 164.250 164.850 166.050 165.750 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 133.950 160.950 136.050 163.050 ;
        RECT 154.950 161.850 157.050 162.750 ;
        RECT 161.400 162.450 162.450 163.950 ;
        RECT 166.950 162.450 169.050 163.050 ;
        RECT 161.400 161.400 169.050 162.450 ;
        RECT 166.950 160.950 169.050 161.400 ;
        RECT 130.950 130.950 133.050 133.050 ;
        RECT 127.950 124.950 130.050 127.050 ;
        RECT 128.400 91.050 129.450 124.950 ;
        RECT 121.950 89.400 126.450 90.450 ;
        RECT 121.950 88.950 124.050 89.400 ;
        RECT 127.950 88.950 130.050 91.050 ;
        RECT 116.400 88.050 117.450 88.950 ;
        RECT 100.950 85.950 103.050 88.050 ;
        RECT 115.950 85.950 118.050 88.050 ;
        RECT 101.400 58.050 102.450 85.950 ;
        RECT 122.400 61.050 123.450 88.950 ;
        RECT 109.950 58.950 112.050 61.050 ;
        RECT 121.950 58.950 124.050 61.050 ;
        RECT 124.950 59.250 127.050 60.150 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 97.950 53.250 100.050 54.150 ;
        RECT 100.950 53.850 103.050 54.750 ;
        RECT 106.950 53.250 109.050 54.150 ;
        RECT 97.950 49.950 100.050 52.050 ;
        RECT 106.950 51.450 109.050 52.050 ;
        RECT 110.400 51.450 111.450 58.950 ;
        RECT 118.950 55.950 121.050 58.050 ;
        RECT 122.250 56.250 123.750 57.150 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 128.250 56.250 130.050 57.150 ;
        RECT 118.950 53.850 120.750 54.750 ;
        RECT 121.950 52.950 124.050 55.050 ;
        RECT 106.950 50.400 111.450 51.450 ;
        RECT 106.950 49.950 109.050 50.400 ;
        RECT 122.400 43.050 123.450 52.950 ;
        RECT 121.950 40.950 124.050 43.050 ;
        RECT 88.950 37.950 91.050 40.050 ;
        RECT 85.950 34.950 88.050 37.050 ;
        RECT 82.950 28.950 85.050 31.050 ;
        RECT 100.950 28.950 103.050 31.050 ;
        RECT 79.950 25.950 82.050 28.050 ;
        RECT 85.950 25.950 88.050 28.050 ;
        RECT 94.950 25.950 97.050 28.050 ;
        RECT 80.400 25.050 81.450 25.950 ;
        RECT 86.400 25.050 87.450 25.950 ;
        RECT 95.400 25.050 96.450 25.950 ;
        RECT 101.400 25.050 102.450 28.950 ;
        RECT 79.950 22.950 82.050 25.050 ;
        RECT 83.250 23.250 84.750 24.150 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 98.250 23.250 99.750 24.150 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 122.400 22.050 123.450 40.950 ;
        RECT 125.400 34.050 126.450 55.950 ;
        RECT 127.950 54.450 130.050 55.050 ;
        RECT 131.400 54.450 132.450 130.950 ;
        RECT 134.400 124.050 135.450 160.950 ;
        RECT 163.950 131.250 166.050 132.150 ;
        RECT 170.400 130.050 171.450 172.950 ;
        RECT 178.950 169.950 181.050 172.050 ;
        RECT 190.950 169.950 193.050 172.050 ;
        RECT 197.400 169.050 198.450 190.950 ;
        RECT 200.400 172.050 201.450 241.950 ;
        RECT 199.950 169.950 202.050 172.050 ;
        RECT 175.950 167.250 178.050 168.150 ;
        RECT 178.950 167.850 181.050 168.750 ;
        RECT 181.950 166.950 184.050 169.050 ;
        RECT 187.950 167.250 190.050 168.150 ;
        RECT 190.950 167.850 193.050 168.750 ;
        RECT 193.950 167.250 195.750 168.150 ;
        RECT 196.950 166.950 199.050 169.050 ;
        RECT 175.950 163.950 178.050 166.050 ;
        RECT 172.950 162.450 175.050 163.050 ;
        RECT 176.400 162.450 177.450 163.950 ;
        RECT 172.950 161.400 177.450 162.450 ;
        RECT 172.950 160.950 175.050 161.400 ;
        RECT 182.400 133.050 183.450 166.950 ;
        RECT 187.950 163.950 190.050 166.050 ;
        RECT 193.950 163.950 196.050 166.050 ;
        RECT 197.250 164.850 199.050 165.750 ;
        RECT 188.400 163.050 189.450 163.950 ;
        RECT 187.950 160.950 190.050 163.050 ;
        RECT 187.950 157.950 190.050 160.050 ;
        RECT 181.950 130.950 184.050 133.050 ;
        RECT 157.950 129.450 160.050 130.050 ;
        RECT 136.950 128.250 139.050 129.150 ;
        RECT 155.400 128.400 160.050 129.450 ;
        RECT 136.950 124.950 139.050 127.050 ;
        RECT 140.250 125.250 141.750 126.150 ;
        RECT 142.950 124.950 145.050 127.050 ;
        RECT 146.250 125.250 148.050 126.150 ;
        RECT 151.950 124.950 154.050 127.050 ;
        RECT 152.400 124.050 153.450 124.950 ;
        RECT 133.950 121.950 136.050 124.050 ;
        RECT 139.950 121.950 142.050 124.050 ;
        RECT 143.250 122.850 144.750 123.750 ;
        RECT 145.950 121.950 148.050 124.050 ;
        RECT 151.950 121.950 154.050 124.050 ;
        RECT 140.400 121.050 141.450 121.950 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 142.950 115.950 145.050 118.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 140.400 94.050 141.450 100.950 ;
        RECT 143.400 97.050 144.450 115.950 ;
        RECT 146.400 100.050 147.450 121.950 ;
        RECT 145.950 97.950 148.050 100.050 ;
        RECT 148.950 97.950 151.050 100.050 ;
        RECT 149.400 97.050 150.450 97.950 ;
        RECT 142.950 94.950 145.050 97.050 ;
        RECT 146.250 95.250 147.750 96.150 ;
        RECT 148.950 94.950 151.050 97.050 ;
        RECT 152.400 94.050 153.450 121.950 ;
        RECT 155.400 115.050 156.450 128.400 ;
        RECT 157.950 127.950 160.050 128.400 ;
        RECT 161.250 128.250 162.750 129.150 ;
        RECT 163.950 127.950 166.050 130.050 ;
        RECT 167.250 128.250 169.050 129.150 ;
        RECT 169.950 127.950 172.050 130.050 ;
        RECT 184.950 128.250 187.050 129.150 ;
        RECT 157.950 125.850 159.750 126.750 ;
        RECT 160.950 124.950 163.050 127.050 ;
        RECT 164.400 121.050 165.450 127.950 ;
        RECT 170.400 127.050 171.450 127.950 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 169.950 124.950 172.050 127.050 ;
        RECT 175.950 125.250 177.750 126.150 ;
        RECT 178.950 124.950 181.050 127.050 ;
        RECT 182.250 125.250 183.750 126.150 ;
        RECT 184.950 124.950 187.050 127.050 ;
        RECT 163.950 118.950 166.050 121.050 ;
        RECT 154.950 112.950 157.050 115.050 ;
        RECT 164.400 97.050 165.450 118.950 ;
        RECT 167.400 117.450 168.450 124.950 ;
        RECT 170.400 121.050 171.450 124.950 ;
        RECT 175.950 121.950 178.050 124.050 ;
        RECT 179.250 122.850 180.750 123.750 ;
        RECT 181.950 121.950 184.050 124.050 ;
        RECT 176.400 121.050 177.450 121.950 ;
        RECT 185.400 121.050 186.450 124.950 ;
        RECT 169.950 118.950 172.050 121.050 ;
        RECT 175.950 118.950 178.050 121.050 ;
        RECT 184.950 118.950 187.050 121.050 ;
        RECT 167.400 116.400 171.450 117.450 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 163.950 94.950 166.050 97.050 ;
        RECT 164.400 94.050 165.450 94.950 ;
        RECT 139.950 91.950 142.050 94.050 ;
        RECT 143.250 92.850 144.750 93.750 ;
        RECT 145.950 91.950 148.050 94.050 ;
        RECT 149.250 92.850 151.050 93.750 ;
        RECT 151.950 91.950 154.050 94.050 ;
        RECT 160.950 92.250 162.750 93.150 ;
        RECT 163.950 91.950 166.050 94.050 ;
        RECT 139.950 89.850 142.050 90.750 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 143.400 55.050 144.450 55.950 ;
        RECT 146.400 55.050 147.450 91.950 ;
        RECT 167.400 91.050 168.450 100.950 ;
        RECT 170.400 94.050 171.450 116.400 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 182.400 100.050 183.450 100.950 ;
        RECT 181.950 97.950 184.050 100.050 ;
        RECT 188.400 97.050 189.450 157.950 ;
        RECT 193.950 154.950 196.050 157.050 ;
        RECT 194.400 124.050 195.450 154.950 ;
        RECT 200.400 133.050 201.450 169.950 ;
        RECT 203.400 157.050 204.450 259.950 ;
        RECT 206.400 259.050 207.450 263.400 ;
        RECT 212.400 262.050 213.450 331.950 ;
        RECT 221.400 322.050 222.450 343.950 ;
        RECT 224.400 340.050 225.450 367.950 ;
        RECT 226.950 340.950 229.050 343.050 ;
        RECT 223.950 337.950 226.050 340.050 ;
        RECT 227.400 334.050 228.450 340.950 ;
        RECT 230.400 339.450 231.450 373.950 ;
        RECT 233.400 373.050 234.450 376.950 ;
        RECT 236.400 376.050 237.450 391.950 ;
        RECT 239.400 388.050 240.450 397.950 ;
        RECT 238.950 385.950 241.050 388.050 ;
        RECT 238.950 383.850 241.050 384.750 ;
        RECT 241.950 383.250 244.050 384.150 ;
        RECT 241.950 379.950 244.050 382.050 ;
        RECT 245.400 379.050 246.450 403.950 ;
        RECT 247.950 396.450 250.050 397.050 ;
        RECT 251.400 396.450 252.450 406.950 ;
        RECT 247.950 395.400 252.450 396.450 ;
        RECT 247.950 394.950 250.050 395.400 ;
        RECT 254.400 391.050 255.450 445.950 ;
        RECT 247.950 388.950 250.050 391.050 ;
        RECT 253.950 388.950 256.050 391.050 ;
        RECT 248.400 384.450 249.450 388.950 ;
        RECT 260.400 385.050 261.450 446.400 ;
        RECT 263.400 406.050 264.450 467.400 ;
        RECT 269.400 457.050 270.450 475.950 ;
        RECT 274.950 469.950 277.050 472.050 ;
        RECT 275.400 457.050 276.450 469.950 ;
        RECT 268.950 454.950 271.050 457.050 ;
        RECT 272.250 455.250 273.750 456.150 ;
        RECT 274.950 454.950 277.050 457.050 ;
        RECT 265.950 451.950 268.050 454.050 ;
        RECT 269.250 452.850 270.750 453.750 ;
        RECT 271.950 451.950 274.050 454.050 ;
        RECT 275.250 452.850 277.050 453.750 ;
        RECT 265.950 449.850 268.050 450.750 ;
        RECT 268.950 417.450 271.050 418.050 ;
        RECT 268.950 416.400 273.450 417.450 ;
        RECT 268.950 415.950 271.050 416.400 ;
        RECT 272.400 415.050 273.450 416.400 ;
        RECT 265.950 413.250 268.050 414.150 ;
        RECT 268.950 413.850 271.050 414.750 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 274.950 413.250 277.050 414.150 ;
        RECT 265.950 409.950 268.050 412.050 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 275.400 409.050 276.450 409.950 ;
        RECT 274.950 406.950 277.050 409.050 ;
        RECT 262.950 403.950 265.050 406.050 ;
        RECT 268.950 403.950 271.050 406.050 ;
        RECT 265.950 397.950 268.050 400.050 ;
        RECT 248.400 383.400 252.450 384.450 ;
        RECT 244.950 376.950 247.050 379.050 ;
        RECT 235.950 373.950 238.050 376.050 ;
        RECT 232.950 370.950 235.050 373.050 ;
        RECT 244.950 352.950 247.050 355.050 ;
        RECT 238.950 346.950 241.050 349.050 ;
        RECT 232.950 344.250 235.050 345.150 ;
        RECT 239.400 343.050 240.450 346.950 ;
        RECT 232.950 340.950 235.050 343.050 ;
        RECT 236.250 341.250 237.750 342.150 ;
        RECT 238.950 340.950 241.050 343.050 ;
        RECT 242.250 341.250 244.050 342.150 ;
        RECT 230.400 338.400 234.450 339.450 ;
        RECT 226.950 331.950 229.050 334.050 ;
        RECT 220.950 319.950 223.050 322.050 ;
        RECT 226.950 313.950 229.050 316.050 ;
        RECT 220.950 310.950 223.050 313.050 ;
        RECT 224.250 311.250 226.050 312.150 ;
        RECT 226.950 311.850 229.050 312.750 ;
        RECT 229.950 311.250 232.050 312.150 ;
        RECT 220.950 308.850 222.750 309.750 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 229.950 307.950 232.050 310.050 ;
        RECT 220.950 295.950 223.050 298.050 ;
        RECT 214.950 272.250 217.050 273.150 ;
        RECT 221.400 271.050 222.450 295.950 ;
        RECT 233.400 291.450 234.450 338.400 ;
        RECT 235.950 337.950 238.050 340.050 ;
        RECT 239.250 338.850 240.750 339.750 ;
        RECT 241.950 337.950 244.050 340.050 ;
        RECT 236.400 337.050 237.450 337.950 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 242.400 334.050 243.450 337.950 ;
        RECT 241.950 331.950 244.050 334.050 ;
        RECT 238.950 319.950 241.050 322.050 ;
        RECT 235.950 316.950 238.050 319.050 ;
        RECT 236.400 292.050 237.450 316.950 ;
        RECT 230.400 290.400 234.450 291.450 ;
        RECT 214.950 268.950 217.050 271.050 ;
        RECT 218.250 269.250 219.750 270.150 ;
        RECT 220.950 268.950 223.050 271.050 ;
        RECT 224.250 269.250 226.050 270.150 ;
        RECT 215.400 265.050 216.450 268.950 ;
        RECT 230.400 268.050 231.450 290.400 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 239.400 273.450 240.450 319.950 ;
        RECT 245.400 310.050 246.450 352.950 ;
        RECT 247.950 349.950 250.050 352.050 ;
        RECT 248.400 313.050 249.450 349.950 ;
        RECT 251.400 313.050 252.450 383.400 ;
        RECT 253.950 382.950 256.050 385.050 ;
        RECT 257.250 383.250 258.750 384.150 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 253.950 380.850 255.750 381.750 ;
        RECT 256.950 379.950 259.050 382.050 ;
        RECT 260.250 380.850 261.750 381.750 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 257.400 378.450 258.450 379.950 ;
        RECT 254.400 377.400 258.450 378.450 ;
        RECT 262.950 377.850 265.050 378.750 ;
        RECT 254.400 370.050 255.450 377.400 ;
        RECT 256.950 373.950 259.050 376.050 ;
        RECT 253.950 367.950 256.050 370.050 ;
        RECT 257.400 352.050 258.450 373.950 ;
        RECT 259.950 372.450 262.050 373.050 ;
        RECT 262.950 372.450 265.050 373.050 ;
        RECT 259.950 371.400 265.050 372.450 ;
        RECT 259.950 370.950 262.050 371.400 ;
        RECT 262.950 370.950 265.050 371.400 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 256.950 349.950 259.050 352.050 ;
        RECT 256.950 343.950 259.050 346.050 ;
        RECT 257.400 343.050 258.450 343.950 ;
        RECT 260.400 343.050 261.450 367.950 ;
        RECT 262.950 352.950 265.050 355.050 ;
        RECT 263.400 343.050 264.450 352.950 ;
        RECT 253.950 341.250 255.750 342.150 ;
        RECT 256.950 340.950 259.050 343.050 ;
        RECT 259.950 340.950 262.050 343.050 ;
        RECT 262.950 340.950 265.050 343.050 ;
        RECT 253.950 337.950 256.050 340.050 ;
        RECT 257.250 338.850 259.050 339.750 ;
        RECT 259.950 338.250 262.050 339.150 ;
        RECT 262.950 338.850 265.050 339.750 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 263.400 334.050 264.450 334.950 ;
        RECT 262.950 331.950 265.050 334.050 ;
        RECT 256.950 328.950 259.050 331.050 ;
        RECT 253.950 313.950 256.050 316.050 ;
        RECT 247.950 310.950 250.050 313.050 ;
        RECT 250.950 310.950 253.050 313.050 ;
        RECT 241.950 308.250 243.750 309.150 ;
        RECT 244.950 307.950 247.050 310.050 ;
        RECT 248.400 309.450 249.450 310.950 ;
        RECT 250.950 309.450 253.050 310.050 ;
        RECT 248.400 308.400 253.050 309.450 ;
        RECT 250.950 307.950 253.050 308.400 ;
        RECT 254.400 307.050 255.450 313.950 ;
        RECT 241.950 304.950 244.050 307.050 ;
        RECT 245.250 305.850 246.750 306.750 ;
        RECT 247.950 304.950 250.050 307.050 ;
        RECT 251.250 305.850 253.050 306.750 ;
        RECT 253.950 304.950 256.050 307.050 ;
        RECT 242.400 304.050 243.450 304.950 ;
        RECT 241.950 301.950 244.050 304.050 ;
        RECT 247.950 302.850 250.050 303.750 ;
        RECT 250.950 301.950 253.050 304.050 ;
        RECT 236.400 272.400 240.450 273.450 ;
        RECT 236.400 271.050 237.450 272.400 ;
        RECT 241.950 272.250 244.050 273.150 ;
        RECT 232.950 269.250 234.750 270.150 ;
        RECT 235.950 268.950 238.050 271.050 ;
        RECT 239.250 269.250 240.750 270.150 ;
        RECT 241.950 268.950 244.050 271.050 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 242.400 268.050 243.450 268.950 ;
        RECT 217.950 265.950 220.050 268.050 ;
        RECT 221.250 266.850 222.750 267.750 ;
        RECT 223.950 265.950 226.050 268.050 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 232.950 265.950 235.050 268.050 ;
        RECT 236.250 266.850 237.750 267.750 ;
        RECT 238.950 265.950 241.050 268.050 ;
        RECT 241.950 265.950 244.050 268.050 ;
        RECT 214.950 262.950 217.050 265.050 ;
        RECT 211.950 259.950 214.050 262.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 214.950 250.950 217.050 253.050 ;
        RECT 205.950 238.950 208.050 241.050 ;
        RECT 206.400 214.050 207.450 238.950 ;
        RECT 211.950 236.850 214.050 237.750 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 215.400 204.450 216.450 250.950 ;
        RECT 218.400 244.050 219.450 265.950 ;
        RECT 226.950 262.950 229.050 265.050 ;
        RECT 223.950 259.950 226.050 262.050 ;
        RECT 217.950 241.950 220.050 244.050 ;
        RECT 217.950 240.450 220.050 241.050 ;
        RECT 217.950 239.400 222.450 240.450 ;
        RECT 217.950 238.950 220.050 239.400 ;
        RECT 217.950 236.850 220.050 237.750 ;
        RECT 221.400 235.050 222.450 239.400 ;
        RECT 220.950 232.950 223.050 235.050 ;
        RECT 212.400 203.400 216.450 204.450 ;
        RECT 212.400 202.050 213.450 203.400 ;
        RECT 211.950 199.950 214.050 202.050 ;
        RECT 215.250 200.250 216.750 201.150 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 211.950 197.850 213.750 198.750 ;
        RECT 214.950 196.950 217.050 199.050 ;
        RECT 218.250 197.850 220.050 198.750 ;
        RECT 215.400 175.050 216.450 196.950 ;
        RECT 214.950 172.950 217.050 175.050 ;
        RECT 205.950 169.950 208.050 172.050 ;
        RECT 214.950 171.450 217.050 172.050 ;
        RECT 214.950 170.400 219.450 171.450 ;
        RECT 214.950 169.950 217.050 170.400 ;
        RECT 206.400 166.050 207.450 169.950 ;
        RECT 211.950 167.250 214.050 168.150 ;
        RECT 214.950 167.850 217.050 168.750 ;
        RECT 205.950 163.950 208.050 166.050 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 212.400 163.050 213.450 163.950 ;
        RECT 218.400 163.050 219.450 170.400 ;
        RECT 211.950 160.950 214.050 163.050 ;
        RECT 217.950 160.950 220.050 163.050 ;
        RECT 202.950 154.950 205.050 157.050 ;
        RECT 199.950 130.950 202.050 133.050 ;
        RECT 205.950 131.250 208.050 132.150 ;
        RECT 214.950 130.950 217.050 133.050 ;
        RECT 199.950 129.450 202.050 130.050 ;
        RECT 197.400 128.400 202.050 129.450 ;
        RECT 193.950 121.950 196.050 124.050 ;
        RECT 172.950 94.950 175.050 97.050 ;
        RECT 178.950 95.250 181.050 96.150 ;
        RECT 181.950 95.850 184.050 96.750 ;
        RECT 184.950 95.250 186.750 96.150 ;
        RECT 187.950 94.950 190.050 97.050 ;
        RECT 169.950 91.950 172.050 94.050 ;
        RECT 160.950 88.950 163.050 91.050 ;
        RECT 164.250 89.850 165.750 90.750 ;
        RECT 166.950 88.950 169.050 91.050 ;
        RECT 170.250 89.850 172.050 90.750 ;
        RECT 166.950 86.850 169.050 87.750 ;
        RECT 173.400 82.050 174.450 94.950 ;
        RECT 178.950 91.950 181.050 94.050 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 188.250 92.850 190.050 93.750 ;
        RECT 179.400 91.050 180.450 91.950 ;
        RECT 178.950 88.950 181.050 91.050 ;
        RECT 197.400 88.050 198.450 128.400 ;
        RECT 199.950 127.950 202.050 128.400 ;
        RECT 203.250 128.250 204.750 129.150 ;
        RECT 205.950 127.950 208.050 130.050 ;
        RECT 209.250 128.250 211.050 129.150 ;
        RECT 211.950 127.950 214.050 130.050 ;
        RECT 199.950 125.850 201.750 126.750 ;
        RECT 202.950 124.950 205.050 127.050 ;
        RECT 208.950 126.450 211.050 127.050 ;
        RECT 212.400 126.450 213.450 127.950 ;
        RECT 208.950 125.400 213.450 126.450 ;
        RECT 208.950 124.950 211.050 125.400 ;
        RECT 199.950 109.950 202.050 112.050 ;
        RECT 196.950 85.950 199.050 88.050 ;
        RECT 184.950 82.950 187.050 85.050 ;
        RECT 166.950 79.950 169.050 82.050 ;
        RECT 172.950 79.950 175.050 82.050 ;
        RECT 151.950 61.950 154.050 64.050 ;
        RECT 127.950 53.400 132.450 54.450 ;
        RECT 127.950 52.950 130.050 53.400 ;
        RECT 139.950 53.250 141.750 54.150 ;
        RECT 142.950 52.950 145.050 55.050 ;
        RECT 145.950 52.950 148.050 55.050 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 124.950 31.950 127.050 34.050 ;
        RECT 128.400 31.050 129.450 52.950 ;
        RECT 139.950 49.950 142.050 52.050 ;
        RECT 143.250 50.850 145.050 51.750 ;
        RECT 145.950 50.250 148.050 51.150 ;
        RECT 148.950 50.850 151.050 51.750 ;
        RECT 145.950 46.950 148.050 49.050 ;
        RECT 146.400 46.050 147.450 46.950 ;
        RECT 145.950 43.950 148.050 46.050 ;
        RECT 152.400 34.050 153.450 61.950 ;
        RECT 160.950 59.250 163.050 60.150 ;
        RECT 167.400 58.050 168.450 79.950 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 157.950 56.250 159.750 57.150 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 164.250 56.250 165.750 57.150 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 155.400 42.450 156.450 55.950 ;
        RECT 157.950 52.950 160.050 55.050 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 167.250 53.850 169.050 54.750 ;
        RECT 181.950 54.450 184.050 55.050 ;
        RECT 179.400 53.400 184.050 54.450 ;
        RECT 158.400 46.050 159.450 52.950 ;
        RECT 157.950 43.950 160.050 46.050 ;
        RECT 179.400 43.050 180.450 53.400 ;
        RECT 181.950 52.950 184.050 53.400 ;
        RECT 181.950 50.850 184.050 51.750 ;
        RECT 185.400 48.450 186.450 82.950 ;
        RECT 187.950 53.250 190.050 54.150 ;
        RECT 200.400 52.050 201.450 109.950 ;
        RECT 208.950 97.950 211.050 100.050 ;
        RECT 202.950 94.950 205.050 97.050 ;
        RECT 206.250 95.250 208.050 96.150 ;
        RECT 208.950 95.850 211.050 96.750 ;
        RECT 211.950 95.250 214.050 96.150 ;
        RECT 202.950 92.850 204.750 93.750 ;
        RECT 205.950 91.950 208.050 94.050 ;
        RECT 211.950 91.950 214.050 94.050 ;
        RECT 206.400 85.050 207.450 91.950 ;
        RECT 212.400 88.050 213.450 91.950 ;
        RECT 211.950 85.950 214.050 88.050 ;
        RECT 205.950 82.950 208.050 85.050 ;
        RECT 208.950 59.250 211.050 60.150 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 206.250 56.250 207.750 57.150 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 212.250 56.250 214.050 57.150 ;
        RECT 202.950 53.850 204.750 54.750 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 211.950 52.950 214.050 55.050 ;
        RECT 212.400 52.050 213.450 52.950 ;
        RECT 187.950 49.950 190.050 52.050 ;
        RECT 191.250 50.250 193.050 51.150 ;
        RECT 199.950 49.950 202.050 52.050 ;
        RECT 211.950 49.950 214.050 52.050 ;
        RECT 182.400 47.400 186.450 48.450 ;
        RECT 155.400 41.400 159.450 42.450 ;
        RECT 136.950 31.950 139.050 34.050 ;
        RECT 151.950 31.950 154.050 34.050 ;
        RECT 127.950 28.950 130.050 31.050 ;
        RECT 128.400 22.050 129.450 28.950 ;
        RECT 137.400 28.050 138.450 31.950 ;
        RECT 130.950 25.950 133.050 28.050 ;
        RECT 133.950 25.950 136.050 28.050 ;
        RECT 136.950 25.950 139.050 28.050 ;
        RECT 131.400 22.050 132.450 25.950 ;
        RECT 64.950 20.400 69.450 21.450 ;
        RECT 64.950 19.950 67.050 20.400 ;
        RECT 70.950 19.950 73.050 22.050 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 80.250 20.850 81.750 21.750 ;
        RECT 82.950 19.950 85.050 22.050 ;
        RECT 86.250 20.850 88.050 21.750 ;
        RECT 94.950 20.850 96.750 21.750 ;
        RECT 97.950 19.950 100.050 22.050 ;
        RECT 101.250 20.850 102.750 21.750 ;
        RECT 103.950 19.950 106.050 22.050 ;
        RECT 118.950 20.250 120.750 21.150 ;
        RECT 121.950 19.950 124.050 22.050 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 127.950 19.950 130.050 22.050 ;
        RECT 130.950 19.950 133.050 22.050 ;
        RECT 10.950 16.950 13.050 19.050 ;
        RECT 14.250 17.850 15.750 18.750 ;
        RECT 16.950 16.950 19.050 19.050 ;
        RECT 20.250 17.850 22.050 18.750 ;
        RECT 22.950 16.950 25.050 19.050 ;
        RECT 25.950 16.950 28.050 19.050 ;
        RECT 29.400 16.050 30.450 19.950 ;
        RECT 35.400 19.050 36.450 19.950 ;
        RECT 125.400 19.050 126.450 19.950 ;
        RECT 134.400 19.050 135.450 25.950 ;
        RECT 152.400 25.050 153.450 31.950 ;
        RECT 158.400 25.050 159.450 41.400 ;
        RECT 160.950 40.950 163.050 43.050 ;
        RECT 178.950 40.950 181.050 43.050 ;
        RECT 136.950 23.850 139.050 24.750 ;
        RECT 139.950 23.250 142.050 24.150 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 155.250 23.250 156.750 24.150 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 140.400 19.050 141.450 19.950 ;
        RECT 143.400 19.050 144.450 22.950 ;
        RECT 161.400 22.050 162.450 40.950 ;
        RECT 169.950 28.950 172.050 31.050 ;
        RECT 151.950 20.850 153.750 21.750 ;
        RECT 154.950 19.950 157.050 22.050 ;
        RECT 158.250 20.850 159.750 21.750 ;
        RECT 160.950 19.950 163.050 22.050 ;
        RECT 170.400 21.450 171.450 28.950 ;
        RECT 175.950 25.950 178.050 28.050 ;
        RECT 182.400 25.050 183.450 47.400 ;
        RECT 190.950 46.950 193.050 49.050 ;
        RECT 184.950 25.950 187.050 28.050 ;
        RECT 172.950 23.250 175.050 24.150 ;
        RECT 175.950 23.850 178.050 24.750 ;
        RECT 178.950 23.250 180.750 24.150 ;
        RECT 181.950 22.950 184.050 25.050 ;
        RECT 185.400 22.050 186.450 25.950 ;
        RECT 191.400 25.050 192.450 46.950 ;
        RECT 200.400 28.050 201.450 49.950 ;
        RECT 215.400 30.450 216.450 130.950 ;
        RECT 218.400 130.050 219.450 160.950 ;
        RECT 224.400 160.050 225.450 259.950 ;
        RECT 227.400 175.050 228.450 262.950 ;
        RECT 239.400 253.050 240.450 265.950 ;
        RECT 238.950 250.950 241.050 253.050 ;
        RECT 245.400 244.050 246.450 268.950 ;
        RECT 235.950 241.950 238.050 244.050 ;
        RECT 244.950 241.950 247.050 244.050 ;
        RECT 251.400 241.050 252.450 301.950 ;
        RECT 257.400 298.050 258.450 328.950 ;
        RECT 263.400 315.450 264.450 331.950 ;
        RECT 266.400 319.050 267.450 397.950 ;
        RECT 269.400 385.050 270.450 403.950 ;
        RECT 268.950 382.950 271.050 385.050 ;
        RECT 271.950 382.950 274.050 385.050 ;
        RECT 268.950 379.950 271.050 382.050 ;
        RECT 269.400 376.050 270.450 379.950 ;
        RECT 268.950 373.950 271.050 376.050 ;
        RECT 272.400 373.050 273.450 382.950 ;
        RECT 275.400 381.450 276.450 406.950 ;
        RECT 278.400 391.050 279.450 493.950 ;
        RECT 287.400 492.450 288.450 523.950 ;
        RECT 290.400 520.050 291.450 523.950 ;
        RECT 296.400 523.050 297.450 523.950 ;
        RECT 295.950 520.950 298.050 523.050 ;
        RECT 289.950 517.950 292.050 520.050 ;
        RECT 290.400 496.050 291.450 517.950 ;
        RECT 298.950 505.950 301.050 508.050 ;
        RECT 289.950 493.950 292.050 496.050 ;
        RECT 284.400 491.400 288.450 492.450 ;
        RECT 284.400 481.050 285.450 491.400 ;
        RECT 286.950 487.950 289.050 490.050 ;
        RECT 292.950 489.450 295.050 490.050 ;
        RECT 290.250 488.250 291.750 489.150 ;
        RECT 292.950 488.400 297.450 489.450 ;
        RECT 292.950 487.950 295.050 488.400 ;
        RECT 286.950 485.850 288.750 486.750 ;
        RECT 289.950 484.950 292.050 487.050 ;
        RECT 293.250 485.850 295.050 486.750 ;
        RECT 290.400 481.050 291.450 484.950 ;
        RECT 283.950 478.950 286.050 481.050 ;
        RECT 289.950 478.950 292.050 481.050 ;
        RECT 283.950 472.950 286.050 475.050 ;
        RECT 284.400 457.050 285.450 472.950 ;
        RECT 289.950 460.950 292.050 463.050 ;
        RECT 290.400 457.050 291.450 460.950 ;
        RECT 296.400 460.050 297.450 488.400 ;
        RECT 295.950 457.950 298.050 460.050 ;
        RECT 283.950 456.450 286.050 457.050 ;
        RECT 281.400 455.400 286.050 456.450 ;
        RECT 281.400 454.050 282.450 455.400 ;
        RECT 283.950 454.950 286.050 455.400 ;
        RECT 287.250 455.250 288.750 456.150 ;
        RECT 289.950 454.950 292.050 457.050 ;
        RECT 280.950 451.950 283.050 454.050 ;
        RECT 283.950 452.850 285.750 453.750 ;
        RECT 286.950 451.950 289.050 454.050 ;
        RECT 290.250 452.850 291.750 453.750 ;
        RECT 292.950 453.450 295.050 454.050 ;
        RECT 292.950 452.400 297.450 453.450 ;
        RECT 292.950 451.950 295.050 452.400 ;
        RECT 292.950 449.850 295.050 450.750 ;
        RECT 296.400 448.050 297.450 452.400 ;
        RECT 295.950 445.950 298.050 448.050 ;
        RECT 295.950 439.950 298.050 442.050 ;
        RECT 286.950 427.950 289.050 430.050 ;
        RECT 287.400 400.050 288.450 427.950 ;
        RECT 289.950 418.950 292.050 421.050 ;
        RECT 290.400 418.050 291.450 418.950 ;
        RECT 296.400 418.050 297.450 439.950 ;
        RECT 299.400 421.050 300.450 505.950 ;
        RECT 302.400 493.050 303.450 523.950 ;
        RECT 305.400 517.050 306.450 550.950 ;
        RECT 307.950 526.950 310.050 529.050 ;
        RECT 304.950 514.950 307.050 517.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 302.400 457.050 303.450 490.950 ;
        RECT 308.400 487.050 309.450 526.950 ;
        RECT 311.400 496.050 312.450 568.950 ;
        RECT 314.400 559.050 315.450 625.950 ;
        RECT 313.950 556.950 316.050 559.050 ;
        RECT 317.400 556.050 318.450 625.950 ;
        RECT 320.400 625.050 321.450 631.950 ;
        RECT 329.400 631.050 330.450 640.950 ;
        RECT 322.950 628.950 325.050 631.050 ;
        RECT 326.250 629.850 328.050 630.750 ;
        RECT 328.950 628.950 331.050 631.050 ;
        RECT 319.950 622.950 322.050 625.050 ;
        RECT 323.400 607.050 324.450 628.950 ;
        RECT 322.950 604.950 325.050 607.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 319.950 596.250 321.750 597.150 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 326.400 595.050 327.450 601.950 ;
        RECT 328.950 595.950 331.050 598.050 ;
        RECT 319.950 592.950 322.050 595.050 ;
        RECT 323.250 593.850 324.750 594.750 ;
        RECT 325.950 592.950 328.050 595.050 ;
        RECT 329.250 593.850 331.050 594.750 ;
        RECT 325.950 590.850 328.050 591.750 ;
        RECT 319.950 562.950 322.050 565.050 ;
        RECT 320.400 562.050 321.450 562.950 ;
        RECT 319.950 559.950 322.050 562.050 ;
        RECT 323.250 560.250 324.750 561.150 ;
        RECT 325.950 559.950 328.050 562.050 ;
        RECT 319.950 557.850 321.750 558.750 ;
        RECT 322.950 556.950 325.050 559.050 ;
        RECT 326.250 557.850 328.050 558.750 ;
        RECT 313.950 553.950 316.050 556.050 ;
        RECT 316.950 553.950 319.050 556.050 ;
        RECT 314.400 552.450 315.450 553.950 ;
        RECT 314.400 551.400 318.450 552.450 ;
        RECT 317.400 529.050 318.450 551.400 ;
        RECT 323.400 532.050 324.450 556.950 ;
        RECT 332.400 544.050 333.450 646.950 ;
        RECT 334.950 634.950 337.050 637.050 ;
        RECT 335.400 628.050 336.450 634.950 ;
        RECT 341.400 633.450 342.450 682.950 ;
        RECT 349.950 668.250 351.750 669.150 ;
        RECT 352.950 667.950 355.050 670.050 ;
        RECT 356.250 668.250 358.050 669.150 ;
        RECT 349.950 664.950 352.050 667.050 ;
        RECT 353.250 665.850 354.750 666.750 ;
        RECT 355.950 666.450 358.050 667.050 ;
        RECT 359.400 666.450 360.450 697.950 ;
        RECT 368.400 688.050 369.450 742.950 ;
        RECT 373.950 740.250 375.750 741.150 ;
        RECT 376.950 739.950 379.050 742.050 ;
        RECT 380.400 739.050 381.450 773.400 ;
        RECT 383.400 772.050 384.450 778.950 ;
        RECT 389.400 775.050 390.450 814.950 ;
        RECT 401.400 814.050 402.450 814.950 ;
        RECT 391.950 812.250 393.750 813.150 ;
        RECT 394.950 811.950 397.050 814.050 ;
        RECT 400.950 811.950 403.050 814.050 ;
        RECT 391.950 808.950 394.050 811.050 ;
        RECT 395.250 809.850 396.750 810.750 ;
        RECT 397.950 808.950 400.050 811.050 ;
        RECT 401.250 809.850 403.050 810.750 ;
        RECT 397.950 806.850 400.050 807.750 ;
        RECT 404.400 804.450 405.450 844.950 ;
        RECT 410.400 841.050 411.450 844.950 ;
        RECT 409.950 838.950 412.050 841.050 ;
        RECT 416.400 835.050 417.450 844.950 ;
        RECT 415.950 832.950 418.050 835.050 ;
        RECT 415.950 829.950 418.050 832.050 ;
        RECT 416.400 814.050 417.450 829.950 ;
        RECT 412.950 812.250 414.750 813.150 ;
        RECT 415.950 811.950 418.050 814.050 ;
        RECT 419.400 811.050 420.450 847.950 ;
        RECT 422.400 835.050 423.450 848.400 ;
        RECT 424.950 847.950 427.050 848.400 ;
        RECT 428.250 848.250 429.750 849.150 ;
        RECT 430.950 847.950 433.050 850.050 ;
        RECT 460.950 848.250 463.050 849.150 ;
        RECT 487.950 847.950 490.050 850.050 ;
        RECT 514.950 847.950 517.050 850.050 ;
        RECT 523.950 847.950 526.050 850.050 ;
        RECT 527.250 848.250 528.750 849.150 ;
        RECT 529.950 847.950 532.050 850.050 ;
        RECT 533.250 848.250 535.050 849.150 ;
        RECT 598.950 848.250 601.050 849.150 ;
        RECT 613.950 847.950 616.050 850.050 ;
        RECT 625.950 849.600 628.050 851.700 ;
        RECT 424.950 845.850 426.750 846.750 ;
        RECT 427.950 844.950 430.050 847.050 ;
        RECT 431.250 845.850 433.050 846.750 ;
        RECT 445.950 844.950 448.050 847.050 ;
        RECT 460.950 844.950 463.050 847.050 ;
        RECT 464.250 845.250 465.750 846.150 ;
        RECT 466.950 844.950 469.050 847.050 ;
        RECT 470.250 845.250 472.050 846.150 ;
        RECT 484.950 845.250 487.050 846.150 ;
        RECT 487.950 845.850 490.050 846.750 ;
        RECT 493.950 845.250 496.050 846.150 ;
        RECT 505.950 845.250 508.050 846.150 ;
        RECT 511.950 845.250 514.050 846.150 ;
        RECT 421.950 832.950 424.050 835.050 ;
        RECT 422.400 814.050 423.450 832.950 ;
        RECT 428.400 820.050 429.450 844.950 ;
        RECT 445.950 842.850 448.050 843.750 ;
        RECT 448.950 842.250 451.050 843.150 ;
        RECT 463.950 841.950 466.050 844.050 ;
        RECT 467.250 842.850 468.750 843.750 ;
        RECT 469.950 841.950 472.050 844.050 ;
        RECT 484.950 841.950 487.050 844.050 ;
        RECT 493.950 841.950 496.050 844.050 ;
        RECT 505.950 841.950 508.050 844.050 ;
        RECT 511.950 843.450 514.050 844.050 ;
        RECT 515.400 843.450 516.450 847.950 ;
        RECT 614.400 847.050 615.450 847.950 ;
        RECT 523.950 845.850 525.750 846.750 ;
        RECT 526.950 844.950 529.050 847.050 ;
        RECT 532.950 844.950 535.050 847.050 ;
        RECT 547.950 844.950 550.050 847.050 ;
        RECT 562.950 846.450 565.050 847.050 ;
        RECT 560.400 845.400 565.050 846.450 ;
        RECT 509.250 842.250 510.750 843.150 ;
        RECT 511.950 842.400 516.450 843.450 ;
        RECT 511.950 841.950 514.050 842.400 ;
        RECT 448.950 838.950 451.050 841.050 ;
        RECT 449.400 832.050 450.450 838.950 ;
        RECT 430.950 829.950 433.050 832.050 ;
        RECT 448.950 829.950 451.050 832.050 ;
        RECT 427.950 817.950 430.050 820.050 ;
        RECT 428.400 814.050 429.450 817.950 ;
        RECT 431.400 817.050 432.450 829.950 ;
        RECT 439.950 820.950 442.050 823.050 ;
        RECT 436.950 817.950 439.050 820.050 ;
        RECT 437.400 817.050 438.450 817.950 ;
        RECT 430.950 814.950 433.050 817.050 ;
        RECT 434.250 815.250 435.750 816.150 ;
        RECT 436.950 814.950 439.050 817.050 ;
        RECT 440.400 814.050 441.450 820.950 ;
        RECT 451.950 817.950 454.050 820.050 ;
        RECT 464.400 817.050 465.450 841.950 ;
        RECT 470.400 841.050 471.450 841.950 ;
        RECT 469.950 838.950 472.050 841.050 ;
        RECT 508.950 838.950 511.050 841.050 ;
        RECT 509.400 829.050 510.450 838.950 ;
        RECT 508.950 826.950 511.050 829.050 ;
        RECT 487.950 817.950 490.050 820.050 ;
        RECT 451.950 815.850 454.050 816.750 ;
        RECT 454.950 815.250 457.050 816.150 ;
        RECT 463.950 814.950 466.050 817.050 ;
        RECT 488.400 814.050 489.450 817.950 ;
        RECT 515.400 817.050 516.450 842.400 ;
        RECT 523.950 841.950 526.050 844.050 ;
        RECT 524.400 819.450 525.450 841.950 ;
        RECT 529.950 820.950 532.050 823.050 ;
        RECT 526.950 819.450 529.050 820.050 ;
        RECT 524.400 818.400 529.050 819.450 ;
        RECT 490.950 814.950 493.050 817.050 ;
        RECT 505.950 814.950 508.050 817.050 ;
        RECT 514.950 814.950 517.050 817.050 ;
        RECT 421.950 811.950 424.050 814.050 ;
        RECT 427.950 811.950 430.050 814.050 ;
        RECT 430.950 812.850 432.750 813.750 ;
        RECT 433.950 811.950 436.050 814.050 ;
        RECT 437.250 812.850 438.750 813.750 ;
        RECT 439.950 811.950 442.050 814.050 ;
        RECT 454.950 811.950 457.050 814.050 ;
        RECT 466.950 812.250 468.750 813.150 ;
        RECT 469.950 811.950 472.050 814.050 ;
        RECT 473.250 812.250 475.050 813.150 ;
        RECT 475.950 811.950 478.050 814.050 ;
        RECT 487.950 811.950 490.050 814.050 ;
        RECT 455.400 811.050 456.450 811.950 ;
        RECT 412.950 808.950 415.050 811.050 ;
        RECT 416.250 809.850 417.750 810.750 ;
        RECT 418.950 808.950 421.050 811.050 ;
        RECT 422.250 809.850 424.050 810.750 ;
        RECT 439.950 809.850 442.050 810.750 ;
        RECT 454.950 808.950 457.050 811.050 ;
        RECT 466.950 808.950 469.050 811.050 ;
        RECT 470.250 809.850 471.750 810.750 ;
        RECT 472.950 808.950 475.050 811.050 ;
        RECT 473.400 808.050 474.450 808.950 ;
        RECT 418.950 806.850 421.050 807.750 ;
        RECT 472.950 805.950 475.050 808.050 ;
        RECT 401.400 803.400 405.450 804.450 ;
        RECT 388.950 772.950 391.050 775.050 ;
        RECT 382.950 769.950 385.050 772.050 ;
        RECT 388.950 770.850 391.050 771.750 ;
        RECT 391.950 770.250 394.050 771.150 ;
        RECT 401.400 769.050 402.450 803.400 ;
        RECT 403.950 776.250 406.050 777.150 ;
        RECT 421.950 775.950 424.050 778.050 ;
        RECT 451.950 777.450 454.050 778.050 ;
        RECT 427.950 776.250 430.050 777.150 ;
        RECT 451.950 776.400 456.450 777.450 ;
        RECT 451.950 775.950 454.050 776.400 ;
        RECT 403.950 772.950 406.050 775.050 ;
        RECT 407.250 773.250 408.750 774.150 ;
        RECT 409.950 772.950 412.050 775.050 ;
        RECT 413.250 773.250 415.050 774.150 ;
        RECT 382.950 766.950 385.050 769.050 ;
        RECT 391.950 766.950 394.050 769.050 ;
        RECT 400.950 766.950 403.050 769.050 ;
        RECT 383.400 742.050 384.450 766.950 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 398.400 748.050 399.450 757.950 ;
        RECT 404.400 754.050 405.450 772.950 ;
        RECT 406.950 769.950 409.050 772.050 ;
        RECT 410.250 770.850 411.750 771.750 ;
        RECT 412.950 769.950 415.050 772.050 ;
        RECT 407.400 769.050 408.450 769.950 ;
        RECT 406.950 766.950 409.050 769.050 ;
        RECT 403.950 751.950 406.050 754.050 ;
        RECT 413.400 748.050 414.450 769.950 ;
        RECT 397.950 745.950 400.050 748.050 ;
        RECT 412.950 745.950 415.050 748.050 ;
        RECT 415.950 745.950 418.050 748.050 ;
        RECT 394.950 743.250 397.050 744.150 ;
        RECT 397.950 743.850 400.050 744.750 ;
        RECT 416.400 742.050 417.450 745.950 ;
        RECT 382.950 741.450 385.050 742.050 ;
        RECT 382.950 740.400 387.450 741.450 ;
        RECT 382.950 739.950 385.050 740.400 ;
        RECT 373.950 736.950 376.050 739.050 ;
        RECT 377.250 737.850 378.750 738.750 ;
        RECT 379.950 736.950 382.050 739.050 ;
        RECT 383.250 737.850 385.050 738.750 ;
        RECT 379.950 734.850 382.050 735.750 ;
        RECT 386.400 735.450 387.450 740.400 ;
        RECT 394.950 739.950 397.050 742.050 ;
        RECT 412.950 740.250 414.750 741.150 ;
        RECT 415.950 739.950 418.050 742.050 ;
        RECT 419.250 740.250 421.050 741.150 ;
        RECT 388.950 736.950 391.050 739.050 ;
        RECT 412.950 736.950 415.050 739.050 ;
        RECT 416.250 737.850 417.750 738.750 ;
        RECT 418.950 736.950 421.050 739.050 ;
        RECT 383.400 734.400 387.450 735.450 ;
        RECT 379.950 730.950 382.050 733.050 ;
        RECT 380.400 709.050 381.450 730.950 ;
        RECT 379.950 706.950 382.050 709.050 ;
        RECT 380.400 706.050 381.450 706.950 ;
        RECT 373.950 703.950 376.050 706.050 ;
        RECT 377.250 704.250 378.750 705.150 ;
        RECT 379.950 703.950 382.050 706.050 ;
        RECT 373.950 701.850 375.750 702.750 ;
        RECT 376.950 700.950 379.050 703.050 ;
        RECT 380.250 701.850 382.050 702.750 ;
        RECT 377.400 691.050 378.450 700.950 ;
        RECT 376.950 688.950 379.050 691.050 ;
        RECT 367.950 685.950 370.050 688.050 ;
        RECT 373.950 676.950 376.050 679.050 ;
        RECT 370.950 673.950 373.050 676.050 ;
        RECT 371.400 670.050 372.450 673.950 ;
        RECT 361.950 667.950 364.050 670.050 ;
        RECT 364.950 667.950 367.050 670.050 ;
        RECT 367.950 668.250 369.750 669.150 ;
        RECT 370.950 667.950 373.050 670.050 ;
        RECT 355.950 665.400 360.450 666.450 ;
        RECT 355.950 664.950 358.050 665.400 ;
        RECT 350.400 664.050 351.450 664.950 ;
        RECT 349.950 661.950 352.050 664.050 ;
        RECT 350.400 661.050 351.450 661.950 ;
        RECT 349.950 658.950 352.050 661.050 ;
        RECT 349.950 652.950 352.050 655.050 ;
        RECT 338.400 632.400 342.450 633.450 ;
        RECT 334.950 625.950 337.050 628.050 ;
        RECT 338.400 616.050 339.450 632.400 ;
        RECT 340.950 629.250 343.050 630.150 ;
        RECT 346.950 629.250 349.050 630.150 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 344.250 626.250 345.750 627.150 ;
        RECT 346.950 625.950 349.050 628.050 ;
        RECT 343.950 622.950 346.050 625.050 ;
        RECT 347.400 616.050 348.450 625.950 ;
        RECT 350.400 625.050 351.450 652.950 ;
        RECT 355.950 649.950 358.050 652.050 ;
        RECT 352.950 637.950 355.050 640.050 ;
        RECT 353.400 628.050 354.450 637.950 ;
        RECT 352.950 625.950 355.050 628.050 ;
        RECT 349.950 622.950 352.050 625.050 ;
        RECT 337.950 613.950 340.050 616.050 ;
        RECT 346.950 613.950 349.050 616.050 ;
        RECT 340.950 601.950 343.050 604.050 ;
        RECT 334.950 597.450 337.050 598.050 ;
        RECT 337.950 597.450 340.050 598.050 ;
        RECT 334.950 596.400 340.050 597.450 ;
        RECT 334.950 595.950 337.050 596.400 ;
        RECT 337.950 595.950 340.050 596.400 ;
        RECT 335.400 558.450 336.450 595.950 ;
        RECT 341.400 595.050 342.450 601.950 ;
        RECT 356.400 601.050 357.450 649.950 ;
        RECT 359.400 634.050 360.450 665.400 ;
        RECT 362.400 649.050 363.450 667.950 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 365.400 646.050 366.450 667.950 ;
        RECT 374.400 667.050 375.450 676.950 ;
        RECT 376.950 667.950 379.050 670.050 ;
        RECT 383.400 669.450 384.450 734.400 ;
        RECT 389.400 730.050 390.450 736.950 ;
        RECT 419.400 736.050 420.450 736.950 ;
        RECT 418.950 733.950 421.050 736.050 ;
        RECT 388.950 727.950 391.050 730.050 ;
        RECT 385.950 703.950 388.050 706.050 ;
        RECT 386.400 700.050 387.450 703.950 ;
        RECT 385.950 697.950 388.050 700.050 ;
        RECT 389.400 685.050 390.450 727.950 ;
        RECT 397.950 709.950 400.050 712.050 ;
        RECT 394.950 701.250 397.050 702.150 ;
        RECT 394.950 697.950 397.050 700.050 ;
        RECT 388.950 682.950 391.050 685.050 ;
        RECT 385.950 676.950 388.050 679.050 ;
        RECT 386.400 670.050 387.450 676.950 ;
        RECT 391.950 673.950 394.050 676.050 ;
        RECT 392.400 670.050 393.450 673.950 ;
        RECT 380.400 668.400 384.450 669.450 ;
        RECT 367.950 664.950 370.050 667.050 ;
        RECT 371.250 665.850 372.750 666.750 ;
        RECT 373.950 664.950 376.050 667.050 ;
        RECT 377.250 665.850 379.050 666.750 ;
        RECT 368.400 652.050 369.450 664.950 ;
        RECT 373.950 662.850 376.050 663.750 ;
        RECT 367.950 649.950 370.050 652.050 ;
        RECT 364.950 643.950 367.050 646.050 ;
        RECT 367.950 637.950 370.050 640.050 ;
        RECT 376.950 637.950 379.050 640.050 ;
        RECT 358.950 631.950 361.050 634.050 ;
        RECT 361.950 632.250 364.050 633.150 ;
        RECT 368.400 631.050 369.450 637.950 ;
        RECT 373.950 634.950 376.050 637.050 ;
        RECT 361.950 628.950 364.050 631.050 ;
        RECT 365.250 629.250 366.750 630.150 ;
        RECT 367.950 628.950 370.050 631.050 ;
        RECT 371.250 629.250 373.050 630.150 ;
        RECT 362.400 622.050 363.450 628.950 ;
        RECT 364.950 625.950 367.050 628.050 ;
        RECT 368.250 626.850 369.750 627.750 ;
        RECT 370.950 625.950 373.050 628.050 ;
        RECT 371.400 625.050 372.450 625.950 ;
        RECT 370.950 622.950 373.050 625.050 ;
        RECT 361.950 619.950 364.050 622.050 ;
        RECT 358.950 616.950 361.050 619.050 ;
        RECT 343.950 598.950 346.050 601.050 ;
        RECT 349.950 598.950 352.050 601.050 ;
        RECT 355.950 598.950 358.050 601.050 ;
        RECT 344.400 598.050 345.450 598.950 ;
        RECT 343.950 595.950 346.050 598.050 ;
        RECT 347.250 596.250 349.050 597.150 ;
        RECT 337.950 593.850 339.750 594.750 ;
        RECT 340.950 592.950 343.050 595.050 ;
        RECT 344.250 593.850 345.750 594.750 ;
        RECT 346.950 592.950 349.050 595.050 ;
        RECT 340.950 590.850 343.050 591.750 ;
        RECT 350.400 565.050 351.450 598.950 ;
        RECT 359.400 583.050 360.450 616.950 ;
        RECT 361.950 613.950 364.050 616.050 ;
        RECT 362.400 598.050 363.450 613.950 ;
        RECT 374.400 612.450 375.450 634.950 ;
        RECT 377.400 619.050 378.450 637.950 ;
        RECT 376.950 616.950 379.050 619.050 ;
        RECT 374.400 611.400 378.450 612.450 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 364.950 598.950 367.050 601.050 ;
        RECT 368.250 599.250 369.750 600.150 ;
        RECT 370.950 598.950 373.050 601.050 ;
        RECT 374.400 598.050 375.450 601.950 ;
        RECT 361.950 595.950 364.050 598.050 ;
        RECT 365.250 596.850 366.750 597.750 ;
        RECT 367.950 595.950 370.050 598.050 ;
        RECT 371.250 596.850 373.050 597.750 ;
        RECT 373.950 595.950 376.050 598.050 ;
        RECT 361.950 593.850 364.050 594.750 ;
        RECT 368.400 589.050 369.450 595.950 ;
        RECT 377.400 595.050 378.450 611.400 ;
        RECT 373.950 592.950 376.050 595.050 ;
        RECT 376.950 592.950 379.050 595.050 ;
        RECT 367.950 586.950 370.050 589.050 ;
        RECT 358.950 580.950 361.050 583.050 ;
        RECT 367.950 580.950 370.050 583.050 ;
        RECT 370.950 580.950 373.050 583.050 ;
        RECT 355.950 571.950 358.050 574.050 ;
        RECT 340.950 563.250 343.050 564.150 ;
        RECT 349.950 562.950 352.050 565.050 ;
        RECT 337.950 560.250 339.750 561.150 ;
        RECT 340.950 559.950 343.050 562.050 ;
        RECT 344.250 560.250 345.750 561.150 ;
        RECT 346.950 559.950 349.050 562.050 ;
        RECT 341.400 559.050 342.450 559.950 ;
        RECT 337.950 558.450 340.050 559.050 ;
        RECT 335.400 557.400 340.050 558.450 ;
        RECT 337.950 556.950 340.050 557.400 ;
        RECT 340.950 556.950 343.050 559.050 ;
        RECT 343.950 556.950 346.050 559.050 ;
        RECT 347.250 557.850 349.050 558.750 ;
        RECT 338.400 550.050 339.450 556.950 ;
        RECT 337.950 547.950 340.050 550.050 ;
        RECT 331.950 541.950 334.050 544.050 ;
        RECT 337.950 535.950 340.050 538.050 ;
        RECT 322.950 529.950 325.050 532.050 ;
        RECT 325.950 529.950 328.050 532.050 ;
        RECT 328.950 529.950 331.050 532.050 ;
        RECT 338.400 531.450 339.450 535.950 ;
        RECT 341.400 535.050 342.450 556.950 ;
        RECT 344.400 556.050 345.450 556.950 ;
        RECT 343.950 553.950 346.050 556.050 ;
        RECT 350.400 555.450 351.450 562.950 ;
        RECT 347.400 554.400 351.450 555.450 ;
        RECT 340.950 532.950 343.050 535.050 ;
        RECT 338.400 530.400 342.450 531.450 ;
        RECT 316.950 526.950 319.050 529.050 ;
        RECT 320.250 527.250 321.750 528.150 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 326.400 526.050 327.450 529.950 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 317.250 524.850 318.750 525.750 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 323.250 524.850 325.050 525.750 ;
        RECT 325.950 523.950 328.050 526.050 ;
        RECT 313.950 521.850 316.050 522.750 ;
        RECT 316.950 508.950 319.050 511.050 ;
        RECT 310.950 493.950 313.050 496.050 ;
        RECT 304.950 485.250 306.750 486.150 ;
        RECT 307.950 484.950 310.050 487.050 ;
        RECT 313.950 484.950 316.050 487.050 ;
        RECT 304.950 481.950 307.050 484.050 ;
        RECT 308.250 482.850 310.050 483.750 ;
        RECT 310.950 482.250 313.050 483.150 ;
        RECT 313.950 482.850 316.050 483.750 ;
        RECT 305.400 472.050 306.450 481.950 ;
        RECT 310.950 480.450 313.050 481.050 ;
        RECT 310.950 479.400 315.450 480.450 ;
        RECT 310.950 478.950 313.050 479.400 ;
        RECT 304.950 469.950 307.050 472.050 ;
        RECT 304.950 460.950 307.050 463.050 ;
        RECT 301.950 454.950 304.050 457.050 ;
        RECT 305.400 430.050 306.450 460.950 ;
        RECT 310.950 457.950 313.050 460.050 ;
        RECT 311.400 454.050 312.450 457.950 ;
        RECT 314.400 457.050 315.450 479.400 ;
        RECT 317.400 463.050 318.450 508.950 ;
        RECT 329.400 493.050 330.450 529.950 ;
        RECT 341.400 529.050 342.450 530.400 ;
        RECT 334.950 528.450 337.050 529.050 ;
        RECT 332.400 527.400 337.050 528.450 ;
        RECT 332.400 523.050 333.450 527.400 ;
        RECT 334.950 526.950 337.050 527.400 ;
        RECT 338.250 527.250 339.750 528.150 ;
        RECT 340.950 526.950 343.050 529.050 ;
        RECT 343.950 526.950 346.050 529.050 ;
        RECT 344.400 526.050 345.450 526.950 ;
        RECT 334.950 524.850 336.750 525.750 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 341.250 524.850 342.750 525.750 ;
        RECT 343.950 523.950 346.050 526.050 ;
        RECT 331.950 520.950 334.050 523.050 ;
        RECT 343.950 521.850 346.050 522.750 ;
        RECT 347.400 522.450 348.450 554.400 ;
        RECT 349.950 529.950 352.050 532.050 ;
        RECT 350.400 526.050 351.450 529.950 ;
        RECT 352.950 526.950 355.050 529.050 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 347.400 521.400 351.450 522.450 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 319.950 489.450 322.050 490.050 ;
        RECT 322.950 489.450 325.050 490.050 ;
        RECT 319.950 488.400 325.050 489.450 ;
        RECT 319.950 487.950 322.050 488.400 ;
        RECT 322.950 487.950 325.050 488.400 ;
        RECT 326.250 488.250 327.750 489.150 ;
        RECT 328.950 487.950 331.050 490.050 ;
        RECT 320.400 466.050 321.450 487.950 ;
        RECT 322.950 485.850 324.750 486.750 ;
        RECT 325.950 484.950 328.050 487.050 ;
        RECT 329.250 485.850 331.050 486.750 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 325.950 466.950 328.050 469.050 ;
        RECT 319.950 463.950 322.050 466.050 ;
        RECT 316.950 460.950 319.050 463.050 ;
        RECT 313.950 454.950 316.050 457.050 ;
        RECT 319.950 456.450 322.050 457.050 ;
        RECT 317.250 455.250 318.750 456.150 ;
        RECT 319.950 455.400 324.450 456.450 ;
        RECT 319.950 454.950 322.050 455.400 ;
        RECT 310.950 451.950 313.050 454.050 ;
        RECT 314.250 452.850 315.750 453.750 ;
        RECT 316.950 451.950 319.050 454.050 ;
        RECT 320.250 452.850 322.050 453.750 ;
        RECT 323.400 451.050 324.450 455.400 ;
        RECT 310.950 449.850 313.050 450.750 ;
        RECT 322.950 448.950 325.050 451.050 ;
        RECT 319.950 433.950 322.050 436.050 ;
        RECT 304.950 427.950 307.050 430.050 ;
        RECT 307.950 421.950 310.050 424.050 ;
        RECT 316.950 421.950 319.050 424.050 ;
        RECT 298.950 418.950 301.050 421.050 ;
        RECT 289.950 415.950 292.050 418.050 ;
        RECT 293.250 416.250 294.750 417.150 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 289.950 413.850 291.750 414.750 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 296.250 413.850 298.050 414.750 ;
        RECT 299.400 412.050 300.450 418.950 ;
        RECT 301.950 415.950 304.050 418.050 ;
        RECT 292.950 409.950 295.050 412.050 ;
        RECT 298.950 409.950 301.050 412.050 ;
        RECT 302.400 411.450 303.450 415.950 ;
        RECT 308.400 415.050 309.450 421.950 ;
        RECT 313.950 416.250 316.050 417.150 ;
        RECT 304.950 413.250 306.750 414.150 ;
        RECT 307.950 412.950 310.050 415.050 ;
        RECT 311.250 413.250 312.750 414.150 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 304.950 411.450 307.050 412.050 ;
        RECT 302.400 410.400 307.050 411.450 ;
        RECT 308.250 410.850 309.750 411.750 ;
        RECT 304.950 409.950 307.050 410.400 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 286.950 397.950 289.050 400.050 ;
        RECT 286.950 391.950 289.050 394.050 ;
        RECT 277.950 388.950 280.050 391.050 ;
        RECT 287.400 385.050 288.450 391.950 ;
        RECT 289.950 388.950 292.050 391.050 ;
        RECT 280.950 382.950 283.050 385.050 ;
        RECT 284.250 383.250 285.750 384.150 ;
        RECT 286.950 382.950 289.050 385.050 ;
        RECT 277.950 381.450 280.050 382.050 ;
        RECT 275.400 380.400 280.050 381.450 ;
        RECT 281.250 380.850 282.750 381.750 ;
        RECT 275.400 373.050 276.450 380.400 ;
        RECT 277.950 379.950 280.050 380.400 ;
        RECT 283.950 379.950 286.050 382.050 ;
        RECT 287.250 380.850 289.050 381.750 ;
        RECT 277.950 377.850 280.050 378.750 ;
        RECT 284.400 378.450 285.450 379.950 ;
        RECT 281.400 377.400 285.450 378.450 ;
        RECT 268.950 370.950 271.050 373.050 ;
        RECT 271.950 370.950 274.050 373.050 ;
        RECT 274.950 370.950 277.050 373.050 ;
        RECT 269.400 340.050 270.450 370.950 ;
        RECT 281.400 370.050 282.450 377.400 ;
        RECT 283.950 370.950 286.050 373.050 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 280.950 367.950 283.050 370.050 ;
        RECT 268.950 337.950 271.050 340.050 ;
        RECT 272.400 334.050 273.450 367.950 ;
        RECT 281.400 367.050 282.450 367.950 ;
        RECT 280.950 364.950 283.050 367.050 ;
        RECT 274.950 349.950 277.050 352.050 ;
        RECT 275.400 346.050 276.450 349.950 ;
        RECT 284.400 348.450 285.450 370.950 ;
        RECT 280.950 347.250 283.050 348.150 ;
        RECT 284.400 347.400 288.450 348.450 ;
        RECT 287.400 346.050 288.450 347.400 ;
        RECT 274.950 343.950 277.050 346.050 ;
        RECT 278.250 344.250 279.750 345.150 ;
        RECT 280.950 343.950 283.050 346.050 ;
        RECT 284.250 344.250 286.050 345.150 ;
        RECT 286.950 343.950 289.050 346.050 ;
        RECT 274.950 341.850 276.750 342.750 ;
        RECT 277.950 340.950 280.050 343.050 ;
        RECT 280.950 340.950 283.050 343.050 ;
        RECT 283.950 342.450 286.050 343.050 ;
        RECT 283.950 341.400 288.450 342.450 ;
        RECT 283.950 340.950 286.050 341.400 ;
        RECT 271.950 331.950 274.050 334.050 ;
        RECT 271.950 328.950 274.050 331.050 ;
        RECT 265.950 316.950 268.050 319.050 ;
        RECT 260.400 314.400 264.450 315.450 ;
        RECT 260.400 313.050 261.450 314.400 ;
        RECT 265.950 313.950 268.050 316.050 ;
        RECT 266.400 313.050 267.450 313.950 ;
        RECT 259.950 310.950 262.050 313.050 ;
        RECT 263.250 311.250 264.750 312.150 ;
        RECT 265.950 310.950 268.050 313.050 ;
        RECT 259.950 308.850 261.750 309.750 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 266.250 308.850 267.750 309.750 ;
        RECT 268.950 309.450 271.050 310.050 ;
        RECT 272.400 309.450 273.450 328.950 ;
        RECT 274.950 325.950 277.050 328.050 ;
        RECT 268.950 308.400 273.450 309.450 ;
        RECT 268.950 307.950 271.050 308.400 ;
        RECT 263.400 307.050 264.450 307.950 ;
        RECT 262.950 304.950 265.050 307.050 ;
        RECT 268.950 305.850 271.050 306.750 ;
        RECT 256.950 295.950 259.050 298.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 253.950 277.950 256.050 280.050 ;
        RECT 254.400 270.450 255.450 277.950 ;
        RECT 256.950 272.250 259.050 273.150 ;
        RECT 263.400 271.050 264.450 289.950 ;
        RECT 256.950 270.450 259.050 271.050 ;
        RECT 254.400 269.400 259.050 270.450 ;
        RECT 256.950 268.950 259.050 269.400 ;
        RECT 260.250 269.250 261.750 270.150 ;
        RECT 262.950 268.950 265.050 271.050 ;
        RECT 266.250 269.250 268.050 270.150 ;
        RECT 257.400 241.050 258.450 268.950 ;
        RECT 259.950 265.950 262.050 268.050 ;
        RECT 263.250 266.850 264.750 267.750 ;
        RECT 265.950 265.950 268.050 268.050 ;
        RECT 260.400 244.050 261.450 265.950 ;
        RECT 266.400 265.050 267.450 265.950 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 272.400 262.050 273.450 308.400 ;
        RECT 275.400 304.050 276.450 325.950 ;
        RECT 281.400 325.050 282.450 340.950 ;
        RECT 287.400 340.050 288.450 341.400 ;
        RECT 283.950 337.950 286.050 340.050 ;
        RECT 286.950 337.950 289.050 340.050 ;
        RECT 284.400 328.050 285.450 337.950 ;
        RECT 283.950 325.950 286.050 328.050 ;
        RECT 280.950 322.950 283.050 325.050 ;
        RECT 290.400 319.050 291.450 388.950 ;
        RECT 277.950 316.950 280.050 319.050 ;
        RECT 289.950 316.950 292.050 319.050 ;
        RECT 274.950 301.950 277.050 304.050 ;
        RECT 274.950 292.950 277.050 295.050 ;
        RECT 275.400 265.050 276.450 292.950 ;
        RECT 278.400 280.050 279.450 316.950 ;
        RECT 283.950 313.950 286.050 316.050 ;
        RECT 280.950 311.250 283.050 312.150 ;
        RECT 283.950 311.850 286.050 312.750 ;
        RECT 286.950 311.250 288.750 312.150 ;
        RECT 289.950 310.950 292.050 313.050 ;
        RECT 280.950 307.950 283.050 310.050 ;
        RECT 286.950 307.950 289.050 310.050 ;
        RECT 290.250 308.850 292.050 309.750 ;
        RECT 286.950 286.950 289.050 289.050 ;
        RECT 277.950 277.950 280.050 280.050 ;
        RECT 277.950 271.950 280.050 274.050 ;
        RECT 283.950 273.450 286.050 274.050 ;
        RECT 287.400 273.450 288.450 286.950 ;
        RECT 289.950 280.950 292.050 283.050 ;
        RECT 281.250 272.250 282.750 273.150 ;
        RECT 283.950 272.400 288.450 273.450 ;
        RECT 283.950 271.950 286.050 272.400 ;
        RECT 277.950 269.850 279.750 270.750 ;
        RECT 280.950 268.950 283.050 271.050 ;
        RECT 284.250 269.850 286.050 270.750 ;
        RECT 274.950 262.950 277.050 265.050 ;
        RECT 271.950 259.950 274.050 262.050 ;
        RECT 281.400 259.050 282.450 268.950 ;
        RECT 280.950 256.950 283.050 259.050 ;
        RECT 277.950 253.950 280.050 256.050 ;
        RECT 268.950 250.950 271.050 253.050 ;
        RECT 259.950 241.950 262.050 244.050 ;
        RECT 232.950 239.250 235.050 240.150 ;
        RECT 235.950 239.850 238.050 240.750 ;
        RECT 238.950 238.950 241.050 241.050 ;
        RECT 244.950 238.950 247.050 241.050 ;
        RECT 248.250 239.250 249.750 240.150 ;
        RECT 250.950 238.950 253.050 241.050 ;
        RECT 256.950 240.450 259.050 241.050 ;
        RECT 254.250 239.250 255.750 240.150 ;
        RECT 256.950 239.400 261.450 240.450 ;
        RECT 256.950 238.950 259.050 239.400 ;
        RECT 232.950 235.950 235.050 238.050 ;
        RECT 233.400 204.450 234.450 235.950 ;
        RECT 230.400 203.400 234.450 204.450 ;
        RECT 230.400 202.050 231.450 203.400 ;
        RECT 229.950 199.950 232.050 202.050 ;
        RECT 235.950 201.450 238.050 202.050 ;
        RECT 239.400 201.450 240.450 238.950 ;
        RECT 244.950 236.850 246.750 237.750 ;
        RECT 247.950 235.950 250.050 238.050 ;
        RECT 251.250 236.850 252.750 237.750 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 257.250 236.850 259.050 237.750 ;
        RECT 254.400 208.050 255.450 235.950 ;
        RECT 253.950 205.950 256.050 208.050 ;
        RECT 260.400 205.050 261.450 239.400 ;
        RECT 265.950 239.250 268.050 240.150 ;
        RECT 265.950 235.950 268.050 238.050 ;
        RECT 266.400 235.050 267.450 235.950 ;
        RECT 265.950 232.950 268.050 235.050 ;
        RECT 269.400 228.450 270.450 250.950 ;
        RECT 274.950 241.950 277.050 244.050 ;
        RECT 266.400 227.400 270.450 228.450 ;
        RECT 262.950 205.950 265.050 208.050 ;
        RECT 256.950 203.250 259.050 204.150 ;
        RECT 259.950 202.950 262.050 205.050 ;
        RECT 233.250 200.250 234.750 201.150 ;
        RECT 235.950 200.400 240.450 201.450 ;
        RECT 235.950 199.950 238.050 200.400 ;
        RECT 229.950 197.850 231.750 198.750 ;
        RECT 232.950 196.950 235.050 199.050 ;
        RECT 236.250 197.850 238.050 198.750 ;
        RECT 232.950 175.950 235.050 178.050 ;
        RECT 226.950 172.950 229.050 175.050 ;
        RECT 227.400 169.050 228.450 172.950 ;
        RECT 229.950 169.950 232.050 172.050 ;
        RECT 233.400 169.050 234.450 175.950 ;
        RECT 226.950 166.950 229.050 169.050 ;
        RECT 230.250 167.850 231.750 168.750 ;
        RECT 232.950 166.950 235.050 169.050 ;
        RECT 226.950 164.850 229.050 165.750 ;
        RECT 229.950 163.950 232.050 166.050 ;
        RECT 232.950 164.850 235.050 165.750 ;
        RECT 223.950 157.950 226.050 160.050 ;
        RECT 217.950 127.950 220.050 130.050 ;
        RECT 220.950 127.950 223.050 130.050 ;
        RECT 221.400 127.050 222.450 127.950 ;
        RECT 220.950 124.950 223.050 127.050 ;
        RECT 217.950 122.250 220.050 123.150 ;
        RECT 220.950 122.850 223.050 123.750 ;
        RECT 217.950 118.950 220.050 121.050 ;
        RECT 217.950 103.950 220.050 106.050 ;
        RECT 218.400 55.050 219.450 103.950 ;
        RECT 230.400 103.050 231.450 163.950 ;
        RECT 239.400 133.050 240.450 200.400 ;
        RECT 250.950 199.950 253.050 202.050 ;
        RECT 254.250 200.250 255.750 201.150 ;
        RECT 256.950 199.950 259.050 202.050 ;
        RECT 260.250 200.250 262.050 201.150 ;
        RECT 250.950 197.850 252.750 198.750 ;
        RECT 253.950 196.950 256.050 199.050 ;
        RECT 259.950 198.450 262.050 199.050 ;
        RECT 263.400 198.450 264.450 205.950 ;
        RECT 259.950 197.400 264.450 198.450 ;
        RECT 259.950 196.950 262.050 197.400 ;
        RECT 241.950 175.950 244.050 178.050 ;
        RECT 238.950 130.950 241.050 133.050 ;
        RECT 239.400 130.050 240.450 130.950 ;
        RECT 232.950 127.950 235.050 130.050 ;
        RECT 236.250 128.250 237.750 129.150 ;
        RECT 238.950 127.950 241.050 130.050 ;
        RECT 232.950 125.850 234.750 126.750 ;
        RECT 235.950 124.950 238.050 127.050 ;
        RECT 239.250 125.850 241.050 126.750 ;
        RECT 242.400 121.050 243.450 175.950 ;
        RECT 244.950 172.950 247.050 175.050 ;
        RECT 245.400 172.050 246.450 172.950 ;
        RECT 244.950 169.950 247.050 172.050 ;
        RECT 244.950 167.850 247.050 168.750 ;
        RECT 247.950 167.250 250.050 168.150 ;
        RECT 266.400 166.050 267.450 227.400 ;
        RECT 268.950 205.950 271.050 208.050 ;
        RECT 269.400 202.050 270.450 205.950 ;
        RECT 275.400 202.050 276.450 241.950 ;
        RECT 278.400 238.050 279.450 253.950 ;
        RECT 287.400 253.050 288.450 272.400 ;
        RECT 290.400 262.050 291.450 280.950 ;
        RECT 293.400 274.050 294.450 409.950 ;
        RECT 295.950 385.950 298.050 388.050 ;
        RECT 307.950 385.950 310.050 388.050 ;
        RECT 296.400 385.050 297.450 385.950 ;
        RECT 295.950 382.950 298.050 385.050 ;
        RECT 299.250 383.250 300.750 384.150 ;
        RECT 301.950 382.950 304.050 385.050 ;
        RECT 295.950 380.850 297.750 381.750 ;
        RECT 298.950 379.950 301.050 382.050 ;
        RECT 302.250 380.850 303.750 381.750 ;
        RECT 304.950 379.950 307.050 382.050 ;
        RECT 299.400 379.050 300.450 379.950 ;
        RECT 298.950 376.950 301.050 379.050 ;
        RECT 304.950 377.850 307.050 378.750 ;
        RECT 295.950 355.950 298.050 358.050 ;
        RECT 296.400 346.050 297.450 355.950 ;
        RECT 308.400 349.050 309.450 385.950 ;
        RECT 301.950 347.250 304.050 348.150 ;
        RECT 307.950 346.950 310.050 349.050 ;
        RECT 295.950 343.950 298.050 346.050 ;
        RECT 299.250 344.250 300.750 345.150 ;
        RECT 301.950 343.950 304.050 346.050 ;
        RECT 305.250 344.250 307.050 345.150 ;
        RECT 295.950 341.850 297.750 342.750 ;
        RECT 298.950 340.950 301.050 343.050 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 299.400 331.050 300.450 340.950 ;
        RECT 305.400 340.050 306.450 340.950 ;
        RECT 304.950 337.950 307.050 340.050 ;
        RECT 298.950 328.950 301.050 331.050 ;
        RECT 295.950 316.950 298.050 319.050 ;
        RECT 296.400 292.050 297.450 316.950 ;
        RECT 299.400 313.050 300.450 328.950 ;
        RECT 308.400 315.450 309.450 346.950 ;
        RECT 311.400 345.450 312.450 409.950 ;
        RECT 314.400 400.050 315.450 412.950 ;
        RECT 313.950 397.950 316.050 400.050 ;
        RECT 317.400 382.050 318.450 421.950 ;
        RECT 320.400 385.050 321.450 433.950 ;
        RECT 323.400 412.050 324.450 448.950 ;
        RECT 326.400 424.050 327.450 466.950 ;
        RECT 329.400 445.050 330.450 481.950 ;
        RECT 332.400 481.050 333.450 520.950 ;
        RECT 340.950 514.950 343.050 517.050 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 334.950 487.950 337.050 490.050 ;
        RECT 335.400 484.050 336.450 487.950 ;
        RECT 334.950 481.950 337.050 484.050 ;
        RECT 331.950 478.950 334.050 481.050 ;
        RECT 335.400 459.450 336.450 481.950 ;
        RECT 338.400 469.050 339.450 490.950 ;
        RECT 341.400 480.450 342.450 514.950 ;
        RECT 346.950 493.950 349.050 496.050 ;
        RECT 347.400 490.050 348.450 493.950 ;
        RECT 346.950 487.950 349.050 490.050 ;
        RECT 343.950 485.250 346.050 486.150 ;
        RECT 346.950 485.850 349.050 486.750 ;
        RECT 343.950 481.950 346.050 484.050 ;
        RECT 341.400 479.400 345.450 480.450 ;
        RECT 337.950 466.950 340.050 469.050 ;
        RECT 332.400 458.400 336.450 459.450 ;
        RECT 332.400 454.050 333.450 458.400 ;
        RECT 334.950 454.950 337.050 457.050 ;
        RECT 338.250 455.250 339.750 456.150 ;
        RECT 340.950 454.950 343.050 457.050 ;
        RECT 331.950 451.950 334.050 454.050 ;
        RECT 335.250 452.850 336.750 453.750 ;
        RECT 337.950 451.950 340.050 454.050 ;
        RECT 341.250 452.850 343.050 453.750 ;
        RECT 331.950 449.850 334.050 450.750 ;
        RECT 328.950 442.950 331.050 445.050 ;
        RECT 338.400 441.450 339.450 451.950 ;
        RECT 338.400 440.400 342.450 441.450 ;
        RECT 334.950 436.950 337.050 439.050 ;
        RECT 328.950 433.950 331.050 436.050 ;
        RECT 325.950 421.950 328.050 424.050 ;
        RECT 325.950 418.950 328.050 421.050 ;
        RECT 322.950 409.950 325.050 412.050 ;
        RECT 319.950 382.950 322.050 385.050 ;
        RECT 313.950 379.950 316.050 382.050 ;
        RECT 316.950 379.950 319.050 382.050 ;
        RECT 319.950 380.250 321.750 381.150 ;
        RECT 322.950 379.950 325.050 382.050 ;
        RECT 314.400 364.050 315.450 379.950 ;
        RECT 326.400 379.050 327.450 418.950 ;
        RECT 329.400 418.050 330.450 433.950 ;
        RECT 328.950 415.950 331.050 418.050 ;
        RECT 331.950 415.950 334.050 418.050 ;
        RECT 328.950 413.250 331.050 414.150 ;
        RECT 331.950 413.850 334.050 414.750 ;
        RECT 328.950 409.950 331.050 412.050 ;
        RECT 331.950 409.950 334.050 412.050 ;
        RECT 328.950 388.950 331.050 391.050 ;
        RECT 329.400 382.050 330.450 388.950 ;
        RECT 328.950 379.950 331.050 382.050 ;
        RECT 316.950 376.950 319.050 379.050 ;
        RECT 319.950 376.950 322.050 379.050 ;
        RECT 323.250 377.850 324.750 378.750 ;
        RECT 325.950 376.950 328.050 379.050 ;
        RECT 329.250 377.850 331.050 378.750 ;
        RECT 313.950 361.950 316.050 364.050 ;
        RECT 317.400 352.050 318.450 376.950 ;
        RECT 320.400 355.050 321.450 376.950 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 325.950 374.850 328.050 375.750 ;
        RECT 319.950 352.950 322.050 355.050 ;
        RECT 316.950 349.950 319.050 352.050 ;
        RECT 320.400 348.450 321.450 352.950 ;
        RECT 323.400 349.050 324.450 373.950 ;
        RECT 332.400 370.050 333.450 409.950 ;
        RECT 335.400 390.450 336.450 436.950 ;
        RECT 337.950 413.250 340.050 414.150 ;
        RECT 337.950 409.950 340.050 412.050 ;
        RECT 338.400 406.050 339.450 409.950 ;
        RECT 337.950 403.950 340.050 406.050 ;
        RECT 335.400 389.400 339.450 390.450 ;
        RECT 334.950 382.950 337.050 385.050 ;
        RECT 335.400 370.050 336.450 382.950 ;
        RECT 338.400 373.050 339.450 389.400 ;
        RECT 341.400 388.050 342.450 440.400 ;
        RECT 344.400 409.050 345.450 479.400 ;
        RECT 346.950 472.950 349.050 475.050 ;
        RECT 347.400 421.050 348.450 472.950 ;
        RECT 350.400 472.050 351.450 521.400 ;
        RECT 353.400 520.050 354.450 526.950 ;
        RECT 356.400 526.050 357.450 571.950 ;
        RECT 358.950 568.950 361.050 571.050 ;
        RECT 359.400 538.050 360.450 568.950 ;
        RECT 361.950 560.250 364.050 561.150 ;
        RECT 368.400 559.050 369.450 580.950 ;
        RECT 371.400 571.050 372.450 580.950 ;
        RECT 370.950 568.950 373.050 571.050 ;
        RECT 361.950 556.950 364.050 559.050 ;
        RECT 365.250 557.250 366.750 558.150 ;
        RECT 367.950 556.950 370.050 559.050 ;
        RECT 371.250 557.250 373.050 558.150 ;
        RECT 364.950 553.950 367.050 556.050 ;
        RECT 368.250 554.850 369.750 555.750 ;
        RECT 370.950 553.950 373.050 556.050 ;
        RECT 365.400 547.050 366.450 553.950 ;
        RECT 364.950 544.950 367.050 547.050 ;
        RECT 358.950 535.950 361.050 538.050 ;
        RECT 364.950 535.950 367.050 538.050 ;
        RECT 365.400 532.050 366.450 535.950 ;
        RECT 358.950 529.950 361.050 532.050 ;
        RECT 364.950 529.950 367.050 532.050 ;
        RECT 359.400 529.050 360.450 529.950 ;
        RECT 358.950 526.950 361.050 529.050 ;
        RECT 362.250 527.250 364.050 528.150 ;
        RECT 364.950 527.850 367.050 528.750 ;
        RECT 367.950 527.250 370.050 528.150 ;
        RECT 355.950 523.950 358.050 526.050 ;
        RECT 358.950 524.850 360.750 525.750 ;
        RECT 361.950 523.950 364.050 526.050 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 352.950 517.950 355.050 520.050 ;
        RECT 352.950 485.250 355.050 486.150 ;
        RECT 352.950 483.450 355.050 484.050 ;
        RECT 356.400 483.450 357.450 523.950 ;
        RECT 362.400 507.450 363.450 523.950 ;
        RECT 359.400 506.400 363.450 507.450 ;
        RECT 359.400 484.050 360.450 506.400 ;
        RECT 361.950 493.950 364.050 496.050 ;
        RECT 362.400 490.050 363.450 493.950 ;
        RECT 368.400 490.050 369.450 523.950 ;
        RECT 361.950 487.950 364.050 490.050 ;
        RECT 365.250 488.250 366.750 489.150 ;
        RECT 367.950 487.950 370.050 490.050 ;
        RECT 370.950 487.950 373.050 490.050 ;
        RECT 361.950 485.850 363.750 486.750 ;
        RECT 364.950 484.950 367.050 487.050 ;
        RECT 368.250 485.850 370.050 486.750 ;
        RECT 352.950 482.400 357.450 483.450 ;
        RECT 352.950 481.950 355.050 482.400 ;
        RECT 358.950 481.950 361.050 484.050 ;
        RECT 355.950 478.950 358.050 481.050 ;
        RECT 349.950 469.950 352.050 472.050 ;
        RECT 352.950 466.950 355.050 469.050 ;
        RECT 353.400 460.050 354.450 466.950 ;
        RECT 352.950 457.950 355.050 460.050 ;
        RECT 353.400 454.050 354.450 457.950 ;
        RECT 356.400 457.050 357.450 478.950 ;
        RECT 365.400 469.050 366.450 484.950 ;
        RECT 371.400 483.450 372.450 487.950 ;
        RECT 368.400 482.400 372.450 483.450 ;
        RECT 364.950 466.950 367.050 469.050 ;
        RECT 361.950 457.950 364.050 460.050 ;
        RECT 355.950 454.950 358.050 457.050 ;
        RECT 359.250 455.250 361.050 456.150 ;
        RECT 361.950 455.850 364.050 456.750 ;
        RECT 364.950 455.250 367.050 456.150 ;
        RECT 352.950 451.950 355.050 454.050 ;
        RECT 355.950 452.850 357.750 453.750 ;
        RECT 358.950 451.950 361.050 454.050 ;
        RECT 361.950 451.950 364.050 454.050 ;
        RECT 364.950 451.950 367.050 454.050 ;
        RECT 346.950 418.950 349.050 421.050 ;
        RECT 349.950 417.450 352.050 418.050 ;
        RECT 347.400 416.400 352.050 417.450 ;
        RECT 355.950 417.450 358.050 418.050 ;
        RECT 343.950 406.950 346.050 409.050 ;
        RECT 347.400 406.050 348.450 416.400 ;
        RECT 349.950 415.950 352.050 416.400 ;
        RECT 353.250 416.250 354.750 417.150 ;
        RECT 355.950 416.400 360.450 417.450 ;
        RECT 355.950 415.950 358.050 416.400 ;
        RECT 349.950 413.850 351.750 414.750 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 356.250 413.850 358.050 414.750 ;
        RECT 359.400 409.050 360.450 416.400 ;
        RECT 362.400 415.050 363.450 451.950 ;
        RECT 365.400 439.050 366.450 451.950 ;
        RECT 364.950 436.950 367.050 439.050 ;
        RECT 364.950 418.950 367.050 421.050 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 358.950 406.950 361.050 409.050 ;
        RECT 346.950 403.950 349.050 406.050 ;
        RECT 346.950 388.950 349.050 391.050 ;
        RECT 361.950 388.950 364.050 391.050 ;
        RECT 347.400 388.050 348.450 388.950 ;
        RECT 340.950 385.950 343.050 388.050 ;
        RECT 346.950 385.950 349.050 388.050 ;
        RECT 352.950 385.950 355.050 388.050 ;
        RECT 341.400 385.050 342.450 385.950 ;
        RECT 340.950 382.950 343.050 385.050 ;
        RECT 344.250 383.250 346.050 384.150 ;
        RECT 346.950 383.850 349.050 384.750 ;
        RECT 349.950 383.250 352.050 384.150 ;
        RECT 340.950 380.850 342.750 381.750 ;
        RECT 343.950 379.950 346.050 382.050 ;
        RECT 349.950 379.950 352.050 382.050 ;
        RECT 344.400 379.050 345.450 379.950 ;
        RECT 343.950 376.950 346.050 379.050 ;
        RECT 350.400 373.050 351.450 379.950 ;
        RECT 353.400 379.050 354.450 385.950 ;
        RECT 355.950 382.950 358.050 385.050 ;
        RECT 352.950 376.950 355.050 379.050 ;
        RECT 337.950 370.950 340.050 373.050 ;
        RECT 349.950 370.950 352.050 373.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 325.950 355.950 328.050 358.050 ;
        RECT 317.400 347.400 321.450 348.450 ;
        RECT 311.400 344.400 315.450 345.450 ;
        RECT 310.950 340.950 313.050 343.050 ;
        RECT 310.950 338.850 313.050 339.750 ;
        RECT 314.400 334.050 315.450 344.400 ;
        RECT 317.400 340.050 318.450 347.400 ;
        RECT 322.950 346.950 325.050 349.050 ;
        RECT 319.950 343.950 322.050 346.050 ;
        RECT 322.950 344.250 325.050 345.150 ;
        RECT 316.950 337.950 319.050 340.050 ;
        RECT 313.950 331.950 316.050 334.050 ;
        RECT 308.400 314.400 312.450 315.450 ;
        RECT 298.950 310.950 301.050 313.050 ;
        RECT 307.950 311.250 310.050 312.150 ;
        RECT 311.400 310.050 312.450 314.400 ;
        RECT 313.950 310.950 316.050 313.050 ;
        RECT 317.250 311.250 319.050 312.150 ;
        RECT 307.950 307.950 310.050 310.050 ;
        RECT 310.950 307.950 313.050 310.050 ;
        RECT 313.950 308.850 315.750 309.750 ;
        RECT 316.950 307.950 319.050 310.050 ;
        RECT 311.400 307.050 312.450 307.950 ;
        RECT 310.950 304.950 313.050 307.050 ;
        RECT 301.950 295.950 304.050 298.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 295.950 280.950 298.050 283.050 ;
        RECT 296.400 274.050 297.450 280.950 ;
        RECT 302.400 274.050 303.450 295.950 ;
        RECT 307.950 289.950 310.050 292.050 ;
        RECT 292.950 271.950 295.050 274.050 ;
        RECT 295.950 271.950 298.050 274.050 ;
        RECT 299.250 272.250 300.750 273.150 ;
        RECT 301.950 271.950 304.050 274.050 ;
        RECT 295.950 269.850 297.750 270.750 ;
        RECT 298.950 268.950 301.050 271.050 ;
        RECT 302.250 269.850 304.050 270.750 ;
        RECT 289.950 259.950 292.050 262.050 ;
        RECT 299.400 253.050 300.450 268.950 ;
        RECT 286.950 250.950 289.050 253.050 ;
        RECT 298.950 250.950 301.050 253.050 ;
        RECT 286.950 245.400 289.050 247.500 ;
        RECT 289.950 245.400 292.050 247.500 ;
        RECT 292.950 245.400 295.050 247.500 ;
        RECT 297.750 245.400 299.850 247.500 ;
        RECT 301.950 245.400 304.050 247.500 ;
        RECT 277.950 235.950 280.050 238.050 ;
        RECT 277.950 233.850 280.050 234.750 ;
        RECT 287.550 231.750 288.750 245.400 ;
        RECT 286.950 229.650 289.050 231.750 ;
        RECT 287.550 225.900 288.750 229.650 ;
        RECT 290.250 228.150 291.450 245.400 ;
        RECT 293.400 231.750 294.600 245.400 ;
        RECT 298.350 239.550 299.550 245.400 ;
        RECT 297.750 237.450 299.850 239.550 ;
        RECT 292.950 229.650 295.050 231.750 ;
        RECT 298.350 228.600 299.550 237.450 ;
        RECT 302.550 236.850 303.750 245.400 ;
        RECT 304.950 241.950 307.050 244.050 ;
        RECT 304.950 239.850 307.050 240.750 ;
        RECT 301.950 234.750 304.050 236.850 ;
        RECT 304.950 235.950 307.050 238.050 ;
        RECT 302.550 228.600 303.750 234.750 ;
        RECT 289.950 226.050 292.050 228.150 ;
        RECT 297.900 226.500 300.000 228.600 ;
        RECT 301.950 226.500 304.050 228.600 ;
        RECT 286.800 223.800 288.900 225.900 ;
        RECT 305.400 223.050 306.450 235.950 ;
        RECT 304.950 220.950 307.050 223.050 ;
        RECT 295.950 203.250 298.050 204.150 ;
        RECT 268.950 199.950 271.050 202.050 ;
        RECT 272.250 200.250 273.750 201.150 ;
        RECT 274.950 199.950 277.050 202.050 ;
        RECT 280.950 199.950 283.050 202.050 ;
        RECT 289.950 199.950 292.050 202.050 ;
        RECT 293.250 200.250 294.750 201.150 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 299.250 200.250 301.050 201.150 ;
        RECT 301.950 199.950 304.050 202.050 ;
        RECT 268.950 197.850 270.750 198.750 ;
        RECT 271.950 196.950 274.050 199.050 ;
        RECT 275.250 197.850 277.050 198.750 ;
        RECT 268.950 184.950 271.050 187.050 ;
        RECT 247.950 163.950 250.050 166.050 ;
        RECT 262.950 164.250 264.750 165.150 ;
        RECT 265.950 163.950 268.050 166.050 ;
        RECT 248.400 133.050 249.450 163.950 ;
        RECT 269.400 163.050 270.450 184.950 ;
        RECT 272.400 169.050 273.450 196.950 ;
        RECT 274.950 169.950 277.050 172.050 ;
        RECT 271.950 166.950 274.050 169.050 ;
        RECT 271.950 165.450 274.050 166.050 ;
        RECT 275.400 165.450 276.450 169.950 ;
        RECT 277.950 166.950 280.050 169.050 ;
        RECT 271.950 164.400 276.450 165.450 ;
        RECT 271.950 163.950 274.050 164.400 ;
        RECT 262.950 160.950 265.050 163.050 ;
        RECT 266.250 161.850 267.750 162.750 ;
        RECT 268.950 160.950 271.050 163.050 ;
        RECT 272.250 161.850 274.050 162.750 ;
        RECT 268.950 158.850 271.050 159.750 ;
        RECT 271.950 148.950 274.050 151.050 ;
        RECT 247.950 130.950 250.050 133.050 ;
        RECT 262.950 131.250 265.050 132.150 ;
        RECT 244.950 127.950 247.050 130.050 ;
        RECT 256.950 127.950 259.050 130.050 ;
        RECT 260.250 128.250 261.750 129.150 ;
        RECT 262.950 127.950 265.050 130.050 ;
        RECT 266.250 128.250 268.050 129.150 ;
        RECT 241.950 118.950 244.050 121.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 226.950 97.950 229.050 100.050 ;
        RECT 227.400 97.050 228.450 97.950 ;
        RECT 226.950 94.950 229.050 97.050 ;
        RECT 223.950 93.450 226.050 94.050 ;
        RECT 221.400 92.400 226.050 93.450 ;
        RECT 221.400 85.050 222.450 92.400 ;
        RECT 223.950 91.950 226.050 92.400 ;
        RECT 227.400 91.050 228.450 94.950 ;
        RECT 229.950 91.950 232.050 94.050 ;
        RECT 233.250 92.250 235.050 93.150 ;
        RECT 238.950 91.950 241.050 94.050 ;
        RECT 223.950 89.850 225.750 90.750 ;
        RECT 226.950 88.950 229.050 91.050 ;
        RECT 230.250 89.850 231.750 90.750 ;
        RECT 232.950 88.950 235.050 91.050 ;
        RECT 226.950 86.850 229.050 87.750 ;
        RECT 220.950 82.950 223.050 85.050 ;
        RECT 220.950 58.950 223.050 61.050 ;
        RECT 217.950 52.950 220.050 55.050 ;
        RECT 221.400 52.050 222.450 58.950 ;
        RECT 239.400 58.050 240.450 91.950 ;
        RECT 245.400 64.050 246.450 127.950 ;
        RECT 256.950 125.850 258.750 126.750 ;
        RECT 259.950 124.950 262.050 127.050 ;
        RECT 260.400 124.050 261.450 124.950 ;
        RECT 259.950 121.950 262.050 124.050 ;
        RECT 263.400 118.050 264.450 127.950 ;
        RECT 265.950 124.950 268.050 127.050 ;
        RECT 272.400 124.050 273.450 148.950 ;
        RECT 275.400 127.050 276.450 164.400 ;
        RECT 278.400 160.050 279.450 166.950 ;
        RECT 281.400 163.050 282.450 199.950 ;
        RECT 289.950 197.850 291.750 198.750 ;
        RECT 292.950 196.950 295.050 199.050 ;
        RECT 298.950 196.950 301.050 199.050 ;
        RECT 299.400 193.050 300.450 196.950 ;
        RECT 298.950 190.950 301.050 193.050 ;
        RECT 302.400 178.050 303.450 199.950 ;
        RECT 308.400 199.050 309.450 289.950 ;
        RECT 316.950 274.950 319.050 277.050 ;
        RECT 317.400 271.050 318.450 274.950 ;
        RECT 316.950 268.950 319.050 271.050 ;
        RECT 316.950 266.850 319.050 267.750 ;
        RECT 310.950 244.950 313.050 247.050 ;
        RECT 313.950 244.950 316.050 247.050 ;
        RECT 316.950 244.950 319.050 247.050 ;
        RECT 311.250 226.050 312.450 244.950 ;
        RECT 314.250 232.350 315.450 244.950 ;
        RECT 313.950 230.250 316.050 232.350 ;
        RECT 314.250 226.050 315.450 230.250 ;
        RECT 317.250 226.050 318.450 244.950 ;
        RECT 320.400 241.050 321.450 343.950 ;
        RECT 322.950 340.950 325.050 343.050 ;
        RECT 323.400 325.050 324.450 340.950 ;
        RECT 326.400 337.050 327.450 355.950 ;
        RECT 331.800 353.100 333.900 355.200 ;
        RECT 332.550 349.350 333.750 353.100 ;
        RECT 334.950 350.850 337.050 352.950 ;
        RECT 328.950 346.950 331.050 349.050 ;
        RECT 331.950 347.250 334.050 349.350 ;
        RECT 325.950 334.950 328.050 337.050 ;
        RECT 322.950 322.950 325.050 325.050 ;
        RECT 322.950 312.450 325.050 313.050 ;
        RECT 326.400 312.450 327.450 334.950 ;
        RECT 329.400 313.050 330.450 346.950 ;
        RECT 332.550 333.600 333.750 347.250 ;
        RECT 335.250 333.600 336.450 350.850 ;
        RECT 342.900 350.400 345.000 352.500 ;
        RECT 346.950 350.400 349.050 352.500 ;
        RECT 337.950 347.250 340.050 349.350 ;
        RECT 338.400 333.600 339.600 347.250 ;
        RECT 343.350 341.550 344.550 350.400 ;
        RECT 347.550 344.250 348.750 350.400 ;
        RECT 346.950 342.150 349.050 344.250 ;
        RECT 342.750 339.450 344.850 341.550 ;
        RECT 343.350 333.600 344.550 339.450 ;
        RECT 347.550 333.600 348.750 342.150 ;
        RECT 349.950 338.250 352.050 339.150 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 331.950 331.500 334.050 333.600 ;
        RECT 334.950 331.500 337.050 333.600 ;
        RECT 337.950 331.500 340.050 333.600 ;
        RECT 342.750 331.500 344.850 333.600 ;
        RECT 346.950 331.500 349.050 333.600 ;
        RECT 349.950 331.950 352.050 334.050 ;
        RECT 340.950 325.950 343.050 328.050 ;
        RECT 334.950 322.950 337.050 325.050 ;
        RECT 322.950 311.400 327.450 312.450 ;
        RECT 322.950 310.950 325.050 311.400 ;
        RECT 328.950 310.950 331.050 313.050 ;
        RECT 322.950 308.850 325.050 309.750 ;
        RECT 331.950 274.950 334.050 277.050 ;
        RECT 322.950 271.950 325.050 274.050 ;
        RECT 328.950 271.950 331.050 274.050 ;
        RECT 323.400 271.050 324.450 271.950 ;
        RECT 329.400 271.050 330.450 271.950 ;
        RECT 322.950 268.950 325.050 271.050 ;
        RECT 328.950 268.950 331.050 271.050 ;
        RECT 322.950 266.850 325.050 267.750 ;
        RECT 325.950 265.950 328.050 268.050 ;
        RECT 328.950 266.850 331.050 267.750 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 322.950 233.850 325.050 234.750 ;
        RECT 310.950 223.950 313.050 226.050 ;
        RECT 313.950 223.950 316.050 226.050 ;
        RECT 316.950 223.950 319.050 226.050 ;
        RECT 316.950 220.950 319.050 223.050 ;
        RECT 310.950 205.950 313.050 208.050 ;
        RECT 311.400 199.050 312.450 205.950 ;
        RECT 307.950 196.950 310.050 199.050 ;
        RECT 310.950 196.950 313.050 199.050 ;
        RECT 310.950 194.850 313.050 195.750 ;
        RECT 313.950 194.250 316.050 195.150 ;
        RECT 313.950 190.950 316.050 193.050 ;
        RECT 313.950 187.950 316.050 190.050 ;
        RECT 301.950 175.950 304.050 178.050 ;
        RECT 310.950 175.950 313.050 178.050 ;
        RECT 311.400 169.050 312.450 175.950 ;
        RECT 304.950 166.950 307.050 169.050 ;
        RECT 308.250 167.250 309.750 168.150 ;
        RECT 310.950 166.950 313.050 169.050 ;
        RECT 283.950 164.250 285.750 165.150 ;
        RECT 286.950 163.950 289.050 166.050 ;
        RECT 290.250 164.250 292.050 165.150 ;
        RECT 301.950 163.950 304.050 166.050 ;
        RECT 305.250 164.850 306.750 165.750 ;
        RECT 307.950 163.950 310.050 166.050 ;
        RECT 311.250 164.850 313.050 165.750 ;
        RECT 280.950 160.950 283.050 163.050 ;
        RECT 283.950 160.950 286.050 163.050 ;
        RECT 287.250 161.850 288.750 162.750 ;
        RECT 289.950 160.950 292.050 163.050 ;
        RECT 292.950 160.950 295.050 163.050 ;
        RECT 301.950 161.850 304.050 162.750 ;
        RECT 284.400 160.050 285.450 160.950 ;
        RECT 277.950 157.950 280.050 160.050 ;
        RECT 283.950 157.950 286.050 160.050 ;
        RECT 277.950 130.950 280.050 133.050 ;
        RECT 283.950 131.250 286.050 132.150 ;
        RECT 278.400 130.050 279.450 130.950 ;
        RECT 277.950 127.950 280.050 130.050 ;
        RECT 281.250 128.250 282.750 129.150 ;
        RECT 283.950 127.950 286.050 130.050 ;
        RECT 287.250 128.250 289.050 129.150 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 277.950 125.850 279.750 126.750 ;
        RECT 280.950 124.950 283.050 127.050 ;
        RECT 286.950 124.950 289.050 127.050 ;
        RECT 281.400 124.050 282.450 124.950 ;
        RECT 271.950 121.950 274.050 124.050 ;
        RECT 280.950 121.950 283.050 124.050 ;
        RECT 265.950 118.950 268.050 121.050 ;
        RECT 262.950 115.950 265.050 118.050 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 248.400 94.050 249.450 97.950 ;
        RECT 250.950 94.950 253.050 97.050 ;
        RECT 254.250 95.250 255.750 96.150 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 259.950 94.950 262.050 97.050 ;
        RECT 247.950 91.950 250.050 94.050 ;
        RECT 251.250 92.850 252.750 93.750 ;
        RECT 253.950 91.950 256.050 94.050 ;
        RECT 257.250 92.850 259.050 93.750 ;
        RECT 247.950 89.850 250.050 90.750 ;
        RECT 244.950 61.950 247.050 64.050 ;
        RECT 254.400 58.050 255.450 91.950 ;
        RECT 256.950 88.950 259.050 91.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 241.950 56.250 244.050 57.150 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 227.400 55.050 228.450 55.950 ;
        RECT 248.400 55.050 249.450 55.950 ;
        RECT 257.400 55.050 258.450 88.950 ;
        RECT 226.950 52.950 229.050 55.050 ;
        RECT 241.950 52.950 244.050 55.050 ;
        RECT 245.250 53.250 246.750 54.150 ;
        RECT 247.950 52.950 250.050 55.050 ;
        RECT 251.250 53.250 253.050 54.150 ;
        RECT 256.950 52.950 259.050 55.050 ;
        RECT 220.950 49.950 223.050 52.050 ;
        RECT 226.950 50.850 229.050 51.750 ;
        RECT 229.950 50.250 232.050 51.150 ;
        RECT 242.400 49.050 243.450 52.950 ;
        RECT 260.400 52.050 261.450 94.950 ;
        RECT 266.400 94.050 267.450 118.950 ;
        RECT 293.400 112.050 294.450 160.950 ;
        RECT 310.950 157.950 313.050 160.050 ;
        RECT 298.950 131.250 301.050 132.150 ;
        RECT 295.950 128.250 297.750 129.150 ;
        RECT 298.950 127.950 301.050 130.050 ;
        RECT 302.250 128.250 303.750 129.150 ;
        RECT 304.950 127.950 307.050 130.050 ;
        RECT 307.950 127.950 310.050 130.050 ;
        RECT 295.950 124.950 298.050 127.050 ;
        RECT 299.400 118.050 300.450 127.950 ;
        RECT 301.950 124.950 304.050 127.050 ;
        RECT 305.250 125.850 307.050 126.750 ;
        RECT 302.400 124.050 303.450 124.950 ;
        RECT 301.950 121.950 304.050 124.050 ;
        RECT 298.950 115.950 301.050 118.050 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 292.950 109.950 295.050 112.050 ;
        RECT 271.950 103.950 274.050 106.050 ;
        RECT 277.950 103.950 280.050 106.050 ;
        RECT 272.400 103.050 273.450 103.950 ;
        RECT 271.950 100.950 274.050 103.050 ;
        RECT 272.400 94.050 273.450 100.950 ;
        RECT 278.400 94.050 279.450 103.950 ;
        RECT 289.950 97.950 292.050 100.050 ;
        RECT 296.400 97.050 297.450 112.950 ;
        RECT 299.400 112.050 300.450 115.950 ;
        RECT 298.950 109.950 301.050 112.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 299.400 97.050 300.450 97.950 ;
        RECT 286.950 95.250 289.050 96.150 ;
        RECT 289.950 95.850 292.050 96.750 ;
        RECT 292.950 95.250 294.750 96.150 ;
        RECT 295.950 94.950 298.050 97.050 ;
        RECT 298.950 94.950 301.050 97.050 ;
        RECT 299.400 94.050 300.450 94.950 ;
        RECT 265.950 91.950 268.050 94.050 ;
        RECT 268.950 92.250 270.750 93.150 ;
        RECT 271.950 91.950 274.050 94.050 ;
        RECT 277.950 91.950 280.050 94.050 ;
        RECT 286.950 91.950 289.050 94.050 ;
        RECT 292.950 91.950 295.050 94.050 ;
        RECT 296.250 92.850 298.050 93.750 ;
        RECT 298.950 91.950 301.050 94.050 ;
        RECT 268.950 88.950 271.050 91.050 ;
        RECT 272.250 89.850 273.750 90.750 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 278.250 89.850 280.050 90.750 ;
        RECT 269.400 88.050 270.450 88.950 ;
        RECT 268.950 85.950 271.050 88.050 ;
        RECT 274.950 86.850 277.050 87.750 ;
        RECT 274.950 82.950 277.050 85.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 262.950 53.250 265.050 54.150 ;
        RECT 265.950 53.850 268.050 54.750 ;
        RECT 271.950 53.250 274.050 54.150 ;
        RECT 244.950 49.950 247.050 52.050 ;
        RECT 248.250 50.850 249.750 51.750 ;
        RECT 250.950 49.950 253.050 52.050 ;
        RECT 259.950 49.950 262.050 52.050 ;
        RECT 262.950 49.950 265.050 52.050 ;
        RECT 271.950 49.950 274.050 52.050 ;
        RECT 229.950 46.950 232.050 49.050 ;
        RECT 241.950 46.950 244.050 49.050 ;
        RECT 245.400 46.050 246.450 49.950 ;
        RECT 244.950 43.950 247.050 46.050 ;
        RECT 212.400 29.400 216.450 30.450 ;
        RECT 196.950 25.950 199.050 28.050 ;
        RECT 199.950 25.950 202.050 28.050 ;
        RECT 200.400 25.050 201.450 25.950 ;
        RECT 212.400 25.050 213.450 29.400 ;
        RECT 238.950 28.950 241.050 31.050 ;
        RECT 239.400 28.050 240.450 28.950 ;
        RECT 214.950 25.950 217.050 28.050 ;
        RECT 238.950 25.950 241.050 28.050 ;
        RECT 259.950 25.950 262.050 28.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 197.250 23.850 198.750 24.750 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 172.950 21.450 175.050 22.050 ;
        RECT 170.400 20.400 175.050 21.450 ;
        RECT 172.950 19.950 175.050 20.400 ;
        RECT 178.950 19.950 181.050 22.050 ;
        RECT 182.250 20.850 184.050 21.750 ;
        RECT 184.950 19.950 187.050 22.050 ;
        RECT 193.950 20.850 196.050 21.750 ;
        RECT 199.950 20.850 202.050 21.750 ;
        RECT 211.950 20.850 214.050 21.750 ;
        RECT 155.400 19.050 156.450 19.950 ;
        RECT 34.950 16.950 37.050 19.050 ;
        RECT 76.950 17.850 79.050 18.750 ;
        RECT 103.950 17.850 106.050 18.750 ;
        RECT 118.950 16.950 121.050 19.050 ;
        RECT 122.250 17.850 123.750 18.750 ;
        RECT 124.950 16.950 127.050 19.050 ;
        RECT 128.250 17.850 130.050 18.750 ;
        RECT 133.950 16.950 136.050 19.050 ;
        RECT 139.950 16.950 142.050 19.050 ;
        RECT 142.950 16.950 145.050 19.050 ;
        RECT 154.950 16.950 157.050 19.050 ;
        RECT 160.950 17.850 163.050 18.750 ;
        RECT 215.400 18.450 216.450 25.950 ;
        RECT 260.400 25.050 261.450 25.950 ;
        RECT 220.950 24.450 223.050 25.050 ;
        RECT 220.950 23.400 225.450 24.450 ;
        RECT 220.950 22.950 223.050 23.400 ;
        RECT 217.950 20.250 220.050 21.150 ;
        RECT 220.950 20.850 223.050 21.750 ;
        RECT 224.400 19.050 225.450 23.400 ;
        RECT 235.950 23.250 238.050 24.150 ;
        RECT 238.950 23.850 241.050 24.750 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 257.250 23.250 258.750 24.150 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 263.400 22.050 264.450 49.950 ;
        RECT 268.950 22.950 271.050 25.050 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 250.950 19.950 253.050 22.050 ;
        RECT 254.250 20.850 255.750 21.750 ;
        RECT 256.950 19.950 259.050 22.050 ;
        RECT 260.250 20.850 262.050 21.750 ;
        RECT 262.950 19.950 265.050 22.050 ;
        RECT 217.950 18.450 220.050 19.050 ;
        RECT 215.400 17.400 220.050 18.450 ;
        RECT 217.950 16.950 220.050 17.400 ;
        RECT 223.950 16.950 226.050 19.050 ;
        RECT 250.950 17.850 253.050 18.750 ;
        RECT 269.400 18.450 270.450 22.950 ;
        RECT 275.400 22.050 276.450 82.950 ;
        RECT 287.400 61.050 288.450 91.950 ;
        RECT 308.400 91.050 309.450 127.950 ;
        RECT 311.400 124.050 312.450 157.950 ;
        RECT 310.950 121.950 313.050 124.050 ;
        RECT 314.400 115.050 315.450 187.950 ;
        RECT 317.400 166.050 318.450 220.950 ;
        RECT 319.950 205.950 322.050 208.050 ;
        RECT 316.950 163.950 319.050 166.050 ;
        RECT 320.400 136.050 321.450 205.950 ;
        RECT 326.400 195.450 327.450 265.950 ;
        RECT 328.950 236.250 331.050 237.150 ;
        RECT 328.950 234.450 331.050 235.050 ;
        RECT 332.400 234.450 333.450 274.950 ;
        RECT 335.400 271.050 336.450 322.950 ;
        RECT 341.400 310.050 342.450 325.950 ;
        RECT 337.950 308.250 339.750 309.150 ;
        RECT 340.950 307.950 343.050 310.050 ;
        RECT 346.950 309.450 349.050 310.050 ;
        RECT 350.400 309.450 351.450 331.950 ;
        RECT 353.400 330.450 354.450 376.950 ;
        RECT 356.400 358.050 357.450 382.950 ;
        RECT 362.400 382.050 363.450 388.950 ;
        RECT 365.400 385.050 366.450 418.950 ;
        RECT 368.400 418.050 369.450 482.400 ;
        RECT 370.950 457.950 373.050 460.050 ;
        RECT 371.400 451.050 372.450 457.950 ;
        RECT 370.950 448.950 373.050 451.050 ;
        RECT 374.400 450.450 375.450 592.950 ;
        RECT 377.400 583.050 378.450 592.950 ;
        RECT 380.400 583.050 381.450 668.400 ;
        RECT 385.950 667.950 388.050 670.050 ;
        RECT 391.950 667.950 394.050 670.050 ;
        RECT 395.250 668.250 397.050 669.150 ;
        RECT 385.950 665.850 387.750 666.750 ;
        RECT 388.950 664.950 391.050 667.050 ;
        RECT 392.250 665.850 393.750 666.750 ;
        RECT 394.950 664.950 397.050 667.050 ;
        RECT 388.950 662.850 391.050 663.750 ;
        RECT 395.400 658.050 396.450 664.950 ;
        RECT 398.400 661.050 399.450 709.950 ;
        RECT 412.950 707.250 415.050 708.150 ;
        RECT 403.950 703.950 406.050 706.050 ;
        RECT 409.950 704.250 411.750 705.150 ;
        RECT 412.950 703.950 415.050 706.050 ;
        RECT 416.250 704.250 417.750 705.150 ;
        RECT 418.950 703.950 421.050 706.050 ;
        RECT 400.950 701.250 403.050 702.150 ;
        RECT 400.950 697.950 403.050 700.050 ;
        RECT 401.400 694.050 402.450 697.950 ;
        RECT 400.950 691.950 403.050 694.050 ;
        RECT 401.400 691.050 402.450 691.950 ;
        RECT 400.950 688.950 403.050 691.050 ;
        RECT 400.950 685.950 403.050 688.050 ;
        RECT 397.950 658.950 400.050 661.050 ;
        RECT 394.950 655.950 397.050 658.050 ;
        RECT 391.950 635.250 394.050 636.150 ;
        RECT 385.950 633.450 388.050 634.050 ;
        RECT 383.400 632.400 388.050 633.450 ;
        RECT 383.400 622.050 384.450 632.400 ;
        RECT 385.950 631.950 388.050 632.400 ;
        RECT 389.250 632.250 390.750 633.150 ;
        RECT 391.950 631.950 394.050 634.050 ;
        RECT 395.250 632.250 397.050 633.150 ;
        RECT 385.950 629.850 387.750 630.750 ;
        RECT 388.950 628.950 391.050 631.050 ;
        RECT 389.400 628.050 390.450 628.950 ;
        RECT 388.950 625.950 391.050 628.050 ;
        RECT 382.950 619.950 385.050 622.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 389.400 600.450 390.450 601.950 ;
        RECT 386.400 599.400 390.450 600.450 ;
        RECT 386.400 598.050 387.450 599.400 ;
        RECT 392.400 598.050 393.450 631.950 ;
        RECT 394.950 628.950 397.050 631.050 ;
        RECT 401.400 622.050 402.450 685.950 ;
        RECT 404.400 646.050 405.450 703.950 ;
        RECT 422.400 703.050 423.450 775.950 ;
        RECT 427.950 772.950 430.050 775.050 ;
        RECT 431.250 773.250 432.750 774.150 ;
        RECT 433.950 772.950 436.050 775.050 ;
        RECT 437.250 773.250 439.050 774.150 ;
        RECT 448.950 773.250 451.050 774.150 ;
        RECT 451.950 773.850 454.050 774.750 ;
        RECT 424.950 754.950 427.050 757.050 ;
        RECT 425.400 736.050 426.450 754.950 ;
        RECT 428.400 748.050 429.450 772.950 ;
        RECT 455.400 772.050 456.450 776.400 ;
        RECT 457.950 773.250 460.050 774.150 ;
        RECT 466.950 773.250 469.050 774.150 ;
        RECT 472.950 773.250 475.050 774.150 ;
        RECT 430.950 769.950 433.050 772.050 ;
        RECT 434.250 770.850 435.750 771.750 ;
        RECT 436.950 769.950 439.050 772.050 ;
        RECT 448.950 769.950 451.050 772.050 ;
        RECT 454.950 769.950 457.050 772.050 ;
        RECT 457.950 769.950 460.050 772.050 ;
        RECT 466.950 769.950 469.050 772.050 ;
        RECT 470.250 770.250 471.750 771.150 ;
        RECT 472.950 769.950 475.050 772.050 ;
        RECT 437.400 769.050 438.450 769.950 ;
        RECT 436.950 766.950 439.050 769.050 ;
        RECT 454.950 763.950 457.050 766.050 ;
        RECT 448.950 751.950 451.050 754.050 ;
        RECT 427.950 745.950 430.050 748.050 ;
        RECT 427.950 743.850 430.050 744.750 ;
        RECT 430.950 743.250 433.050 744.150 ;
        RECT 445.950 742.950 448.050 745.050 ;
        RECT 430.950 739.950 433.050 742.050 ;
        RECT 442.950 739.950 445.050 742.050 ;
        RECT 446.400 739.050 447.450 742.950 ;
        RECT 449.400 742.050 450.450 751.950 ;
        RECT 448.950 739.950 451.050 742.050 ;
        RECT 452.250 740.250 454.050 741.150 ;
        RECT 430.950 736.950 433.050 739.050 ;
        RECT 442.950 737.850 444.750 738.750 ;
        RECT 445.950 736.950 448.050 739.050 ;
        RECT 449.250 737.850 450.750 738.750 ;
        RECT 451.950 738.450 454.050 739.050 ;
        RECT 455.400 738.450 456.450 763.950 ;
        RECT 458.400 751.050 459.450 769.950 ;
        RECT 469.950 766.950 472.050 769.050 ;
        RECT 473.400 751.050 474.450 769.950 ;
        RECT 457.950 748.950 460.050 751.050 ;
        RECT 466.950 748.950 469.050 751.050 ;
        RECT 472.950 748.950 475.050 751.050 ;
        RECT 467.400 742.050 468.450 748.950 ;
        RECT 476.400 748.050 477.450 811.950 ;
        RECT 491.400 811.050 492.450 814.950 ;
        RECT 493.950 811.950 496.050 814.050 ;
        RECT 497.250 812.250 499.050 813.150 ;
        RECT 499.950 811.950 502.050 814.050 ;
        RECT 487.950 809.850 489.750 810.750 ;
        RECT 490.950 808.950 493.050 811.050 ;
        RECT 494.250 809.850 495.750 810.750 ;
        RECT 496.950 808.950 499.050 811.050 ;
        RECT 490.950 806.850 493.050 807.750 ;
        RECT 490.950 774.450 493.050 775.050 ;
        RECT 488.400 773.400 493.050 774.450 ;
        RECT 475.950 745.950 478.050 748.050 ;
        RECT 484.950 745.950 487.050 748.050 ;
        RECT 469.950 742.950 472.050 745.050 ;
        RECT 475.950 744.450 478.050 745.050 ;
        RECT 473.250 743.250 474.750 744.150 ;
        RECT 475.950 743.400 480.450 744.450 ;
        RECT 475.950 742.950 478.050 743.400 ;
        RECT 466.950 739.950 469.050 742.050 ;
        RECT 470.250 740.850 471.750 741.750 ;
        RECT 472.950 739.950 475.050 742.050 ;
        RECT 476.250 740.850 478.050 741.750 ;
        RECT 451.950 737.400 456.450 738.450 ;
        RECT 466.950 737.850 469.050 738.750 ;
        RECT 473.400 738.450 474.450 739.950 ;
        RECT 470.400 737.400 474.450 738.450 ;
        RECT 451.950 736.950 454.050 737.400 ;
        RECT 424.950 733.950 427.050 736.050 ;
        RECT 409.950 700.950 412.050 703.050 ;
        RECT 415.950 700.950 418.050 703.050 ;
        RECT 419.250 701.850 421.050 702.750 ;
        RECT 421.950 700.950 424.050 703.050 ;
        RECT 410.400 700.050 411.450 700.950 ;
        RECT 416.400 700.050 417.450 700.950 ;
        RECT 409.950 697.950 412.050 700.050 ;
        RECT 415.950 697.950 418.050 700.050 ;
        RECT 416.400 697.050 417.450 697.950 ;
        RECT 415.950 694.950 418.050 697.050 ;
        RECT 412.950 682.950 415.050 685.050 ;
        RECT 424.950 682.950 427.050 685.050 ;
        RECT 413.400 676.050 414.450 682.950 ;
        RECT 406.950 673.950 409.050 676.050 ;
        RECT 412.950 673.950 415.050 676.050 ;
        RECT 407.400 667.050 408.450 673.950 ;
        RECT 425.400 673.050 426.450 682.950 ;
        RECT 431.400 679.050 432.450 736.950 ;
        RECT 445.950 734.850 448.050 735.750 ;
        RECT 470.400 727.050 471.450 737.400 ;
        RECT 475.950 736.950 478.050 739.050 ;
        RECT 476.400 735.450 477.450 736.950 ;
        RECT 473.400 734.400 477.450 735.450 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 469.950 706.950 472.050 709.050 ;
        RECT 442.950 703.950 445.050 706.050 ;
        RECT 454.950 703.950 457.050 706.050 ;
        RECT 433.950 701.250 436.050 702.150 ;
        RECT 439.950 701.250 442.050 702.150 ;
        RECT 433.950 697.950 436.050 700.050 ;
        RECT 439.950 699.450 442.050 700.050 ;
        RECT 443.400 699.450 444.450 703.950 ;
        RECT 455.400 703.050 456.450 703.950 ;
        RECT 451.950 701.250 453.750 702.150 ;
        RECT 454.950 700.950 457.050 703.050 ;
        RECT 458.250 701.250 459.750 702.150 ;
        RECT 460.950 700.950 463.050 703.050 ;
        RECT 464.250 701.250 466.050 702.150 ;
        RECT 437.250 698.250 438.750 699.150 ;
        RECT 439.950 698.400 444.450 699.450 ;
        RECT 439.950 697.950 442.050 698.400 ;
        RECT 451.950 697.950 454.050 700.050 ;
        RECT 455.250 698.850 456.750 699.750 ;
        RECT 457.950 697.950 460.050 700.050 ;
        RECT 461.250 698.850 462.750 699.750 ;
        RECT 463.950 697.950 466.050 700.050 ;
        RECT 434.400 688.050 435.450 697.950 ;
        RECT 436.950 694.950 439.050 697.050 ;
        RECT 437.400 694.050 438.450 694.950 ;
        RECT 436.950 691.950 439.050 694.050 ;
        RECT 452.400 688.050 453.450 697.950 ;
        RECT 458.400 696.450 459.450 697.950 ;
        RECT 455.400 695.400 459.450 696.450 ;
        RECT 433.950 685.950 436.050 688.050 ;
        RECT 451.950 685.950 454.050 688.050 ;
        RECT 430.950 676.950 433.050 679.050 ;
        RECT 436.950 676.950 439.050 679.050 ;
        RECT 427.950 673.950 430.050 676.050 ;
        RECT 409.950 671.250 412.050 672.150 ;
        RECT 412.950 671.850 415.050 672.750 ;
        RECT 424.950 672.450 427.050 673.050 ;
        RECT 422.400 671.400 427.050 672.450 ;
        RECT 428.250 671.850 429.750 672.750 ;
        RECT 409.950 667.950 412.050 670.050 ;
        RECT 412.950 667.950 415.050 670.050 ;
        RECT 406.950 664.950 409.050 667.050 ;
        RECT 409.950 652.950 412.050 655.050 ;
        RECT 403.950 643.950 406.050 646.050 ;
        RECT 406.950 637.950 409.050 640.050 ;
        RECT 407.400 634.050 408.450 637.950 ;
        RECT 406.950 631.950 409.050 634.050 ;
        RECT 406.950 628.950 409.050 631.050 ;
        RECT 403.950 626.250 406.050 627.150 ;
        RECT 406.950 626.850 409.050 627.750 ;
        RECT 403.950 622.950 406.050 625.050 ;
        RECT 400.950 619.950 403.050 622.050 ;
        RECT 404.400 619.050 405.450 622.950 ;
        RECT 406.950 619.950 409.050 622.050 ;
        RECT 403.950 616.950 406.050 619.050 ;
        RECT 394.950 598.950 397.050 601.050 ;
        RECT 400.950 598.950 403.050 601.050 ;
        RECT 395.400 598.050 396.450 598.950 ;
        RECT 401.400 598.050 402.450 598.950 ;
        RECT 382.950 596.250 384.750 597.150 ;
        RECT 385.950 595.950 388.050 598.050 ;
        RECT 389.250 596.250 391.050 597.150 ;
        RECT 391.950 595.950 394.050 598.050 ;
        RECT 394.950 595.950 397.050 598.050 ;
        RECT 397.950 596.250 399.750 597.150 ;
        RECT 400.950 595.950 403.050 598.050 ;
        RECT 404.250 596.250 406.050 597.150 ;
        RECT 382.950 592.950 385.050 595.050 ;
        RECT 386.250 593.850 387.750 594.750 ;
        RECT 388.950 592.950 391.050 595.050 ;
        RECT 391.950 592.950 394.050 595.050 ;
        RECT 394.950 594.450 397.050 595.050 ;
        RECT 397.950 594.450 400.050 595.050 ;
        RECT 394.950 593.400 400.050 594.450 ;
        RECT 401.250 593.850 402.750 594.750 ;
        RECT 394.950 592.950 397.050 593.400 ;
        RECT 397.950 592.950 400.050 593.400 ;
        RECT 403.950 592.950 406.050 595.050 ;
        RECT 388.950 589.950 391.050 592.050 ;
        RECT 376.950 580.950 379.050 583.050 ;
        RECT 379.950 580.950 382.050 583.050 ;
        RECT 385.950 562.950 388.050 565.050 ;
        RECT 386.400 562.050 387.450 562.950 ;
        RECT 379.950 561.450 382.050 562.050 ;
        RECT 377.400 560.400 382.050 561.450 ;
        RECT 377.400 550.050 378.450 560.400 ;
        RECT 379.950 559.950 382.050 560.400 ;
        RECT 383.250 560.250 384.750 561.150 ;
        RECT 385.950 559.950 388.050 562.050 ;
        RECT 379.950 557.850 381.750 558.750 ;
        RECT 382.950 556.950 385.050 559.050 ;
        RECT 386.250 557.850 388.050 558.750 ;
        RECT 389.400 553.050 390.450 589.950 ;
        RECT 392.400 589.050 393.450 592.950 ;
        RECT 391.950 586.950 394.050 589.050 ;
        RECT 391.950 580.950 394.050 583.050 ;
        RECT 388.950 550.950 391.050 553.050 ;
        RECT 376.950 547.950 379.050 550.050 ;
        RECT 376.950 544.950 379.050 547.050 ;
        RECT 377.400 469.050 378.450 544.950 ;
        RECT 388.950 541.950 391.050 544.050 ;
        RECT 389.400 529.050 390.450 541.950 ;
        RECT 379.950 526.950 382.050 529.050 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 388.950 526.950 391.050 529.050 ;
        RECT 379.950 524.850 382.050 525.750 ;
        RECT 382.950 524.250 385.050 525.150 ;
        RECT 382.950 520.950 385.050 523.050 ;
        RECT 386.400 493.050 387.450 526.950 ;
        RECT 388.950 524.850 391.050 525.750 ;
        RECT 392.400 499.050 393.450 580.950 ;
        RECT 395.400 550.050 396.450 592.950 ;
        RECT 400.950 586.950 403.050 589.050 ;
        RECT 397.950 580.950 400.050 583.050 ;
        RECT 398.400 571.050 399.450 580.950 ;
        RECT 397.950 568.950 400.050 571.050 ;
        RECT 401.400 559.050 402.450 586.950 ;
        RECT 407.400 570.450 408.450 619.950 ;
        RECT 410.400 574.050 411.450 652.950 ;
        RECT 413.400 619.050 414.450 667.950 ;
        RECT 422.400 636.450 423.450 671.400 ;
        RECT 424.950 670.950 427.050 671.400 ;
        RECT 430.950 670.950 433.050 673.050 ;
        RECT 424.950 668.850 427.050 669.750 ;
        RECT 430.950 668.850 433.050 669.750 ;
        RECT 419.400 635.400 423.450 636.450 ;
        RECT 415.950 631.950 418.050 634.050 ;
        RECT 412.950 616.950 415.050 619.050 ;
        RECT 416.400 598.050 417.450 631.950 ;
        RECT 419.400 630.450 420.450 635.400 ;
        RECT 424.950 635.250 427.050 636.150 ;
        RECT 433.950 634.950 436.050 637.050 ;
        RECT 421.950 632.250 423.750 633.150 ;
        RECT 424.950 631.950 427.050 634.050 ;
        RECT 428.250 632.250 429.750 633.150 ;
        RECT 430.950 631.950 433.050 634.050 ;
        RECT 421.950 630.450 424.050 631.050 ;
        RECT 427.950 630.450 430.050 631.050 ;
        RECT 419.400 629.400 424.050 630.450 ;
        RECT 421.950 628.950 424.050 629.400 ;
        RECT 425.400 629.400 430.050 630.450 ;
        RECT 431.250 629.850 433.050 630.750 ;
        RECT 425.400 616.050 426.450 629.400 ;
        RECT 427.950 628.950 430.050 629.400 ;
        RECT 434.400 625.050 435.450 634.950 ;
        RECT 437.400 631.050 438.450 676.950 ;
        RECT 451.950 673.950 454.050 676.050 ;
        RECT 448.950 670.950 451.050 673.050 ;
        RECT 439.950 667.950 442.050 670.050 ;
        RECT 442.950 668.250 444.750 669.150 ;
        RECT 445.950 667.950 448.050 670.050 ;
        RECT 440.400 652.050 441.450 667.950 ;
        RECT 449.400 667.050 450.450 670.950 ;
        RECT 452.400 670.050 453.450 673.950 ;
        RECT 451.950 667.950 454.050 670.050 ;
        RECT 442.950 664.950 445.050 667.050 ;
        RECT 446.250 665.850 447.750 666.750 ;
        RECT 448.950 664.950 451.050 667.050 ;
        RECT 452.250 665.850 454.050 666.750 ;
        RECT 439.950 649.950 442.050 652.050 ;
        RECT 443.400 643.050 444.450 664.950 ;
        RECT 448.950 662.850 451.050 663.750 ;
        RECT 455.400 655.050 456.450 695.400 ;
        RECT 466.950 676.950 469.050 679.050 ;
        RECT 467.400 670.050 468.450 676.950 ;
        RECT 470.400 676.050 471.450 706.950 ;
        RECT 473.400 706.050 474.450 734.400 ;
        RECT 475.950 730.950 478.050 733.050 ;
        RECT 472.950 703.950 475.050 706.050 ;
        RECT 469.950 673.950 472.050 676.050 ;
        RECT 463.950 668.250 465.750 669.150 ;
        RECT 466.950 667.950 469.050 670.050 ;
        RECT 470.400 667.050 471.450 673.950 ;
        RECT 473.400 670.050 474.450 703.950 ;
        RECT 476.400 700.050 477.450 730.950 ;
        RECT 479.400 712.050 480.450 743.400 ;
        RECT 478.950 709.950 481.050 712.050 ;
        RECT 485.400 709.050 486.450 745.950 ;
        RECT 488.400 742.050 489.450 773.400 ;
        RECT 490.950 772.950 493.050 773.400 ;
        RECT 490.950 770.850 493.050 771.750 ;
        RECT 493.950 770.250 496.050 771.150 ;
        RECT 493.950 766.950 496.050 769.050 ;
        RECT 490.950 751.950 493.050 754.050 ;
        RECT 491.400 745.050 492.450 751.950 ;
        RECT 497.400 748.050 498.450 808.950 ;
        RECT 500.400 808.050 501.450 811.950 ;
        RECT 506.400 810.450 507.450 814.950 ;
        RECT 508.950 812.250 510.750 813.150 ;
        RECT 511.950 811.950 514.050 814.050 ;
        RECT 515.250 812.250 517.050 813.150 ;
        RECT 508.950 810.450 511.050 811.050 ;
        RECT 506.400 809.400 511.050 810.450 ;
        RECT 512.250 809.850 513.750 810.750 ;
        RECT 508.950 808.950 511.050 809.400 ;
        RECT 514.950 808.950 517.050 811.050 ;
        RECT 499.950 805.950 502.050 808.050 ;
        RECT 524.400 790.050 525.450 818.400 ;
        RECT 526.950 817.950 529.050 818.400 ;
        RECT 530.400 817.050 531.450 820.950 ;
        RECT 533.400 820.050 534.450 844.950 ;
        RECT 547.950 842.850 550.050 843.750 ;
        RECT 550.950 842.250 553.050 843.150 ;
        RECT 550.950 838.950 553.050 841.050 ;
        RECT 541.950 835.950 544.050 838.050 ;
        RECT 532.950 817.950 535.050 820.050 ;
        RECT 526.950 815.850 528.750 816.750 ;
        RECT 529.950 814.950 532.050 817.050 ;
        RECT 535.950 815.250 538.050 816.150 ;
        RECT 538.950 814.950 541.050 817.050 ;
        RECT 529.950 812.850 532.050 813.750 ;
        RECT 535.950 811.950 538.050 814.050 ;
        RECT 523.950 787.950 526.050 790.050 ;
        RECT 532.950 781.950 535.050 784.050 ;
        RECT 533.400 778.050 534.450 781.950 ;
        RECT 526.950 776.250 529.050 777.150 ;
        RECT 532.950 775.950 535.050 778.050 ;
        RECT 533.400 775.050 534.450 775.950 ;
        RECT 505.950 773.250 508.050 774.150 ;
        RECT 511.950 773.250 514.050 774.150 ;
        RECT 526.950 772.950 529.050 775.050 ;
        RECT 530.250 773.250 531.750 774.150 ;
        RECT 532.950 772.950 535.050 775.050 ;
        RECT 536.250 773.250 538.050 774.150 ;
        RECT 505.950 769.950 508.050 772.050 ;
        RECT 509.250 770.250 510.750 771.150 ;
        RECT 511.950 769.950 514.050 772.050 ;
        RECT 506.400 769.050 507.450 769.950 ;
        RECT 505.950 766.950 508.050 769.050 ;
        RECT 508.950 766.950 511.050 769.050 ;
        RECT 509.400 753.450 510.450 766.950 ;
        RECT 506.400 752.400 510.450 753.450 ;
        RECT 496.950 745.950 499.050 748.050 ;
        RECT 506.400 745.050 507.450 752.400 ;
        RECT 512.400 751.050 513.450 769.950 ;
        RECT 527.400 769.050 528.450 772.950 ;
        RECT 529.950 769.950 532.050 772.050 ;
        RECT 533.250 770.850 534.750 771.750 ;
        RECT 535.950 771.450 538.050 772.050 ;
        RECT 539.400 771.450 540.450 814.950 ;
        RECT 535.950 770.400 540.450 771.450 ;
        RECT 535.950 769.950 538.050 770.400 ;
        RECT 526.950 766.950 529.050 769.050 ;
        RECT 508.950 748.950 511.050 751.050 ;
        RECT 511.950 748.950 514.050 751.050 ;
        RECT 526.950 748.950 529.050 751.050 ;
        RECT 509.400 745.050 510.450 748.950 ;
        RECT 527.400 748.050 528.450 748.950 ;
        RECT 530.400 748.050 531.450 769.950 ;
        RECT 532.950 766.950 535.050 769.050 ;
        RECT 514.950 745.950 517.050 748.050 ;
        RECT 523.950 745.950 526.050 748.050 ;
        RECT 526.950 745.950 529.050 748.050 ;
        RECT 529.950 745.950 532.050 748.050 ;
        RECT 490.950 742.950 493.050 745.050 ;
        RECT 494.250 743.250 495.750 744.150 ;
        RECT 496.950 742.950 499.050 745.050 ;
        RECT 505.950 742.950 508.050 745.050 ;
        RECT 508.950 742.950 511.050 745.050 ;
        RECT 512.250 743.250 514.050 744.150 ;
        RECT 514.950 743.850 517.050 744.750 ;
        RECT 517.950 743.250 520.050 744.150 ;
        RECT 506.400 742.050 507.450 742.950 ;
        RECT 487.950 739.950 490.050 742.050 ;
        RECT 491.250 740.850 492.750 741.750 ;
        RECT 493.950 739.950 496.050 742.050 ;
        RECT 497.250 740.850 499.050 741.750 ;
        RECT 505.950 739.950 508.050 742.050 ;
        RECT 508.950 740.850 510.750 741.750 ;
        RECT 511.950 739.950 514.050 742.050 ;
        RECT 514.950 739.950 517.050 742.050 ;
        RECT 517.950 739.950 520.050 742.050 ;
        RECT 487.950 737.850 490.050 738.750 ;
        RECT 494.400 733.050 495.450 739.950 ;
        RECT 515.400 736.050 516.450 739.950 ;
        RECT 514.950 733.950 517.050 736.050 ;
        RECT 493.950 730.950 496.050 733.050 ;
        RECT 496.950 727.950 499.050 730.050 ;
        RECT 484.950 706.950 487.050 709.050 ;
        RECT 485.400 706.050 486.450 706.950 ;
        RECT 497.400 706.050 498.450 727.950 ;
        RECT 514.950 718.950 517.050 721.050 ;
        RECT 508.950 715.950 511.050 718.050 ;
        RECT 502.950 707.250 505.050 708.150 ;
        RECT 478.950 703.950 481.050 706.050 ;
        RECT 482.250 704.250 483.750 705.150 ;
        RECT 484.950 703.950 487.050 706.050 ;
        RECT 496.950 703.950 499.050 706.050 ;
        RECT 500.250 704.250 501.750 705.150 ;
        RECT 502.950 703.950 505.050 706.050 ;
        RECT 506.250 704.250 508.050 705.150 ;
        RECT 478.950 701.850 480.750 702.750 ;
        RECT 481.950 700.950 484.050 703.050 ;
        RECT 485.250 701.850 487.050 702.750 ;
        RECT 487.950 700.950 490.050 703.050 ;
        RECT 496.950 701.850 498.750 702.750 ;
        RECT 499.950 700.950 502.050 703.050 ;
        RECT 475.950 697.950 478.050 700.050 ;
        RECT 475.950 694.950 478.050 697.050 ;
        RECT 472.950 667.950 475.050 670.050 ;
        RECT 463.950 664.950 466.050 667.050 ;
        RECT 467.250 665.850 468.750 666.750 ;
        RECT 469.950 664.950 472.050 667.050 ;
        RECT 473.250 665.850 475.050 666.750 ;
        RECT 454.950 652.950 457.050 655.050 ;
        RECT 448.950 649.950 451.050 652.050 ;
        RECT 454.950 649.950 457.050 652.050 ;
        RECT 442.950 640.950 445.050 643.050 ;
        RECT 449.400 634.050 450.450 649.950 ;
        RECT 451.950 634.950 454.050 637.050 ;
        RECT 442.950 631.950 445.050 634.050 ;
        RECT 446.250 632.250 447.750 633.150 ;
        RECT 448.950 631.950 451.050 634.050 ;
        RECT 436.950 628.950 439.050 631.050 ;
        RECT 442.950 629.850 444.750 630.750 ;
        RECT 445.950 628.950 448.050 631.050 ;
        RECT 449.250 629.850 451.050 630.750 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 433.950 622.950 436.050 625.050 ;
        RECT 427.950 619.950 430.050 622.050 ;
        RECT 424.950 613.950 427.050 616.050 ;
        RECT 425.400 613.050 426.450 613.950 ;
        RECT 424.950 610.950 427.050 613.050 ;
        RECT 421.950 604.950 424.050 607.050 ;
        RECT 422.400 601.050 423.450 604.950 ;
        RECT 421.950 598.950 424.050 601.050 ;
        RECT 422.400 598.050 423.450 598.950 ;
        RECT 412.950 595.950 415.050 598.050 ;
        RECT 415.950 595.950 418.050 598.050 ;
        RECT 421.950 595.950 424.050 598.050 ;
        RECT 425.250 596.250 427.050 597.150 ;
        RECT 413.400 595.050 414.450 595.950 ;
        RECT 412.950 592.950 415.050 595.050 ;
        RECT 415.950 593.850 417.750 594.750 ;
        RECT 418.950 592.950 421.050 595.050 ;
        RECT 422.250 593.850 423.750 594.750 ;
        RECT 424.950 592.950 427.050 595.050 ;
        RECT 413.400 591.450 414.450 592.950 ;
        RECT 413.400 590.400 417.450 591.450 ;
        RECT 418.950 590.850 421.050 591.750 ;
        RECT 412.950 577.950 415.050 580.050 ;
        RECT 409.950 571.950 412.050 574.050 ;
        RECT 407.400 569.400 411.450 570.450 ;
        RECT 403.950 565.950 406.050 568.050 ;
        RECT 404.400 562.050 405.450 565.950 ;
        RECT 403.950 559.950 406.050 562.050 ;
        RECT 406.950 560.250 409.050 561.150 ;
        RECT 397.950 557.250 399.750 558.150 ;
        RECT 400.950 556.950 403.050 559.050 ;
        RECT 404.250 557.250 405.750 558.150 ;
        RECT 406.950 556.950 409.050 559.050 ;
        RECT 397.950 553.950 400.050 556.050 ;
        RECT 401.250 554.850 402.750 555.750 ;
        RECT 403.950 553.950 406.050 556.050 ;
        RECT 406.950 553.950 409.050 556.050 ;
        RECT 394.950 547.950 397.050 550.050 ;
        RECT 398.400 546.450 399.450 553.950 ;
        RECT 404.400 553.050 405.450 553.950 ;
        RECT 403.950 550.950 406.050 553.050 ;
        RECT 395.400 545.400 399.450 546.450 ;
        RECT 391.950 496.950 394.050 499.050 ;
        RECT 385.950 490.950 388.050 493.050 ;
        RECT 382.950 488.250 385.050 489.150 ;
        RECT 382.950 484.950 385.050 487.050 ;
        RECT 386.250 485.250 387.750 486.150 ;
        RECT 388.950 484.950 391.050 487.050 ;
        RECT 392.250 485.250 394.050 486.150 ;
        RECT 383.400 478.050 384.450 484.950 ;
        RECT 385.950 481.950 388.050 484.050 ;
        RECT 389.250 482.850 390.750 483.750 ;
        RECT 391.950 481.950 394.050 484.050 ;
        RECT 382.950 475.950 385.050 478.050 ;
        RECT 392.400 475.050 393.450 481.950 ;
        RECT 391.950 472.950 394.050 475.050 ;
        RECT 388.950 469.950 391.050 472.050 ;
        RECT 376.950 466.950 379.050 469.050 ;
        RECT 385.950 466.950 388.050 469.050 ;
        RECT 376.950 463.950 379.050 466.050 ;
        RECT 377.400 457.050 378.450 463.950 ;
        RECT 386.400 460.050 387.450 466.950 ;
        RECT 382.950 457.950 385.050 460.050 ;
        RECT 385.950 457.950 388.050 460.050 ;
        RECT 376.950 454.950 379.050 457.050 ;
        RECT 380.250 455.250 382.050 456.150 ;
        RECT 382.950 455.850 385.050 456.750 ;
        RECT 385.950 455.250 388.050 456.150 ;
        RECT 376.950 452.850 378.750 453.750 ;
        RECT 379.950 451.950 382.050 454.050 ;
        RECT 385.950 451.950 388.050 454.050 ;
        RECT 374.400 449.400 378.450 450.450 ;
        RECT 367.950 415.950 370.050 418.050 ;
        RECT 367.950 413.250 370.050 414.150 ;
        RECT 373.950 413.250 376.050 414.150 ;
        RECT 367.950 409.950 370.050 412.050 ;
        RECT 371.250 410.250 372.750 411.150 ;
        RECT 373.950 409.950 376.050 412.050 ;
        RECT 367.950 406.950 370.050 409.050 ;
        RECT 370.950 406.950 373.050 409.050 ;
        RECT 364.950 382.950 367.050 385.050 ;
        RECT 358.950 380.250 360.750 381.150 ;
        RECT 361.950 379.950 364.050 382.050 ;
        RECT 365.250 380.250 367.050 381.150 ;
        RECT 358.950 376.950 361.050 379.050 ;
        RECT 362.250 377.850 363.750 378.750 ;
        RECT 364.950 376.950 367.050 379.050 ;
        RECT 368.400 376.050 369.450 406.950 ;
        RECT 371.400 406.050 372.450 406.950 ;
        RECT 374.400 406.050 375.450 409.950 ;
        RECT 370.950 403.950 373.050 406.050 ;
        RECT 373.950 403.950 376.050 406.050 ;
        RECT 371.400 379.050 372.450 403.950 ;
        RECT 374.400 382.050 375.450 403.950 ;
        RECT 377.400 394.050 378.450 449.400 ;
        RECT 379.950 448.950 382.050 451.050 ;
        RECT 376.950 391.950 379.050 394.050 ;
        RECT 380.400 390.450 381.450 448.950 ;
        RECT 386.400 424.050 387.450 451.950 ;
        RECT 389.400 451.050 390.450 469.950 ;
        RECT 395.400 466.050 396.450 545.400 ;
        RECT 397.950 524.250 399.750 525.150 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 404.250 524.250 406.050 525.150 ;
        RECT 407.400 523.050 408.450 553.950 ;
        RECT 410.400 547.050 411.450 569.400 ;
        RECT 409.950 544.950 412.050 547.050 ;
        RECT 409.950 541.950 412.050 544.050 ;
        RECT 410.400 526.050 411.450 541.950 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 397.950 520.950 400.050 523.050 ;
        RECT 401.250 521.850 402.750 522.750 ;
        RECT 403.950 520.950 406.050 523.050 ;
        RECT 406.950 520.950 409.050 523.050 ;
        RECT 398.400 505.050 399.450 520.950 ;
        RECT 397.950 502.950 400.050 505.050 ;
        RECT 413.400 502.050 414.450 577.950 ;
        RECT 412.950 499.950 415.050 502.050 ;
        RECT 412.950 496.950 415.050 499.050 ;
        RECT 400.950 493.950 403.050 496.050 ;
        RECT 397.950 490.950 400.050 493.050 ;
        RECT 398.400 481.050 399.450 490.950 ;
        RECT 397.950 478.950 400.050 481.050 ;
        RECT 397.950 475.950 400.050 478.050 ;
        RECT 394.950 463.950 397.050 466.050 ;
        RECT 395.400 463.050 396.450 463.950 ;
        RECT 394.950 460.950 397.050 463.050 ;
        RECT 398.400 457.050 399.450 475.950 ;
        RECT 401.400 463.050 402.450 493.950 ;
        RECT 406.950 487.950 409.050 490.050 ;
        RECT 407.400 487.050 408.450 487.950 ;
        RECT 413.400 487.050 414.450 496.950 ;
        RECT 416.400 493.050 417.450 590.400 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 418.950 559.950 421.050 562.050 ;
        RECT 419.400 553.050 420.450 559.950 ;
        RECT 422.400 559.050 423.450 568.950 ;
        RECT 425.400 565.050 426.450 592.950 ;
        RECT 424.950 562.950 427.050 565.050 ;
        RECT 425.400 559.050 426.450 562.950 ;
        RECT 421.950 556.950 424.050 559.050 ;
        RECT 424.950 556.950 427.050 559.050 ;
        RECT 421.950 554.850 424.050 555.750 ;
        RECT 424.950 554.250 427.050 555.150 ;
        RECT 418.950 550.950 421.050 553.050 ;
        RECT 424.950 550.950 427.050 553.050 ;
        RECT 428.400 529.050 429.450 619.950 ;
        RECT 431.400 607.050 432.450 622.950 ;
        RECT 430.950 604.950 433.050 607.050 ;
        RECT 430.950 601.950 433.050 604.050 ;
        RECT 431.400 592.050 432.450 601.950 ;
        RECT 437.400 600.450 438.450 628.950 ;
        RECT 442.950 616.950 445.050 619.050 ;
        RECT 434.400 599.400 438.450 600.450 ;
        RECT 430.950 589.950 433.050 592.050 ;
        RECT 434.400 576.450 435.450 599.400 ;
        RECT 443.400 598.050 444.450 616.950 ;
        RECT 446.400 610.050 447.450 628.950 ;
        RECT 445.950 607.950 448.050 610.050 ;
        RECT 452.400 606.450 453.450 634.950 ;
        RECT 455.400 628.050 456.450 649.950 ;
        RECT 460.950 630.450 463.050 631.050 ;
        RECT 458.400 629.400 463.050 630.450 ;
        RECT 464.400 630.450 465.450 664.950 ;
        RECT 469.950 662.850 472.050 663.750 ;
        RECT 472.950 655.950 475.050 658.050 ;
        RECT 466.950 630.450 469.050 631.050 ;
        RECT 464.400 629.400 469.050 630.450 ;
        RECT 454.950 625.950 457.050 628.050 ;
        RECT 458.400 616.050 459.450 629.400 ;
        RECT 460.950 628.950 463.050 629.400 ;
        RECT 466.950 628.950 469.050 629.400 ;
        RECT 470.250 629.250 472.050 630.150 ;
        RECT 460.950 626.850 463.050 627.750 ;
        RECT 463.950 626.250 466.050 627.150 ;
        RECT 466.950 626.850 468.750 627.750 ;
        RECT 469.950 625.950 472.050 628.050 ;
        RECT 463.950 624.450 466.050 625.050 ;
        RECT 466.950 624.450 469.050 625.050 ;
        RECT 463.950 623.400 469.050 624.450 ;
        RECT 463.950 622.950 466.050 623.400 ;
        RECT 466.950 622.950 469.050 623.400 ;
        RECT 460.950 616.950 463.050 619.050 ;
        RECT 457.950 613.950 460.050 616.050 ;
        RECT 449.400 605.400 453.450 606.450 ;
        RECT 449.400 604.050 450.450 605.400 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 461.400 603.450 462.450 616.950 ;
        RECT 458.400 602.400 462.450 603.450 ;
        RECT 436.950 595.950 439.050 598.050 ;
        RECT 442.950 595.950 445.050 598.050 ;
        RECT 446.250 596.250 448.050 597.150 ;
        RECT 448.950 595.950 451.050 598.050 ;
        RECT 436.950 593.850 438.750 594.750 ;
        RECT 439.950 592.950 442.050 595.050 ;
        RECT 443.250 593.850 444.750 594.750 ;
        RECT 445.950 592.950 448.050 595.050 ;
        RECT 439.950 590.850 442.050 591.750 ;
        RECT 442.950 589.950 445.050 592.050 ;
        RECT 443.400 583.050 444.450 589.950 ;
        RECT 449.400 589.050 450.450 595.950 ;
        RECT 455.400 595.050 456.450 601.950 ;
        RECT 454.950 592.950 457.050 595.050 ;
        RECT 458.400 592.050 459.450 602.400 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 460.950 599.250 463.050 600.150 ;
        RECT 463.950 599.850 466.050 600.750 ;
        RECT 460.950 595.950 463.050 598.050 ;
        RECT 457.950 589.950 460.050 592.050 ;
        RECT 448.950 586.950 451.050 589.050 ;
        RECT 448.950 583.950 451.050 586.050 ;
        RECT 451.950 583.950 454.050 586.050 ;
        RECT 442.950 580.950 445.050 583.050 ;
        RECT 431.400 575.400 435.450 576.450 ;
        RECT 431.400 529.050 432.450 575.400 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 436.950 560.250 439.050 561.150 ;
        RECT 443.400 559.050 444.450 568.950 ;
        RECT 436.950 556.950 439.050 559.050 ;
        RECT 440.250 557.250 441.750 558.150 ;
        RECT 442.950 556.950 445.050 559.050 ;
        RECT 446.250 557.250 448.050 558.150 ;
        RECT 449.400 556.050 450.450 583.950 ;
        RECT 439.950 553.950 442.050 556.050 ;
        RECT 443.250 554.850 444.750 555.750 ;
        RECT 445.950 553.950 448.050 556.050 ;
        RECT 448.950 553.950 451.050 556.050 ;
        RECT 446.400 553.050 447.450 553.950 ;
        RECT 445.950 550.950 448.050 553.050 ;
        RECT 439.950 547.950 442.050 550.050 ;
        RECT 433.950 535.950 436.050 538.050 ;
        RECT 421.950 526.950 424.050 529.050 ;
        RECT 425.250 527.250 426.750 528.150 ;
        RECT 427.950 526.950 430.050 529.050 ;
        RECT 430.950 526.950 433.050 529.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 422.250 524.850 423.750 525.750 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 428.250 524.850 430.050 525.750 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 425.400 523.050 426.450 523.950 ;
        RECT 418.950 521.850 421.050 522.750 ;
        RECT 424.950 520.950 427.050 523.050 ;
        RECT 427.950 520.950 430.050 523.050 ;
        RECT 428.400 508.050 429.450 520.950 ;
        RECT 427.950 505.950 430.050 508.050 ;
        RECT 418.950 499.950 421.050 502.050 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 419.400 489.450 420.450 499.950 ;
        RECT 431.400 496.050 432.450 523.950 ;
        RECT 430.950 493.950 433.050 496.050 ;
        RECT 424.950 491.250 427.050 492.150 ;
        RECT 431.400 490.050 432.450 493.950 ;
        RECT 416.400 488.400 420.450 489.450 ;
        RECT 403.950 485.250 405.750 486.150 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 412.950 484.950 415.050 487.050 ;
        RECT 403.950 481.950 406.050 484.050 ;
        RECT 407.250 482.850 409.050 483.750 ;
        RECT 409.950 482.250 412.050 483.150 ;
        RECT 412.950 482.850 415.050 483.750 ;
        RECT 409.950 478.950 412.050 481.050 ;
        RECT 416.400 480.450 417.450 488.400 ;
        RECT 421.950 488.250 423.750 489.150 ;
        RECT 424.950 487.950 427.050 490.050 ;
        RECT 428.250 488.250 429.750 489.150 ;
        RECT 430.950 487.950 433.050 490.050 ;
        RECT 425.400 487.050 426.450 487.950 ;
        RECT 418.950 484.950 421.050 487.050 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 427.950 484.950 430.050 487.050 ;
        RECT 431.250 485.850 433.050 486.750 ;
        RECT 419.400 484.050 420.450 484.950 ;
        RECT 418.950 481.950 421.050 484.050 ;
        RECT 424.950 481.950 427.050 484.050 ;
        RECT 416.400 479.400 420.450 480.450 ;
        RECT 403.950 466.950 406.050 469.050 ;
        RECT 412.950 466.950 415.050 469.050 ;
        RECT 400.950 460.950 403.050 463.050 ;
        RECT 404.400 457.050 405.450 466.950 ;
        RECT 397.950 454.950 400.050 457.050 ;
        RECT 401.250 455.250 402.750 456.150 ;
        RECT 403.950 454.950 406.050 457.050 ;
        RECT 407.250 455.250 408.750 456.150 ;
        RECT 409.950 454.950 412.050 457.050 ;
        RECT 397.950 452.850 399.750 453.750 ;
        RECT 400.950 451.950 403.050 454.050 ;
        RECT 404.250 452.850 405.750 453.750 ;
        RECT 406.950 451.950 409.050 454.050 ;
        RECT 410.250 452.850 412.050 453.750 ;
        RECT 401.400 451.050 402.450 451.950 ;
        RECT 388.950 448.950 391.050 451.050 ;
        RECT 400.950 448.950 403.050 451.050 ;
        RECT 403.950 448.950 406.050 451.050 ;
        RECT 388.950 436.950 391.050 439.050 ;
        RECT 385.950 421.950 388.050 424.050 ;
        RECT 386.400 411.450 387.450 421.950 ;
        RECT 389.400 418.050 390.450 436.950 ;
        RECT 394.950 419.250 397.050 420.150 ;
        RECT 401.400 418.050 402.450 448.950 ;
        RECT 388.950 415.950 391.050 418.050 ;
        RECT 392.250 416.250 393.750 417.150 ;
        RECT 394.950 415.950 397.050 418.050 ;
        RECT 398.250 416.250 400.050 417.150 ;
        RECT 400.950 415.950 403.050 418.050 ;
        RECT 388.950 413.850 390.750 414.750 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 392.400 411.450 393.450 412.950 ;
        RECT 386.400 410.400 393.450 411.450 ;
        RECT 395.400 393.450 396.450 415.950 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 404.400 412.050 405.450 448.950 ;
        RECT 407.400 448.050 408.450 451.950 ;
        RECT 406.950 445.950 409.050 448.050 ;
        RECT 406.950 442.950 409.050 445.050 ;
        RECT 403.950 409.950 406.050 412.050 ;
        RECT 397.950 406.950 400.050 409.050 ;
        RECT 392.400 392.400 396.450 393.450 ;
        RECT 392.400 391.050 393.450 392.400 ;
        RECT 377.400 389.400 381.450 390.450 ;
        RECT 373.950 379.950 376.050 382.050 ;
        RECT 370.950 376.950 373.050 379.050 ;
        RECT 373.950 376.950 376.050 379.050 ;
        RECT 364.950 373.950 367.050 376.050 ;
        RECT 367.950 373.950 370.050 376.050 ;
        RECT 355.950 355.950 358.050 358.050 ;
        RECT 355.950 352.950 358.050 355.050 ;
        RECT 358.950 352.950 361.050 355.050 ;
        RECT 361.950 352.950 364.050 355.050 ;
        RECT 356.250 334.050 357.450 352.950 ;
        RECT 359.250 348.750 360.450 352.950 ;
        RECT 358.950 346.650 361.050 348.750 ;
        RECT 359.250 334.050 360.450 346.650 ;
        RECT 362.250 334.050 363.450 352.950 ;
        RECT 365.400 339.450 366.450 373.950 ;
        RECT 374.400 373.050 375.450 376.950 ;
        RECT 373.950 370.950 376.050 373.050 ;
        RECT 377.400 355.050 378.450 389.400 ;
        RECT 385.950 388.950 388.050 391.050 ;
        RECT 391.950 388.950 394.050 391.050 ;
        RECT 394.950 388.950 397.050 391.050 ;
        RECT 382.950 385.950 385.050 388.050 ;
        RECT 383.400 382.050 384.450 385.950 ;
        RECT 386.400 385.050 387.450 388.950 ;
        RECT 385.950 382.950 388.050 385.050 ;
        RECT 389.250 383.250 390.750 384.150 ;
        RECT 391.950 382.950 394.050 385.050 ;
        RECT 382.950 379.950 385.050 382.050 ;
        RECT 386.250 380.850 387.750 381.750 ;
        RECT 388.950 379.950 391.050 382.050 ;
        RECT 392.250 380.850 394.050 381.750 ;
        RECT 382.950 377.850 385.050 378.750 ;
        RECT 389.400 373.050 390.450 379.950 ;
        RECT 388.950 370.950 391.050 373.050 ;
        RECT 382.950 361.950 385.050 364.050 ;
        RECT 376.950 352.950 379.050 355.050 ;
        RECT 373.950 345.450 376.050 346.050 ;
        RECT 367.950 344.250 370.050 345.150 ;
        RECT 371.400 344.400 376.050 345.450 ;
        RECT 365.400 338.400 369.450 339.450 ;
        RECT 355.950 331.950 358.050 334.050 ;
        RECT 358.950 331.950 361.050 334.050 ;
        RECT 361.950 331.950 364.050 334.050 ;
        RECT 353.400 329.400 357.450 330.450 ;
        RECT 352.950 311.250 355.050 312.150 ;
        RECT 346.950 308.400 351.450 309.450 ;
        RECT 346.950 307.950 349.050 308.400 ;
        RECT 337.950 304.950 340.050 307.050 ;
        RECT 341.250 305.850 342.750 306.750 ;
        RECT 343.950 304.950 346.050 307.050 ;
        RECT 347.250 305.850 349.050 306.750 ;
        RECT 338.400 295.050 339.450 304.950 ;
        RECT 343.950 302.850 346.050 303.750 ;
        RECT 343.950 298.950 346.050 301.050 ;
        RECT 337.950 292.950 340.050 295.050 ;
        RECT 337.950 271.950 340.050 274.050 ;
        RECT 340.950 272.250 343.050 273.150 ;
        RECT 334.950 268.950 337.050 271.050 ;
        RECT 335.400 256.050 336.450 268.950 ;
        RECT 334.950 253.950 337.050 256.050 ;
        RECT 338.400 249.450 339.450 271.950 ;
        RECT 340.950 268.950 343.050 271.050 ;
        RECT 344.400 264.450 345.450 298.950 ;
        RECT 350.400 292.050 351.450 308.400 ;
        RECT 352.950 307.950 355.050 310.050 ;
        RECT 353.400 304.050 354.450 307.950 ;
        RECT 352.950 301.950 355.050 304.050 ;
        RECT 356.400 301.050 357.450 329.400 ;
        RECT 364.950 322.950 367.050 325.050 ;
        RECT 361.950 313.950 364.050 316.050 ;
        RECT 355.950 298.950 358.050 301.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 362.400 286.050 363.450 313.950 ;
        RECT 365.400 310.050 366.450 322.950 ;
        RECT 364.950 307.950 367.050 310.050 ;
        RECT 364.950 305.850 367.050 306.750 ;
        RECT 368.400 294.450 369.450 338.400 ;
        RECT 371.400 310.050 372.450 344.400 ;
        RECT 373.950 343.950 376.050 344.400 ;
        RECT 373.950 341.850 376.050 342.750 ;
        RECT 377.400 328.050 378.450 352.950 ;
        RECT 383.400 328.050 384.450 361.950 ;
        RECT 395.400 360.450 396.450 388.950 ;
        RECT 392.400 359.400 396.450 360.450 ;
        RECT 388.950 341.250 391.050 342.150 ;
        RECT 388.950 337.950 391.050 340.050 ;
        RECT 389.400 334.050 390.450 337.950 ;
        RECT 392.400 336.450 393.450 359.400 ;
        RECT 398.400 346.050 399.450 406.950 ;
        RECT 404.400 387.450 405.450 409.950 ;
        RECT 407.400 388.050 408.450 442.950 ;
        RECT 413.400 421.050 414.450 466.950 ;
        RECT 415.950 460.950 418.050 463.050 ;
        RECT 416.400 457.050 417.450 460.950 ;
        RECT 415.950 454.950 418.050 457.050 ;
        RECT 419.400 450.450 420.450 479.400 ;
        RECT 421.950 455.250 424.050 456.150 ;
        RECT 421.950 453.450 424.050 454.050 ;
        RECT 425.400 453.450 426.450 481.950 ;
        RECT 428.400 481.050 429.450 484.950 ;
        RECT 427.950 478.950 430.050 481.050 ;
        RECT 430.950 477.450 433.050 478.050 ;
        RECT 428.400 476.400 433.050 477.450 ;
        RECT 428.400 472.050 429.450 476.400 ;
        RECT 430.950 475.950 433.050 476.400 ;
        RECT 427.950 469.950 430.050 472.050 ;
        RECT 430.950 460.950 433.050 463.050 ;
        RECT 431.400 460.050 432.450 460.950 ;
        RECT 430.950 457.950 433.050 460.050 ;
        RECT 427.950 454.950 430.050 457.050 ;
        RECT 431.250 455.850 433.050 456.750 ;
        RECT 421.950 452.400 426.450 453.450 ;
        RECT 427.950 452.850 430.050 453.750 ;
        RECT 421.950 451.950 424.050 452.400 ;
        RECT 430.950 451.950 433.050 454.050 ;
        RECT 419.400 449.400 423.450 450.450 ;
        RECT 415.950 427.950 418.050 430.050 ;
        RECT 412.950 418.950 415.050 421.050 ;
        RECT 412.950 415.950 415.050 418.050 ;
        RECT 409.950 413.250 412.050 414.150 ;
        RECT 412.950 413.850 415.050 414.750 ;
        RECT 409.950 409.950 412.050 412.050 ;
        RECT 416.400 411.450 417.450 427.950 ;
        RECT 418.950 413.250 421.050 414.150 ;
        RECT 418.950 411.450 421.050 412.050 ;
        RECT 416.400 410.400 421.050 411.450 ;
        RECT 418.950 409.950 421.050 410.400 ;
        RECT 410.400 406.050 411.450 409.950 ;
        RECT 422.400 408.450 423.450 449.400 ;
        RECT 427.950 430.950 430.050 433.050 ;
        RECT 424.950 418.950 427.050 421.050 ;
        RECT 425.400 415.050 426.450 418.950 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 424.950 409.950 427.050 412.050 ;
        RECT 419.400 407.400 423.450 408.450 ;
        RECT 409.950 403.950 412.050 406.050 ;
        RECT 401.400 386.400 405.450 387.450 ;
        RECT 401.400 385.050 402.450 386.400 ;
        RECT 406.950 385.950 409.050 388.050 ;
        RECT 415.950 385.950 418.050 388.050 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 404.250 383.250 405.750 384.150 ;
        RECT 406.950 382.950 409.050 385.050 ;
        RECT 400.950 380.850 402.750 381.750 ;
        RECT 403.950 379.950 406.050 382.050 ;
        RECT 407.250 380.850 408.750 381.750 ;
        RECT 409.950 381.450 412.050 382.050 ;
        RECT 409.950 380.400 414.450 381.450 ;
        RECT 409.950 379.950 412.050 380.400 ;
        RECT 404.400 373.050 405.450 379.950 ;
        RECT 406.950 376.950 409.050 379.050 ;
        RECT 409.950 377.850 412.050 378.750 ;
        RECT 403.950 370.950 406.050 373.050 ;
        RECT 397.950 343.950 400.050 346.050 ;
        RECT 407.400 345.450 408.450 376.950 ;
        RECT 413.400 376.050 414.450 380.400 ;
        RECT 412.950 373.950 415.050 376.050 ;
        RECT 416.400 367.050 417.450 385.950 ;
        RECT 415.950 364.950 418.050 367.050 ;
        RECT 419.400 346.050 420.450 407.400 ;
        RECT 421.950 403.950 424.050 406.050 ;
        RECT 422.400 391.050 423.450 403.950 ;
        RECT 421.950 388.950 424.050 391.050 ;
        RECT 425.400 387.450 426.450 409.950 ;
        RECT 422.400 386.400 426.450 387.450 ;
        RECT 428.400 387.450 429.450 430.950 ;
        RECT 431.400 430.050 432.450 451.950 ;
        RECT 434.400 445.050 435.450 535.950 ;
        RECT 440.400 528.450 441.450 547.950 ;
        RECT 448.950 529.950 451.050 532.050 ;
        RECT 449.400 529.050 450.450 529.950 ;
        RECT 442.950 528.450 445.050 529.050 ;
        RECT 440.400 527.400 445.050 528.450 ;
        RECT 436.950 493.950 439.050 496.050 ;
        RECT 437.400 487.050 438.450 493.950 ;
        RECT 440.400 490.050 441.450 527.400 ;
        RECT 442.950 526.950 445.050 527.400 ;
        RECT 448.950 526.950 451.050 529.050 ;
        RECT 442.950 524.850 445.050 525.750 ;
        RECT 448.950 524.850 451.050 525.750 ;
        RECT 452.400 520.050 453.450 583.950 ;
        RECT 461.400 565.050 462.450 595.950 ;
        RECT 467.400 577.050 468.450 622.950 ;
        RECT 470.400 619.050 471.450 625.950 ;
        RECT 473.400 619.050 474.450 655.950 ;
        RECT 469.950 616.950 472.050 619.050 ;
        RECT 472.950 616.950 475.050 619.050 ;
        RECT 472.950 607.950 475.050 610.050 ;
        RECT 469.950 604.950 472.050 607.050 ;
        RECT 470.400 577.050 471.450 604.950 ;
        RECT 466.950 574.950 469.050 577.050 ;
        RECT 469.950 574.950 472.050 577.050 ;
        RECT 466.950 568.950 469.050 571.050 ;
        RECT 460.950 562.950 463.050 565.050 ;
        RECT 454.950 559.950 457.050 562.050 ;
        RECT 458.250 560.250 459.750 561.150 ;
        RECT 460.950 559.950 463.050 562.050 ;
        RECT 454.950 557.850 456.750 558.750 ;
        RECT 457.950 556.950 460.050 559.050 ;
        RECT 461.250 557.850 463.050 558.750 ;
        RECT 454.950 553.950 457.050 556.050 ;
        RECT 455.400 532.050 456.450 553.950 ;
        RECT 458.400 532.050 459.450 556.950 ;
        RECT 467.400 556.050 468.450 568.950 ;
        RECT 466.950 553.950 469.050 556.050 ;
        RECT 469.950 550.950 472.050 553.050 ;
        RECT 460.950 547.950 463.050 550.050 ;
        RECT 461.400 541.050 462.450 547.950 ;
        RECT 460.950 538.950 463.050 541.050 ;
        RECT 463.950 538.950 466.050 541.050 ;
        RECT 454.950 529.950 457.050 532.050 ;
        RECT 457.950 529.950 460.050 532.050 ;
        RECT 451.950 517.950 454.050 520.050 ;
        RECT 455.400 499.050 456.450 529.950 ;
        RECT 457.950 526.950 460.050 529.050 ;
        RECT 458.400 526.050 459.450 526.950 ;
        RECT 464.400 526.050 465.450 538.950 ;
        RECT 457.950 523.950 460.050 526.050 ;
        RECT 460.950 524.250 462.750 525.150 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 467.250 524.250 469.050 525.150 ;
        RECT 458.400 522.450 459.450 523.950 ;
        RECT 460.950 522.450 463.050 523.050 ;
        RECT 458.400 521.400 463.050 522.450 ;
        RECT 464.250 521.850 465.750 522.750 ;
        RECT 460.950 520.950 463.050 521.400 ;
        RECT 466.950 520.950 469.050 523.050 ;
        RECT 467.400 520.050 468.450 520.950 ;
        RECT 457.950 517.950 460.050 520.050 ;
        RECT 466.950 517.950 469.050 520.050 ;
        RECT 454.950 496.950 457.050 499.050 ;
        RECT 445.950 491.250 448.050 492.150 ;
        RECT 439.950 487.950 442.050 490.050 ;
        RECT 442.950 488.250 444.750 489.150 ;
        RECT 445.950 487.950 448.050 490.050 ;
        RECT 451.950 489.450 454.050 490.050 ;
        RECT 449.250 488.250 450.750 489.150 ;
        RECT 451.950 488.400 456.450 489.450 ;
        RECT 451.950 487.950 454.050 488.400 ;
        RECT 436.950 484.950 439.050 487.050 ;
        RECT 440.400 486.450 441.450 487.950 ;
        RECT 442.950 486.450 445.050 487.050 ;
        RECT 440.400 485.400 445.050 486.450 ;
        RECT 442.950 484.950 445.050 485.400 ;
        RECT 446.400 484.050 447.450 487.950 ;
        RECT 448.950 484.950 451.050 487.050 ;
        RECT 452.250 485.850 454.050 486.750 ;
        RECT 439.950 481.950 442.050 484.050 ;
        RECT 445.950 481.950 448.050 484.050 ;
        RECT 440.400 478.050 441.450 481.950 ;
        RECT 449.400 480.450 450.450 484.950 ;
        RECT 451.950 481.950 454.050 484.050 ;
        RECT 446.400 479.400 450.450 480.450 ;
        RECT 436.950 475.950 439.050 478.050 ;
        RECT 439.950 475.950 442.050 478.050 ;
        RECT 433.950 442.950 436.050 445.050 ;
        RECT 433.950 430.950 436.050 433.050 ;
        RECT 430.950 427.950 433.050 430.050 ;
        RECT 434.400 415.050 435.450 430.950 ;
        RECT 437.400 421.050 438.450 475.950 ;
        RECT 439.950 460.950 442.050 463.050 ;
        RECT 440.400 457.050 441.450 460.950 ;
        RECT 446.400 460.050 447.450 479.400 ;
        RECT 442.950 457.950 445.050 460.050 ;
        RECT 445.950 457.950 448.050 460.050 ;
        RECT 439.950 454.950 442.050 457.050 ;
        RECT 443.250 455.850 444.750 456.750 ;
        RECT 445.950 456.450 448.050 457.050 ;
        RECT 445.950 455.400 450.450 456.450 ;
        RECT 445.950 454.950 448.050 455.400 ;
        RECT 439.950 452.850 442.050 453.750 ;
        RECT 445.950 452.850 448.050 453.750 ;
        RECT 445.950 436.950 448.050 439.050 ;
        RECT 436.950 418.950 439.050 421.050 ;
        RECT 439.950 416.250 442.050 417.150 ;
        RECT 430.950 413.250 432.750 414.150 ;
        RECT 433.950 412.950 436.050 415.050 ;
        RECT 437.250 413.250 438.750 414.150 ;
        RECT 430.950 409.950 433.050 412.050 ;
        RECT 434.250 410.850 435.750 411.750 ;
        RECT 436.950 409.950 439.050 412.050 ;
        RECT 431.400 409.050 432.450 409.950 ;
        RECT 430.950 406.950 433.050 409.050 ;
        RECT 436.950 406.950 439.050 409.050 ;
        RECT 430.950 387.450 433.050 388.050 ;
        RECT 428.400 386.400 433.050 387.450 ;
        RECT 422.400 382.050 423.450 386.400 ;
        RECT 430.950 385.950 433.050 386.400 ;
        RECT 424.950 382.950 427.050 385.050 ;
        RECT 428.250 383.250 430.050 384.150 ;
        RECT 430.950 383.850 433.050 384.750 ;
        RECT 433.950 383.250 436.050 384.150 ;
        RECT 421.950 379.950 424.050 382.050 ;
        RECT 424.950 380.850 426.750 381.750 ;
        RECT 427.950 379.950 430.050 382.050 ;
        RECT 430.950 379.950 433.050 382.050 ;
        RECT 433.950 381.450 436.050 382.050 ;
        RECT 437.400 381.450 438.450 406.950 ;
        RECT 439.950 400.950 442.050 403.050 ;
        RECT 440.400 382.050 441.450 400.950 ;
        RECT 446.400 391.050 447.450 436.950 ;
        RECT 449.400 418.050 450.450 455.400 ;
        RECT 448.950 415.950 451.050 418.050 ;
        RECT 448.950 406.950 451.050 409.050 ;
        RECT 449.400 391.050 450.450 406.950 ;
        RECT 445.950 388.950 448.050 391.050 ;
        RECT 448.950 388.950 451.050 391.050 ;
        RECT 449.400 388.050 450.450 388.950 ;
        RECT 448.950 385.950 451.050 388.050 ;
        RECT 445.950 383.250 448.050 384.150 ;
        RECT 448.950 383.850 451.050 384.750 ;
        RECT 433.950 380.400 438.450 381.450 ;
        RECT 433.950 379.950 436.050 380.400 ;
        RECT 439.950 379.950 442.050 382.050 ;
        RECT 445.950 379.950 448.050 382.050 ;
        RECT 452.400 381.450 453.450 481.950 ;
        RECT 455.400 481.050 456.450 488.400 ;
        RECT 458.400 484.050 459.450 517.950 ;
        RECT 463.950 508.950 466.050 511.050 ;
        RECT 460.950 490.950 463.050 493.050 ;
        RECT 457.950 481.950 460.050 484.050 ;
        RECT 454.950 478.950 457.050 481.050 ;
        RECT 454.950 466.950 457.050 469.050 ;
        RECT 455.400 424.050 456.450 466.950 ;
        RECT 461.400 457.050 462.450 490.950 ;
        RECT 464.400 478.050 465.450 508.950 ;
        RECT 470.400 502.050 471.450 550.950 ;
        RECT 473.400 511.050 474.450 607.950 ;
        RECT 476.400 604.050 477.450 694.950 ;
        RECT 482.400 685.050 483.450 700.950 ;
        RECT 488.400 697.050 489.450 700.950 ;
        RECT 487.950 694.950 490.050 697.050 ;
        RECT 503.400 694.050 504.450 703.950 ;
        RECT 505.950 702.450 508.050 703.050 ;
        RECT 509.400 702.450 510.450 715.950 ;
        RECT 511.950 706.950 514.050 709.050 ;
        RECT 512.400 703.050 513.450 706.950 ;
        RECT 505.950 701.400 510.450 702.450 ;
        RECT 505.950 700.950 508.050 701.400 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 502.950 691.950 505.050 694.050 ;
        RECT 493.950 688.950 496.050 691.050 ;
        RECT 481.950 682.950 484.050 685.050 ;
        RECT 482.400 682.050 483.450 682.950 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 481.950 673.950 484.050 676.050 ;
        RECT 481.950 671.850 484.050 672.750 ;
        RECT 484.950 671.250 487.050 672.150 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 485.400 631.050 486.450 667.950 ;
        RECT 488.400 631.050 489.450 679.950 ;
        RECT 481.950 630.450 484.050 631.050 ;
        RECT 479.400 629.400 484.050 630.450 ;
        RECT 479.400 616.050 480.450 629.400 ;
        RECT 481.950 628.950 484.050 629.400 ;
        RECT 484.950 628.950 487.050 631.050 ;
        RECT 487.950 628.950 490.050 631.050 ;
        RECT 491.250 629.250 493.050 630.150 ;
        RECT 481.950 626.850 484.050 627.750 ;
        RECT 484.950 626.250 487.050 627.150 ;
        RECT 487.950 626.850 489.750 627.750 ;
        RECT 490.950 625.950 493.050 628.050 ;
        RECT 484.950 622.950 487.050 625.050 ;
        RECT 481.950 616.950 484.050 619.050 ;
        RECT 484.950 616.950 487.050 619.050 ;
        RECT 478.950 613.950 481.050 616.050 ;
        RECT 482.400 612.450 483.450 616.950 ;
        RECT 479.400 611.400 483.450 612.450 ;
        RECT 475.950 601.950 478.050 604.050 ;
        RECT 479.400 598.050 480.450 611.400 ;
        RECT 481.950 607.950 484.050 610.050 ;
        RECT 475.950 596.250 477.750 597.150 ;
        RECT 478.950 595.950 481.050 598.050 ;
        RECT 482.400 595.050 483.450 607.950 ;
        RECT 485.400 598.050 486.450 616.950 ;
        RECT 490.950 613.950 493.050 616.050 ;
        RECT 487.950 598.950 490.050 601.050 ;
        RECT 491.400 600.450 492.450 613.950 ;
        RECT 494.400 607.050 495.450 688.950 ;
        RECT 496.950 673.950 499.050 676.050 ;
        RECT 497.400 673.050 498.450 673.950 ;
        RECT 496.950 670.950 499.050 673.050 ;
        RECT 500.250 671.250 501.750 672.150 ;
        RECT 502.950 670.950 505.050 673.050 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 506.400 670.050 507.450 670.950 ;
        RECT 496.950 668.850 498.750 669.750 ;
        RECT 499.950 667.950 502.050 670.050 ;
        RECT 503.250 668.850 504.750 669.750 ;
        RECT 505.950 667.950 508.050 670.050 ;
        RECT 500.400 667.050 501.450 667.950 ;
        RECT 499.950 664.950 502.050 667.050 ;
        RECT 505.950 665.850 508.050 666.750 ;
        RECT 499.950 658.950 502.050 661.050 ;
        RECT 496.950 640.950 499.050 643.050 ;
        RECT 497.400 615.450 498.450 640.950 ;
        RECT 500.400 625.050 501.450 658.950 ;
        RECT 511.950 632.250 514.050 633.150 ;
        RECT 502.950 629.250 504.750 630.150 ;
        RECT 505.950 628.950 508.050 631.050 ;
        RECT 509.250 629.250 510.750 630.150 ;
        RECT 511.950 628.950 514.050 631.050 ;
        RECT 502.950 625.950 505.050 628.050 ;
        RECT 506.250 626.850 507.750 627.750 ;
        RECT 508.950 625.950 511.050 628.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 505.950 622.950 508.050 625.050 ;
        RECT 497.400 614.400 501.450 615.450 ;
        RECT 500.400 613.050 501.450 614.400 ;
        RECT 496.950 610.950 499.050 613.050 ;
        RECT 499.950 610.950 502.050 613.050 ;
        RECT 493.950 604.950 496.050 607.050 ;
        RECT 497.400 604.050 498.450 610.950 ;
        RECT 499.950 607.950 502.050 610.050 ;
        RECT 500.400 604.050 501.450 607.950 ;
        RECT 502.950 604.950 505.050 607.050 ;
        RECT 496.950 601.950 499.050 604.050 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 491.400 599.400 495.450 600.450 ;
        RECT 484.950 595.950 487.050 598.050 ;
        RECT 488.400 595.050 489.450 598.950 ;
        RECT 490.950 595.950 493.050 598.050 ;
        RECT 475.950 592.950 478.050 595.050 ;
        RECT 479.250 593.850 480.750 594.750 ;
        RECT 481.950 592.950 484.050 595.050 ;
        RECT 485.250 593.850 487.050 594.750 ;
        RECT 487.950 592.950 490.050 595.050 ;
        RECT 476.400 538.050 477.450 592.950 ;
        RECT 481.950 590.850 484.050 591.750 ;
        RECT 484.950 580.950 487.050 583.050 ;
        RECT 485.400 577.050 486.450 580.950 ;
        RECT 484.950 574.950 487.050 577.050 ;
        RECT 487.950 574.950 490.050 577.050 ;
        RECT 478.950 562.950 481.050 565.050 ;
        RECT 479.400 562.050 480.450 562.950 ;
        RECT 478.950 559.950 481.050 562.050 ;
        RECT 482.250 560.250 483.750 561.150 ;
        RECT 484.950 559.950 487.050 562.050 ;
        RECT 478.950 557.850 480.750 558.750 ;
        RECT 481.950 556.950 484.050 559.050 ;
        RECT 485.250 557.850 487.050 558.750 ;
        RECT 488.400 547.050 489.450 574.950 ;
        RECT 491.400 549.450 492.450 595.950 ;
        RECT 494.400 574.050 495.450 599.400 ;
        RECT 496.950 599.250 499.050 600.150 ;
        RECT 499.950 599.850 502.050 600.750 ;
        RECT 496.950 595.950 499.050 598.050 ;
        RECT 493.950 571.950 496.050 574.050 ;
        RECT 499.950 571.950 502.050 574.050 ;
        RECT 493.950 562.950 496.050 565.050 ;
        RECT 494.400 553.050 495.450 562.950 ;
        RECT 496.950 559.950 499.050 562.050 ;
        RECT 497.400 559.050 498.450 559.950 ;
        RECT 500.400 559.050 501.450 571.950 ;
        RECT 503.400 571.050 504.450 604.950 ;
        RECT 506.400 577.050 507.450 622.950 ;
        RECT 509.400 616.050 510.450 625.950 ;
        RECT 515.400 616.050 516.450 718.950 ;
        RECT 518.400 715.050 519.450 739.950 ;
        RECT 517.950 712.950 520.050 715.050 ;
        RECT 520.950 712.950 523.050 715.050 ;
        RECT 521.400 706.050 522.450 712.950 ;
        RECT 520.950 703.950 523.050 706.050 ;
        RECT 521.400 703.050 522.450 703.950 ;
        RECT 524.400 703.050 525.450 745.950 ;
        RECT 526.950 743.850 528.750 744.750 ;
        RECT 529.950 744.450 532.050 745.050 ;
        RECT 533.400 744.450 534.450 766.950 ;
        RECT 529.950 743.400 534.450 744.450 ;
        RECT 529.950 742.950 532.050 743.400 ;
        RECT 529.950 740.850 532.050 741.750 ;
        RECT 526.950 736.950 529.050 739.050 ;
        RECT 527.400 703.050 528.450 736.950 ;
        RECT 533.400 730.050 534.450 743.400 ;
        RECT 535.950 743.250 538.050 744.150 ;
        RECT 535.950 739.950 538.050 742.050 ;
        RECT 536.400 739.050 537.450 739.950 ;
        RECT 535.950 736.950 538.050 739.050 ;
        RECT 542.400 736.050 543.450 835.950 ;
        RECT 560.400 832.050 561.450 845.400 ;
        RECT 562.950 844.950 565.050 845.400 ;
        RECT 577.950 844.950 580.050 847.050 ;
        RECT 589.950 845.250 591.750 846.150 ;
        RECT 592.950 844.950 595.050 847.050 ;
        RECT 596.250 845.250 597.750 846.150 ;
        RECT 598.950 844.950 601.050 847.050 ;
        RECT 613.950 844.950 616.050 847.050 ;
        RECT 562.950 842.850 565.050 843.750 ;
        RECT 565.950 842.250 568.050 843.150 ;
        RECT 574.950 842.250 577.050 843.150 ;
        RECT 577.950 842.850 580.050 843.750 ;
        RECT 589.950 841.950 592.050 844.050 ;
        RECT 593.250 842.850 594.750 843.750 ;
        RECT 595.950 841.950 598.050 844.050 ;
        RECT 590.400 841.050 591.450 841.950 ;
        RECT 565.950 838.950 568.050 841.050 ;
        RECT 574.950 838.950 577.050 841.050 ;
        RECT 589.950 840.450 592.050 841.050 ;
        RECT 589.950 839.400 594.450 840.450 ;
        RECT 589.950 838.950 592.050 839.400 ;
        RECT 566.400 838.050 567.450 838.950 ;
        RECT 565.950 835.950 568.050 838.050 ;
        RECT 556.950 829.950 559.050 832.050 ;
        RECT 559.950 829.950 562.050 832.050 ;
        RECT 557.400 814.050 558.450 829.950 ;
        RECT 560.400 817.050 561.450 829.950 ;
        RECT 568.950 826.950 571.050 829.050 ;
        RECT 562.950 823.950 565.050 826.050 ;
        RECT 565.950 823.950 568.050 826.050 ;
        RECT 559.950 814.950 562.050 817.050 ;
        RECT 550.950 812.250 552.750 813.150 ;
        RECT 553.950 811.950 556.050 814.050 ;
        RECT 556.950 811.950 559.050 814.050 ;
        RECT 559.950 811.950 562.050 814.050 ;
        RECT 550.950 808.950 553.050 811.050 ;
        RECT 554.250 809.850 555.750 810.750 ;
        RECT 556.950 808.950 559.050 811.050 ;
        RECT 560.250 809.850 562.050 810.750 ;
        RECT 556.950 806.850 559.050 807.750 ;
        RECT 544.950 778.950 547.050 781.050 ;
        RECT 545.400 778.050 546.450 778.950 ;
        RECT 544.950 775.950 547.050 778.050 ;
        RECT 550.950 777.450 553.050 778.050 ;
        RECT 553.950 777.450 556.050 778.050 ;
        RECT 548.250 776.250 549.750 777.150 ;
        RECT 550.950 776.400 556.050 777.450 ;
        RECT 550.950 775.950 553.050 776.400 ;
        RECT 553.950 775.950 556.050 776.400 ;
        RECT 544.950 773.850 546.750 774.750 ;
        RECT 547.950 772.950 550.050 775.050 ;
        RECT 551.250 773.850 553.050 774.750 ;
        RECT 548.400 772.050 549.450 772.950 ;
        RECT 547.950 769.950 550.050 772.050 ;
        RECT 554.400 748.050 555.450 775.950 ;
        RECT 556.950 763.950 559.050 766.050 ;
        RECT 553.950 745.950 556.050 748.050 ;
        RECT 557.400 745.050 558.450 763.950 ;
        RECT 550.950 744.450 553.050 745.050 ;
        RECT 548.400 743.400 553.050 744.450 ;
        RECT 554.250 743.850 555.750 744.750 ;
        RECT 535.950 733.950 538.050 736.050 ;
        RECT 541.950 733.950 544.050 736.050 ;
        RECT 532.950 727.950 535.050 730.050 ;
        RECT 517.950 701.250 519.750 702.150 ;
        RECT 520.950 700.950 523.050 703.050 ;
        RECT 523.950 700.950 526.050 703.050 ;
        RECT 526.950 702.450 529.050 703.050 ;
        RECT 526.950 701.400 531.450 702.450 ;
        RECT 526.950 700.950 529.050 701.400 ;
        RECT 530.400 700.050 531.450 701.400 ;
        RECT 517.950 697.950 520.050 700.050 ;
        RECT 521.250 698.850 523.050 699.750 ;
        RECT 523.950 698.250 526.050 699.150 ;
        RECT 526.950 698.850 529.050 699.750 ;
        RECT 529.950 697.950 532.050 700.050 ;
        RECT 518.400 697.050 519.450 697.950 ;
        RECT 517.950 694.950 520.050 697.050 ;
        RECT 523.950 694.950 526.050 697.050 ;
        RECT 517.950 676.950 520.050 679.050 ;
        RECT 520.950 676.950 523.050 679.050 ;
        RECT 518.400 631.050 519.450 676.950 ;
        RECT 521.400 673.050 522.450 676.950 ;
        RECT 526.950 673.950 529.050 676.050 ;
        RECT 520.950 670.950 523.050 673.050 ;
        RECT 520.950 668.850 523.050 669.750 ;
        RECT 523.950 668.250 526.050 669.150 ;
        RECT 523.950 666.450 526.050 667.050 ;
        RECT 527.400 666.450 528.450 673.950 ;
        RECT 529.950 670.950 532.050 673.050 ;
        RECT 529.950 668.850 532.050 669.750 ;
        RECT 532.950 667.950 535.050 670.050 ;
        RECT 523.950 665.400 528.450 666.450 ;
        RECT 523.950 664.950 526.050 665.400 ;
        RECT 527.400 661.050 528.450 665.400 ;
        RECT 526.950 658.950 529.050 661.050 ;
        RECT 517.950 628.950 520.050 631.050 ;
        RECT 523.950 628.950 526.050 631.050 ;
        RECT 529.950 628.950 532.050 631.050 ;
        RECT 520.950 622.950 523.050 625.050 ;
        RECT 508.950 613.950 511.050 616.050 ;
        RECT 514.950 613.950 517.050 616.050 ;
        RECT 508.950 610.950 511.050 613.050 ;
        RECT 505.950 574.950 508.050 577.050 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 509.400 568.050 510.450 610.950 ;
        RECT 521.400 601.050 522.450 622.950 ;
        RECT 524.400 619.050 525.450 628.950 ;
        RECT 526.950 626.250 529.050 627.150 ;
        RECT 529.950 626.850 532.050 627.750 ;
        RECT 533.400 625.050 534.450 667.950 ;
        RECT 536.400 637.050 537.450 733.950 ;
        RECT 548.400 712.050 549.450 743.400 ;
        RECT 550.950 742.950 553.050 743.400 ;
        RECT 556.950 742.950 559.050 745.050 ;
        RECT 550.950 740.850 553.050 741.750 ;
        RECT 556.950 740.850 559.050 741.750 ;
        RECT 556.950 730.950 559.050 733.050 ;
        RECT 550.950 727.950 553.050 730.050 ;
        RECT 547.950 709.950 550.050 712.050 ;
        RECT 538.950 706.950 541.050 709.050 ;
        RECT 544.950 707.250 547.050 708.150 ;
        RECT 539.400 706.050 540.450 706.950 ;
        RECT 538.950 703.950 541.050 706.050 ;
        RECT 542.250 704.250 543.750 705.150 ;
        RECT 544.950 703.950 547.050 706.050 ;
        RECT 548.250 704.250 550.050 705.150 ;
        RECT 545.400 703.050 546.450 703.950 ;
        RECT 538.950 701.850 540.750 702.750 ;
        RECT 541.950 700.950 544.050 703.050 ;
        RECT 544.950 700.950 547.050 703.050 ;
        RECT 547.950 700.950 550.050 703.050 ;
        RECT 542.400 700.050 543.450 700.950 ;
        RECT 541.950 697.950 544.050 700.050 ;
        RECT 545.400 697.050 546.450 700.950 ;
        RECT 544.950 694.950 547.050 697.050 ;
        RECT 547.950 688.950 550.050 691.050 ;
        RECT 548.400 679.050 549.450 688.950 ;
        RECT 547.950 676.950 550.050 679.050 ;
        RECT 538.950 670.950 541.050 673.050 ;
        RECT 544.950 670.950 547.050 673.050 ;
        RECT 539.400 667.050 540.450 670.950 ;
        RECT 545.400 670.050 546.450 670.950 ;
        RECT 541.950 668.250 543.750 669.150 ;
        RECT 544.950 667.950 547.050 670.050 ;
        RECT 548.250 668.250 550.050 669.150 ;
        RECT 538.950 664.950 541.050 667.050 ;
        RECT 541.950 664.950 544.050 667.050 ;
        RECT 545.250 665.850 546.750 666.750 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 542.400 661.050 543.450 664.950 ;
        RECT 544.950 661.950 547.050 664.050 ;
        RECT 541.950 658.950 544.050 661.050 ;
        RECT 545.400 658.050 546.450 661.950 ;
        RECT 544.950 655.950 547.050 658.050 ;
        RECT 538.950 637.950 541.050 640.050 ;
        RECT 535.950 634.950 538.050 637.050 ;
        RECT 526.950 622.950 529.050 625.050 ;
        RECT 532.950 622.950 535.050 625.050 ;
        RECT 523.950 616.950 526.050 619.050 ;
        RECT 523.950 613.950 526.050 616.050 ;
        RECT 514.950 598.950 517.050 601.050 ;
        RECT 518.250 599.250 519.750 600.150 ;
        RECT 520.950 598.950 523.050 601.050 ;
        RECT 511.950 595.950 514.050 598.050 ;
        RECT 515.250 596.850 516.750 597.750 ;
        RECT 517.950 595.950 520.050 598.050 ;
        RECT 521.250 596.850 523.050 597.750 ;
        RECT 511.950 593.850 514.050 594.750 ;
        RECT 518.400 592.050 519.450 595.950 ;
        RECT 524.400 594.450 525.450 613.950 ;
        RECT 532.950 607.950 535.050 610.050 ;
        RECT 533.400 598.050 534.450 607.950 ;
        RECT 536.400 607.050 537.450 634.950 ;
        RECT 539.400 630.450 540.450 637.950 ;
        RECT 544.950 635.250 547.050 636.150 ;
        RECT 551.400 634.050 552.450 727.950 ;
        RECT 553.950 721.950 556.050 724.050 ;
        RECT 554.400 673.050 555.450 721.950 ;
        RECT 557.400 699.450 558.450 730.950 ;
        RECT 563.400 706.050 564.450 823.950 ;
        RECT 566.400 808.050 567.450 823.950 ;
        RECT 569.400 814.050 570.450 826.950 ;
        RECT 575.400 820.050 576.450 838.950 ;
        RECT 593.400 829.050 594.450 839.400 ;
        RECT 596.400 835.050 597.450 841.950 ;
        RECT 599.400 841.050 600.450 844.950 ;
        RECT 610.950 842.250 613.050 843.150 ;
        RECT 613.950 842.850 616.050 843.750 ;
        RECT 622.950 843.450 625.050 844.050 ;
        RECT 620.400 842.400 625.050 843.450 ;
        RECT 598.950 838.950 601.050 841.050 ;
        RECT 610.950 838.950 613.050 841.050 ;
        RECT 595.950 832.950 598.050 835.050 ;
        RECT 595.950 829.950 598.050 832.050 ;
        RECT 592.950 826.950 595.050 829.050 ;
        RECT 596.400 826.050 597.450 829.950 ;
        RECT 577.950 823.950 580.050 826.050 ;
        RECT 592.950 823.950 595.050 826.050 ;
        RECT 595.950 823.950 598.050 826.050 ;
        RECT 578.400 820.050 579.450 823.950 ;
        RECT 586.950 820.950 589.050 823.050 ;
        RECT 574.950 817.950 577.050 820.050 ;
        RECT 577.950 817.950 580.050 820.050 ;
        RECT 571.950 814.950 574.050 817.050 ;
        RECT 575.250 815.250 577.050 816.150 ;
        RECT 577.950 815.850 580.050 816.750 ;
        RECT 580.950 815.250 583.050 816.150 ;
        RECT 583.950 814.950 586.050 817.050 ;
        RECT 568.950 811.950 571.050 814.050 ;
        RECT 571.950 812.850 573.750 813.750 ;
        RECT 574.950 811.950 577.050 814.050 ;
        RECT 577.950 811.950 580.050 814.050 ;
        RECT 580.950 813.450 583.050 814.050 ;
        RECT 584.400 813.450 585.450 814.950 ;
        RECT 580.950 812.400 585.450 813.450 ;
        RECT 580.950 811.950 583.050 812.400 ;
        RECT 565.950 805.950 568.050 808.050 ;
        RECT 565.950 775.950 568.050 778.050 ;
        RECT 571.950 777.450 574.050 778.050 ;
        RECT 569.250 776.250 570.750 777.150 ;
        RECT 571.950 776.400 576.450 777.450 ;
        RECT 571.950 775.950 574.050 776.400 ;
        RECT 565.950 773.850 567.750 774.750 ;
        RECT 568.950 772.950 571.050 775.050 ;
        RECT 572.250 773.850 574.050 774.750 ;
        RECT 575.400 757.050 576.450 776.400 ;
        RECT 574.950 754.950 577.050 757.050 ;
        RECT 575.400 751.050 576.450 754.950 ;
        RECT 565.950 748.950 568.050 751.050 ;
        RECT 574.950 748.950 577.050 751.050 ;
        RECT 578.400 750.450 579.450 811.950 ;
        RECT 581.400 811.050 582.450 811.950 ;
        RECT 580.950 808.950 583.050 811.050 ;
        RECT 583.950 808.950 586.050 811.050 ;
        RECT 587.400 810.450 588.450 820.950 ;
        RECT 593.400 814.050 594.450 823.950 ;
        RECT 589.950 812.250 591.750 813.150 ;
        RECT 592.950 811.950 595.050 814.050 ;
        RECT 596.250 812.250 598.050 813.150 ;
        RECT 589.950 810.450 592.050 811.050 ;
        RECT 587.400 809.400 592.050 810.450 ;
        RECT 593.250 809.850 594.750 810.750 ;
        RECT 589.950 808.950 592.050 809.400 ;
        RECT 595.950 808.950 598.050 811.050 ;
        RECT 584.400 775.050 585.450 808.950 ;
        RECT 596.400 790.050 597.450 808.950 ;
        RECT 599.400 808.050 600.450 838.950 ;
        RECT 620.400 838.050 621.450 842.400 ;
        RECT 622.950 841.950 625.050 842.400 ;
        RECT 622.950 839.850 625.050 840.750 ;
        RECT 619.950 835.950 622.050 838.050 ;
        RECT 626.550 837.600 627.750 849.600 ;
        RECT 634.950 845.250 637.050 846.150 ;
        RECT 640.950 845.250 643.050 846.150 ;
        RECT 634.950 841.950 637.050 844.050 ;
        RECT 640.950 841.950 643.050 844.050 ;
        RECT 635.400 841.050 636.450 841.950 ;
        RECT 634.950 838.950 637.050 841.050 ;
        RECT 647.400 837.600 648.600 854.400 ;
        RECT 817.950 853.950 820.050 856.050 ;
        RECT 868.950 853.950 871.050 856.050 ;
        RECT 724.950 850.950 727.050 853.050 ;
        RECT 745.950 850.950 748.050 853.050 ;
        RECT 667.950 848.250 670.050 849.150 ;
        RECT 725.400 847.050 726.450 850.950 ;
        RECT 733.950 847.950 736.050 850.050 ;
        RECT 739.950 848.250 742.050 849.150 ;
        RECT 667.950 844.950 670.050 847.050 ;
        RECT 671.250 845.250 672.750 846.150 ;
        RECT 673.950 844.950 676.050 847.050 ;
        RECT 677.250 845.250 679.050 846.150 ;
        RECT 682.950 844.950 685.050 847.050 ;
        RECT 688.950 846.450 691.050 847.050 ;
        RECT 686.400 845.400 691.050 846.450 ;
        RECT 670.950 841.950 673.050 844.050 ;
        RECT 674.250 842.850 675.750 843.750 ;
        RECT 625.950 835.500 628.050 837.600 ;
        RECT 646.950 835.500 649.050 837.600 ;
        RECT 679.950 826.950 682.050 829.050 ;
        RECT 664.950 820.950 667.050 823.050 ;
        RECT 646.950 817.950 649.050 820.050 ;
        RECT 655.950 817.950 658.050 820.050 ;
        RECT 613.950 814.950 616.050 817.050 ;
        RECT 619.950 816.450 622.050 817.050 ;
        RECT 622.950 816.450 625.050 817.050 ;
        RECT 617.250 815.250 618.750 816.150 ;
        RECT 619.950 815.400 625.050 816.450 ;
        RECT 619.950 814.950 622.050 815.400 ;
        RECT 622.950 814.950 625.050 815.400 ;
        RECT 610.950 813.450 613.050 814.050 ;
        RECT 608.400 812.400 613.050 813.450 ;
        RECT 614.250 812.850 615.750 813.750 ;
        RECT 598.950 805.950 601.050 808.050 ;
        RECT 608.400 805.050 609.450 812.400 ;
        RECT 610.950 811.950 613.050 812.400 ;
        RECT 616.950 811.950 619.050 814.050 ;
        RECT 620.250 812.850 622.050 813.750 ;
        RECT 623.400 811.050 624.450 814.950 ;
        RECT 631.950 812.250 633.750 813.150 ;
        RECT 634.950 811.950 637.050 814.050 ;
        RECT 638.250 812.250 640.050 813.150 ;
        RECT 610.950 809.850 613.050 810.750 ;
        RECT 622.950 808.950 625.050 811.050 ;
        RECT 631.950 808.950 634.050 811.050 ;
        RECT 635.250 809.850 636.750 810.750 ;
        RECT 637.950 808.950 640.050 811.050 ;
        RECT 647.400 810.450 648.450 817.950 ;
        RECT 649.950 812.250 651.750 813.150 ;
        RECT 652.950 811.950 655.050 814.050 ;
        RECT 656.400 811.050 657.450 817.950 ;
        RECT 658.950 813.450 661.050 814.050 ;
        RECT 658.950 812.400 663.450 813.450 ;
        RECT 658.950 811.950 661.050 812.400 ;
        RECT 662.400 811.050 663.450 812.400 ;
        RECT 649.950 810.450 652.050 811.050 ;
        RECT 647.400 809.400 652.050 810.450 ;
        RECT 653.250 809.850 654.750 810.750 ;
        RECT 649.950 808.950 652.050 809.400 ;
        RECT 655.950 808.950 658.050 811.050 ;
        RECT 659.250 809.850 661.050 810.750 ;
        RECT 661.950 808.950 664.050 811.050 ;
        RECT 619.950 805.950 622.050 808.050 ;
        RECT 607.950 802.950 610.050 805.050 ;
        RECT 610.950 802.950 613.050 805.050 ;
        RECT 595.950 787.950 598.050 790.050 ;
        RECT 592.950 778.950 595.050 781.050 ;
        RECT 595.950 778.950 598.050 781.050 ;
        RECT 604.950 779.250 607.050 780.150 ;
        RECT 593.400 778.050 594.450 778.950 ;
        RECT 586.950 775.950 589.050 778.050 ;
        RECT 590.250 776.250 591.750 777.150 ;
        RECT 592.950 775.950 595.050 778.050 ;
        RECT 583.950 772.950 586.050 775.050 ;
        RECT 586.950 773.850 588.750 774.750 ;
        RECT 589.950 772.950 592.050 775.050 ;
        RECT 593.250 773.850 595.050 774.750 ;
        RECT 586.950 763.950 589.050 766.050 ;
        RECT 578.400 749.400 582.450 750.450 ;
        RECT 566.400 738.450 567.450 748.950 ;
        RECT 577.950 745.950 580.050 748.050 ;
        RECT 578.400 742.050 579.450 745.950 ;
        RECT 568.950 740.250 570.750 741.150 ;
        RECT 571.950 739.950 574.050 742.050 ;
        RECT 577.950 739.950 580.050 742.050 ;
        RECT 568.950 738.450 571.050 739.050 ;
        RECT 566.400 737.400 571.050 738.450 ;
        RECT 572.250 737.850 573.750 738.750 ;
        RECT 568.950 736.950 571.050 737.400 ;
        RECT 574.950 736.950 577.050 739.050 ;
        RECT 578.250 737.850 580.050 738.750 ;
        RECT 569.400 721.050 570.450 736.950 ;
        RECT 574.950 734.850 577.050 735.750 ;
        RECT 581.400 724.050 582.450 749.400 ;
        RECT 587.400 741.450 588.450 763.950 ;
        RECT 590.400 760.050 591.450 772.950 ;
        RECT 589.950 757.950 592.050 760.050 ;
        RECT 592.950 745.950 595.050 748.050 ;
        RECT 589.950 743.250 592.050 744.150 ;
        RECT 592.950 743.850 595.050 744.750 ;
        RECT 589.950 741.450 592.050 742.050 ;
        RECT 587.400 740.400 592.050 741.450 ;
        RECT 589.950 739.950 592.050 740.400 ;
        RECT 580.950 721.950 583.050 724.050 ;
        RECT 568.950 718.950 571.050 721.050 ;
        RECT 586.950 715.950 589.050 718.050 ;
        RECT 571.950 706.950 574.050 709.050 ;
        RECT 580.950 707.250 583.050 708.150 ;
        RECT 562.950 703.950 565.050 706.050 ;
        RECT 568.950 703.950 571.050 706.050 ;
        RECT 569.400 703.050 570.450 703.950 ;
        RECT 559.950 701.250 561.750 702.150 ;
        RECT 562.950 700.950 565.050 703.050 ;
        RECT 568.950 700.950 571.050 703.050 ;
        RECT 559.950 699.450 562.050 700.050 ;
        RECT 557.400 698.400 562.050 699.450 ;
        RECT 563.250 698.850 565.050 699.750 ;
        RECT 559.950 697.950 562.050 698.400 ;
        RECT 565.950 698.250 568.050 699.150 ;
        RECT 568.950 698.850 571.050 699.750 ;
        RECT 572.400 697.050 573.450 706.950 ;
        RECT 587.400 706.050 588.450 715.950 ;
        RECT 574.950 703.950 577.050 706.050 ;
        RECT 577.950 704.250 579.750 705.150 ;
        RECT 580.950 703.950 583.050 706.050 ;
        RECT 584.250 704.250 585.750 705.150 ;
        RECT 586.950 703.950 589.050 706.050 ;
        RECT 559.950 694.950 562.050 697.050 ;
        RECT 565.950 694.950 568.050 697.050 ;
        RECT 571.950 694.950 574.050 697.050 ;
        RECT 556.950 688.950 559.050 691.050 ;
        RECT 553.950 670.950 556.050 673.050 ;
        RECT 554.400 667.050 555.450 670.950 ;
        RECT 553.950 664.950 556.050 667.050 ;
        RECT 541.950 632.250 543.750 633.150 ;
        RECT 544.950 631.950 547.050 634.050 ;
        RECT 548.250 632.250 549.750 633.150 ;
        RECT 550.950 631.950 553.050 634.050 ;
        RECT 541.950 630.450 544.050 631.050 ;
        RECT 539.400 629.400 544.050 630.450 ;
        RECT 541.950 628.950 544.050 629.400 ;
        RECT 545.400 628.050 546.450 631.950 ;
        RECT 547.950 628.950 550.050 631.050 ;
        RECT 551.250 629.850 553.050 630.750 ;
        RECT 538.950 625.950 541.050 628.050 ;
        RECT 544.950 625.950 547.050 628.050 ;
        RECT 535.950 604.950 538.050 607.050 ;
        RECT 529.950 596.250 531.750 597.150 ;
        RECT 532.950 595.950 535.050 598.050 ;
        RECT 536.250 596.250 538.050 597.150 ;
        RECT 521.400 593.400 525.450 594.450 ;
        RECT 517.950 589.950 520.050 592.050 ;
        RECT 502.950 565.950 505.050 568.050 ;
        RECT 508.950 565.950 511.050 568.050 ;
        RECT 503.400 562.050 504.450 565.950 ;
        RECT 505.950 562.950 508.050 565.050 ;
        RECT 511.950 563.250 514.050 564.150 ;
        RECT 502.950 559.950 505.050 562.050 ;
        RECT 496.950 556.950 499.050 559.050 ;
        RECT 499.950 556.950 502.050 559.050 ;
        RECT 496.950 554.850 499.050 555.750 ;
        RECT 499.950 554.250 502.050 555.150 ;
        RECT 493.950 550.950 496.050 553.050 ;
        RECT 499.950 550.950 502.050 553.050 ;
        RECT 491.400 548.400 495.450 549.450 ;
        RECT 487.950 544.950 490.050 547.050 ;
        RECT 490.950 544.950 493.050 547.050 ;
        RECT 475.950 535.950 478.050 538.050 ;
        RECT 478.950 526.950 481.050 529.050 ;
        RECT 475.950 523.950 478.050 526.050 ;
        RECT 479.400 523.050 480.450 526.950 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 485.250 524.250 487.050 525.150 ;
        RECT 487.950 523.950 490.050 526.050 ;
        RECT 475.950 521.850 477.750 522.750 ;
        RECT 478.950 520.950 481.050 523.050 ;
        RECT 482.250 521.850 483.750 522.750 ;
        RECT 484.950 520.950 487.050 523.050 ;
        RECT 488.400 520.050 489.450 523.950 ;
        RECT 478.950 518.850 481.050 519.750 ;
        RECT 487.950 517.950 490.050 520.050 ;
        RECT 491.400 516.450 492.450 544.950 ;
        RECT 488.400 515.400 492.450 516.450 ;
        RECT 472.950 508.950 475.050 511.050 ;
        RECT 466.950 499.950 469.050 502.050 ;
        RECT 469.950 499.950 472.050 502.050 ;
        RECT 478.950 499.950 481.050 502.050 ;
        RECT 484.950 499.950 487.050 502.050 ;
        RECT 467.400 490.050 468.450 499.950 ;
        RECT 472.950 496.950 475.050 499.050 ;
        RECT 473.400 492.450 474.450 496.950 ;
        RECT 473.400 491.400 477.450 492.450 ;
        RECT 466.950 487.950 469.050 490.050 ;
        RECT 470.250 488.250 471.750 489.150 ;
        RECT 472.950 487.950 475.050 490.050 ;
        RECT 466.950 485.850 468.750 486.750 ;
        RECT 469.950 484.950 472.050 487.050 ;
        RECT 473.250 485.850 475.050 486.750 ;
        RECT 463.950 475.950 466.050 478.050 ;
        RECT 470.400 475.050 471.450 484.950 ;
        RECT 463.950 472.950 466.050 475.050 ;
        RECT 469.950 472.950 472.050 475.050 ;
        RECT 460.950 454.950 463.050 457.050 ;
        RECT 464.400 454.050 465.450 472.950 ;
        RECT 472.950 460.950 475.050 463.050 ;
        RECT 469.950 454.950 472.050 457.050 ;
        RECT 460.950 452.250 462.750 453.150 ;
        RECT 463.950 451.950 466.050 454.050 ;
        RECT 467.250 452.250 469.050 453.150 ;
        RECT 460.950 448.950 463.050 451.050 ;
        RECT 464.250 449.850 465.750 450.750 ;
        RECT 466.950 448.950 469.050 451.050 ;
        RECT 467.400 448.050 468.450 448.950 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 470.400 439.050 471.450 454.950 ;
        RECT 473.400 448.050 474.450 460.950 ;
        RECT 472.950 445.950 475.050 448.050 ;
        RECT 469.950 436.950 472.050 439.050 ;
        RECT 469.950 430.950 472.050 433.050 ;
        RECT 454.950 421.950 457.050 424.050 ;
        RECT 466.950 421.950 469.050 424.050 ;
        RECT 460.950 419.250 463.050 420.150 ;
        RECT 467.400 418.050 468.450 421.950 ;
        RECT 454.950 415.950 457.050 418.050 ;
        RECT 458.250 416.250 459.750 417.150 ;
        RECT 460.950 415.950 463.050 418.050 ;
        RECT 464.250 416.250 466.050 417.150 ;
        RECT 466.950 415.950 469.050 418.050 ;
        RECT 454.950 413.850 456.750 414.750 ;
        RECT 457.950 412.950 460.050 415.050 ;
        RECT 463.950 412.950 466.050 415.050 ;
        RECT 454.950 409.950 457.050 412.050 ;
        RECT 455.400 382.050 456.450 409.950 ;
        RECT 458.400 403.050 459.450 412.950 ;
        RECT 464.400 412.050 465.450 412.950 ;
        RECT 470.400 412.050 471.450 430.950 ;
        RECT 476.400 421.050 477.450 491.400 ;
        RECT 479.400 475.050 480.450 499.950 ;
        RECT 485.400 490.050 486.450 499.950 ;
        RECT 488.400 490.050 489.450 515.400 ;
        RECT 494.400 502.050 495.450 548.400 ;
        RECT 499.950 524.250 501.750 525.150 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 506.400 525.450 507.450 562.950 ;
        RECT 508.950 560.250 510.750 561.150 ;
        RECT 511.950 559.950 514.050 562.050 ;
        RECT 515.250 560.250 516.750 561.150 ;
        RECT 517.950 559.950 520.050 562.050 ;
        RECT 514.950 556.950 517.050 559.050 ;
        RECT 518.250 557.850 520.050 558.750 ;
        RECT 508.950 529.950 511.050 532.050 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 509.400 529.050 510.450 529.950 ;
        RECT 508.950 526.950 511.050 529.050 ;
        RECT 508.950 525.450 511.050 526.050 ;
        RECT 506.400 524.400 511.050 525.450 ;
        RECT 508.950 523.950 511.050 524.400 ;
        RECT 499.950 520.950 502.050 523.050 ;
        RECT 503.250 521.850 504.750 522.750 ;
        RECT 505.950 520.950 508.050 523.050 ;
        RECT 509.250 521.850 511.050 522.750 ;
        RECT 512.400 520.050 513.450 529.950 ;
        RECT 514.950 526.950 517.050 529.050 ;
        RECT 521.400 528.450 522.450 593.400 ;
        RECT 529.950 592.950 532.050 595.050 ;
        RECT 533.250 593.850 534.750 594.750 ;
        RECT 535.950 592.950 538.050 595.050 ;
        RECT 523.950 586.950 526.050 589.050 ;
        RECT 524.400 532.050 525.450 586.950 ;
        RECT 526.950 571.950 529.050 574.050 ;
        RECT 527.400 532.050 528.450 571.950 ;
        RECT 532.950 562.950 535.050 565.050 ;
        RECT 533.400 559.050 534.450 562.950 ;
        RECT 535.950 559.950 538.050 562.050 ;
        RECT 532.950 556.950 535.050 559.050 ;
        RECT 529.950 554.250 532.050 555.150 ;
        RECT 532.950 554.850 535.050 555.750 ;
        RECT 529.950 550.950 532.050 553.050 ;
        RECT 532.950 550.950 535.050 553.050 ;
        RECT 530.400 538.050 531.450 550.950 ;
        RECT 529.950 535.950 532.050 538.050 ;
        RECT 523.950 529.950 526.050 532.050 ;
        RECT 526.950 529.950 529.050 532.050 ;
        RECT 530.400 529.050 531.450 535.950 ;
        RECT 533.400 535.050 534.450 550.950 ;
        RECT 532.950 532.950 535.050 535.050 ;
        RECT 523.950 528.450 526.050 529.050 ;
        RECT 521.400 527.400 526.050 528.450 ;
        RECT 523.950 526.950 526.050 527.400 ;
        RECT 527.250 527.250 528.750 528.150 ;
        RECT 529.950 526.950 532.050 529.050 ;
        RECT 499.950 517.950 502.050 520.050 ;
        RECT 502.950 517.950 505.050 520.050 ;
        RECT 505.950 518.850 508.050 519.750 ;
        RECT 511.950 517.950 514.050 520.050 ;
        RECT 493.950 499.950 496.050 502.050 ;
        RECT 496.950 496.950 499.050 499.050 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 494.400 490.050 495.450 490.950 ;
        RECT 484.950 487.950 487.050 490.050 ;
        RECT 487.950 487.950 490.050 490.050 ;
        RECT 491.250 488.250 492.750 489.150 ;
        RECT 493.950 487.950 496.050 490.050 ;
        RECT 487.950 485.850 489.750 486.750 ;
        RECT 490.950 484.950 493.050 487.050 ;
        RECT 494.250 485.850 496.050 486.750 ;
        RECT 478.950 472.950 481.050 475.050 ;
        RECT 491.400 472.050 492.450 484.950 ;
        RECT 490.950 469.950 493.050 472.050 ;
        RECT 481.950 466.950 484.050 469.050 ;
        RECT 482.400 457.050 483.450 466.950 ;
        RECT 490.950 460.950 493.050 463.050 ;
        RECT 487.950 457.950 490.050 460.050 ;
        RECT 481.950 454.950 484.050 457.050 ;
        RECT 481.950 452.850 484.050 453.750 ;
        RECT 484.950 452.250 487.050 453.150 ;
        RECT 484.950 450.450 487.050 451.050 ;
        RECT 488.400 450.450 489.450 457.950 ;
        RECT 491.400 457.050 492.450 460.950 ;
        RECT 490.950 454.950 493.050 457.050 ;
        RECT 490.950 452.850 493.050 453.750 ;
        RECT 484.950 449.400 489.450 450.450 ;
        RECT 484.950 448.950 487.050 449.400 ;
        RECT 493.950 439.950 496.050 442.050 ;
        RECT 494.400 427.050 495.450 439.950 ;
        RECT 493.950 424.950 496.050 427.050 ;
        RECT 475.950 418.950 478.050 421.050 ;
        RECT 478.950 418.950 481.050 421.050 ;
        RECT 484.950 418.950 487.050 421.050 ;
        RECT 487.950 418.950 490.050 421.050 ;
        RECT 479.400 418.050 480.450 418.950 ;
        RECT 472.950 415.950 475.050 418.050 ;
        RECT 476.250 416.250 477.750 417.150 ;
        RECT 478.950 415.950 481.050 418.050 ;
        RECT 481.950 415.950 484.050 418.050 ;
        RECT 472.950 413.850 474.750 414.750 ;
        RECT 475.950 412.950 478.050 415.050 ;
        RECT 479.250 413.850 481.050 414.750 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 469.950 409.950 472.050 412.050 ;
        RECT 457.950 400.950 460.050 403.050 ;
        RECT 476.400 400.050 477.450 412.950 ;
        RECT 475.950 397.950 478.050 400.050 ;
        RECT 478.950 388.950 481.050 391.050 ;
        RECT 458.400 386.400 468.450 387.450 ;
        RECT 458.400 385.050 459.450 386.400 ;
        RECT 467.400 385.050 468.450 386.400 ;
        RECT 475.950 385.950 478.050 388.050 ;
        RECT 457.950 382.950 460.050 385.050 ;
        RECT 461.250 383.250 462.750 384.150 ;
        RECT 463.950 382.950 466.050 385.050 ;
        RECT 466.950 382.950 469.050 385.050 ;
        RECT 472.950 382.950 475.050 385.050 ;
        RECT 449.400 380.400 453.450 381.450 ;
        RECT 421.950 376.950 424.050 379.050 ;
        RECT 407.400 344.400 411.450 345.450 ;
        RECT 410.400 343.050 411.450 344.400 ;
        RECT 415.950 344.250 418.050 345.150 ;
        RECT 418.950 343.950 421.050 346.050 ;
        RECT 394.950 341.250 397.050 342.150 ;
        RECT 406.950 341.250 408.750 342.150 ;
        RECT 409.950 340.950 412.050 343.050 ;
        RECT 413.250 341.250 414.750 342.150 ;
        RECT 415.950 340.950 418.050 343.050 ;
        RECT 394.950 337.950 397.050 340.050 ;
        RECT 406.950 337.950 409.050 340.050 ;
        RECT 410.250 338.850 411.750 339.750 ;
        RECT 412.950 337.950 415.050 340.050 ;
        RECT 415.950 337.950 418.050 340.050 ;
        RECT 407.400 337.050 408.450 337.950 ;
        RECT 392.400 335.400 396.450 336.450 ;
        RECT 388.950 331.950 391.050 334.050 ;
        RECT 376.950 325.950 379.050 328.050 ;
        RECT 382.950 325.950 385.050 328.050 ;
        RECT 373.950 317.400 376.050 319.500 ;
        RECT 376.950 317.400 379.050 319.500 ;
        RECT 379.950 317.400 382.050 319.500 ;
        RECT 384.750 317.400 386.850 319.500 ;
        RECT 388.950 317.400 391.050 319.500 ;
        RECT 370.950 307.950 373.050 310.050 ;
        RECT 374.550 303.750 375.750 317.400 ;
        RECT 373.950 301.650 376.050 303.750 ;
        RECT 374.550 297.900 375.750 301.650 ;
        RECT 377.250 300.150 378.450 317.400 ;
        RECT 380.400 303.750 381.600 317.400 ;
        RECT 385.350 311.550 386.550 317.400 ;
        RECT 384.750 309.450 386.850 311.550 ;
        RECT 379.950 301.650 382.050 303.750 ;
        RECT 385.350 300.600 386.550 309.450 ;
        RECT 389.550 308.850 390.750 317.400 ;
        RECT 391.950 316.950 394.050 319.050 ;
        RECT 392.400 316.050 393.450 316.950 ;
        RECT 391.950 313.950 394.050 316.050 ;
        RECT 391.950 311.850 394.050 312.750 ;
        RECT 388.950 306.750 391.050 308.850 ;
        RECT 391.950 307.950 394.050 310.050 ;
        RECT 389.550 300.600 390.750 306.750 ;
        RECT 376.950 298.050 379.050 300.150 ;
        RECT 384.900 298.500 387.000 300.600 ;
        RECT 388.950 298.500 391.050 300.600 ;
        RECT 373.800 295.800 375.900 297.900 ;
        RECT 392.400 295.050 393.450 307.950 ;
        RECT 368.400 293.400 372.450 294.450 ;
        RECT 361.950 283.950 364.050 286.050 ;
        RECT 349.800 281.100 351.900 283.200 ;
        RECT 350.550 277.350 351.750 281.100 ;
        RECT 352.950 278.850 355.050 280.950 ;
        RECT 349.950 275.250 352.050 277.350 ;
        RECT 328.950 233.400 333.450 234.450 ;
        RECT 335.400 248.400 339.450 249.450 ;
        RECT 341.400 263.400 345.450 264.450 ;
        RECT 328.950 232.950 331.050 233.400 ;
        RECT 335.400 208.050 336.450 248.400 ;
        RECT 337.950 244.950 340.050 247.050 ;
        RECT 338.400 238.050 339.450 244.950 ;
        RECT 337.950 235.950 340.050 238.050 ;
        RECT 334.950 205.950 337.050 208.050 ;
        RECT 334.950 203.250 337.050 204.150 ;
        RECT 328.950 199.950 331.050 202.050 ;
        RECT 332.250 200.250 333.750 201.150 ;
        RECT 334.950 199.950 337.050 202.050 ;
        RECT 338.250 200.250 340.050 201.150 ;
        RECT 328.950 197.850 330.750 198.750 ;
        RECT 331.950 196.950 334.050 199.050 ;
        RECT 337.950 196.950 340.050 199.050 ;
        RECT 332.400 196.050 333.450 196.950 ;
        RECT 326.400 194.400 330.450 195.450 ;
        RECT 325.950 166.950 328.050 169.050 ;
        RECT 326.400 166.050 327.450 166.950 ;
        RECT 322.950 164.250 324.750 165.150 ;
        RECT 325.950 163.950 328.050 166.050 ;
        RECT 329.400 163.050 330.450 194.400 ;
        RECT 331.950 193.950 334.050 196.050 ;
        RECT 338.400 172.050 339.450 196.950 ;
        RECT 341.400 190.050 342.450 263.400 ;
        RECT 350.550 261.600 351.750 275.250 ;
        RECT 353.250 261.600 354.450 278.850 ;
        RECT 360.900 278.400 363.000 280.500 ;
        RECT 364.950 278.400 367.050 280.500 ;
        RECT 355.950 275.250 358.050 277.350 ;
        RECT 356.400 261.600 357.600 275.250 ;
        RECT 361.350 269.550 362.550 278.400 ;
        RECT 365.550 272.250 366.750 278.400 ;
        RECT 364.950 270.150 367.050 272.250 ;
        RECT 360.750 267.450 362.850 269.550 ;
        RECT 361.350 261.600 362.550 267.450 ;
        RECT 365.550 261.600 366.750 270.150 ;
        RECT 367.950 266.250 370.050 267.150 ;
        RECT 367.950 262.950 370.050 265.050 ;
        RECT 349.950 259.500 352.050 261.600 ;
        RECT 352.950 259.500 355.050 261.600 ;
        RECT 355.950 259.500 358.050 261.600 ;
        RECT 360.750 259.500 362.850 261.600 ;
        RECT 364.950 259.500 367.050 261.600 ;
        RECT 371.400 256.050 372.450 293.400 ;
        RECT 391.950 292.950 394.050 295.050 ;
        RECT 388.950 289.950 391.050 292.050 ;
        RECT 382.950 283.950 385.050 286.050 ;
        RECT 373.950 280.950 376.050 283.050 ;
        RECT 376.950 280.950 379.050 283.050 ;
        RECT 379.950 280.950 382.050 283.050 ;
        RECT 374.250 262.050 375.450 280.950 ;
        RECT 377.250 276.750 378.450 280.950 ;
        RECT 376.950 274.650 379.050 276.750 ;
        RECT 377.250 262.050 378.450 274.650 ;
        RECT 380.250 262.050 381.450 280.950 ;
        RECT 383.400 265.050 384.450 283.950 ;
        RECT 385.950 272.250 388.050 273.150 ;
        RECT 382.950 262.950 385.050 265.050 ;
        RECT 373.950 259.950 376.050 262.050 ;
        RECT 376.950 259.950 379.050 262.050 ;
        RECT 379.950 259.950 382.050 262.050 ;
        RECT 385.950 259.950 388.050 262.050 ;
        RECT 358.950 253.950 361.050 256.050 ;
        RECT 370.950 253.950 373.050 256.050 ;
        RECT 349.950 241.950 352.050 244.050 ;
        RECT 350.400 241.050 351.450 241.950 ;
        RECT 343.950 238.950 346.050 241.050 ;
        RECT 347.250 239.250 348.750 240.150 ;
        RECT 349.950 238.950 352.050 241.050 ;
        RECT 343.950 236.850 345.750 237.750 ;
        RECT 346.950 235.950 349.050 238.050 ;
        RECT 350.250 236.850 351.750 237.750 ;
        RECT 352.950 235.950 355.050 238.050 ;
        RECT 352.950 233.850 355.050 234.750 ;
        RECT 359.400 231.450 360.450 253.950 ;
        RECT 376.950 250.950 379.050 253.050 ;
        RECT 373.950 244.950 376.050 247.050 ;
        RECT 361.950 238.950 364.050 241.050 ;
        RECT 362.400 234.450 363.450 238.950 ;
        RECT 364.950 236.250 366.750 237.150 ;
        RECT 367.950 235.950 370.050 238.050 ;
        RECT 371.250 236.250 373.050 237.150 ;
        RECT 364.950 234.450 367.050 235.050 ;
        RECT 362.400 233.400 367.050 234.450 ;
        RECT 368.250 233.850 369.750 234.750 ;
        RECT 370.950 234.450 373.050 235.050 ;
        RECT 374.400 234.450 375.450 244.950 ;
        RECT 364.950 232.950 367.050 233.400 ;
        RECT 370.950 233.400 375.450 234.450 ;
        RECT 370.950 232.950 373.050 233.400 ;
        RECT 365.400 232.050 366.450 232.950 ;
        RECT 359.400 230.400 363.450 231.450 ;
        RECT 343.950 214.950 346.050 217.050 ;
        RECT 344.400 202.050 345.450 214.950 ;
        RECT 355.950 203.250 358.050 204.150 ;
        RECT 343.950 199.950 346.050 202.050 ;
        RECT 349.950 201.450 352.050 202.050 ;
        RECT 347.400 200.400 352.050 201.450 ;
        RECT 347.400 193.050 348.450 200.400 ;
        RECT 349.950 199.950 352.050 200.400 ;
        RECT 353.250 200.250 354.750 201.150 ;
        RECT 355.950 199.950 358.050 202.050 ;
        RECT 359.250 200.250 361.050 201.150 ;
        RECT 349.950 197.850 351.750 198.750 ;
        RECT 352.950 196.950 355.050 199.050 ;
        RECT 353.400 196.050 354.450 196.950 ;
        RECT 352.950 193.950 355.050 196.050 ;
        RECT 346.950 190.950 349.050 193.050 ;
        RECT 349.950 190.950 352.050 193.050 ;
        RECT 340.950 187.950 343.050 190.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 331.950 169.950 334.050 172.050 ;
        RECT 337.950 169.950 340.050 172.050 ;
        RECT 332.400 166.050 333.450 169.950 ;
        RECT 347.400 169.050 348.450 178.950 ;
        RECT 346.950 166.950 349.050 169.050 ;
        RECT 347.400 166.050 348.450 166.950 ;
        RECT 350.400 166.050 351.450 190.950 ;
        RECT 353.400 190.050 354.450 193.950 ;
        RECT 352.950 187.950 355.050 190.050 ;
        RECT 356.400 187.050 357.450 199.950 ;
        RECT 358.950 196.950 361.050 199.050 ;
        RECT 355.950 184.950 358.050 187.050 ;
        RECT 355.950 166.950 358.050 169.050 ;
        RECT 331.950 163.950 334.050 166.050 ;
        RECT 340.950 163.950 343.050 166.050 ;
        RECT 343.950 164.250 345.750 165.150 ;
        RECT 346.950 163.950 349.050 166.050 ;
        RECT 349.950 163.950 352.050 166.050 ;
        RECT 352.950 163.950 355.050 166.050 ;
        RECT 322.950 160.950 325.050 163.050 ;
        RECT 326.250 161.850 327.750 162.750 ;
        RECT 328.950 160.950 331.050 163.050 ;
        RECT 332.250 161.850 334.050 162.750 ;
        RECT 328.950 158.850 331.050 159.750 ;
        RECT 334.950 136.950 337.050 139.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 319.950 127.950 322.050 130.050 ;
        RECT 325.950 128.250 328.050 129.150 ;
        RECT 320.400 127.050 321.450 127.950 ;
        RECT 316.950 125.250 318.750 126.150 ;
        RECT 319.950 124.950 322.050 127.050 ;
        RECT 323.250 125.250 324.750 126.150 ;
        RECT 325.950 124.950 328.050 127.050 ;
        RECT 316.950 121.950 319.050 124.050 ;
        RECT 320.250 122.850 321.750 123.750 ;
        RECT 322.950 121.950 325.050 124.050 ;
        RECT 317.400 121.050 318.450 121.950 ;
        RECT 316.950 118.950 319.050 121.050 ;
        RECT 313.950 112.950 316.050 115.050 ;
        RECT 326.400 103.050 327.450 124.950 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 313.950 97.950 316.050 100.050 ;
        RECT 316.950 97.950 319.050 100.050 ;
        RECT 317.400 97.050 318.450 97.950 ;
        RECT 310.950 94.950 313.050 97.050 ;
        RECT 314.250 95.850 315.750 96.750 ;
        RECT 316.950 94.950 319.050 97.050 ;
        RECT 310.950 92.850 313.050 93.750 ;
        RECT 316.950 92.850 319.050 93.750 ;
        RECT 326.400 93.450 327.450 100.950 ;
        RECT 328.950 95.250 331.050 96.150 ;
        RECT 328.950 93.450 331.050 94.050 ;
        RECT 326.400 92.400 331.050 93.450 ;
        RECT 328.950 91.950 331.050 92.400 ;
        RECT 307.950 88.950 310.050 91.050 ;
        RECT 325.950 85.950 328.050 88.050 ;
        RECT 310.950 73.950 313.050 76.050 ;
        RECT 286.950 58.950 289.050 61.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 278.400 51.450 279.450 55.950 ;
        RECT 280.950 53.250 283.050 54.150 ;
        RECT 286.950 53.250 289.050 54.150 ;
        RECT 280.950 51.450 283.050 52.050 ;
        RECT 278.400 50.400 283.050 51.450 ;
        RECT 280.950 49.950 283.050 50.400 ;
        RECT 284.250 50.250 285.750 51.150 ;
        RECT 286.950 49.950 289.050 52.050 ;
        RECT 283.950 46.950 286.050 49.050 ;
        RECT 299.400 48.450 300.450 55.950 ;
        RECT 304.950 52.950 307.050 55.050 ;
        RECT 301.950 50.250 304.050 51.150 ;
        RECT 304.950 50.850 307.050 51.750 ;
        RECT 301.950 48.450 304.050 49.050 ;
        RECT 299.400 47.400 304.050 48.450 ;
        RECT 301.950 46.950 304.050 47.400 ;
        RECT 284.400 28.050 285.450 46.950 ;
        RECT 283.950 25.950 286.050 28.050 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 287.400 22.050 288.450 22.950 ;
        RECT 271.950 20.250 273.750 21.150 ;
        RECT 274.950 19.950 277.050 22.050 ;
        RECT 278.250 20.250 280.050 21.150 ;
        RECT 286.950 19.950 289.050 22.050 ;
        RECT 292.950 19.950 295.050 22.050 ;
        RECT 296.250 20.250 298.050 21.150 ;
        RECT 311.400 19.050 312.450 73.950 ;
        RECT 319.950 56.250 322.050 57.150 ;
        RECT 326.400 55.050 327.450 85.950 ;
        RECT 332.400 57.450 333.450 133.950 ;
        RECT 335.400 123.450 336.450 136.950 ;
        RECT 341.400 133.050 342.450 163.950 ;
        RECT 350.400 163.050 351.450 163.950 ;
        RECT 343.950 160.950 346.050 163.050 ;
        RECT 347.250 161.850 348.750 162.750 ;
        RECT 349.950 160.950 352.050 163.050 ;
        RECT 353.250 161.850 355.050 162.750 ;
        RECT 344.400 139.050 345.450 160.950 ;
        RECT 349.950 158.850 352.050 159.750 ;
        RECT 343.950 136.950 346.050 139.050 ;
        RECT 343.950 133.950 346.050 136.050 ;
        RECT 340.950 130.950 343.050 133.050 ;
        RECT 344.400 130.050 345.450 133.950 ;
        RECT 343.950 129.450 346.050 130.050 ;
        RECT 341.400 128.400 346.050 129.450 ;
        RECT 337.950 125.250 340.050 126.150 ;
        RECT 337.950 123.450 340.050 124.050 ;
        RECT 335.400 122.400 340.050 123.450 ;
        RECT 337.950 121.950 340.050 122.400 ;
        RECT 338.400 100.050 339.450 121.950 ;
        RECT 337.950 97.950 340.050 100.050 ;
        RECT 341.400 97.050 342.450 128.400 ;
        RECT 343.950 127.950 346.050 128.400 ;
        RECT 343.950 125.850 346.050 126.750 ;
        RECT 346.950 125.250 349.050 126.150 ;
        RECT 346.950 121.950 349.050 124.050 ;
        RECT 347.400 121.050 348.450 121.950 ;
        RECT 346.950 118.950 349.050 121.050 ;
        RECT 356.400 106.050 357.450 166.950 ;
        RECT 359.400 166.050 360.450 196.950 ;
        RECT 358.950 163.950 361.050 166.050 ;
        RECT 362.400 159.450 363.450 230.400 ;
        RECT 364.950 229.950 367.050 232.050 ;
        RECT 377.400 231.450 378.450 250.950 ;
        RECT 379.950 241.950 382.050 244.050 ;
        RECT 374.400 230.400 378.450 231.450 ;
        RECT 370.950 198.450 373.050 199.050 ;
        RECT 374.400 198.450 375.450 230.400 ;
        RECT 380.400 222.450 381.450 241.950 ;
        RECT 386.400 238.050 387.450 259.950 ;
        RECT 389.400 259.050 390.450 289.950 ;
        RECT 392.400 277.050 393.450 292.950 ;
        RECT 391.950 274.950 394.050 277.050 ;
        RECT 392.400 274.050 393.450 274.950 ;
        RECT 391.950 271.950 394.050 274.050 ;
        RECT 391.950 269.850 394.050 270.750 ;
        RECT 395.400 268.050 396.450 335.400 ;
        RECT 406.950 334.950 409.050 337.050 ;
        RECT 406.950 331.950 409.050 334.050 ;
        RECT 397.950 316.950 400.050 319.050 ;
        RECT 400.950 316.950 403.050 319.050 ;
        RECT 403.950 316.950 406.050 319.050 ;
        RECT 398.250 298.050 399.450 316.950 ;
        RECT 401.250 304.350 402.450 316.950 ;
        RECT 400.950 302.250 403.050 304.350 ;
        RECT 401.250 298.050 402.450 302.250 ;
        RECT 404.250 298.050 405.450 316.950 ;
        RECT 397.950 295.950 400.050 298.050 ;
        RECT 400.950 295.950 403.050 298.050 ;
        RECT 403.950 295.950 406.050 298.050 ;
        RECT 407.400 292.050 408.450 331.950 ;
        RECT 413.400 316.050 414.450 337.950 ;
        RECT 416.400 331.050 417.450 337.950 ;
        RECT 415.950 328.950 418.050 331.050 ;
        RECT 412.950 313.950 415.050 316.050 ;
        RECT 415.950 308.250 418.050 309.150 ;
        RECT 409.950 305.850 412.050 306.750 ;
        RECT 415.950 304.950 418.050 307.050 ;
        RECT 416.400 295.050 417.450 304.950 ;
        RECT 415.950 292.950 418.050 295.050 ;
        RECT 406.950 289.950 409.050 292.050 ;
        RECT 403.950 283.950 406.050 286.050 ;
        RECT 404.400 274.050 405.450 283.950 ;
        RECT 419.400 283.050 420.450 343.950 ;
        RECT 422.400 283.050 423.450 376.950 ;
        RECT 424.950 358.950 427.050 361.050 ;
        RECT 425.400 343.050 426.450 358.950 ;
        RECT 431.400 343.050 432.450 379.950 ;
        RECT 446.400 349.050 447.450 379.950 ;
        RECT 445.950 346.950 448.050 349.050 ;
        RECT 436.950 344.250 439.050 345.150 ;
        RECT 424.950 340.950 427.050 343.050 ;
        RECT 427.950 341.250 429.750 342.150 ;
        RECT 430.950 340.950 433.050 343.050 ;
        RECT 434.250 341.250 435.750 342.150 ;
        RECT 436.950 340.950 439.050 343.050 ;
        RECT 427.950 337.950 430.050 340.050 ;
        RECT 431.250 338.850 432.750 339.750 ;
        RECT 433.950 337.950 436.050 340.050 ;
        RECT 428.400 334.050 429.450 337.950 ;
        RECT 437.400 337.050 438.450 340.950 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 427.950 331.950 430.050 334.050 ;
        RECT 433.950 316.950 436.050 319.050 ;
        RECT 427.950 313.950 430.050 316.050 ;
        RECT 428.400 313.050 429.450 313.950 ;
        RECT 434.400 313.050 435.450 316.950 ;
        RECT 437.400 316.050 438.450 334.950 ;
        RECT 439.950 331.950 442.050 334.050 ;
        RECT 436.950 313.950 439.050 316.050 ;
        RECT 427.950 312.450 430.050 313.050 ;
        RECT 425.400 311.400 430.050 312.450 ;
        RECT 425.400 304.050 426.450 311.400 ;
        RECT 427.950 310.950 430.050 311.400 ;
        RECT 431.250 311.250 432.750 312.150 ;
        RECT 433.950 310.950 436.050 313.050 ;
        RECT 427.950 308.850 429.750 309.750 ;
        RECT 430.950 307.950 433.050 310.050 ;
        RECT 434.250 308.850 435.750 309.750 ;
        RECT 436.950 307.950 439.050 310.050 ;
        RECT 436.950 305.850 439.050 306.750 ;
        RECT 424.950 301.950 427.050 304.050 ;
        RECT 436.950 298.950 439.050 301.050 ;
        RECT 418.950 280.950 421.050 283.050 ;
        RECT 421.950 280.950 424.050 283.050 ;
        RECT 412.950 274.950 415.050 277.050 ;
        RECT 403.950 273.450 406.050 274.050 ;
        RECT 401.400 272.400 406.050 273.450 ;
        RECT 409.950 273.450 412.050 274.050 ;
        RECT 413.400 273.450 414.450 274.950 ;
        RECT 394.950 265.950 397.050 268.050 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 388.950 238.950 391.050 241.050 ;
        RECT 394.950 240.450 397.050 241.050 ;
        RECT 392.250 239.250 393.750 240.150 ;
        RECT 394.950 239.400 399.450 240.450 ;
        RECT 394.950 238.950 397.050 239.400 ;
        RECT 385.950 235.950 388.050 238.050 ;
        RECT 389.250 236.850 390.750 237.750 ;
        RECT 391.950 235.950 394.050 238.050 ;
        RECT 395.250 236.850 397.050 237.750 ;
        RECT 385.950 233.850 388.050 234.750 ;
        RECT 370.950 197.400 375.450 198.450 ;
        RECT 370.950 196.950 373.050 197.400 ;
        RECT 367.950 194.250 370.050 195.150 ;
        RECT 370.950 194.850 373.050 195.750 ;
        RECT 367.950 190.950 370.050 193.050 ;
        RECT 374.400 178.050 375.450 197.400 ;
        RECT 377.400 221.400 381.450 222.450 ;
        RECT 377.400 186.450 378.450 221.400 ;
        RECT 379.950 217.950 382.050 220.050 ;
        RECT 380.400 193.050 381.450 217.950 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 382.950 208.950 385.050 211.050 ;
        RECT 383.400 196.050 384.450 208.950 ;
        RECT 389.400 204.450 390.450 211.950 ;
        RECT 392.400 211.050 393.450 235.950 ;
        RECT 398.400 229.050 399.450 239.400 ;
        RECT 397.950 226.950 400.050 229.050 ;
        RECT 391.950 208.950 394.050 211.050 ;
        RECT 386.400 203.400 390.450 204.450 ;
        RECT 386.400 198.450 387.450 203.400 ;
        RECT 394.950 202.950 397.050 205.050 ;
        RECT 388.950 200.250 391.050 201.150 ;
        RECT 395.400 199.050 396.450 202.950 ;
        RECT 401.400 199.050 402.450 272.400 ;
        RECT 403.950 271.950 406.050 272.400 ;
        RECT 407.250 272.250 408.750 273.150 ;
        RECT 409.950 272.400 414.450 273.450 ;
        RECT 409.950 271.950 412.050 272.400 ;
        RECT 403.950 269.850 405.750 270.750 ;
        RECT 406.950 268.950 409.050 271.050 ;
        RECT 410.250 269.850 412.050 270.750 ;
        RECT 403.950 262.950 406.050 265.050 ;
        RECT 388.950 198.450 391.050 199.050 ;
        RECT 386.400 197.400 391.050 198.450 ;
        RECT 388.950 196.950 391.050 197.400 ;
        RECT 392.250 197.250 393.750 198.150 ;
        RECT 394.950 196.950 397.050 199.050 ;
        RECT 398.250 197.250 400.050 198.150 ;
        RECT 400.950 196.950 403.050 199.050 ;
        RECT 382.950 193.950 385.050 196.050 ;
        RECT 391.950 193.950 394.050 196.050 ;
        RECT 395.250 194.850 396.750 195.750 ;
        RECT 397.950 193.950 400.050 196.050 ;
        RECT 379.950 190.950 382.050 193.050 ;
        RECT 377.400 185.400 381.450 186.450 ;
        RECT 376.950 181.950 379.050 184.050 ;
        RECT 373.950 175.950 376.050 178.050 ;
        RECT 364.950 169.950 367.050 172.050 ;
        RECT 365.400 166.050 366.450 169.950 ;
        RECT 374.400 169.050 375.450 175.950 ;
        RECT 367.950 166.950 370.050 169.050 ;
        RECT 371.250 167.250 372.750 168.150 ;
        RECT 373.950 166.950 376.050 169.050 ;
        RECT 364.950 163.950 367.050 166.050 ;
        RECT 368.250 164.850 369.750 165.750 ;
        RECT 370.950 163.950 373.050 166.050 ;
        RECT 374.250 164.850 376.050 165.750 ;
        RECT 364.950 161.850 367.050 162.750 ;
        RECT 362.400 158.400 366.450 159.450 ;
        RECT 361.950 154.950 364.050 157.050 ;
        RECT 362.400 127.050 363.450 154.950 ;
        RECT 361.950 124.950 364.050 127.050 ;
        RECT 365.400 124.050 366.450 158.400 ;
        RECT 377.400 157.050 378.450 181.950 ;
        RECT 380.400 166.050 381.450 185.400 ;
        RECT 382.950 169.950 385.050 172.050 ;
        RECT 379.950 163.950 382.050 166.050 ;
        RECT 383.400 162.450 384.450 169.950 ;
        RECT 388.950 166.950 391.050 169.050 ;
        RECT 389.400 166.050 390.450 166.950 ;
        RECT 385.950 164.250 387.750 165.150 ;
        RECT 388.950 163.950 391.050 166.050 ;
        RECT 394.950 163.950 397.050 166.050 ;
        RECT 385.950 162.450 388.050 163.050 ;
        RECT 383.400 161.400 388.050 162.450 ;
        RECT 389.250 161.850 390.750 162.750 ;
        RECT 376.950 154.950 379.050 157.050 ;
        RECT 383.400 136.050 384.450 161.400 ;
        RECT 385.950 160.950 388.050 161.400 ;
        RECT 391.950 160.950 394.050 163.050 ;
        RECT 395.250 161.850 397.050 162.750 ;
        RECT 391.950 158.850 394.050 159.750 ;
        RECT 382.950 133.950 385.050 136.050 ;
        RECT 376.950 127.950 379.050 130.050 ;
        RECT 382.950 129.450 385.050 130.050 ;
        RECT 380.250 128.250 381.750 129.150 ;
        RECT 382.950 128.400 387.450 129.450 ;
        RECT 382.950 127.950 385.050 128.400 ;
        RECT 386.400 127.050 387.450 128.400 ;
        RECT 394.950 127.950 397.050 130.050 ;
        RECT 395.400 127.050 396.450 127.950 ;
        RECT 376.950 125.850 378.750 126.750 ;
        RECT 379.950 124.950 382.050 127.050 ;
        RECT 383.250 125.850 385.050 126.750 ;
        RECT 385.950 124.950 388.050 127.050 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 358.950 122.250 361.050 123.150 ;
        RECT 361.950 122.850 364.050 123.750 ;
        RECT 364.950 121.950 367.050 124.050 ;
        RECT 358.950 118.950 361.050 121.050 ;
        RECT 355.950 103.950 358.050 106.050 ;
        RECT 334.950 94.950 337.050 97.050 ;
        RECT 338.250 95.850 340.050 96.750 ;
        RECT 340.950 94.950 343.050 97.050 ;
        RECT 346.950 96.450 349.050 97.050 ;
        RECT 344.400 95.400 349.050 96.450 ;
        RECT 334.950 92.850 337.050 93.750 ;
        RECT 344.400 76.050 345.450 95.400 ;
        RECT 346.950 94.950 349.050 95.400 ;
        RECT 355.950 96.450 358.050 97.050 ;
        RECT 359.400 96.450 360.450 118.950 ;
        RECT 364.950 112.950 367.050 115.050 ;
        RECT 355.950 95.400 360.450 96.450 ;
        RECT 355.950 94.950 358.050 95.400 ;
        RECT 346.950 92.850 349.050 93.750 ;
        RECT 352.950 92.250 355.050 93.150 ;
        RECT 355.950 92.850 358.050 93.750 ;
        RECT 352.950 88.950 355.050 91.050 ;
        RECT 365.400 90.450 366.450 112.950 ;
        RECT 367.950 92.250 369.750 93.150 ;
        RECT 370.950 91.950 373.050 94.050 ;
        RECT 374.250 92.250 376.050 93.150 ;
        RECT 367.950 90.450 370.050 91.050 ;
        RECT 365.400 89.400 370.050 90.450 ;
        RECT 371.250 89.850 372.750 90.750 ;
        RECT 367.950 88.950 370.050 89.400 ;
        RECT 373.950 88.950 376.050 91.050 ;
        RECT 349.950 79.950 352.050 82.050 ;
        RECT 343.950 73.950 346.050 76.050 ;
        RECT 337.950 61.950 340.050 64.050 ;
        RECT 332.400 56.400 336.450 57.450 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 323.250 53.250 324.750 54.150 ;
        RECT 325.950 52.950 328.050 55.050 ;
        RECT 329.250 53.250 331.050 54.150 ;
        RECT 331.950 52.950 334.050 55.050 ;
        RECT 322.950 49.950 325.050 52.050 ;
        RECT 326.250 50.850 327.750 51.750 ;
        RECT 328.950 51.450 331.050 52.050 ;
        RECT 332.400 51.450 333.450 52.950 ;
        RECT 328.950 50.400 333.450 51.450 ;
        RECT 328.950 49.950 331.050 50.400 ;
        RECT 323.400 25.050 324.450 49.950 ;
        RECT 325.950 28.950 328.050 31.050 ;
        RECT 326.400 28.050 327.450 28.950 ;
        RECT 325.950 25.950 328.050 28.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 317.400 22.050 318.450 22.950 ;
        RECT 313.950 20.250 315.750 21.150 ;
        RECT 316.950 19.950 319.050 22.050 ;
        RECT 322.950 21.450 325.050 22.050 ;
        RECT 326.400 21.450 327.450 25.950 ;
        RECT 331.950 24.450 334.050 25.050 ;
        RECT 335.400 24.450 336.450 56.400 ;
        RECT 338.400 28.050 339.450 61.950 ;
        RECT 350.400 55.050 351.450 79.950 ;
        RECT 352.950 58.950 355.050 61.050 ;
        RECT 340.950 53.250 342.750 54.150 ;
        RECT 343.950 52.950 346.050 55.050 ;
        RECT 349.950 52.950 352.050 55.050 ;
        RECT 340.950 49.950 343.050 52.050 ;
        RECT 344.250 50.850 346.050 51.750 ;
        RECT 346.950 50.250 349.050 51.150 ;
        RECT 349.950 50.850 352.050 51.750 ;
        RECT 353.400 49.050 354.450 58.950 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 368.400 52.050 369.450 88.950 ;
        RECT 374.400 85.050 375.450 88.950 ;
        RECT 373.950 82.950 376.050 85.050 ;
        RECT 380.400 64.050 381.450 124.950 ;
        RECT 394.950 122.850 397.050 123.750 ;
        RECT 398.400 115.050 399.450 193.950 ;
        RECT 401.400 166.050 402.450 196.950 ;
        RECT 404.400 181.050 405.450 262.950 ;
        RECT 407.400 262.050 408.450 268.950 ;
        RECT 413.400 265.050 414.450 272.400 ;
        RECT 415.950 271.950 418.050 274.050 ;
        RECT 412.950 262.950 415.050 265.050 ;
        RECT 406.950 259.950 409.050 262.050 ;
        RECT 407.400 244.050 408.450 259.950 ;
        RECT 406.950 241.950 409.050 244.050 ;
        RECT 416.400 241.050 417.450 271.950 ;
        RECT 419.400 271.050 420.450 280.950 ;
        RECT 421.950 277.950 424.050 280.050 ;
        RECT 418.950 268.950 421.050 271.050 ;
        RECT 422.400 265.050 423.450 277.950 ;
        RECT 430.950 275.250 433.050 276.150 ;
        RECT 424.950 271.950 427.050 274.050 ;
        RECT 428.250 272.250 429.750 273.150 ;
        RECT 434.250 272.250 436.050 273.150 ;
        RECT 424.950 269.850 426.750 270.750 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 433.950 268.950 436.050 271.050 ;
        RECT 434.400 268.050 435.450 268.950 ;
        RECT 433.950 265.950 436.050 268.050 ;
        RECT 421.950 262.950 424.050 265.050 ;
        RECT 437.400 262.050 438.450 298.950 ;
        RECT 436.950 259.950 439.050 262.050 ;
        RECT 421.950 256.950 424.050 259.050 ;
        RECT 436.950 256.950 439.050 259.050 ;
        RECT 418.950 241.950 421.050 244.050 ;
        RECT 415.950 238.950 418.050 241.050 ;
        RECT 406.950 236.250 408.750 237.150 ;
        RECT 409.950 235.950 412.050 238.050 ;
        RECT 413.250 236.250 415.050 237.150 ;
        RECT 406.950 232.950 409.050 235.050 ;
        RECT 410.250 233.850 411.750 234.750 ;
        RECT 412.950 232.950 415.050 235.050 ;
        RECT 413.400 232.050 414.450 232.950 ;
        RECT 419.400 232.050 420.450 241.950 ;
        RECT 412.950 229.950 415.050 232.050 ;
        RECT 418.950 229.950 421.050 232.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 410.400 199.050 411.450 211.950 ;
        RECT 413.400 200.400 420.450 201.450 ;
        RECT 413.400 199.050 414.450 200.400 ;
        RECT 409.950 196.950 412.050 199.050 ;
        RECT 412.950 196.950 415.050 199.050 ;
        RECT 416.250 197.250 418.050 198.150 ;
        RECT 406.950 194.850 409.050 195.750 ;
        RECT 409.950 194.250 412.050 195.150 ;
        RECT 412.950 194.850 414.750 195.750 ;
        RECT 415.950 193.950 418.050 196.050 ;
        RECT 409.950 190.950 412.050 193.050 ;
        RECT 415.950 190.950 418.050 193.050 ;
        RECT 410.400 184.050 411.450 190.950 ;
        RECT 409.950 181.950 412.050 184.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 413.400 169.050 414.450 178.950 ;
        RECT 406.950 167.850 409.050 168.750 ;
        RECT 409.950 167.250 412.050 168.150 ;
        RECT 412.950 166.950 415.050 169.050 ;
        RECT 400.950 163.950 403.050 166.050 ;
        RECT 409.950 163.950 412.050 166.050 ;
        RECT 413.400 130.050 414.450 166.950 ;
        RECT 416.400 166.050 417.450 190.950 ;
        RECT 419.400 184.050 420.450 200.400 ;
        RECT 422.400 196.050 423.450 256.950 ;
        RECT 433.950 247.950 436.050 250.050 ;
        RECT 427.950 244.950 430.050 247.050 ;
        RECT 428.400 241.050 429.450 244.950 ;
        RECT 434.400 241.050 435.450 247.950 ;
        RECT 424.950 238.950 427.050 241.050 ;
        RECT 427.950 238.950 430.050 241.050 ;
        RECT 431.250 239.250 432.750 240.150 ;
        RECT 433.950 238.950 436.050 241.050 ;
        RECT 425.400 238.050 426.450 238.950 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 428.250 236.850 429.750 237.750 ;
        RECT 430.950 235.950 433.050 238.050 ;
        RECT 434.250 236.850 436.050 237.750 ;
        RECT 424.950 233.850 427.050 234.750 ;
        RECT 427.950 226.950 430.050 229.050 ;
        RECT 424.950 208.950 427.050 211.050 ;
        RECT 425.400 196.050 426.450 208.950 ;
        RECT 428.400 208.050 429.450 226.950 ;
        RECT 431.400 211.050 432.450 235.950 ;
        RECT 437.400 232.050 438.450 256.950 ;
        RECT 436.950 229.950 439.050 232.050 ;
        RECT 440.400 214.050 441.450 331.950 ;
        RECT 449.400 301.050 450.450 380.400 ;
        RECT 454.950 379.950 457.050 382.050 ;
        RECT 457.950 380.850 459.750 381.750 ;
        RECT 460.950 379.950 463.050 382.050 ;
        RECT 464.250 380.850 465.750 381.750 ;
        RECT 466.950 381.450 469.050 382.050 ;
        RECT 466.950 380.400 471.450 381.450 ;
        RECT 466.950 379.950 469.050 380.400 ;
        RECT 461.400 370.050 462.450 379.950 ;
        RECT 466.950 377.850 469.050 378.750 ;
        RECT 460.950 367.950 463.050 370.050 ;
        RECT 451.950 361.950 454.050 364.050 ;
        RECT 452.400 346.050 453.450 361.950 ;
        RECT 463.950 355.950 466.050 358.050 ;
        RECT 457.950 346.950 460.050 349.050 ;
        RECT 458.400 346.050 459.450 346.950 ;
        RECT 451.950 343.950 454.050 346.050 ;
        RECT 455.250 344.250 456.750 345.150 ;
        RECT 457.950 343.950 460.050 346.050 ;
        RECT 451.950 341.850 453.750 342.750 ;
        RECT 454.950 340.950 457.050 343.050 ;
        RECT 458.250 341.850 460.050 342.750 ;
        RECT 454.950 337.950 457.050 340.050 ;
        RECT 455.400 322.050 456.450 337.950 ;
        RECT 454.950 319.950 457.050 322.050 ;
        RECT 451.950 308.250 453.750 309.150 ;
        RECT 454.950 307.950 457.050 310.050 ;
        RECT 458.250 308.250 460.050 309.150 ;
        RECT 451.950 304.950 454.050 307.050 ;
        RECT 455.250 305.850 456.750 306.750 ;
        RECT 457.950 304.950 460.050 307.050 ;
        RECT 448.950 298.950 451.050 301.050 ;
        RECT 452.400 297.450 453.450 304.950 ;
        RECT 458.400 304.050 459.450 304.950 ;
        RECT 457.950 301.950 460.050 304.050 ;
        RECT 458.400 301.050 459.450 301.950 ;
        RECT 457.950 298.950 460.050 301.050 ;
        RECT 449.400 296.400 453.450 297.450 ;
        RECT 449.400 280.050 450.450 296.400 ;
        RECT 451.950 289.950 454.050 292.050 ;
        RECT 448.950 277.950 451.050 280.050 ;
        RECT 445.950 272.250 448.050 273.150 ;
        RECT 452.400 271.050 453.450 289.950 ;
        RECT 445.950 268.950 448.050 271.050 ;
        RECT 449.250 269.250 450.750 270.150 ;
        RECT 451.950 268.950 454.050 271.050 ;
        RECT 455.250 269.250 457.050 270.150 ;
        RECT 448.950 265.950 451.050 268.050 ;
        RECT 452.250 266.850 453.750 267.750 ;
        RECT 454.950 265.950 457.050 268.050 ;
        RECT 449.400 265.050 450.450 265.950 ;
        RECT 455.400 265.050 456.450 265.950 ;
        RECT 448.950 262.950 451.050 265.050 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 448.950 244.950 451.050 247.050 ;
        RECT 449.400 241.050 450.450 244.950 ;
        RECT 458.400 244.050 459.450 298.950 ;
        RECT 460.950 292.950 463.050 295.050 ;
        RECT 461.400 264.450 462.450 292.950 ;
        RECT 464.400 274.050 465.450 355.950 ;
        RECT 470.400 346.050 471.450 380.400 ;
        RECT 473.400 379.050 474.450 382.950 ;
        RECT 472.950 376.950 475.050 379.050 ;
        RECT 476.400 376.050 477.450 385.950 ;
        RECT 479.400 385.050 480.450 388.950 ;
        RECT 482.400 388.050 483.450 415.950 ;
        RECT 485.400 412.050 486.450 418.950 ;
        RECT 484.950 409.950 487.050 412.050 ;
        RECT 488.400 409.050 489.450 418.950 ;
        RECT 497.400 418.050 498.450 496.950 ;
        RECT 500.400 484.050 501.450 517.950 ;
        RECT 503.400 505.050 504.450 517.950 ;
        RECT 511.950 514.950 514.050 517.050 ;
        RECT 512.400 505.050 513.450 514.950 ;
        RECT 502.950 502.950 505.050 505.050 ;
        RECT 511.950 502.950 514.050 505.050 ;
        RECT 508.950 487.950 511.050 490.050 ;
        RECT 505.950 484.950 508.050 487.050 ;
        RECT 499.950 481.950 502.050 484.050 ;
        RECT 502.950 482.250 505.050 483.150 ;
        RECT 505.950 482.850 508.050 483.750 ;
        RECT 502.950 478.950 505.050 481.050 ;
        RECT 502.950 472.950 505.050 475.050 ;
        RECT 499.950 466.950 502.050 469.050 ;
        RECT 500.400 460.050 501.450 466.950 ;
        RECT 499.950 457.950 502.050 460.050 ;
        RECT 503.400 457.050 504.450 472.950 ;
        RECT 509.400 463.050 510.450 487.950 ;
        RECT 508.950 460.950 511.050 463.050 ;
        RECT 499.950 455.850 501.750 456.750 ;
        RECT 502.950 454.950 505.050 457.050 ;
        RECT 505.950 454.950 508.050 457.050 ;
        RECT 508.950 455.250 511.050 456.150 ;
        RECT 502.950 452.850 505.050 453.750 ;
        RECT 506.400 442.050 507.450 454.950 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 508.950 448.950 511.050 451.050 ;
        RECT 505.950 439.950 508.050 442.050 ;
        RECT 493.950 416.250 496.050 417.150 ;
        RECT 496.950 415.950 499.050 418.050 ;
        RECT 505.950 415.950 508.050 418.050 ;
        RECT 497.250 413.250 498.750 414.150 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 503.250 413.250 505.050 414.150 ;
        RECT 496.950 409.950 499.050 412.050 ;
        RECT 500.250 410.850 501.750 411.750 ;
        RECT 502.950 409.950 505.050 412.050 ;
        RECT 503.400 409.050 504.450 409.950 ;
        RECT 487.950 406.950 490.050 409.050 ;
        RECT 502.950 406.950 505.050 409.050 ;
        RECT 493.950 400.950 496.050 403.050 ;
        RECT 496.950 400.950 499.050 403.050 ;
        RECT 484.950 388.950 487.050 391.050 ;
        RECT 481.950 385.950 484.050 388.050 ;
        RECT 478.950 382.950 481.050 385.050 ;
        RECT 485.400 382.050 486.450 388.950 ;
        RECT 490.950 382.950 493.050 385.050 ;
        RECT 478.950 379.950 481.050 382.050 ;
        RECT 481.950 380.250 483.750 381.150 ;
        RECT 484.950 379.950 487.050 382.050 ;
        RECT 488.250 380.250 490.050 381.150 ;
        RECT 475.950 373.950 478.050 376.050 ;
        RECT 479.400 373.050 480.450 379.950 ;
        RECT 491.400 379.050 492.450 382.950 ;
        RECT 481.950 376.950 484.050 379.050 ;
        RECT 485.250 377.850 486.750 378.750 ;
        RECT 487.950 376.950 490.050 379.050 ;
        RECT 490.950 376.950 493.050 379.050 ;
        RECT 481.950 373.950 484.050 376.050 ;
        RECT 478.950 370.950 481.050 373.050 ;
        RECT 478.950 361.950 481.050 364.050 ;
        RECT 479.400 355.050 480.450 361.950 ;
        RECT 478.950 352.950 481.050 355.050 ;
        RECT 475.950 349.950 478.050 352.050 ;
        RECT 478.950 349.950 481.050 352.050 ;
        RECT 476.400 346.050 477.450 349.950 ;
        RECT 469.950 345.450 472.050 346.050 ;
        RECT 467.400 344.400 472.050 345.450 ;
        RECT 467.400 337.050 468.450 344.400 ;
        RECT 469.950 343.950 472.050 344.400 ;
        RECT 473.250 344.250 474.750 345.150 ;
        RECT 475.950 343.950 478.050 346.050 ;
        RECT 469.950 341.850 471.750 342.750 ;
        RECT 472.950 340.950 475.050 343.050 ;
        RECT 476.250 341.850 478.050 342.750 ;
        RECT 473.400 337.050 474.450 340.950 ;
        RECT 479.400 340.050 480.450 349.950 ;
        RECT 482.400 340.050 483.450 373.950 ;
        RECT 494.400 370.050 495.450 400.950 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 487.950 358.950 490.050 361.050 ;
        RECT 484.950 352.950 487.050 355.050 ;
        RECT 478.950 337.950 481.050 340.050 ;
        RECT 481.950 337.950 484.050 340.050 ;
        RECT 466.950 334.950 469.050 337.050 ;
        RECT 472.950 334.950 475.050 337.050 ;
        RECT 478.950 336.450 481.050 337.050 ;
        RECT 481.950 336.450 484.050 337.050 ;
        RECT 478.950 335.400 484.050 336.450 ;
        RECT 478.950 334.950 481.050 335.400 ;
        RECT 481.950 334.950 484.050 335.400 ;
        RECT 469.950 325.950 472.050 328.050 ;
        RECT 470.400 310.050 471.450 325.950 ;
        RECT 475.950 313.950 478.050 316.050 ;
        RECT 466.950 308.250 468.750 309.150 ;
        RECT 469.950 307.950 472.050 310.050 ;
        RECT 473.250 308.250 475.050 309.150 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 470.250 305.850 471.750 306.750 ;
        RECT 472.950 306.450 475.050 307.050 ;
        RECT 476.400 306.450 477.450 313.950 ;
        RECT 485.400 310.050 486.450 352.950 ;
        RECT 488.400 346.050 489.450 358.950 ;
        RECT 497.400 346.050 498.450 400.950 ;
        RECT 506.400 400.050 507.450 415.950 ;
        RECT 509.400 403.050 510.450 448.950 ;
        RECT 512.400 418.050 513.450 502.950 ;
        RECT 515.400 478.050 516.450 526.950 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 524.250 524.850 525.750 525.750 ;
        RECT 526.950 523.950 529.050 526.050 ;
        RECT 530.250 524.850 532.050 525.750 ;
        RECT 517.950 520.950 520.050 523.050 ;
        RECT 520.950 521.850 523.050 522.750 ;
        RECT 523.950 520.950 526.050 523.050 ;
        RECT 518.400 514.050 519.450 520.950 ;
        RECT 524.400 517.050 525.450 520.950 ;
        RECT 523.950 514.950 526.050 517.050 ;
        RECT 517.950 511.950 520.050 514.050 ;
        RECT 533.400 508.050 534.450 532.950 ;
        RECT 532.950 505.950 535.050 508.050 ;
        RECT 536.400 499.050 537.450 559.950 ;
        RECT 539.400 519.450 540.450 625.950 ;
        RECT 548.400 625.050 549.450 628.950 ;
        RECT 541.950 622.950 544.050 625.050 ;
        RECT 547.950 622.950 550.050 625.050 ;
        RECT 542.400 553.050 543.450 622.950 ;
        RECT 557.400 613.050 558.450 688.950 ;
        RECT 560.400 628.050 561.450 694.950 ;
        RECT 566.400 694.050 567.450 694.950 ;
        RECT 565.950 691.950 568.050 694.050 ;
        RECT 571.950 682.950 574.050 685.050 ;
        RECT 572.400 676.050 573.450 682.950 ;
        RECT 571.950 673.950 574.050 676.050 ;
        RECT 562.950 671.250 565.050 672.150 ;
        RECT 568.950 670.950 571.050 673.050 ;
        RECT 572.250 671.850 574.050 672.750 ;
        RECT 562.950 667.950 565.050 670.050 ;
        RECT 568.950 668.850 571.050 669.750 ;
        RECT 571.950 667.950 574.050 670.050 ;
        RECT 565.950 635.250 568.050 636.150 ;
        RECT 572.400 634.050 573.450 667.950 ;
        RECT 562.950 632.250 564.750 633.150 ;
        RECT 565.950 631.950 568.050 634.050 ;
        RECT 569.250 632.250 570.750 633.150 ;
        RECT 571.950 631.950 574.050 634.050 ;
        RECT 575.400 631.050 576.450 703.950 ;
        RECT 577.950 700.950 580.050 703.050 ;
        RECT 577.950 699.450 580.050 700.050 ;
        RECT 581.400 699.450 582.450 703.950 ;
        RECT 583.950 700.950 586.050 703.050 ;
        RECT 587.250 701.850 589.050 702.750 ;
        RECT 577.950 698.400 582.450 699.450 ;
        RECT 577.950 697.950 580.050 698.400 ;
        RECT 578.400 670.050 579.450 697.950 ;
        RECT 584.400 697.050 585.450 700.950 ;
        RECT 583.950 694.950 586.050 697.050 ;
        RECT 584.400 694.050 585.450 694.950 ;
        RECT 583.950 691.950 586.050 694.050 ;
        RECT 590.400 691.050 591.450 739.950 ;
        RECT 596.400 730.050 597.450 778.950 ;
        RECT 611.400 778.050 612.450 802.950 ;
        RECT 601.950 776.250 603.750 777.150 ;
        RECT 604.950 775.950 607.050 778.050 ;
        RECT 608.250 776.250 609.750 777.150 ;
        RECT 610.950 775.950 613.050 778.050 ;
        RECT 598.950 772.950 601.050 775.050 ;
        RECT 601.950 774.450 604.050 775.050 ;
        RECT 601.950 773.400 606.450 774.450 ;
        RECT 601.950 772.950 604.050 773.400 ;
        RECT 599.400 763.050 600.450 772.950 ;
        RECT 601.950 769.950 604.050 772.050 ;
        RECT 602.400 769.050 603.450 769.950 ;
        RECT 601.950 766.950 604.050 769.050 ;
        RECT 598.950 760.950 601.050 763.050 ;
        RECT 601.950 745.950 604.050 748.050 ;
        RECT 602.400 742.050 603.450 745.950 ;
        RECT 601.950 739.950 604.050 742.050 ;
        RECT 605.400 739.050 606.450 773.400 ;
        RECT 607.950 772.950 610.050 775.050 ;
        RECT 611.250 773.850 613.050 774.750 ;
        RECT 613.950 757.950 616.050 760.050 ;
        RECT 607.950 742.950 610.050 745.050 ;
        RECT 608.400 742.050 609.450 742.950 ;
        RECT 607.950 739.950 610.050 742.050 ;
        RECT 611.250 740.250 613.050 741.150 ;
        RECT 601.950 737.850 603.750 738.750 ;
        RECT 604.950 736.950 607.050 739.050 ;
        RECT 608.250 737.850 609.750 738.750 ;
        RECT 610.950 736.950 613.050 739.050 ;
        RECT 604.950 734.850 607.050 735.750 ;
        RECT 595.950 727.950 598.050 730.050 ;
        RECT 592.950 718.950 595.050 721.050 ;
        RECT 593.400 706.050 594.450 718.950 ;
        RECT 592.950 703.950 595.050 706.050 ;
        RECT 589.950 688.950 592.050 691.050 ;
        RECT 589.950 682.950 592.050 685.050 ;
        RECT 583.950 673.950 586.050 676.050 ;
        RECT 584.400 670.050 585.450 673.950 ;
        RECT 577.950 667.950 580.050 670.050 ;
        RECT 580.950 668.250 582.750 669.150 ;
        RECT 583.950 667.950 586.050 670.050 ;
        RECT 587.250 668.250 589.050 669.150 ;
        RECT 580.950 664.950 583.050 667.050 ;
        RECT 584.250 665.850 585.750 666.750 ;
        RECT 586.950 666.450 589.050 667.050 ;
        RECT 590.400 666.450 591.450 682.950 ;
        RECT 586.950 665.400 591.450 666.450 ;
        RECT 586.950 664.950 589.050 665.400 ;
        RECT 586.950 637.950 589.050 640.050 ;
        RECT 587.400 634.050 588.450 637.950 ;
        RECT 596.400 637.050 597.450 727.950 ;
        RECT 601.950 707.250 604.050 708.150 ;
        RECT 598.950 704.250 600.750 705.150 ;
        RECT 601.950 703.950 604.050 706.050 ;
        RECT 607.950 705.450 610.050 706.050 ;
        RECT 605.250 704.250 606.750 705.150 ;
        RECT 607.950 704.400 612.450 705.450 ;
        RECT 607.950 703.950 610.050 704.400 ;
        RECT 598.950 700.950 601.050 703.050 ;
        RECT 604.950 700.950 607.050 703.050 ;
        RECT 608.250 701.850 610.050 702.750 ;
        RECT 599.400 700.050 600.450 700.950 ;
        RECT 598.950 697.950 601.050 700.050 ;
        RECT 595.950 634.950 598.050 637.050 ;
        RECT 586.950 631.950 589.050 634.050 ;
        RECT 592.950 633.450 595.050 634.050 ;
        RECT 590.250 632.250 591.750 633.150 ;
        RECT 592.950 632.400 597.450 633.450 ;
        RECT 592.950 631.950 595.050 632.400 ;
        RECT 562.950 630.450 565.050 631.050 ;
        RECT 562.950 629.400 567.450 630.450 ;
        RECT 562.950 628.950 565.050 629.400 ;
        RECT 559.950 625.950 562.050 628.050 ;
        RECT 544.950 610.950 547.050 613.050 ;
        RECT 556.950 610.950 559.050 613.050 ;
        RECT 559.950 610.950 562.050 613.050 ;
        RECT 545.400 571.050 546.450 610.950 ;
        RECT 556.950 607.950 559.050 610.050 ;
        RECT 557.400 601.050 558.450 607.950 ;
        RECT 560.400 604.050 561.450 610.950 ;
        RECT 566.400 607.050 567.450 629.400 ;
        RECT 568.950 628.950 571.050 631.050 ;
        RECT 572.250 629.850 574.050 630.750 ;
        RECT 574.950 628.950 577.050 631.050 ;
        RECT 586.950 629.850 588.750 630.750 ;
        RECT 589.950 628.950 592.050 631.050 ;
        RECT 593.250 629.850 595.050 630.750 ;
        RECT 596.400 628.050 597.450 632.400 ;
        RECT 595.950 625.950 598.050 628.050 ;
        RECT 599.400 625.050 600.450 697.950 ;
        RECT 605.400 691.050 606.450 700.950 ;
        RECT 611.400 697.050 612.450 704.400 ;
        RECT 610.950 694.950 613.050 697.050 ;
        RECT 604.950 688.950 607.050 691.050 ;
        RECT 601.950 673.950 604.050 676.050 ;
        RECT 602.400 673.050 603.450 673.950 ;
        RECT 601.950 670.950 604.050 673.050 ;
        RECT 601.950 668.850 604.050 669.750 ;
        RECT 605.400 667.050 606.450 688.950 ;
        RECT 614.400 679.050 615.450 757.950 ;
        RECT 620.400 754.050 621.450 805.950 ;
        RECT 632.400 805.050 633.450 808.950 ;
        RECT 655.950 806.850 658.050 807.750 ;
        RECT 631.950 802.950 634.050 805.050 ;
        RECT 640.950 799.950 643.050 802.050 ;
        RECT 625.950 776.250 628.050 777.150 ;
        RECT 637.950 775.950 640.050 778.050 ;
        RECT 625.950 772.950 628.050 775.050 ;
        RECT 629.250 773.250 630.750 774.150 ;
        RECT 631.950 772.950 634.050 775.050 ;
        RECT 635.250 773.250 637.050 774.150 ;
        RECT 626.400 769.050 627.450 772.950 ;
        RECT 638.400 772.050 639.450 775.950 ;
        RECT 628.950 769.950 631.050 772.050 ;
        RECT 632.250 770.850 633.750 771.750 ;
        RECT 634.950 769.950 637.050 772.050 ;
        RECT 637.950 769.950 640.050 772.050 ;
        RECT 625.950 766.950 628.050 769.050 ;
        RECT 619.950 751.950 622.050 754.050 ;
        RECT 619.950 745.950 622.050 748.050 ;
        RECT 616.950 742.950 619.050 745.050 ;
        RECT 617.400 739.050 618.450 742.950 ;
        RECT 620.400 741.450 621.450 745.950 ;
        RECT 626.400 745.050 627.450 766.950 ;
        RECT 635.400 757.050 636.450 769.950 ;
        RECT 634.950 754.950 637.050 757.050 ;
        RECT 634.950 751.950 637.050 754.050 ;
        RECT 625.950 742.950 628.050 745.050 ;
        RECT 622.950 741.450 625.050 742.050 ;
        RECT 620.400 740.400 625.050 741.450 ;
        RECT 616.950 736.950 619.050 739.050 ;
        RECT 620.400 735.450 621.450 740.400 ;
        RECT 622.950 739.950 625.050 740.400 ;
        RECT 628.950 739.950 631.050 742.050 ;
        RECT 632.250 740.250 634.050 741.150 ;
        RECT 622.950 737.850 624.750 738.750 ;
        RECT 625.950 736.950 628.050 739.050 ;
        RECT 629.250 737.850 630.750 738.750 ;
        RECT 631.950 736.950 634.050 739.050 ;
        RECT 617.400 734.400 621.450 735.450 ;
        RECT 625.950 734.850 628.050 735.750 ;
        RECT 617.400 682.050 618.450 734.400 ;
        RECT 622.950 712.950 625.050 715.050 ;
        RECT 623.400 703.050 624.450 712.950 ;
        RECT 625.950 703.950 628.050 706.050 ;
        RECT 626.400 703.050 627.450 703.950 ;
        RECT 622.950 700.950 625.050 703.050 ;
        RECT 625.950 700.950 628.050 703.050 ;
        RECT 619.950 698.250 622.050 699.150 ;
        RECT 622.950 698.850 625.050 699.750 ;
        RECT 626.400 697.050 627.450 700.950 ;
        RECT 619.950 694.950 622.050 697.050 ;
        RECT 625.950 694.950 628.050 697.050 ;
        RECT 635.400 691.050 636.450 751.950 ;
        RECT 641.400 745.050 642.450 799.950 ;
        RECT 661.950 781.950 664.050 784.050 ;
        RECT 655.950 776.250 658.050 777.150 ;
        RECT 643.950 772.950 646.050 775.050 ;
        RECT 646.950 773.250 648.750 774.150 ;
        RECT 649.950 772.950 652.050 775.050 ;
        RECT 653.250 773.250 654.750 774.150 ;
        RECT 655.950 772.950 658.050 775.050 ;
        RECT 644.400 765.450 645.450 772.950 ;
        RECT 656.400 772.050 657.450 772.950 ;
        RECT 646.950 769.950 649.050 772.050 ;
        RECT 650.250 770.850 651.750 771.750 ;
        RECT 652.950 769.950 655.050 772.050 ;
        RECT 655.950 769.950 658.050 772.050 ;
        RECT 647.400 769.050 648.450 769.950 ;
        RECT 646.950 766.950 649.050 769.050 ;
        RECT 644.400 764.400 648.450 765.450 ;
        RECT 647.400 745.050 648.450 764.400 ;
        RECT 658.950 760.950 661.050 763.050 ;
        RECT 655.950 745.950 658.050 748.050 ;
        RECT 656.400 745.050 657.450 745.950 ;
        RECT 640.950 742.950 643.050 745.050 ;
        RECT 643.950 742.950 646.050 745.050 ;
        RECT 646.950 742.950 649.050 745.050 ;
        RECT 655.950 744.450 658.050 745.050 ;
        RECT 653.400 743.400 658.050 744.450 ;
        RECT 640.950 733.950 643.050 736.050 ;
        RECT 641.400 733.050 642.450 733.950 ;
        RECT 640.950 730.950 643.050 733.050 ;
        RECT 641.400 709.050 642.450 730.950 ;
        RECT 640.950 706.950 643.050 709.050 ;
        RECT 641.400 706.050 642.450 706.950 ;
        RECT 640.950 703.950 643.050 706.050 ;
        RECT 644.400 703.050 645.450 742.950 ;
        RECT 646.950 740.850 649.050 741.750 ;
        RECT 649.950 740.250 652.050 741.150 ;
        RECT 653.400 739.050 654.450 743.400 ;
        RECT 655.950 742.950 658.050 743.400 ;
        RECT 655.950 740.850 658.050 741.750 ;
        RECT 649.950 736.950 652.050 739.050 ;
        RECT 652.950 736.950 655.050 739.050 ;
        RECT 655.950 736.950 658.050 739.050 ;
        RECT 650.400 724.050 651.450 736.950 ;
        RECT 649.950 721.950 652.050 724.050 ;
        RECT 637.950 701.250 640.050 702.150 ;
        RECT 640.950 701.850 643.050 702.750 ;
        RECT 643.950 700.950 646.050 703.050 ;
        RECT 646.950 701.250 649.050 702.150 ;
        RECT 649.950 700.950 652.050 703.050 ;
        RECT 637.950 697.950 640.050 700.050 ;
        RECT 646.950 697.950 649.050 700.050 ;
        RECT 638.400 694.050 639.450 697.950 ;
        RECT 637.950 691.950 640.050 694.050 ;
        RECT 634.950 688.950 637.050 691.050 ;
        RECT 634.950 685.950 637.050 688.050 ;
        RECT 616.950 679.950 619.050 682.050 ;
        RECT 607.950 676.950 610.050 679.050 ;
        RECT 613.950 676.950 616.050 679.050 ;
        RECT 608.400 673.050 609.450 676.950 ;
        RECT 617.400 676.050 618.450 679.950 ;
        RECT 616.950 673.950 619.050 676.050 ;
        RECT 617.400 673.050 618.450 673.950 ;
        RECT 607.950 670.950 610.050 673.050 ;
        RECT 616.950 670.950 619.050 673.050 ;
        RECT 625.950 672.450 628.050 673.050 ;
        RECT 625.950 671.400 630.450 672.450 ;
        RECT 625.950 670.950 628.050 671.400 ;
        RECT 607.950 668.850 610.050 669.750 ;
        RECT 616.950 668.850 619.050 669.750 ;
        RECT 622.950 668.250 625.050 669.150 ;
        RECT 625.950 668.850 628.050 669.750 ;
        RECT 604.950 664.950 607.050 667.050 ;
        RECT 622.950 664.950 625.050 667.050 ;
        RECT 605.400 639.450 606.450 664.950 ;
        RECT 623.400 664.050 624.450 664.950 ;
        RECT 622.950 661.950 625.050 664.050 ;
        RECT 605.400 638.400 609.450 639.450 ;
        RECT 604.950 634.950 607.050 637.050 ;
        RECT 598.950 622.950 601.050 625.050 ;
        RECT 580.950 610.950 583.050 613.050 ;
        RECT 568.950 607.950 571.050 610.050 ;
        RECT 565.950 604.950 568.050 607.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 550.950 599.250 553.050 600.150 ;
        RECT 556.950 598.950 559.050 601.050 ;
        RECT 560.250 599.850 562.050 600.750 ;
        RECT 562.950 598.950 565.050 601.050 ;
        RECT 550.950 595.950 553.050 598.050 ;
        RECT 556.950 596.850 559.050 597.750 ;
        RECT 551.400 595.050 552.450 595.950 ;
        RECT 550.950 592.950 553.050 595.050 ;
        RECT 556.950 589.950 559.050 592.050 ;
        RECT 544.950 568.950 547.050 571.050 ;
        RECT 545.400 556.050 546.450 568.950 ;
        RECT 557.400 562.050 558.450 589.950 ;
        RECT 556.950 559.950 559.050 562.050 ;
        RECT 547.950 557.250 550.050 558.150 ;
        RECT 553.950 557.250 556.050 558.150 ;
        RECT 544.950 553.950 547.050 556.050 ;
        RECT 547.950 553.950 550.050 556.050 ;
        RECT 551.250 554.250 552.750 555.150 ;
        RECT 553.950 553.950 556.050 556.050 ;
        RECT 541.950 550.950 544.050 553.050 ;
        RECT 544.950 541.950 547.050 544.050 ;
        RECT 541.950 535.950 544.050 538.050 ;
        RECT 542.400 526.050 543.450 535.950 ;
        RECT 545.400 529.050 546.450 541.950 ;
        RECT 548.400 535.050 549.450 553.950 ;
        RECT 550.950 550.950 553.050 553.050 ;
        RECT 551.400 547.050 552.450 550.950 ;
        RECT 550.950 544.950 553.050 547.050 ;
        RECT 550.950 541.950 553.050 544.050 ;
        RECT 547.950 532.950 550.050 535.050 ;
        RECT 551.400 529.050 552.450 541.950 ;
        RECT 553.950 529.950 556.050 532.050 ;
        RECT 544.950 526.950 547.050 529.050 ;
        RECT 548.250 527.250 549.750 528.150 ;
        RECT 550.950 526.950 553.050 529.050 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 545.250 524.850 546.750 525.750 ;
        RECT 547.950 523.950 550.050 526.050 ;
        RECT 551.250 524.850 553.050 525.750 ;
        RECT 541.950 521.850 544.050 522.750 ;
        RECT 539.400 518.400 543.450 519.450 ;
        RECT 535.950 496.950 538.050 499.050 ;
        RECT 542.400 493.050 543.450 518.400 ;
        RECT 550.950 517.950 553.050 520.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 526.950 491.250 529.050 492.150 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 514.950 475.950 517.050 478.050 ;
        RECT 515.400 469.050 516.450 475.950 ;
        RECT 514.950 466.950 517.050 469.050 ;
        RECT 518.400 451.050 519.450 490.950 ;
        RECT 551.400 490.050 552.450 517.950 ;
        RECT 554.400 514.050 555.450 529.950 ;
        RECT 553.950 511.950 556.050 514.050 ;
        RECT 553.950 508.950 556.050 511.050 ;
        RECT 520.950 487.950 523.050 490.050 ;
        RECT 524.250 488.250 525.750 489.150 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 530.250 488.250 532.050 489.150 ;
        RECT 550.950 487.950 553.050 490.050 ;
        RECT 520.950 485.850 522.750 486.750 ;
        RECT 523.950 484.950 526.050 487.050 ;
        RECT 520.950 469.950 523.050 472.050 ;
        RECT 517.950 448.950 520.050 451.050 ;
        RECT 514.950 442.950 517.050 445.050 ;
        RECT 515.400 418.050 516.450 442.950 ;
        RECT 521.400 421.050 522.450 469.950 ;
        RECT 524.400 457.050 525.450 484.950 ;
        RECT 527.400 475.050 528.450 487.950 ;
        RECT 529.950 484.950 532.050 487.050 ;
        RECT 538.950 484.950 541.050 487.050 ;
        RECT 544.950 484.950 547.050 487.050 ;
        RECT 548.250 485.250 550.050 486.150 ;
        RECT 554.400 484.050 555.450 508.950 ;
        RECT 529.950 481.950 532.050 484.050 ;
        RECT 538.950 482.850 541.050 483.750 ;
        RECT 541.950 482.250 544.050 483.150 ;
        RECT 544.950 482.850 546.750 483.750 ;
        RECT 547.950 481.950 550.050 484.050 ;
        RECT 553.950 481.950 556.050 484.050 ;
        RECT 526.950 472.950 529.050 475.050 ;
        RECT 530.400 471.450 531.450 481.950 ;
        RECT 532.950 478.950 535.050 481.050 ;
        RECT 541.950 478.950 544.050 481.050 ;
        RECT 553.950 478.950 556.050 481.050 ;
        RECT 527.400 470.400 531.450 471.450 ;
        RECT 527.400 457.050 528.450 470.400 ;
        RECT 533.400 457.050 534.450 478.950 ;
        RECT 542.400 475.050 543.450 478.950 ;
        RECT 541.950 472.950 544.050 475.050 ;
        RECT 554.400 469.050 555.450 478.950 ;
        RECT 553.950 466.950 556.050 469.050 ;
        RECT 547.950 457.950 550.050 460.050 ;
        RECT 548.400 457.050 549.450 457.950 ;
        RECT 554.400 457.050 555.450 466.950 ;
        RECT 523.950 454.950 526.050 457.050 ;
        RECT 526.950 454.950 529.050 457.050 ;
        RECT 530.250 455.250 531.750 456.150 ;
        RECT 532.950 454.950 535.050 457.050 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 547.950 454.950 550.050 457.050 ;
        RECT 551.250 455.250 552.750 456.150 ;
        RECT 553.950 454.950 556.050 457.050 ;
        RECT 524.400 454.050 525.450 454.950 ;
        RECT 545.400 454.050 546.450 454.950 ;
        RECT 523.950 451.950 526.050 454.050 ;
        RECT 527.250 452.850 528.750 453.750 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 533.250 452.850 535.050 453.750 ;
        RECT 544.950 451.950 547.050 454.050 ;
        RECT 548.250 452.850 549.750 453.750 ;
        RECT 550.950 451.950 553.050 454.050 ;
        RECT 554.250 452.850 556.050 453.750 ;
        RECT 530.400 451.050 531.450 451.950 ;
        RECT 551.400 451.050 552.450 451.950 ;
        RECT 523.950 449.850 526.050 450.750 ;
        RECT 526.950 448.950 529.050 451.050 ;
        RECT 529.950 448.950 532.050 451.050 ;
        RECT 544.950 449.850 547.050 450.750 ;
        RECT 550.950 448.950 553.050 451.050 ;
        RECT 527.400 423.450 528.450 448.950 ;
        RECT 557.400 427.050 558.450 559.950 ;
        RECT 559.950 556.950 562.050 559.050 ;
        RECT 560.400 550.050 561.450 556.950 ;
        RECT 559.950 547.950 562.050 550.050 ;
        RECT 563.400 531.450 564.450 598.950 ;
        RECT 566.400 589.050 567.450 604.950 ;
        RECT 569.400 594.450 570.450 607.950 ;
        RECT 571.950 596.250 573.750 597.150 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 578.250 596.250 580.050 597.150 ;
        RECT 571.950 594.450 574.050 595.050 ;
        RECT 569.400 593.400 574.050 594.450 ;
        RECT 575.250 593.850 576.750 594.750 ;
        RECT 577.950 594.450 580.050 595.050 ;
        RECT 581.400 594.450 582.450 610.950 ;
        RECT 583.950 604.950 586.050 607.050 ;
        RECT 571.950 592.950 574.050 593.400 ;
        RECT 577.950 593.400 582.450 594.450 ;
        RECT 577.950 592.950 580.050 593.400 ;
        RECT 577.950 589.950 580.050 592.050 ;
        RECT 565.950 586.950 568.050 589.050 ;
        RECT 571.950 574.950 574.050 577.050 ;
        RECT 572.400 562.050 573.450 574.950 ;
        RECT 574.950 562.950 577.050 565.050 ;
        RECT 565.950 559.950 568.050 562.050 ;
        RECT 569.250 560.250 570.750 561.150 ;
        RECT 571.950 559.950 574.050 562.050 ;
        RECT 565.950 557.850 567.750 558.750 ;
        RECT 568.950 556.950 571.050 559.050 ;
        RECT 572.250 557.850 574.050 558.750 ;
        RECT 569.400 552.450 570.450 556.950 ;
        RECT 566.400 551.400 570.450 552.450 ;
        RECT 566.400 538.050 567.450 551.400 ;
        RECT 575.400 550.050 576.450 562.950 ;
        RECT 568.950 547.950 571.050 550.050 ;
        RECT 574.950 547.950 577.050 550.050 ;
        RECT 565.950 535.950 568.050 538.050 ;
        RECT 560.400 530.400 564.450 531.450 ;
        RECT 556.950 424.950 559.050 427.050 ;
        RECT 560.400 423.450 561.450 530.400 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 562.950 524.850 565.050 525.750 ;
        RECT 565.950 524.250 568.050 525.150 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 569.400 520.050 570.450 547.950 ;
        RECT 571.950 528.450 574.050 529.050 ;
        RECT 571.950 527.400 576.450 528.450 ;
        RECT 571.950 526.950 574.050 527.400 ;
        RECT 575.400 526.050 576.450 527.400 ;
        RECT 571.950 524.850 574.050 525.750 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 568.950 517.950 571.050 520.050 ;
        RECT 562.950 488.250 565.050 489.150 ;
        RECT 569.400 487.050 570.450 517.950 ;
        RECT 575.400 511.050 576.450 523.950 ;
        RECT 574.950 508.950 577.050 511.050 ;
        RECT 562.950 484.950 565.050 487.050 ;
        RECT 566.250 485.250 567.750 486.150 ;
        RECT 568.950 484.950 571.050 487.050 ;
        RECT 572.250 485.250 574.050 486.150 ;
        RECT 574.950 484.950 577.050 487.050 ;
        RECT 563.400 460.050 564.450 484.950 ;
        RECT 575.400 484.050 576.450 484.950 ;
        RECT 565.950 481.950 568.050 484.050 ;
        RECT 569.250 482.850 570.750 483.750 ;
        RECT 571.950 483.450 574.050 484.050 ;
        RECT 574.950 483.450 577.050 484.050 ;
        RECT 571.950 482.400 577.050 483.450 ;
        RECT 571.950 481.950 574.050 482.400 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 566.400 475.050 567.450 481.950 ;
        RECT 565.950 472.950 568.050 475.050 ;
        RECT 568.950 472.950 571.050 475.050 ;
        RECT 562.950 457.950 565.050 460.050 ;
        RECT 565.950 455.250 568.050 456.150 ;
        RECT 565.950 451.950 568.050 454.050 ;
        RECT 527.400 422.400 531.450 423.450 ;
        RECT 560.400 422.400 564.450 423.450 ;
        RECT 520.950 418.950 523.050 421.050 ;
        RECT 526.950 418.950 529.050 421.050 ;
        RECT 511.950 415.950 514.050 418.050 ;
        RECT 514.950 415.950 517.050 418.050 ;
        RECT 517.950 417.450 520.050 418.050 ;
        RECT 517.950 416.400 522.450 417.450 ;
        RECT 517.950 415.950 520.050 416.400 ;
        RECT 514.950 413.250 517.050 414.150 ;
        RECT 517.950 413.850 520.050 414.750 ;
        RECT 514.950 409.950 517.050 412.050 ;
        RECT 511.950 406.950 514.050 409.050 ;
        RECT 508.950 400.950 511.050 403.050 ;
        RECT 499.950 397.950 502.050 400.050 ;
        RECT 505.950 397.950 508.050 400.050 ;
        RECT 500.400 373.050 501.450 397.950 ;
        RECT 505.950 382.950 508.050 385.050 ;
        RECT 506.400 382.050 507.450 382.950 ;
        RECT 512.400 382.050 513.450 406.950 ;
        RECT 517.950 403.950 520.050 406.050 ;
        RECT 502.950 380.250 504.750 381.150 ;
        RECT 505.950 379.950 508.050 382.050 ;
        RECT 511.950 379.950 514.050 382.050 ;
        RECT 502.950 376.950 505.050 379.050 ;
        RECT 506.250 377.850 507.750 378.750 ;
        RECT 508.950 376.950 511.050 379.050 ;
        RECT 512.250 377.850 514.050 378.750 ;
        RECT 514.950 376.950 517.050 379.050 ;
        RECT 502.950 373.950 505.050 376.050 ;
        RECT 508.950 374.850 511.050 375.750 ;
        RECT 499.950 370.950 502.050 373.050 ;
        RECT 499.950 352.950 502.050 355.050 ;
        RECT 487.950 343.950 490.050 346.050 ;
        RECT 490.950 345.450 493.050 346.050 ;
        RECT 493.950 345.450 496.050 346.050 ;
        RECT 490.950 344.400 496.050 345.450 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 493.950 343.950 496.050 344.400 ;
        RECT 496.950 343.950 499.050 346.050 ;
        RECT 500.400 343.050 501.450 352.950 ;
        RECT 490.950 341.250 492.750 342.150 ;
        RECT 499.950 340.950 502.050 343.050 ;
        RECT 490.950 337.950 493.050 340.050 ;
        RECT 494.250 338.850 496.050 339.750 ;
        RECT 496.950 338.250 499.050 339.150 ;
        RECT 499.950 338.850 502.050 339.750 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 497.400 334.050 498.450 334.950 ;
        RECT 496.950 331.950 499.050 334.050 ;
        RECT 503.400 328.050 504.450 373.950 ;
        RECT 515.400 370.050 516.450 376.950 ;
        RECT 514.950 367.950 517.050 370.050 ;
        RECT 508.950 364.950 511.050 367.050 ;
        RECT 505.950 352.950 508.050 355.050 ;
        RECT 506.400 349.050 507.450 352.950 ;
        RECT 505.950 346.950 508.050 349.050 ;
        RECT 509.400 346.050 510.450 364.950 ;
        RECT 518.400 358.050 519.450 403.950 ;
        RECT 521.400 403.050 522.450 416.400 ;
        RECT 523.950 413.250 526.050 414.150 ;
        RECT 527.400 412.050 528.450 418.950 ;
        RECT 523.950 411.450 526.050 412.050 ;
        RECT 526.950 411.450 529.050 412.050 ;
        RECT 523.950 410.400 529.050 411.450 ;
        RECT 523.950 409.950 526.050 410.400 ;
        RECT 526.950 409.950 529.050 410.400 ;
        RECT 523.950 406.950 526.050 409.050 ;
        RECT 520.950 400.950 523.050 403.050 ;
        RECT 520.950 397.950 523.050 400.050 ;
        RECT 521.400 385.050 522.450 397.950 ;
        RECT 520.950 382.950 523.050 385.050 ;
        RECT 520.950 380.850 523.050 381.750 ;
        RECT 520.950 370.950 523.050 373.050 ;
        RECT 517.950 355.950 520.050 358.050 ;
        RECT 517.950 352.950 520.050 355.050 ;
        RECT 505.950 343.950 508.050 346.050 ;
        RECT 508.950 343.950 511.050 346.050 ;
        RECT 502.950 325.950 505.050 328.050 ;
        RECT 496.950 316.950 499.050 319.050 ;
        RECT 490.950 313.950 493.050 316.050 ;
        RECT 491.250 311.850 492.750 312.750 ;
        RECT 484.950 307.950 487.050 310.050 ;
        RECT 487.950 308.850 490.050 309.750 ;
        RECT 490.950 307.950 493.050 310.050 ;
        RECT 493.950 308.850 496.050 309.750 ;
        RECT 472.950 305.400 477.450 306.450 ;
        RECT 472.950 304.950 475.050 305.400 ;
        RECT 478.950 304.950 481.050 307.050 ;
        RECT 467.400 274.050 468.450 304.950 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 472.950 280.950 475.050 283.050 ;
        RECT 463.950 271.950 466.050 274.050 ;
        RECT 466.950 271.950 469.050 274.050 ;
        RECT 463.950 269.250 466.050 270.150 ;
        RECT 469.950 269.250 472.050 270.150 ;
        RECT 467.250 266.250 468.750 267.150 ;
        RECT 469.950 265.950 472.050 268.050 ;
        RECT 461.400 263.400 465.450 264.450 ;
        RECT 460.950 259.950 463.050 262.050 ;
        RECT 454.950 241.950 457.050 244.050 ;
        RECT 457.950 241.950 460.050 244.050 ;
        RECT 455.400 241.050 456.450 241.950 ;
        RECT 448.950 238.950 451.050 241.050 ;
        RECT 452.250 239.250 453.750 240.150 ;
        RECT 454.950 238.950 457.050 241.050 ;
        RECT 461.400 240.450 462.450 259.950 ;
        RECT 458.400 239.400 462.450 240.450 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 449.250 236.850 450.750 237.750 ;
        RECT 451.950 235.950 454.050 238.050 ;
        RECT 455.250 236.850 457.050 237.750 ;
        RECT 445.950 233.850 448.050 234.750 ;
        RECT 445.950 229.950 448.050 232.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 430.950 208.950 433.050 211.050 ;
        RECT 427.950 205.950 430.050 208.050 ;
        RECT 436.950 205.950 439.050 208.050 ;
        RECT 437.400 205.050 438.450 205.950 ;
        RECT 427.950 202.950 430.050 205.050 ;
        RECT 436.950 202.950 439.050 205.050 ;
        RECT 421.950 193.950 424.050 196.050 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 428.400 193.050 429.450 202.950 ;
        RECT 430.950 200.250 433.050 201.150 ;
        RECT 437.400 199.050 438.450 202.950 ;
        RECT 430.950 196.950 433.050 199.050 ;
        RECT 434.250 197.250 435.750 198.150 ;
        RECT 436.950 196.950 439.050 199.050 ;
        RECT 440.250 197.250 442.050 198.150 ;
        RECT 446.400 196.050 447.450 229.950 ;
        RECT 452.400 229.050 453.450 235.950 ;
        RECT 451.950 226.950 454.050 229.050 ;
        RECT 454.950 205.950 457.050 208.050 ;
        RECT 448.950 202.950 451.050 205.050 ;
        RECT 433.950 193.950 436.050 196.050 ;
        RECT 437.250 194.850 438.750 195.750 ;
        RECT 439.950 193.950 442.050 196.050 ;
        RECT 445.950 193.950 448.050 196.050 ;
        RECT 424.950 190.950 427.050 193.050 ;
        RECT 427.950 190.950 430.050 193.050 ;
        RECT 418.950 181.950 421.050 184.050 ;
        RECT 425.400 172.050 426.450 190.950 ;
        RECT 424.950 169.950 427.050 172.050 ;
        RECT 440.400 171.450 441.450 193.950 ;
        RECT 449.400 180.450 450.450 202.950 ;
        RECT 455.400 201.450 456.450 205.950 ;
        RECT 458.400 205.050 459.450 239.400 ;
        RECT 460.950 236.250 463.050 237.150 ;
        RECT 460.950 234.450 463.050 235.050 ;
        RECT 464.400 234.450 465.450 263.400 ;
        RECT 466.950 262.950 469.050 265.050 ;
        RECT 470.400 252.450 471.450 265.950 ;
        RECT 467.400 251.400 471.450 252.450 ;
        RECT 467.400 241.050 468.450 251.400 ;
        RECT 473.400 249.450 474.450 280.950 ;
        RECT 476.400 259.050 477.450 289.950 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 479.400 253.050 480.450 304.950 ;
        RECT 487.950 295.950 490.050 298.050 ;
        RECT 485.250 269.250 487.050 270.150 ;
        RECT 481.950 266.850 483.750 267.750 ;
        RECT 484.950 265.950 487.050 268.050 ;
        RECT 478.950 250.950 481.050 253.050 ;
        RECT 485.400 250.050 486.450 265.950 ;
        RECT 488.400 259.050 489.450 295.950 ;
        RECT 491.400 271.050 492.450 307.950 ;
        RECT 497.400 307.050 498.450 316.950 ;
        RECT 502.950 313.950 505.050 316.050 ;
        RECT 496.950 304.950 499.050 307.050 ;
        RECT 496.950 271.950 499.050 274.050 ;
        RECT 490.950 268.950 493.050 271.050 ;
        RECT 494.250 269.250 496.050 270.150 ;
        RECT 490.950 266.850 492.750 267.750 ;
        RECT 493.950 265.950 496.050 268.050 ;
        RECT 494.400 262.050 495.450 265.950 ;
        RECT 493.950 259.950 496.050 262.050 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 497.400 253.050 498.450 271.950 ;
        RECT 503.400 268.050 504.450 313.950 ;
        RECT 506.400 277.050 507.450 343.950 ;
        RECT 508.950 341.250 511.050 342.150 ;
        RECT 514.950 341.250 517.050 342.150 ;
        RECT 508.950 337.950 511.050 340.050 ;
        RECT 514.950 339.450 517.050 340.050 ;
        RECT 518.400 339.450 519.450 352.950 ;
        RECT 521.400 349.050 522.450 370.950 ;
        RECT 520.950 346.950 523.050 349.050 ;
        RECT 512.250 338.250 513.750 339.150 ;
        RECT 514.950 338.400 519.450 339.450 ;
        RECT 514.950 337.950 517.050 338.400 ;
        RECT 509.400 334.050 510.450 337.950 ;
        RECT 511.950 334.950 514.050 337.050 ;
        RECT 508.950 331.950 511.050 334.050 ;
        RECT 512.400 328.050 513.450 334.950 ;
        RECT 508.950 325.950 511.050 328.050 ;
        RECT 511.950 325.950 514.050 328.050 ;
        RECT 509.400 313.050 510.450 325.950 ;
        RECT 514.950 322.950 517.050 325.050 ;
        RECT 508.950 310.950 511.050 313.050 ;
        RECT 508.950 308.850 511.050 309.750 ;
        RECT 511.950 308.250 514.050 309.150 ;
        RECT 511.950 304.950 514.050 307.050 ;
        RECT 505.950 274.950 508.050 277.050 ;
        RECT 512.400 274.050 513.450 304.950 ;
        RECT 505.950 271.950 508.050 274.050 ;
        RECT 511.950 271.950 514.050 274.050 ;
        RECT 502.950 265.950 505.050 268.050 ;
        RECT 496.950 250.950 499.050 253.050 ;
        RECT 470.400 248.400 474.450 249.450 ;
        RECT 466.950 238.950 469.050 241.050 ;
        RECT 460.950 233.400 465.450 234.450 ;
        RECT 466.950 233.850 469.050 234.750 ;
        RECT 460.950 232.950 463.050 233.400 ;
        RECT 466.950 229.950 469.050 232.050 ;
        RECT 467.400 211.050 468.450 229.950 ;
        RECT 470.400 229.050 471.450 248.400 ;
        RECT 481.950 247.950 484.050 250.050 ;
        RECT 484.950 247.950 487.050 250.050 ;
        RECT 472.950 244.950 475.050 247.050 ;
        RECT 475.950 244.950 478.050 247.050 ;
        RECT 478.950 244.950 481.050 247.050 ;
        RECT 469.950 226.950 472.050 229.050 ;
        RECT 473.550 226.050 474.750 244.950 ;
        RECT 476.550 232.350 477.750 244.950 ;
        RECT 475.950 230.250 478.050 232.350 ;
        RECT 476.550 226.050 477.750 230.250 ;
        RECT 479.550 226.050 480.750 244.950 ;
        RECT 472.950 223.950 475.050 226.050 ;
        RECT 475.950 223.950 478.050 226.050 ;
        RECT 478.950 223.950 481.050 226.050 ;
        RECT 482.400 213.450 483.450 247.950 ;
        RECT 484.950 244.950 487.050 247.050 ;
        RECT 487.950 245.400 490.050 247.500 ;
        RECT 492.150 245.400 494.250 247.500 ;
        RECT 496.950 245.400 499.050 247.500 ;
        RECT 499.950 245.400 502.050 247.500 ;
        RECT 502.950 245.400 505.050 247.500 ;
        RECT 485.400 244.050 486.450 244.950 ;
        RECT 484.950 241.950 487.050 244.050 ;
        RECT 484.950 239.850 487.050 240.750 ;
        RECT 488.250 236.850 489.450 245.400 ;
        RECT 492.450 239.550 493.650 245.400 ;
        RECT 492.150 237.450 494.250 239.550 ;
        RECT 487.950 234.750 490.050 236.850 ;
        RECT 488.250 228.600 489.450 234.750 ;
        RECT 492.450 228.600 493.650 237.450 ;
        RECT 497.400 231.750 498.600 245.400 ;
        RECT 496.950 229.650 499.050 231.750 ;
        RECT 487.950 226.500 490.050 228.600 ;
        RECT 492.000 226.500 494.100 228.600 ;
        RECT 500.550 228.150 501.750 245.400 ;
        RECT 503.250 231.750 504.450 245.400 ;
        RECT 502.950 229.650 505.050 231.750 ;
        RECT 499.950 226.050 502.050 228.150 ;
        RECT 503.250 225.900 504.450 229.650 ;
        RECT 506.400 228.450 507.450 271.950 ;
        RECT 508.950 268.950 511.050 271.050 ;
        RECT 508.950 266.850 511.050 267.750 ;
        RECT 511.950 266.250 514.050 267.150 ;
        RECT 508.950 262.950 511.050 265.050 ;
        RECT 511.950 262.950 514.050 265.050 ;
        RECT 509.400 231.450 510.450 262.950 ;
        RECT 512.400 256.050 513.450 262.950 ;
        RECT 511.950 253.950 514.050 256.050 ;
        RECT 511.950 237.450 514.050 238.050 ;
        RECT 515.400 237.450 516.450 322.950 ;
        RECT 521.400 319.050 522.450 346.950 ;
        RECT 524.400 340.050 525.450 406.950 ;
        RECT 530.400 400.050 531.450 422.400 ;
        RECT 547.950 418.950 550.050 421.050 ;
        RECT 553.950 419.250 556.050 420.150 ;
        RECT 559.950 418.950 562.050 421.050 ;
        RECT 532.950 413.250 535.050 414.150 ;
        RECT 538.950 413.250 541.050 414.150 ;
        RECT 532.950 409.950 535.050 412.050 ;
        RECT 536.250 410.250 537.750 411.150 ;
        RECT 538.950 409.950 541.050 412.050 ;
        RECT 533.400 403.050 534.450 409.950 ;
        RECT 535.950 406.950 538.050 409.050 ;
        RECT 538.950 403.950 541.050 406.050 ;
        RECT 532.950 400.950 535.050 403.050 ;
        RECT 529.950 397.950 532.050 400.050 ;
        RECT 535.950 397.950 538.050 400.050 ;
        RECT 529.950 384.450 532.050 385.050 ;
        RECT 529.950 383.400 534.450 384.450 ;
        RECT 529.950 382.950 532.050 383.400 ;
        RECT 526.950 380.250 529.050 381.150 ;
        RECT 529.950 380.850 532.050 381.750 ;
        RECT 526.950 376.950 529.050 379.050 ;
        RECT 527.400 376.050 528.450 376.950 ;
        RECT 526.950 373.950 529.050 376.050 ;
        RECT 526.950 355.950 529.050 358.050 ;
        RECT 523.950 337.950 526.050 340.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 520.950 316.950 523.050 319.050 ;
        RECT 517.950 310.950 520.050 313.050 ;
        RECT 517.950 308.850 520.050 309.750 ;
        RECT 517.950 295.950 520.050 298.050 ;
        RECT 511.950 236.400 516.450 237.450 ;
        RECT 511.950 235.950 514.050 236.400 ;
        RECT 511.950 233.850 514.050 234.750 ;
        RECT 514.950 232.950 517.050 235.050 ;
        RECT 509.400 230.400 513.450 231.450 ;
        RECT 506.400 227.400 510.450 228.450 ;
        RECT 503.100 223.800 505.200 225.900 ;
        RECT 487.950 220.950 490.050 223.050 ;
        RECT 490.950 220.950 493.050 223.050 ;
        RECT 482.400 212.400 486.450 213.450 ;
        RECT 466.950 208.950 469.050 211.050 ;
        RECT 457.950 202.950 460.050 205.050 ;
        RECT 478.950 202.950 481.050 205.050 ;
        RECT 451.950 200.250 454.050 201.150 ;
        RECT 455.400 200.400 459.450 201.450 ;
        RECT 458.400 199.050 459.450 200.400 ;
        RECT 472.950 200.250 475.050 201.150 ;
        RECT 479.400 199.050 480.450 202.950 ;
        RECT 451.950 196.950 454.050 199.050 ;
        RECT 455.250 197.250 456.750 198.150 ;
        RECT 457.950 196.950 460.050 199.050 ;
        RECT 461.250 197.250 463.050 198.150 ;
        RECT 472.950 196.950 475.050 199.050 ;
        RECT 476.250 197.250 477.750 198.150 ;
        RECT 478.950 196.950 481.050 199.050 ;
        RECT 482.250 197.250 484.050 198.150 ;
        RECT 454.950 193.950 457.050 196.050 ;
        RECT 458.250 194.850 459.750 195.750 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 469.950 193.950 472.050 196.050 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 479.250 194.850 480.750 195.750 ;
        RECT 454.950 190.950 457.050 193.050 ;
        RECT 446.400 179.400 453.450 180.450 ;
        RECT 437.400 170.400 441.450 171.450 ;
        RECT 425.250 167.850 426.750 168.750 ;
        RECT 427.950 168.450 430.050 169.050 ;
        RECT 427.950 167.400 432.450 168.450 ;
        RECT 427.950 166.950 430.050 167.400 ;
        RECT 415.950 163.950 418.050 166.050 ;
        RECT 421.950 164.850 424.050 165.750 ;
        RECT 427.950 164.850 430.050 165.750 ;
        RECT 431.400 157.050 432.450 167.400 ;
        RECT 433.950 166.950 436.050 169.050 ;
        RECT 430.950 154.950 433.050 157.050 ;
        RECT 434.400 130.050 435.450 166.950 ;
        RECT 437.400 148.050 438.450 170.400 ;
        RECT 442.950 169.950 445.050 172.050 ;
        RECT 446.400 169.050 447.450 179.400 ;
        RECT 439.950 166.950 442.050 169.050 ;
        RECT 443.250 167.850 444.750 168.750 ;
        RECT 445.950 166.950 448.050 169.050 ;
        RECT 439.950 164.850 442.050 165.750 ;
        RECT 445.950 164.850 448.050 165.750 ;
        RECT 445.950 160.950 448.050 163.050 ;
        RECT 436.950 145.950 439.050 148.050 ;
        RECT 446.400 142.050 447.450 160.950 ;
        RECT 445.950 139.950 448.050 142.050 ;
        RECT 439.950 130.950 442.050 133.050 ;
        RECT 440.400 130.050 441.450 130.950 ;
        RECT 412.950 129.450 415.050 130.050 ;
        RECT 410.400 128.400 415.050 129.450 ;
        RECT 418.950 129.450 421.050 130.050 ;
        RECT 400.950 125.250 403.050 126.150 ;
        RECT 410.400 124.050 411.450 128.400 ;
        RECT 412.950 127.950 415.050 128.400 ;
        RECT 416.250 128.250 417.750 129.150 ;
        RECT 418.950 128.400 423.450 129.450 ;
        RECT 418.950 127.950 421.050 128.400 ;
        RECT 412.950 125.850 414.750 126.750 ;
        RECT 415.950 124.950 418.050 127.050 ;
        RECT 419.250 125.850 421.050 126.750 ;
        RECT 400.950 121.950 403.050 124.050 ;
        RECT 404.250 122.250 406.050 123.150 ;
        RECT 409.950 121.950 412.050 124.050 ;
        RECT 403.950 118.950 406.050 121.050 ;
        RECT 404.400 118.050 405.450 118.950 ;
        RECT 422.400 118.050 423.450 128.400 ;
        RECT 427.950 127.950 430.050 130.050 ;
        RECT 433.950 127.950 436.050 130.050 ;
        RECT 437.250 128.250 438.750 129.150 ;
        RECT 439.950 127.950 442.050 130.050 ;
        RECT 403.950 115.950 406.050 118.050 ;
        RECT 421.950 115.950 424.050 118.050 ;
        RECT 397.950 112.950 400.050 115.050 ;
        RECT 409.950 97.950 412.050 100.050 ;
        RECT 428.400 97.050 429.450 127.950 ;
        RECT 452.400 127.050 453.450 179.400 ;
        RECT 455.400 127.050 456.450 190.950 ;
        RECT 457.950 169.950 460.050 172.050 ;
        RECT 458.400 169.050 459.450 169.950 ;
        RECT 461.400 169.050 462.450 193.950 ;
        RECT 457.950 166.950 460.050 169.050 ;
        RECT 460.950 166.950 463.050 169.050 ;
        RECT 466.950 166.950 469.050 169.050 ;
        RECT 457.950 164.850 460.050 165.750 ;
        RECT 463.950 164.250 466.050 165.150 ;
        RECT 466.950 164.850 469.050 165.750 ;
        RECT 463.950 160.950 466.050 163.050 ;
        RECT 470.400 160.050 471.450 193.950 ;
        RECT 476.400 184.050 477.450 193.950 ;
        RECT 478.950 184.950 481.050 187.050 ;
        RECT 475.950 181.950 478.050 184.050 ;
        RECT 472.950 172.950 475.050 175.050 ;
        RECT 473.400 163.050 474.450 172.950 ;
        RECT 472.950 160.950 475.050 163.050 ;
        RECT 469.950 157.950 472.050 160.050 ;
        RECT 466.950 130.950 469.050 133.050 ;
        RECT 433.950 125.850 435.750 126.750 ;
        RECT 436.950 124.950 439.050 127.050 ;
        RECT 440.250 125.850 442.050 126.750 ;
        RECT 451.950 124.950 454.050 127.050 ;
        RECT 454.950 124.950 457.050 127.050 ;
        RECT 457.950 124.950 460.050 127.050 ;
        RECT 430.950 97.950 433.050 100.050 ;
        RECT 406.950 96.450 409.050 97.050 ;
        RECT 404.400 95.400 409.050 96.450 ;
        RECT 410.250 95.850 411.750 96.750 ;
        RECT 412.950 96.450 415.050 97.050 ;
        RECT 421.950 96.450 424.050 97.050 ;
        RECT 388.950 92.250 390.750 93.150 ;
        RECT 391.950 91.950 394.050 94.050 ;
        RECT 395.250 92.250 397.050 93.150 ;
        RECT 388.950 88.950 391.050 91.050 ;
        RECT 392.250 89.850 393.750 90.750 ;
        RECT 394.950 88.950 397.050 91.050 ;
        RECT 389.400 82.050 390.450 88.950 ;
        RECT 388.950 79.950 391.050 82.050 ;
        RECT 395.400 79.050 396.450 88.950 ;
        RECT 404.400 82.050 405.450 95.400 ;
        RECT 406.950 94.950 409.050 95.400 ;
        RECT 412.950 95.400 417.450 96.450 ;
        RECT 412.950 94.950 415.050 95.400 ;
        RECT 406.950 92.850 409.050 93.750 ;
        RECT 409.950 91.950 412.050 94.050 ;
        RECT 412.950 92.850 415.050 93.750 ;
        RECT 403.950 79.950 406.050 82.050 ;
        RECT 394.950 76.950 397.050 79.050 ;
        RECT 388.950 64.950 391.050 67.050 ;
        RECT 379.950 61.950 382.050 64.050 ;
        RECT 382.950 59.250 385.050 60.150 ;
        RECT 376.950 57.450 379.050 58.050 ;
        RECT 374.400 56.400 379.050 57.450 ;
        RECT 361.950 50.850 364.050 51.750 ;
        RECT 364.950 50.250 367.050 51.150 ;
        RECT 367.950 49.950 370.050 52.050 ;
        RECT 346.950 46.950 349.050 49.050 ;
        RECT 352.950 46.950 355.050 49.050 ;
        RECT 364.950 46.950 367.050 49.050 ;
        RECT 355.950 43.950 358.050 46.050 ;
        RECT 337.950 25.950 340.050 28.050 ;
        RECT 331.950 23.400 336.450 24.450 ;
        RECT 331.950 22.950 334.050 23.400 ;
        RECT 349.950 22.950 352.050 25.050 ;
        RECT 322.950 20.400 327.450 21.450 ;
        RECT 331.950 20.850 334.050 21.750 ;
        RECT 337.950 20.850 340.050 21.750 ;
        RECT 322.950 19.950 325.050 20.400 ;
        RECT 271.950 18.450 274.050 19.050 ;
        RECT 269.400 17.400 274.050 18.450 ;
        RECT 275.250 17.850 276.750 18.750 ;
        RECT 271.950 16.950 274.050 17.400 ;
        RECT 277.950 16.950 280.050 19.050 ;
        RECT 286.950 17.850 288.750 18.750 ;
        RECT 289.950 16.950 292.050 19.050 ;
        RECT 293.250 17.850 294.750 18.750 ;
        RECT 295.950 16.950 298.050 19.050 ;
        RECT 310.950 16.950 313.050 19.050 ;
        RECT 313.950 16.950 316.050 19.050 ;
        RECT 317.250 17.850 318.750 18.750 ;
        RECT 319.950 16.950 322.050 19.050 ;
        RECT 323.250 17.850 325.050 18.750 ;
        RECT 350.400 18.450 351.450 22.950 ;
        RECT 356.400 22.050 357.450 43.950 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 374.400 24.450 375.450 56.400 ;
        RECT 376.950 55.950 379.050 56.400 ;
        RECT 380.250 56.250 381.750 57.150 ;
        RECT 382.950 55.950 385.050 58.050 ;
        RECT 386.250 56.250 388.050 57.150 ;
        RECT 376.950 53.850 378.750 54.750 ;
        RECT 379.950 52.950 382.050 55.050 ;
        RECT 385.950 54.450 388.050 55.050 ;
        RECT 389.400 54.450 390.450 64.950 ;
        RECT 395.400 61.050 396.450 76.950 ;
        RECT 397.950 67.950 400.050 70.050 ;
        RECT 394.950 58.950 397.050 61.050 ;
        RECT 398.400 55.050 399.450 67.950 ;
        RECT 406.950 58.950 409.050 61.050 ;
        RECT 403.950 56.250 406.050 57.150 ;
        RECT 385.950 53.400 390.450 54.450 ;
        RECT 385.950 52.950 388.050 53.400 ;
        RECT 394.950 53.250 396.750 54.150 ;
        RECT 397.950 52.950 400.050 55.050 ;
        RECT 401.250 53.250 402.750 54.150 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 386.400 49.050 387.450 52.950 ;
        RECT 404.400 52.050 405.450 52.950 ;
        RECT 394.950 49.950 397.050 52.050 ;
        RECT 398.250 50.850 399.750 51.750 ;
        RECT 400.950 49.950 403.050 52.050 ;
        RECT 403.950 49.950 406.050 52.050 ;
        RECT 385.950 46.950 388.050 49.050 ;
        RECT 395.400 46.050 396.450 49.950 ;
        RECT 394.950 43.950 397.050 46.050 ;
        RECT 407.400 31.050 408.450 58.950 ;
        RECT 410.400 55.050 411.450 91.950 ;
        RECT 416.400 79.050 417.450 95.400 ;
        RECT 419.400 95.400 424.050 96.450 ;
        RECT 419.400 88.050 420.450 95.400 ;
        RECT 421.950 94.950 424.050 95.400 ;
        RECT 425.250 95.250 426.750 96.150 ;
        RECT 427.950 94.950 430.050 97.050 ;
        RECT 431.400 94.050 432.450 97.950 ;
        RECT 421.950 92.850 423.750 93.750 ;
        RECT 424.950 91.950 427.050 94.050 ;
        RECT 428.250 92.850 429.750 93.750 ;
        RECT 430.950 91.950 433.050 94.050 ;
        RECT 430.950 89.850 433.050 90.750 ;
        RECT 418.950 85.950 421.050 88.050 ;
        RECT 415.950 76.950 418.050 79.050 ;
        RECT 418.950 76.950 421.050 79.050 ;
        RECT 419.400 55.050 420.450 76.950 ;
        RECT 437.400 70.050 438.450 124.950 ;
        RECT 451.950 122.250 454.050 123.150 ;
        RECT 454.950 122.850 457.050 123.750 ;
        RECT 451.950 118.950 454.050 121.050 ;
        RECT 452.400 117.450 453.450 118.950 ;
        RECT 449.400 116.400 453.450 117.450 ;
        RECT 449.400 94.050 450.450 116.400 ;
        RECT 454.950 94.950 457.050 97.050 ;
        RECT 445.950 92.250 447.750 93.150 ;
        RECT 448.950 91.950 451.050 94.050 ;
        RECT 452.250 92.250 454.050 93.150 ;
        RECT 445.950 88.950 448.050 91.050 ;
        RECT 449.250 89.850 450.750 90.750 ;
        RECT 451.950 88.950 454.050 91.050 ;
        RECT 445.950 79.950 448.050 82.050 ;
        RECT 436.950 67.950 439.050 70.050 ;
        RECT 424.950 61.950 427.050 64.050 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 418.950 52.950 421.050 55.050 ;
        RECT 412.950 49.950 415.050 52.050 ;
        RECT 418.950 50.850 421.050 51.750 ;
        RECT 421.950 50.250 424.050 51.150 ;
        RECT 376.950 28.950 379.050 31.050 ;
        RECT 406.950 28.950 409.050 31.050 ;
        RECT 377.400 25.050 378.450 28.950 ;
        RECT 397.950 25.950 400.050 28.050 ;
        RECT 371.400 23.400 375.450 24.450 ;
        RECT 352.950 20.250 354.750 21.150 ;
        RECT 355.950 19.950 358.050 22.050 ;
        RECT 359.250 20.250 361.050 21.150 ;
        RECT 367.950 20.850 370.050 21.750 ;
        RECT 371.400 19.050 372.450 23.400 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 395.250 23.250 397.050 24.150 ;
        RECT 397.950 23.850 400.050 24.750 ;
        RECT 400.950 23.250 403.050 24.150 ;
        RECT 407.400 22.050 408.450 28.950 ;
        RECT 413.400 25.050 414.450 49.950 ;
        RECT 425.400 49.050 426.450 61.950 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 431.400 52.050 432.450 55.950 ;
        RECT 433.950 53.250 436.050 54.150 ;
        RECT 439.950 53.250 442.050 54.150 ;
        RECT 430.950 49.950 433.050 52.050 ;
        RECT 433.950 49.950 436.050 52.050 ;
        RECT 437.250 50.250 438.750 51.150 ;
        RECT 439.950 49.950 442.050 52.050 ;
        RECT 434.400 49.050 435.450 49.950 ;
        RECT 421.950 48.450 424.050 49.050 ;
        RECT 424.950 48.450 427.050 49.050 ;
        RECT 421.950 47.400 427.050 48.450 ;
        RECT 421.950 46.950 424.050 47.400 ;
        RECT 424.950 46.950 427.050 47.400 ;
        RECT 433.950 46.950 436.050 49.050 ;
        RECT 436.950 46.950 439.050 49.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 421.950 24.450 424.050 25.050 ;
        RECT 421.950 23.400 426.450 24.450 ;
        RECT 421.950 22.950 424.050 23.400 ;
        RECT 425.400 22.050 426.450 23.400 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 437.400 22.050 438.450 22.950 ;
        RECT 373.950 20.250 376.050 21.150 ;
        RECT 376.950 20.850 379.050 21.750 ;
        RECT 391.950 20.850 393.750 21.750 ;
        RECT 394.950 19.950 397.050 22.050 ;
        RECT 400.950 19.950 403.050 22.050 ;
        RECT 406.950 19.950 409.050 22.050 ;
        RECT 412.950 20.850 415.050 21.750 ;
        RECT 415.950 20.250 418.050 21.150 ;
        RECT 421.950 20.850 424.050 21.750 ;
        RECT 424.950 19.950 427.050 22.050 ;
        RECT 433.950 20.250 435.750 21.150 ;
        RECT 436.950 19.950 439.050 22.050 ;
        RECT 440.250 20.250 442.050 21.150 ;
        RECT 352.950 18.450 355.050 19.050 ;
        RECT 350.400 17.400 355.050 18.450 ;
        RECT 356.250 17.850 357.750 18.750 ;
        RECT 352.950 16.950 355.050 17.400 ;
        RECT 358.950 16.950 361.050 19.050 ;
        RECT 370.950 18.450 373.050 19.050 ;
        RECT 373.950 18.450 376.050 19.050 ;
        RECT 370.950 17.400 376.050 18.450 ;
        RECT 370.950 16.950 373.050 17.400 ;
        RECT 373.950 16.950 376.050 17.400 ;
        RECT 415.950 16.950 418.050 19.050 ;
        RECT 433.950 16.950 436.050 19.050 ;
        RECT 437.250 17.850 438.750 18.750 ;
        RECT 439.950 16.950 442.050 19.050 ;
        RECT 119.400 16.050 120.450 16.950 ;
        RECT 278.400 16.050 279.450 16.950 ;
        RECT 314.400 16.050 315.450 16.950 ;
        RECT 416.400 16.050 417.450 16.950 ;
        RECT 434.400 16.050 435.450 16.950 ;
        RECT 446.400 16.050 447.450 79.950 ;
        RECT 451.950 52.950 454.050 55.050 ;
        RECT 448.950 50.250 451.050 51.150 ;
        RECT 451.950 50.850 454.050 51.750 ;
        RECT 448.950 46.950 451.050 49.050 ;
        RECT 449.400 19.050 450.450 46.950 ;
        RECT 455.400 28.050 456.450 94.950 ;
        RECT 458.400 61.050 459.450 124.950 ;
        RECT 467.400 121.050 468.450 130.950 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 469.950 122.850 472.050 123.750 ;
        RECT 472.950 122.250 475.050 123.150 ;
        RECT 466.950 118.950 469.050 121.050 ;
        RECT 472.950 118.950 475.050 121.050 ;
        RECT 463.950 97.950 466.050 100.050 ;
        RECT 460.950 95.250 463.050 96.150 ;
        RECT 463.950 95.850 466.050 96.750 ;
        RECT 466.950 95.250 468.750 96.150 ;
        RECT 469.950 94.950 472.050 97.050 ;
        RECT 472.950 94.950 475.050 97.050 ;
        RECT 460.950 91.950 463.050 94.050 ;
        RECT 466.950 91.950 469.050 94.050 ;
        RECT 470.250 92.850 472.050 93.750 ;
        RECT 463.950 85.950 466.050 88.050 ;
        RECT 457.950 58.950 460.050 61.050 ;
        RECT 464.400 51.450 465.450 85.950 ;
        RECT 473.400 82.050 474.450 94.950 ;
        RECT 476.400 94.050 477.450 124.950 ;
        RECT 479.400 100.050 480.450 184.950 ;
        RECT 485.400 172.050 486.450 212.400 ;
        RECT 488.400 172.050 489.450 220.950 ;
        RECT 491.400 193.050 492.450 220.950 ;
        RECT 493.950 208.950 496.050 211.050 ;
        RECT 494.400 199.050 495.450 208.950 ;
        RECT 509.400 199.050 510.450 227.400 ;
        RECT 493.950 196.950 496.050 199.050 ;
        RECT 508.950 196.950 511.050 199.050 ;
        RECT 512.400 196.050 513.450 230.400 ;
        RECT 515.400 226.050 516.450 232.950 ;
        RECT 514.950 223.950 517.050 226.050 ;
        RECT 493.950 194.850 496.050 195.750 ;
        RECT 496.950 194.250 499.050 195.150 ;
        RECT 505.950 194.250 508.050 195.150 ;
        RECT 508.950 194.850 511.050 195.750 ;
        RECT 511.950 193.950 514.050 196.050 ;
        RECT 490.950 190.950 493.050 193.050 ;
        RECT 496.950 190.950 499.050 193.050 ;
        RECT 505.950 190.950 508.050 193.050 ;
        RECT 506.400 187.050 507.450 190.950 ;
        RECT 505.950 184.950 508.050 187.050 ;
        RECT 515.400 181.050 516.450 223.950 ;
        RECT 518.400 220.050 519.450 295.950 ;
        RECT 524.400 289.050 525.450 334.950 ;
        RECT 527.400 331.050 528.450 355.950 ;
        RECT 533.400 343.050 534.450 383.400 ;
        RECT 536.400 373.050 537.450 397.950 ;
        RECT 539.400 375.450 540.450 403.950 ;
        RECT 544.950 400.950 547.050 403.050 ;
        RECT 545.400 382.050 546.450 400.950 ;
        RECT 548.400 385.050 549.450 418.950 ;
        RECT 560.400 418.050 561.450 418.950 ;
        RECT 550.950 416.250 552.750 417.150 ;
        RECT 553.950 415.950 556.050 418.050 ;
        RECT 557.250 416.250 558.750 417.150 ;
        RECT 559.950 415.950 562.050 418.050 ;
        RECT 563.400 415.050 564.450 422.400 ;
        RECT 556.950 412.950 559.050 415.050 ;
        RECT 560.250 413.850 562.050 414.750 ;
        RECT 562.950 412.950 565.050 415.050 ;
        RECT 550.950 406.950 553.050 409.050 ;
        RECT 547.950 382.950 550.050 385.050 ;
        RECT 541.950 380.250 543.750 381.150 ;
        RECT 544.950 379.950 547.050 382.050 ;
        RECT 548.250 380.250 550.050 381.150 ;
        RECT 541.950 376.950 544.050 379.050 ;
        RECT 545.250 377.850 546.750 378.750 ;
        RECT 547.950 376.950 550.050 379.050 ;
        RECT 539.400 374.400 543.450 375.450 ;
        RECT 535.950 370.950 538.050 373.050 ;
        RECT 536.400 346.050 537.450 370.950 ;
        RECT 535.950 343.950 538.050 346.050 ;
        RECT 538.950 344.250 541.050 345.150 ;
        RECT 529.950 341.250 531.750 342.150 ;
        RECT 532.950 340.950 535.050 343.050 ;
        RECT 536.250 341.250 537.750 342.150 ;
        RECT 538.950 340.950 541.050 343.050 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 533.250 338.850 534.750 339.750 ;
        RECT 535.950 337.950 538.050 340.050 ;
        RECT 526.950 328.950 529.050 331.050 ;
        RECT 539.400 328.050 540.450 340.950 ;
        RECT 538.950 325.950 541.050 328.050 ;
        RECT 529.950 313.950 532.050 316.050 ;
        RECT 535.950 313.950 538.050 316.050 ;
        RECT 536.400 313.050 537.450 313.950 ;
        RECT 526.950 311.250 529.050 312.150 ;
        RECT 529.950 311.850 532.050 312.750 ;
        RECT 532.950 311.250 534.750 312.150 ;
        RECT 535.950 310.950 538.050 313.050 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 536.250 308.850 538.050 309.750 ;
        RECT 542.400 307.050 543.450 374.400 ;
        RECT 548.400 373.050 549.450 376.950 ;
        RECT 551.400 376.050 552.450 406.950 ;
        RECT 553.950 400.950 556.050 403.050 ;
        RECT 550.950 373.950 553.050 376.050 ;
        RECT 547.950 370.950 550.050 373.050 ;
        RECT 550.950 358.950 553.050 361.050 ;
        RECT 544.950 355.950 547.050 358.050 ;
        RECT 547.950 355.950 550.050 358.050 ;
        RECT 545.400 340.050 546.450 355.950 ;
        RECT 544.950 337.950 547.050 340.050 ;
        RECT 548.400 337.050 549.450 355.950 ;
        RECT 551.400 346.050 552.450 358.950 ;
        RECT 554.400 358.050 555.450 400.950 ;
        RECT 563.400 388.050 564.450 412.950 ;
        RECT 565.950 409.950 568.050 412.050 ;
        RECT 556.950 385.950 559.050 388.050 ;
        RECT 562.950 385.950 565.050 388.050 ;
        RECT 557.400 384.450 558.450 385.950 ;
        RECT 566.400 385.050 567.450 409.950 ;
        RECT 569.400 406.050 570.450 472.950 ;
        RECT 574.950 457.950 577.050 460.050 ;
        RECT 571.950 454.950 574.050 457.050 ;
        RECT 575.250 455.850 577.050 456.750 ;
        RECT 571.950 452.850 574.050 453.750 ;
        RECT 574.950 451.950 577.050 454.050 ;
        RECT 575.400 450.450 576.450 451.950 ;
        RECT 572.400 449.400 576.450 450.450 ;
        RECT 572.400 442.050 573.450 449.400 ;
        RECT 571.950 439.950 574.050 442.050 ;
        RECT 574.950 433.950 577.050 436.050 ;
        RECT 575.400 420.450 576.450 433.950 ;
        RECT 578.400 424.050 579.450 589.950 ;
        RECT 584.400 574.050 585.450 604.950 ;
        RECT 589.950 598.950 592.050 601.050 ;
        RECT 595.950 598.950 598.050 601.050 ;
        RECT 599.250 599.250 600.750 600.150 ;
        RECT 601.950 598.950 604.050 601.050 ;
        RECT 583.950 571.950 586.050 574.050 ;
        RECT 586.950 565.950 589.050 568.050 ;
        RECT 587.400 559.050 588.450 565.950 ;
        RECT 586.950 556.950 589.050 559.050 ;
        RECT 583.950 554.250 586.050 555.150 ;
        RECT 586.950 554.850 589.050 555.750 ;
        RECT 583.950 550.950 586.050 553.050 ;
        RECT 584.400 547.050 585.450 550.950 ;
        RECT 583.950 544.950 586.050 547.050 ;
        RECT 583.950 541.950 586.050 544.050 ;
        RECT 580.950 538.950 583.050 541.050 ;
        RECT 581.400 529.050 582.450 538.950 ;
        RECT 584.400 532.050 585.450 541.950 ;
        RECT 583.950 529.950 586.050 532.050 ;
        RECT 580.950 526.950 583.050 529.050 ;
        RECT 584.250 527.850 585.750 528.750 ;
        RECT 586.950 526.950 589.050 529.050 ;
        RECT 580.950 524.850 583.050 525.750 ;
        RECT 586.950 524.850 589.050 525.750 ;
        RECT 586.950 505.950 589.050 508.050 ;
        RECT 583.950 484.950 586.050 487.050 ;
        RECT 580.950 482.250 583.050 483.150 ;
        RECT 583.950 482.850 586.050 483.750 ;
        RECT 587.400 481.050 588.450 505.950 ;
        RECT 580.950 478.950 583.050 481.050 ;
        RECT 586.950 478.950 589.050 481.050 ;
        RECT 581.400 463.050 582.450 478.950 ;
        RECT 586.950 475.950 589.050 478.050 ;
        RECT 580.950 460.950 583.050 463.050 ;
        RECT 580.950 454.950 583.050 457.050 ;
        RECT 583.950 454.950 586.050 457.050 ;
        RECT 581.400 448.050 582.450 454.950 ;
        RECT 584.400 451.050 585.450 454.950 ;
        RECT 583.950 448.950 586.050 451.050 ;
        RECT 580.950 445.950 583.050 448.050 ;
        RECT 577.950 421.950 580.050 424.050 ;
        RECT 580.950 421.950 583.050 424.050 ;
        RECT 575.400 419.400 579.450 420.450 ;
        RECT 578.400 418.050 579.450 419.400 ;
        RECT 571.950 415.950 574.050 418.050 ;
        RECT 575.250 416.250 576.750 417.150 ;
        RECT 577.950 415.950 580.050 418.050 ;
        RECT 571.950 413.850 573.750 414.750 ;
        RECT 574.950 412.950 577.050 415.050 ;
        RECT 578.250 413.850 580.050 414.750 ;
        RECT 568.950 403.950 571.050 406.050 ;
        RECT 575.400 397.050 576.450 412.950 ;
        RECT 574.950 394.950 577.050 397.050 ;
        RECT 574.950 391.950 577.050 394.050 ;
        RECT 571.950 385.950 574.050 388.050 ;
        RECT 572.400 385.050 573.450 385.950 ;
        RECT 559.950 384.450 562.050 385.050 ;
        RECT 557.400 383.400 562.050 384.450 ;
        RECT 559.950 382.950 562.050 383.400 ;
        RECT 563.250 383.250 564.750 384.150 ;
        RECT 565.950 382.950 568.050 385.050 ;
        RECT 569.250 383.250 570.750 384.150 ;
        RECT 571.950 382.950 574.050 385.050 ;
        RECT 559.950 380.850 561.750 381.750 ;
        RECT 562.950 379.950 565.050 382.050 ;
        RECT 566.250 380.850 567.750 381.750 ;
        RECT 568.950 379.950 571.050 382.050 ;
        RECT 572.250 380.850 574.050 381.750 ;
        RECT 563.400 379.050 564.450 379.950 ;
        RECT 559.950 376.950 562.050 379.050 ;
        RECT 562.950 376.950 565.050 379.050 ;
        RECT 568.950 376.950 571.050 379.050 ;
        RECT 553.950 355.950 556.050 358.050 ;
        RECT 550.950 343.950 553.050 346.050 ;
        RECT 556.950 345.450 559.050 346.050 ;
        RECT 560.400 345.450 561.450 376.950 ;
        RECT 565.950 370.950 568.050 373.050 ;
        RECT 562.950 352.950 565.050 355.050 ;
        RECT 554.250 344.250 555.750 345.150 ;
        RECT 556.950 344.400 561.450 345.450 ;
        RECT 556.950 343.950 559.050 344.400 ;
        RECT 550.950 341.850 552.750 342.750 ;
        RECT 553.950 340.950 556.050 343.050 ;
        RECT 557.250 341.850 559.050 342.750 ;
        RECT 559.950 340.950 562.050 343.050 ;
        RECT 554.400 340.050 555.450 340.950 ;
        RECT 550.950 337.950 553.050 340.050 ;
        RECT 553.950 337.950 556.050 340.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 547.950 331.950 550.050 334.050 ;
        RECT 544.950 310.950 547.050 313.050 ;
        RECT 541.950 304.950 544.050 307.050 ;
        RECT 538.950 301.950 541.050 304.050 ;
        RECT 523.950 286.950 526.050 289.050 ;
        RECT 529.950 286.950 532.050 289.050 ;
        RECT 524.400 280.050 525.450 286.950 ;
        RECT 523.950 277.950 526.050 280.050 ;
        RECT 530.400 271.050 531.450 286.950 ;
        RECT 535.950 271.950 538.050 274.050 ;
        RECT 520.950 269.250 522.750 270.150 ;
        RECT 523.950 268.950 526.050 271.050 ;
        RECT 527.250 269.250 528.750 270.150 ;
        RECT 529.950 268.950 532.050 271.050 ;
        RECT 533.250 269.250 535.050 270.150 ;
        RECT 520.950 265.950 523.050 268.050 ;
        RECT 524.250 266.850 525.750 267.750 ;
        RECT 526.950 265.950 529.050 268.050 ;
        RECT 530.250 266.850 531.750 267.750 ;
        RECT 532.950 265.950 535.050 268.050 ;
        RECT 521.400 262.050 522.450 265.950 ;
        RECT 520.950 259.950 523.050 262.050 ;
        RECT 520.950 253.950 523.050 256.050 ;
        RECT 521.400 235.050 522.450 253.950 ;
        RECT 523.950 239.250 526.050 240.150 ;
        RECT 523.950 235.950 526.050 238.050 ;
        RECT 520.950 232.950 523.050 235.050 ;
        RECT 520.950 229.950 523.050 232.050 ;
        RECT 517.950 217.950 520.050 220.050 ;
        RECT 517.950 205.950 520.050 208.050 ;
        RECT 518.400 196.050 519.450 205.950 ;
        RECT 517.950 193.950 520.050 196.050 ;
        RECT 517.950 190.950 520.050 193.050 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 505.950 172.950 508.050 175.050 ;
        RECT 506.400 172.050 507.450 172.950 ;
        RECT 484.950 169.950 487.050 172.050 ;
        RECT 487.950 169.950 490.050 172.050 ;
        RECT 505.950 169.950 508.050 172.050 ;
        RECT 508.950 169.950 511.050 172.050 ;
        RECT 514.950 169.950 517.050 172.050 ;
        RECT 509.400 169.050 510.450 169.950 ;
        RECT 485.250 167.850 486.750 168.750 ;
        RECT 487.950 168.450 490.050 169.050 ;
        RECT 487.950 167.400 492.450 168.450 ;
        RECT 487.950 166.950 490.050 167.400 ;
        RECT 481.950 164.850 484.050 165.750 ;
        RECT 484.950 163.950 487.050 166.050 ;
        RECT 487.950 164.850 490.050 165.750 ;
        RECT 478.950 97.950 481.050 100.050 ;
        RECT 485.400 96.450 486.450 163.950 ;
        RECT 491.400 160.050 492.450 167.400 ;
        RECT 496.950 166.950 499.050 169.050 ;
        RECT 502.950 168.450 505.050 169.050 ;
        RECT 500.400 167.400 505.050 168.450 ;
        RECT 506.250 167.850 507.750 168.750 ;
        RECT 490.950 157.950 493.050 160.050 ;
        RECT 487.950 136.950 490.050 139.050 ;
        RECT 488.400 130.050 489.450 136.950 ;
        RECT 487.950 127.950 490.050 130.050 ;
        RECT 491.250 128.250 492.750 129.150 ;
        RECT 493.950 127.950 496.050 130.050 ;
        RECT 487.950 125.850 489.750 126.750 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 494.250 125.850 496.050 126.750 ;
        RECT 491.400 118.050 492.450 124.950 ;
        RECT 490.950 115.950 493.050 118.050 ;
        RECT 497.400 97.050 498.450 166.950 ;
        RECT 500.400 157.050 501.450 167.400 ;
        RECT 502.950 166.950 505.050 167.400 ;
        RECT 508.950 166.950 511.050 169.050 ;
        RECT 502.950 164.850 505.050 165.750 ;
        RECT 508.950 164.850 511.050 165.750 ;
        RECT 499.950 154.950 502.050 157.050 ;
        RECT 500.400 121.050 501.450 154.950 ;
        RECT 515.400 154.050 516.450 169.950 ;
        RECT 514.950 151.950 517.050 154.050 ;
        RECT 508.950 125.250 511.050 126.150 ;
        RECT 514.950 125.250 517.050 126.150 ;
        RECT 508.950 121.950 511.050 124.050 ;
        RECT 512.250 122.250 513.750 123.150 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 499.950 118.950 502.050 121.050 ;
        RECT 511.950 118.950 514.050 121.050 ;
        RECT 515.400 118.050 516.450 121.950 ;
        RECT 514.950 115.950 517.050 118.050 ;
        RECT 505.950 97.950 508.050 100.050 ;
        RECT 511.950 97.950 514.050 100.050 ;
        RECT 482.400 95.400 486.450 96.450 ;
        RECT 475.950 91.950 478.050 94.050 ;
        RECT 472.950 79.950 475.050 82.050 ;
        RECT 476.400 70.050 477.450 91.950 ;
        RECT 475.950 67.950 478.050 70.050 ;
        RECT 469.950 61.950 472.050 64.050 ;
        RECT 470.400 55.050 471.450 61.950 ;
        RECT 482.400 61.050 483.450 95.400 ;
        RECT 490.950 94.950 493.050 97.050 ;
        RECT 496.950 94.950 499.050 97.050 ;
        RECT 484.950 92.250 486.750 93.150 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 491.400 91.050 492.450 94.950 ;
        RECT 493.950 91.950 496.050 94.050 ;
        RECT 484.950 88.950 487.050 91.050 ;
        RECT 488.250 89.850 489.750 90.750 ;
        RECT 490.950 88.950 493.050 91.050 ;
        RECT 494.250 89.850 496.050 90.750 ;
        RECT 490.950 86.850 493.050 87.750 ;
        RECT 487.950 82.950 490.050 85.050 ;
        RECT 481.950 58.950 484.050 61.050 ;
        RECT 472.950 55.950 475.050 58.050 ;
        RECT 473.400 55.050 474.450 55.950 ;
        RECT 488.400 55.050 489.450 82.950 ;
        RECT 497.400 64.050 498.450 94.950 ;
        RECT 506.400 94.050 507.450 97.950 ;
        RECT 499.950 91.950 502.050 94.050 ;
        RECT 502.950 92.250 504.750 93.150 ;
        RECT 505.950 91.950 508.050 94.050 ;
        RECT 509.250 92.250 511.050 93.150 ;
        RECT 496.950 61.950 499.050 64.050 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 494.400 55.050 495.450 55.950 ;
        RECT 466.950 53.250 468.750 54.150 ;
        RECT 469.950 52.950 472.050 55.050 ;
        RECT 472.950 52.950 475.050 55.050 ;
        RECT 475.950 52.950 478.050 55.050 ;
        RECT 487.950 52.950 490.050 55.050 ;
        RECT 493.950 52.950 496.050 55.050 ;
        RECT 497.250 53.250 499.050 54.150 ;
        RECT 466.950 51.450 469.050 52.050 ;
        RECT 464.400 50.400 469.050 51.450 ;
        RECT 470.250 50.850 472.050 51.750 ;
        RECT 466.950 49.950 469.050 50.400 ;
        RECT 472.950 50.250 475.050 51.150 ;
        RECT 475.950 50.850 478.050 51.750 ;
        RECT 487.950 50.850 490.050 51.750 ;
        RECT 490.950 50.250 493.050 51.150 ;
        RECT 493.950 50.850 495.750 51.750 ;
        RECT 496.950 49.950 499.050 52.050 ;
        RECT 472.950 46.950 475.050 49.050 ;
        RECT 490.950 46.950 493.050 49.050 ;
        RECT 497.400 33.450 498.450 49.950 ;
        RECT 500.400 49.050 501.450 91.950 ;
        RECT 502.950 88.950 505.050 91.050 ;
        RECT 506.250 89.850 507.750 90.750 ;
        RECT 508.950 90.450 511.050 91.050 ;
        RECT 512.400 90.450 513.450 97.950 ;
        RECT 508.950 89.400 513.450 90.450 ;
        RECT 508.950 88.950 511.050 89.400 ;
        RECT 503.400 85.050 504.450 88.950 ;
        RECT 502.950 82.950 505.050 85.050 ;
        RECT 511.950 58.950 514.050 61.050 ;
        RECT 512.400 55.050 513.450 58.950 ;
        RECT 518.400 55.050 519.450 190.950 ;
        RECT 521.400 181.050 522.450 229.950 ;
        RECT 524.400 208.050 525.450 235.950 ;
        RECT 527.400 232.050 528.450 265.950 ;
        RECT 533.400 253.050 534.450 265.950 ;
        RECT 532.950 250.950 535.050 253.050 ;
        RECT 532.950 241.950 535.050 244.050 ;
        RECT 529.950 238.950 532.050 241.050 ;
        RECT 530.400 232.050 531.450 238.950 ;
        RECT 526.950 229.950 529.050 232.050 ;
        RECT 529.950 229.950 532.050 232.050 ;
        RECT 526.950 226.950 529.050 229.050 ;
        RECT 523.950 205.950 526.050 208.050 ;
        RECT 523.950 197.250 526.050 198.150 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 175.950 526.050 178.050 ;
        RECT 524.400 172.050 525.450 175.950 ;
        RECT 523.950 169.950 526.050 172.050 ;
        RECT 520.950 167.250 523.050 168.150 ;
        RECT 523.950 167.850 526.050 168.750 ;
        RECT 520.950 163.950 523.050 166.050 ;
        RECT 521.400 130.050 522.450 163.950 ;
        RECT 527.400 151.050 528.450 226.950 ;
        RECT 529.950 220.950 532.050 223.050 ;
        RECT 530.400 217.050 531.450 220.950 ;
        RECT 529.950 214.950 532.050 217.050 ;
        RECT 529.950 197.250 532.050 198.150 ;
        RECT 529.950 193.950 532.050 196.050 ;
        RECT 533.400 175.050 534.450 241.950 ;
        RECT 536.400 190.050 537.450 271.950 ;
        RECT 539.400 244.050 540.450 301.950 ;
        RECT 545.400 294.450 546.450 310.950 ;
        RECT 548.400 304.050 549.450 331.950 ;
        RECT 551.400 316.050 552.450 337.950 ;
        RECT 550.950 313.950 553.050 316.050 ;
        RECT 553.950 312.450 556.050 313.050 ;
        RECT 551.400 311.400 556.050 312.450 ;
        RECT 547.950 301.950 550.050 304.050 ;
        RECT 551.400 301.050 552.450 311.400 ;
        RECT 553.950 310.950 556.050 311.400 ;
        RECT 557.250 311.250 559.050 312.150 ;
        RECT 553.950 308.850 555.750 309.750 ;
        RECT 556.950 304.950 559.050 307.050 ;
        RECT 550.950 298.950 553.050 301.050 ;
        RECT 557.400 298.050 558.450 304.950 ;
        RECT 556.950 295.950 559.050 298.050 ;
        RECT 542.400 293.400 546.450 294.450 ;
        RECT 542.400 286.050 543.450 293.400 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 541.950 283.950 544.050 286.050 ;
        RECT 541.950 274.950 544.050 277.050 ;
        RECT 542.400 268.050 543.450 274.950 ;
        RECT 541.950 265.950 544.050 268.050 ;
        RECT 545.400 265.050 546.450 289.950 ;
        RECT 553.950 283.950 556.050 286.050 ;
        RECT 547.950 272.250 550.050 273.150 ;
        RECT 554.400 271.050 555.450 283.950 ;
        RECT 547.950 268.950 550.050 271.050 ;
        RECT 551.250 269.250 552.750 270.150 ;
        RECT 553.950 268.950 556.050 271.050 ;
        RECT 557.250 269.250 559.050 270.150 ;
        RECT 548.400 265.050 549.450 268.950 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 554.250 266.850 555.750 267.750 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 544.950 262.950 547.050 265.050 ;
        RECT 547.950 262.950 550.050 265.050 ;
        RECT 548.400 262.050 549.450 262.950 ;
        RECT 547.950 259.950 550.050 262.050 ;
        RECT 544.950 256.950 547.050 259.050 ;
        RECT 545.400 244.050 546.450 256.950 ;
        RECT 551.400 253.050 552.450 265.950 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 550.950 250.950 553.050 253.050 ;
        RECT 538.950 241.950 541.050 244.050 ;
        RECT 544.950 241.950 547.050 244.050 ;
        RECT 550.950 241.950 553.050 244.050 ;
        RECT 538.950 238.950 541.050 241.050 ;
        RECT 542.250 239.250 544.050 240.150 ;
        RECT 544.950 239.850 547.050 240.750 ;
        RECT 547.950 239.250 550.050 240.150 ;
        RECT 538.950 236.850 540.750 237.750 ;
        RECT 541.950 235.950 544.050 238.050 ;
        RECT 547.950 235.950 550.050 238.050 ;
        RECT 542.400 235.050 543.450 235.950 ;
        RECT 541.950 232.950 544.050 235.050 ;
        RECT 538.950 229.950 541.050 232.050 ;
        RECT 535.950 187.950 538.050 190.050 ;
        RECT 539.400 178.050 540.450 229.950 ;
        RECT 548.400 211.050 549.450 235.950 ;
        RECT 551.400 235.050 552.450 241.950 ;
        RECT 554.400 238.050 555.450 256.950 ;
        RECT 560.400 250.050 561.450 340.950 ;
        RECT 559.950 247.950 562.050 250.050 ;
        RECT 563.400 247.050 564.450 352.950 ;
        RECT 566.400 337.050 567.450 370.950 ;
        RECT 569.400 346.050 570.450 376.950 ;
        RECT 571.950 373.950 574.050 376.050 ;
        RECT 572.400 364.050 573.450 373.950 ;
        RECT 571.950 361.950 574.050 364.050 ;
        RECT 568.950 343.950 571.050 346.050 ;
        RECT 568.950 341.250 571.050 342.150 ;
        RECT 568.950 337.950 571.050 340.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 569.400 331.050 570.450 337.950 ;
        RECT 568.950 328.950 571.050 331.050 ;
        RECT 572.400 328.050 573.450 361.950 ;
        RECT 575.400 346.050 576.450 391.950 ;
        RECT 577.950 385.950 580.050 388.050 ;
        RECT 578.400 382.050 579.450 385.950 ;
        RECT 577.950 379.950 580.050 382.050 ;
        RECT 577.950 376.950 580.050 379.050 ;
        RECT 578.400 352.050 579.450 376.950 ;
        RECT 577.950 349.950 580.050 352.050 ;
        RECT 574.950 343.950 577.050 346.050 ;
        RECT 574.950 341.250 577.050 342.150 ;
        RECT 574.950 337.950 577.050 340.050 ;
        RECT 575.400 337.050 576.450 337.950 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 565.950 325.950 568.050 328.050 ;
        RECT 571.950 325.950 574.050 328.050 ;
        RECT 566.400 307.050 567.450 325.950 ;
        RECT 575.400 313.050 576.450 334.950 ;
        RECT 578.400 333.450 579.450 349.950 ;
        RECT 581.400 336.450 582.450 421.950 ;
        RECT 587.400 406.050 588.450 475.950 ;
        RECT 590.400 472.050 591.450 598.950 ;
        RECT 592.950 595.950 595.050 598.050 ;
        RECT 596.250 596.850 597.750 597.750 ;
        RECT 598.950 595.950 601.050 598.050 ;
        RECT 602.250 596.850 604.050 597.750 ;
        RECT 605.400 595.050 606.450 634.950 ;
        RECT 608.400 634.050 609.450 638.400 ;
        RECT 613.950 634.950 616.050 637.050 ;
        RECT 614.400 634.050 615.450 634.950 ;
        RECT 607.950 631.950 610.050 634.050 ;
        RECT 611.250 632.250 612.750 633.150 ;
        RECT 613.950 631.950 616.050 634.050 ;
        RECT 619.950 631.950 622.050 634.050 ;
        RECT 607.950 629.850 609.750 630.750 ;
        RECT 610.950 628.950 613.050 631.050 ;
        RECT 614.250 629.850 616.050 630.750 ;
        RECT 607.950 625.950 610.050 628.050 ;
        RECT 592.950 593.850 595.050 594.750 ;
        RECT 598.950 592.950 601.050 595.050 ;
        RECT 604.950 592.950 607.050 595.050 ;
        RECT 599.400 552.450 600.450 592.950 ;
        RECT 601.950 556.950 604.050 559.050 ;
        RECT 601.950 554.850 604.050 555.750 ;
        RECT 604.950 554.250 607.050 555.150 ;
        RECT 604.950 552.450 607.050 553.050 ;
        RECT 608.400 552.450 609.450 625.950 ;
        RECT 611.400 601.050 612.450 628.950 ;
        RECT 620.400 610.050 621.450 631.950 ;
        RECT 623.400 616.050 624.450 661.950 ;
        RECT 629.400 640.050 630.450 671.400 ;
        RECT 635.400 646.050 636.450 685.950 ;
        RECT 647.400 682.050 648.450 697.950 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 637.950 670.950 640.050 673.050 ;
        RECT 634.950 643.950 637.050 646.050 ;
        RECT 625.950 637.950 628.050 640.050 ;
        RECT 628.950 637.950 631.050 640.050 ;
        RECT 626.400 634.050 627.450 637.950 ;
        RECT 625.950 631.950 628.050 634.050 ;
        RECT 631.950 633.450 634.050 634.050 ;
        RECT 635.400 633.450 636.450 643.950 ;
        RECT 629.250 632.250 630.750 633.150 ;
        RECT 631.950 632.400 636.450 633.450 ;
        RECT 631.950 631.950 634.050 632.400 ;
        RECT 625.950 629.850 627.750 630.750 ;
        RECT 628.950 628.950 631.050 631.050 ;
        RECT 632.250 629.850 634.050 630.750 ;
        RECT 635.400 628.050 636.450 632.400 ;
        RECT 628.950 625.950 631.050 628.050 ;
        RECT 634.950 625.950 637.050 628.050 ;
        RECT 622.950 613.950 625.050 616.050 ;
        RECT 613.950 607.950 616.050 610.050 ;
        RECT 619.950 607.950 622.050 610.050 ;
        RECT 625.950 607.950 628.050 610.050 ;
        RECT 614.400 601.050 615.450 607.950 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 620.400 604.050 621.450 604.950 ;
        RECT 619.950 601.950 622.050 604.050 ;
        RECT 610.950 598.950 613.050 601.050 ;
        RECT 613.950 598.950 616.050 601.050 ;
        RECT 617.250 599.250 619.050 600.150 ;
        RECT 619.950 599.850 622.050 600.750 ;
        RECT 622.950 599.250 625.050 600.150 ;
        RECT 613.950 596.850 615.750 597.750 ;
        RECT 616.950 595.950 619.050 598.050 ;
        RECT 622.950 597.450 625.050 598.050 ;
        RECT 626.400 597.450 627.450 607.950 ;
        RECT 622.950 596.400 627.450 597.450 ;
        RECT 622.950 595.950 625.050 596.400 ;
        RECT 629.400 592.050 630.450 625.950 ;
        RECT 638.400 607.050 639.450 670.950 ;
        RECT 640.950 668.250 642.750 669.150 ;
        RECT 643.950 667.950 646.050 670.050 ;
        RECT 647.250 668.250 649.050 669.150 ;
        RECT 640.950 664.950 643.050 667.050 ;
        RECT 644.250 665.850 645.750 666.750 ;
        RECT 646.950 664.950 649.050 667.050 ;
        RECT 647.400 661.050 648.450 664.950 ;
        RECT 650.400 661.050 651.450 700.950 ;
        RECT 652.950 667.950 655.050 670.050 ;
        RECT 640.950 658.950 643.050 661.050 ;
        RECT 646.950 658.950 649.050 661.050 ;
        RECT 649.950 658.950 652.050 661.050 ;
        RECT 641.400 658.050 642.450 658.950 ;
        RECT 640.950 655.950 643.050 658.050 ;
        RECT 637.950 604.950 640.050 607.050 ;
        RECT 631.950 596.250 633.750 597.150 ;
        RECT 634.950 595.950 637.050 598.050 ;
        RECT 638.250 596.250 640.050 597.150 ;
        RECT 631.950 592.950 634.050 595.050 ;
        RECT 635.250 593.850 636.750 594.750 ;
        RECT 637.950 592.950 640.050 595.050 ;
        RECT 632.400 592.050 633.450 592.950 ;
        RECT 628.950 589.950 631.050 592.050 ;
        RECT 631.950 589.950 634.050 592.050 ;
        RECT 638.400 577.050 639.450 592.950 ;
        RECT 637.950 574.950 640.050 577.050 ;
        RECT 613.950 567.300 616.050 569.400 ;
        RECT 614.550 563.700 615.750 567.300 ;
        RECT 634.950 566.400 637.050 568.500 ;
        RECT 613.950 561.600 616.050 563.700 ;
        RECT 610.950 553.950 613.050 556.050 ;
        RECT 599.400 551.400 603.450 552.450 ;
        RECT 598.950 544.950 601.050 547.050 ;
        RECT 595.950 541.950 598.050 544.050 ;
        RECT 596.400 523.050 597.450 541.950 ;
        RECT 599.400 529.050 600.450 544.950 ;
        RECT 598.950 526.950 601.050 529.050 ;
        RECT 595.950 520.950 598.050 523.050 ;
        RECT 598.950 505.950 601.050 508.050 ;
        RECT 595.950 495.300 598.050 497.400 ;
        RECT 596.550 491.700 597.750 495.300 ;
        RECT 592.950 487.950 595.050 490.050 ;
        RECT 595.950 489.600 598.050 491.700 ;
        RECT 593.400 487.050 594.450 487.950 ;
        RECT 592.950 484.950 595.050 487.050 ;
        RECT 593.400 484.050 594.450 484.950 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 592.950 479.850 595.050 480.750 ;
        RECT 596.550 477.600 597.750 489.600 ;
        RECT 595.950 475.500 598.050 477.600 ;
        RECT 599.400 475.050 600.450 505.950 ;
        RECT 602.400 505.050 603.450 551.400 ;
        RECT 604.950 551.400 609.450 552.450 ;
        RECT 610.950 551.850 613.050 552.750 ;
        RECT 604.950 550.950 607.050 551.400 ;
        RECT 605.400 544.050 606.450 550.950 ;
        RECT 614.550 549.600 615.750 561.600 ;
        RECT 619.950 556.950 622.050 559.050 ;
        RECT 622.950 557.250 625.050 558.150 ;
        RECT 628.950 557.250 631.050 558.150 ;
        RECT 620.400 550.050 621.450 556.950 ;
        RECT 622.950 553.950 625.050 556.050 ;
        RECT 628.950 553.950 631.050 556.050 ;
        RECT 631.950 553.950 634.050 556.050 ;
        RECT 613.950 547.500 616.050 549.600 ;
        RECT 619.950 547.950 622.050 550.050 ;
        RECT 604.950 541.950 607.050 544.050 ;
        RECT 623.400 541.050 624.450 553.950 ;
        RECT 622.950 538.950 625.050 541.050 ;
        RECT 629.400 538.050 630.450 553.950 ;
        RECT 628.950 535.950 631.050 538.050 ;
        RECT 628.950 532.950 631.050 535.050 ;
        RECT 607.950 529.950 610.050 532.050 ;
        RECT 622.950 529.950 625.050 532.050 ;
        RECT 608.400 529.050 609.450 529.950 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 613.950 528.450 616.050 529.050 ;
        RECT 611.250 527.250 612.750 528.150 ;
        RECT 613.950 527.400 618.450 528.450 ;
        RECT 622.950 527.850 625.050 528.750 ;
        RECT 613.950 526.950 616.050 527.400 ;
        RECT 617.400 526.050 618.450 527.400 ;
        RECT 625.950 527.250 628.050 528.150 ;
        RECT 604.950 523.950 607.050 526.050 ;
        RECT 608.250 524.850 609.750 525.750 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 614.250 524.850 616.050 525.750 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 604.950 521.850 607.050 522.750 ;
        RECT 611.400 522.450 612.450 523.950 ;
        RECT 608.400 521.400 612.450 522.450 ;
        RECT 601.950 502.950 604.050 505.050 ;
        RECT 601.950 487.950 604.050 490.050 ;
        RECT 598.950 472.950 601.050 475.050 ;
        RECT 589.950 469.950 592.050 472.050 ;
        RECT 595.950 469.950 598.050 472.050 ;
        RECT 589.950 454.950 592.050 457.050 ;
        RECT 589.950 452.850 592.050 453.750 ;
        RECT 592.950 452.250 595.050 453.150 ;
        RECT 592.950 448.950 595.050 451.050 ;
        RECT 593.400 448.050 594.450 448.950 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 596.400 421.050 597.450 469.950 ;
        RECT 598.950 457.950 601.050 460.050 ;
        RECT 599.400 457.050 600.450 457.950 ;
        RECT 598.950 454.950 601.050 457.050 ;
        RECT 598.950 452.850 601.050 453.750 ;
        RECT 602.400 436.050 603.450 487.950 ;
        RECT 604.950 485.250 607.050 486.150 ;
        RECT 604.950 481.950 607.050 484.050 ;
        RECT 605.400 475.050 606.450 481.950 ;
        RECT 604.950 472.950 607.050 475.050 ;
        RECT 608.400 460.050 609.450 521.400 ;
        RECT 611.400 520.050 612.450 521.400 ;
        RECT 625.950 520.950 628.050 523.050 ;
        RECT 610.950 517.950 613.050 520.050 ;
        RECT 622.950 499.950 625.050 502.050 ;
        RECT 619.950 496.950 622.050 499.050 ;
        RECT 616.950 494.400 619.050 496.500 ;
        RECT 610.950 485.250 613.050 486.150 ;
        RECT 613.950 484.950 616.050 487.050 ;
        RECT 610.950 481.950 613.050 484.050 ;
        RECT 611.400 478.050 612.450 481.950 ;
        RECT 610.950 475.950 613.050 478.050 ;
        RECT 610.950 466.950 613.050 469.050 ;
        RECT 611.400 460.050 612.450 466.950 ;
        RECT 614.400 460.050 615.450 484.950 ;
        RECT 617.400 477.600 618.600 494.400 ;
        RECT 616.950 475.500 619.050 477.600 ;
        RECT 607.950 457.950 610.050 460.050 ;
        RECT 610.950 457.950 613.050 460.050 ;
        RECT 613.950 457.950 616.050 460.050 ;
        RECT 604.950 456.450 607.050 457.050 ;
        RECT 607.950 456.450 610.050 457.050 ;
        RECT 604.950 455.400 610.050 456.450 ;
        RECT 611.250 455.850 612.750 456.750 ;
        RECT 613.950 456.450 616.050 457.050 ;
        RECT 604.950 454.950 607.050 455.400 ;
        RECT 607.950 454.950 610.050 455.400 ;
        RECT 613.950 455.400 618.450 456.450 ;
        RECT 613.950 454.950 616.050 455.400 ;
        RECT 601.950 433.950 604.050 436.050 ;
        RECT 601.950 430.950 604.050 433.050 ;
        RECT 589.950 418.950 592.050 421.050 ;
        RECT 595.950 418.950 598.050 421.050 ;
        RECT 598.950 418.950 601.050 421.050 ;
        RECT 586.950 403.950 589.050 406.050 ;
        RECT 586.950 385.950 589.050 388.050 ;
        RECT 590.400 385.050 591.450 418.950 ;
        RECT 599.400 418.050 600.450 418.950 ;
        RECT 602.400 418.050 603.450 430.950 ;
        RECT 598.950 415.950 601.050 418.050 ;
        RECT 601.950 415.950 604.050 418.050 ;
        RECT 592.950 413.250 594.750 414.150 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 592.950 409.950 595.050 412.050 ;
        RECT 596.250 410.850 598.050 411.750 ;
        RECT 593.400 397.050 594.450 409.950 ;
        RECT 599.400 403.050 600.450 415.950 ;
        RECT 598.950 400.950 601.050 403.050 ;
        RECT 595.950 397.950 598.050 400.050 ;
        RECT 592.950 394.950 595.050 397.050 ;
        RECT 583.950 382.950 586.050 385.050 ;
        RECT 587.250 383.850 588.750 384.750 ;
        RECT 589.950 382.950 592.050 385.050 ;
        RECT 583.950 380.850 586.050 381.750 ;
        RECT 586.950 379.950 589.050 382.050 ;
        RECT 589.950 380.850 592.050 381.750 ;
        RECT 583.950 340.950 586.050 343.050 ;
        RECT 583.950 338.850 586.050 339.750 ;
        RECT 581.400 335.400 585.450 336.450 ;
        RECT 578.400 332.400 582.450 333.450 ;
        RECT 568.950 310.950 571.050 313.050 ;
        RECT 574.950 310.950 577.050 313.050 ;
        RECT 569.400 310.050 570.450 310.950 ;
        RECT 568.950 307.950 571.050 310.050 ;
        RECT 574.950 307.950 577.050 310.050 ;
        RECT 578.250 308.250 580.050 309.150 ;
        RECT 565.950 304.950 568.050 307.050 ;
        RECT 568.950 305.850 570.750 306.750 ;
        RECT 571.950 304.950 574.050 307.050 ;
        RECT 575.250 305.850 576.750 306.750 ;
        RECT 577.950 306.450 580.050 307.050 ;
        RECT 581.400 306.450 582.450 332.400 ;
        RECT 577.950 305.400 582.450 306.450 ;
        RECT 577.950 304.950 580.050 305.400 ;
        RECT 565.950 301.950 568.050 304.050 ;
        RECT 571.950 302.850 574.050 303.750 ;
        RECT 566.400 268.050 567.450 301.950 ;
        RECT 568.950 280.950 571.050 283.050 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 566.400 262.050 567.450 265.950 ;
        RECT 565.950 259.950 568.050 262.050 ;
        RECT 562.950 244.950 565.050 247.050 ;
        RECT 562.950 241.950 565.050 244.050 ;
        RECT 563.400 241.050 564.450 241.950 ;
        RECT 556.950 238.950 559.050 241.050 ;
        RECT 560.250 239.250 561.750 240.150 ;
        RECT 562.950 238.950 565.050 241.050 ;
        RECT 553.950 235.950 556.050 238.050 ;
        RECT 556.950 236.850 558.750 237.750 ;
        RECT 559.950 235.950 562.050 238.050 ;
        RECT 563.250 236.850 564.750 237.750 ;
        RECT 565.950 235.950 568.050 238.050 ;
        RECT 550.950 232.950 553.050 235.050 ;
        RECT 560.400 232.050 561.450 235.950 ;
        RECT 565.950 233.850 568.050 234.750 ;
        RECT 559.950 229.950 562.050 232.050 ;
        RECT 569.400 214.050 570.450 280.950 ;
        RECT 577.950 274.950 580.050 277.050 ;
        RECT 571.950 272.250 574.050 273.150 ;
        RECT 578.400 271.050 579.450 274.950 ;
        RECT 571.950 268.950 574.050 271.050 ;
        RECT 575.250 269.250 576.750 270.150 ;
        RECT 577.950 268.950 580.050 271.050 ;
        RECT 581.250 269.250 583.050 270.150 ;
        RECT 572.400 265.050 573.450 268.950 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 578.250 266.850 579.750 267.750 ;
        RECT 580.950 265.950 583.050 268.050 ;
        RECT 581.400 265.050 582.450 265.950 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 580.950 264.450 583.050 265.050 ;
        RECT 578.400 263.400 583.050 264.450 ;
        RECT 578.400 229.050 579.450 263.400 ;
        RECT 580.950 262.950 583.050 263.400 ;
        RECT 584.400 256.050 585.450 335.400 ;
        RECT 587.400 301.050 588.450 379.950 ;
        RECT 589.950 373.950 592.050 376.050 ;
        RECT 590.400 309.450 591.450 373.950 ;
        RECT 592.950 349.950 595.050 352.050 ;
        RECT 596.400 351.450 597.450 397.950 ;
        RECT 598.950 383.250 601.050 384.150 ;
        RECT 598.950 379.950 601.050 382.050 ;
        RECT 599.400 355.050 600.450 379.950 ;
        RECT 602.400 373.050 603.450 415.950 ;
        RECT 605.400 379.050 606.450 454.950 ;
        RECT 607.950 452.850 610.050 453.750 ;
        RECT 613.950 452.850 616.050 453.750 ;
        RECT 617.400 448.050 618.450 455.400 ;
        RECT 616.950 445.950 619.050 448.050 ;
        RECT 607.950 416.250 610.050 417.150 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 611.250 413.250 612.750 414.150 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 617.250 413.250 619.050 414.150 ;
        RECT 608.400 406.050 609.450 412.950 ;
        RECT 610.950 409.950 613.050 412.050 ;
        RECT 614.250 410.850 615.750 411.750 ;
        RECT 616.950 409.950 619.050 412.050 ;
        RECT 611.400 409.050 612.450 409.950 ;
        RECT 617.400 409.050 618.450 409.950 ;
        RECT 610.950 406.950 613.050 409.050 ;
        RECT 616.950 406.950 619.050 409.050 ;
        RECT 620.400 406.050 621.450 496.950 ;
        RECT 623.400 457.050 624.450 499.950 ;
        RECT 626.400 469.050 627.450 520.950 ;
        RECT 629.400 487.050 630.450 532.950 ;
        RECT 632.400 532.050 633.450 553.950 ;
        RECT 635.400 549.600 636.600 566.400 ;
        RECT 634.950 547.500 637.050 549.600 ;
        RECT 638.400 534.450 639.450 574.950 ;
        RECT 641.400 535.050 642.450 655.950 ;
        RECT 653.400 633.450 654.450 667.950 ;
        RECT 656.400 664.050 657.450 736.950 ;
        RECT 659.400 673.050 660.450 760.950 ;
        RECT 662.400 742.050 663.450 781.950 ;
        RECT 661.950 739.950 664.050 742.050 ;
        RECT 662.400 709.050 663.450 739.950 ;
        RECT 665.400 733.050 666.450 820.950 ;
        RECT 673.950 817.950 676.050 820.050 ;
        RECT 680.400 817.050 681.450 826.950 ;
        RECT 683.400 826.050 684.450 844.950 ;
        RECT 686.400 841.050 687.450 845.400 ;
        RECT 688.950 844.950 691.050 845.400 ;
        RECT 724.950 844.950 727.050 847.050 ;
        RECT 688.950 842.850 691.050 843.750 ;
        RECT 709.950 842.850 712.050 843.750 ;
        RECT 724.950 842.850 727.050 843.750 ;
        RECT 727.950 842.250 730.050 843.150 ;
        RECT 685.950 838.950 688.050 841.050 ;
        RECT 721.950 838.950 724.050 841.050 ;
        RECT 727.950 838.950 730.050 841.050 ;
        RECT 686.400 829.050 687.450 838.950 ;
        RECT 685.950 826.950 688.050 829.050 ;
        RECT 682.950 823.950 685.050 826.050 ;
        RECT 706.950 823.950 709.050 826.050 ;
        RECT 691.950 819.450 694.050 820.050 ;
        RECT 689.400 818.400 694.050 819.450 ;
        RECT 689.400 817.050 690.450 818.400 ;
        RECT 691.950 817.950 694.050 818.400 ;
        RECT 707.400 817.050 708.450 823.950 ;
        RECT 712.950 817.950 715.050 820.050 ;
        RECT 713.400 817.050 714.450 817.950 ;
        RECT 670.950 815.250 673.050 816.150 ;
        RECT 673.950 815.850 676.050 816.750 ;
        RECT 676.950 815.250 678.750 816.150 ;
        RECT 679.950 814.950 682.050 817.050 ;
        RECT 688.950 814.950 691.050 817.050 ;
        RECT 691.950 815.850 694.050 816.750 ;
        RECT 694.950 815.250 697.050 816.150 ;
        RECT 706.950 814.950 709.050 817.050 ;
        RECT 710.250 815.250 711.750 816.150 ;
        RECT 712.950 814.950 715.050 817.050 ;
        RECT 722.400 816.450 723.450 838.950 ;
        RECT 727.950 821.400 730.050 823.500 ;
        RECT 724.950 818.250 727.050 819.150 ;
        RECT 724.950 816.450 727.050 817.050 ;
        RECT 722.400 815.400 727.050 816.450 ;
        RECT 724.950 814.950 727.050 815.400 ;
        RECT 670.950 811.950 673.050 814.050 ;
        RECT 676.950 811.950 679.050 814.050 ;
        RECT 680.250 812.850 682.050 813.750 ;
        RECT 694.950 811.950 697.050 814.050 ;
        RECT 706.950 812.850 708.750 813.750 ;
        RECT 709.950 811.950 712.050 814.050 ;
        RECT 713.250 812.850 714.750 813.750 ;
        RECT 715.950 813.450 718.050 814.050 ;
        RECT 715.950 812.400 720.450 813.450 ;
        RECT 715.950 811.950 718.050 812.400 ;
        RECT 671.400 805.050 672.450 811.950 ;
        RECT 677.400 811.050 678.450 811.950 ;
        RECT 710.400 811.050 711.450 811.950 ;
        RECT 676.950 808.950 679.050 811.050 ;
        RECT 682.950 808.950 685.050 811.050 ;
        RECT 709.950 808.950 712.050 811.050 ;
        RECT 715.950 809.850 718.050 810.750 ;
        RECT 670.950 802.950 673.050 805.050 ;
        RECT 670.950 772.950 673.050 775.050 ;
        RECT 667.950 770.250 670.050 771.150 ;
        RECT 670.950 770.850 673.050 771.750 ;
        RECT 679.950 769.950 682.050 772.050 ;
        RECT 667.950 766.950 670.050 769.050 ;
        RECT 667.950 745.950 670.050 748.050 ;
        RECT 667.950 743.850 669.750 744.750 ;
        RECT 670.950 744.450 673.050 745.050 ;
        RECT 673.950 744.450 676.050 745.050 ;
        RECT 670.950 743.400 676.050 744.450 ;
        RECT 670.950 742.950 673.050 743.400 ;
        RECT 673.950 742.950 676.050 743.400 ;
        RECT 676.950 743.250 679.050 744.150 ;
        RECT 670.950 740.850 673.050 741.750 ;
        RECT 664.950 730.950 667.050 733.050 ;
        RECT 674.400 724.050 675.450 742.950 ;
        RECT 676.950 741.450 679.050 742.050 ;
        RECT 680.400 741.450 681.450 769.950 ;
        RECT 676.950 740.400 681.450 741.450 ;
        RECT 676.950 739.950 679.050 740.400 ;
        RECT 683.400 739.050 684.450 808.950 ;
        RECT 719.400 807.450 720.450 812.400 ;
        RECT 716.400 806.400 720.450 807.450 ;
        RECT 700.950 787.950 703.050 790.050 ;
        RECT 685.950 778.950 688.050 781.050 ;
        RECT 691.950 779.250 694.050 780.150 ;
        RECT 686.400 778.050 687.450 778.950 ;
        RECT 685.950 775.950 688.050 778.050 ;
        RECT 689.250 776.250 690.750 777.150 ;
        RECT 691.950 775.950 694.050 778.050 ;
        RECT 695.250 776.250 697.050 777.150 ;
        RECT 685.950 773.850 687.750 774.750 ;
        RECT 688.950 772.950 691.050 775.050 ;
        RECT 689.400 772.050 690.450 772.950 ;
        RECT 688.950 769.950 691.050 772.050 ;
        RECT 692.400 769.050 693.450 775.950 ;
        RECT 694.950 772.950 697.050 775.050 ;
        RECT 697.950 769.950 700.050 772.050 ;
        RECT 691.950 766.950 694.050 769.050 ;
        RECT 698.400 757.050 699.450 769.950 ;
        RECT 691.950 754.950 694.050 757.050 ;
        RECT 697.950 754.950 700.050 757.050 ;
        RECT 692.400 748.050 693.450 754.950 ;
        RECT 688.950 745.950 691.050 748.050 ;
        RECT 691.950 745.950 694.050 748.050 ;
        RECT 689.400 745.050 690.450 745.950 ;
        RECT 688.950 742.950 691.050 745.050 ;
        RECT 692.250 743.850 693.750 744.750 ;
        RECT 694.950 742.950 697.050 745.050 ;
        RECT 688.950 740.850 691.050 741.750 ;
        RECT 694.950 740.850 697.050 741.750 ;
        RECT 701.400 741.450 702.450 787.950 ;
        RECT 703.950 772.950 706.050 775.050 ;
        RECT 709.950 772.950 712.050 775.050 ;
        RECT 713.250 773.250 715.050 774.150 ;
        RECT 703.950 770.850 706.050 771.750 ;
        RECT 706.950 770.250 709.050 771.150 ;
        RECT 709.950 770.850 711.750 771.750 ;
        RECT 712.950 771.450 715.050 772.050 ;
        RECT 716.400 771.450 717.450 806.400 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 712.950 770.400 717.450 771.450 ;
        RECT 712.950 769.950 715.050 770.400 ;
        RECT 706.950 766.950 709.050 769.050 ;
        RECT 712.950 766.950 715.050 769.050 ;
        RECT 706.950 754.950 709.050 757.050 ;
        RECT 698.400 740.400 702.450 741.450 ;
        RECT 682.950 736.950 685.050 739.050 ;
        RECT 691.950 736.950 694.050 739.050 ;
        RECT 692.400 727.050 693.450 736.950 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 673.950 721.950 676.050 724.050 ;
        RECT 688.950 721.950 691.050 724.050 ;
        RECT 661.950 706.950 664.050 709.050 ;
        RECT 667.950 707.250 670.050 708.150 ;
        RECT 673.950 706.950 676.050 709.050 ;
        RECT 682.950 707.250 685.050 708.150 ;
        RECT 661.950 703.950 664.050 706.050 ;
        RECT 665.250 704.250 666.750 705.150 ;
        RECT 667.950 703.950 670.050 706.050 ;
        RECT 671.250 704.250 673.050 705.150 ;
        RECT 661.950 701.850 663.750 702.750 ;
        RECT 664.950 700.950 667.050 703.050 ;
        RECT 668.400 697.050 669.450 703.950 ;
        RECT 670.950 700.950 673.050 703.050 ;
        RECT 667.950 694.950 670.050 697.050 ;
        RECT 671.400 682.050 672.450 700.950 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 670.950 676.950 673.050 679.050 ;
        RECT 658.950 670.950 661.050 673.050 ;
        RECT 661.950 670.950 664.050 673.050 ;
        RECT 667.950 672.450 670.050 673.050 ;
        RECT 671.400 672.450 672.450 676.950 ;
        RECT 665.250 671.250 666.750 672.150 ;
        RECT 667.950 671.400 672.450 672.450 ;
        RECT 667.950 670.950 670.050 671.400 ;
        RECT 658.950 667.950 661.050 670.050 ;
        RECT 662.250 668.850 663.750 669.750 ;
        RECT 664.950 667.950 667.050 670.050 ;
        RECT 668.250 668.850 670.050 669.750 ;
        RECT 665.400 667.050 666.450 667.950 ;
        RECT 658.950 665.850 661.050 666.750 ;
        RECT 664.950 664.950 667.050 667.050 ;
        RECT 655.950 661.950 658.050 664.050 ;
        RECT 671.400 648.450 672.450 671.400 ;
        RECT 674.400 667.050 675.450 706.950 ;
        RECT 689.400 706.050 690.450 721.950 ;
        RECT 679.950 704.250 681.750 705.150 ;
        RECT 682.950 703.950 685.050 706.050 ;
        RECT 686.250 704.250 687.750 705.150 ;
        RECT 688.950 703.950 691.050 706.050 ;
        RECT 679.950 700.950 682.050 703.050 ;
        RECT 679.950 688.950 682.050 691.050 ;
        RECT 680.400 670.050 681.450 688.950 ;
        RECT 683.400 688.050 684.450 703.950 ;
        RECT 685.950 700.950 688.050 703.050 ;
        RECT 689.250 701.850 691.050 702.750 ;
        RECT 686.400 700.050 687.450 700.950 ;
        RECT 685.950 697.950 688.050 700.050 ;
        RECT 688.950 694.950 691.050 697.050 ;
        RECT 682.950 685.950 685.050 688.050 ;
        RECT 676.950 668.250 678.750 669.150 ;
        RECT 679.950 667.950 682.050 670.050 ;
        RECT 683.250 668.250 685.050 669.150 ;
        RECT 673.950 664.950 676.050 667.050 ;
        RECT 676.950 664.950 679.050 667.050 ;
        RECT 680.250 665.850 681.750 666.750 ;
        RECT 682.950 664.950 685.050 667.050 ;
        RECT 671.400 647.400 675.450 648.450 ;
        RECT 643.950 632.250 646.050 633.150 ;
        RECT 653.400 632.400 657.450 633.450 ;
        RECT 643.950 628.950 646.050 631.050 ;
        RECT 647.250 629.250 648.750 630.150 ;
        RECT 649.950 628.950 652.050 631.050 ;
        RECT 653.250 629.250 655.050 630.150 ;
        RECT 644.400 619.050 645.450 628.950 ;
        RECT 646.950 625.950 649.050 628.050 ;
        RECT 650.250 626.850 651.750 627.750 ;
        RECT 652.950 627.450 655.050 628.050 ;
        RECT 656.400 627.450 657.450 632.400 ;
        RECT 664.950 629.250 667.050 630.150 ;
        RECT 670.950 628.950 673.050 631.050 ;
        RECT 652.950 626.400 657.450 627.450 ;
        RECT 652.950 625.950 655.050 626.400 ;
        RECT 656.400 625.050 657.450 626.400 ;
        RECT 658.950 625.950 661.050 628.050 ;
        RECT 661.950 626.250 663.750 627.150 ;
        RECT 664.950 625.950 667.050 628.050 ;
        RECT 670.950 626.850 673.050 627.750 ;
        RECT 655.950 622.950 658.050 625.050 ;
        RECT 659.400 619.050 660.450 625.950 ;
        RECT 661.950 622.950 664.050 625.050 ;
        RECT 674.400 622.050 675.450 647.400 ;
        RECT 683.400 646.050 684.450 664.950 ;
        RECT 689.400 652.050 690.450 694.950 ;
        RECT 692.400 655.050 693.450 724.950 ;
        RECT 698.400 693.450 699.450 740.400 ;
        RECT 703.950 709.950 706.050 712.050 ;
        RECT 704.400 703.050 705.450 709.950 ;
        RECT 703.950 700.950 706.050 703.050 ;
        RECT 700.950 698.250 703.050 699.150 ;
        RECT 703.950 698.850 706.050 699.750 ;
        RECT 700.950 694.950 703.050 697.050 ;
        RECT 698.400 692.400 702.450 693.450 ;
        RECT 701.400 670.050 702.450 692.400 ;
        RECT 697.950 668.250 699.750 669.150 ;
        RECT 700.950 667.950 703.050 670.050 ;
        RECT 704.250 668.250 706.050 669.150 ;
        RECT 697.950 664.950 700.050 667.050 ;
        RECT 701.250 665.850 702.750 666.750 ;
        RECT 703.950 664.950 706.050 667.050 ;
        RECT 698.400 660.450 699.450 664.950 ;
        RECT 704.400 661.050 705.450 664.950 ;
        RECT 698.400 659.400 702.450 660.450 ;
        RECT 691.950 652.950 694.050 655.050 ;
        RECT 697.950 652.950 700.050 655.050 ;
        RECT 688.950 649.950 691.050 652.050 ;
        RECT 682.950 643.950 685.050 646.050 ;
        RECT 689.400 634.050 690.450 649.950 ;
        RECT 691.950 643.950 694.050 646.050 ;
        RECT 682.950 631.950 685.050 634.050 ;
        RECT 685.950 632.250 688.050 633.150 ;
        RECT 688.950 631.950 691.050 634.050 ;
        RECT 673.950 619.950 676.050 622.050 ;
        RECT 643.950 616.950 646.050 619.050 ;
        RECT 649.950 616.950 652.050 619.050 ;
        RECT 658.950 616.950 661.050 619.050 ;
        RECT 643.950 613.950 646.050 616.050 ;
        RECT 644.400 540.450 645.450 613.950 ;
        RECT 650.400 601.050 651.450 616.950 ;
        RECT 655.950 604.950 658.050 607.050 ;
        RECT 656.400 601.050 657.450 604.950 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 653.250 599.250 654.750 600.150 ;
        RECT 655.950 598.950 658.050 601.050 ;
        RECT 670.950 600.450 673.050 601.050 ;
        RECT 668.400 599.400 673.050 600.450 ;
        RECT 649.950 596.850 651.750 597.750 ;
        RECT 652.950 595.950 655.050 598.050 ;
        RECT 656.250 596.850 657.750 597.750 ;
        RECT 658.950 595.950 661.050 598.050 ;
        RECT 664.950 595.950 667.050 598.050 ;
        RECT 658.950 593.850 661.050 594.750 ;
        RECT 661.950 583.950 664.050 586.050 ;
        RECT 649.950 580.950 652.050 583.050 ;
        RECT 655.950 580.950 658.050 583.050 ;
        RECT 644.400 539.400 648.450 540.450 ;
        RECT 643.950 535.950 646.050 538.050 ;
        RECT 635.400 533.400 639.450 534.450 ;
        RECT 631.950 529.950 634.050 532.050 ;
        RECT 632.400 499.050 633.450 529.950 ;
        RECT 631.950 496.950 634.050 499.050 ;
        RECT 635.400 490.050 636.450 533.400 ;
        RECT 640.950 532.950 643.050 535.050 ;
        RECT 644.400 529.050 645.450 535.950 ;
        RECT 647.400 529.050 648.450 539.400 ;
        RECT 650.400 534.450 651.450 580.950 ;
        RECT 656.400 559.050 657.450 580.950 ;
        RECT 662.400 559.050 663.450 583.950 ;
        RECT 665.400 562.050 666.450 595.950 ;
        RECT 664.950 559.950 667.050 562.050 ;
        RECT 652.950 557.250 654.750 558.150 ;
        RECT 655.950 556.950 658.050 559.050 ;
        RECT 659.250 557.250 660.750 558.150 ;
        RECT 661.950 556.950 664.050 559.050 ;
        RECT 665.250 557.250 667.050 558.150 ;
        RECT 668.400 556.050 669.450 599.400 ;
        RECT 670.950 598.950 673.050 599.400 ;
        RECT 674.250 599.250 675.750 600.150 ;
        RECT 676.950 598.950 679.050 601.050 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 680.400 598.050 681.450 598.950 ;
        RECT 670.950 596.850 672.750 597.750 ;
        RECT 673.950 595.950 676.050 598.050 ;
        RECT 677.250 596.850 678.750 597.750 ;
        RECT 679.950 595.950 682.050 598.050 ;
        RECT 670.950 586.950 673.050 589.050 ;
        RECT 671.400 561.450 672.450 586.950 ;
        RECT 674.400 565.050 675.450 595.950 ;
        RECT 679.950 593.850 682.050 594.750 ;
        RECT 683.400 588.450 684.450 631.950 ;
        RECT 692.400 631.050 693.450 643.950 ;
        RECT 685.950 628.950 688.050 631.050 ;
        RECT 689.250 629.250 690.750 630.150 ;
        RECT 691.950 628.950 694.050 631.050 ;
        RECT 695.250 629.250 697.050 630.150 ;
        RECT 686.400 619.050 687.450 628.950 ;
        RECT 688.950 625.950 691.050 628.050 ;
        RECT 692.250 626.850 693.750 627.750 ;
        RECT 694.950 625.950 697.050 628.050 ;
        RECT 685.950 616.950 688.050 619.050 ;
        RECT 689.400 603.450 690.450 625.950 ;
        RECT 695.400 625.050 696.450 625.950 ;
        RECT 698.400 625.050 699.450 652.950 ;
        RECT 701.400 628.050 702.450 659.400 ;
        RECT 703.950 658.950 706.050 661.050 ;
        RECT 707.400 636.450 708.450 754.950 ;
        RECT 713.400 745.050 714.450 766.950 ;
        RECT 719.400 745.050 720.450 802.950 ;
        RECT 725.400 802.050 726.450 814.950 ;
        RECT 728.550 809.400 729.750 821.400 ;
        RECT 727.950 807.300 730.050 809.400 ;
        RECT 728.550 803.700 729.750 807.300 ;
        RECT 724.950 799.950 727.050 802.050 ;
        RECT 727.950 801.600 730.050 803.700 ;
        RECT 724.950 773.250 727.050 774.150 ;
        RECT 730.950 773.250 733.050 774.150 ;
        RECT 724.950 769.950 727.050 772.050 ;
        RECT 728.250 770.250 729.750 771.150 ;
        RECT 730.950 769.950 733.050 772.050 ;
        RECT 725.400 766.050 726.450 769.950 ;
        RECT 727.950 766.950 730.050 769.050 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 728.400 763.050 729.450 766.950 ;
        RECT 727.950 760.950 730.050 763.050 ;
        RECT 734.400 757.050 735.450 847.950 ;
        RECT 746.400 847.050 747.450 850.950 ;
        RECT 764.250 848.250 765.750 849.150 ;
        RECT 779.250 848.250 780.750 849.150 ;
        RECT 796.950 847.950 799.050 850.050 ;
        RECT 802.950 848.250 805.050 849.150 ;
        RECT 797.400 847.050 798.450 847.950 ;
        RECT 818.400 847.050 819.450 853.950 ;
        RECT 833.250 848.250 834.750 849.150 ;
        RECT 739.950 844.950 742.050 847.050 ;
        RECT 743.250 845.250 744.750 846.150 ;
        RECT 745.950 844.950 748.050 847.050 ;
        RECT 749.250 845.250 751.050 846.150 ;
        RECT 760.950 845.850 762.750 846.750 ;
        RECT 763.950 844.950 766.050 847.050 ;
        RECT 767.250 845.850 769.050 846.750 ;
        RECT 775.950 845.850 777.750 846.750 ;
        RECT 778.950 844.950 781.050 847.050 ;
        RECT 782.250 845.850 784.050 846.750 ;
        RECT 793.950 845.250 795.750 846.150 ;
        RECT 796.950 844.950 799.050 847.050 ;
        RECT 800.250 845.250 801.750 846.150 ;
        RECT 802.950 844.950 805.050 847.050 ;
        RECT 817.950 844.950 820.050 847.050 ;
        RECT 829.950 845.850 831.750 846.750 ;
        RECT 832.950 844.950 835.050 847.050 ;
        RECT 836.250 845.850 838.050 846.750 ;
        RECT 850.950 844.950 853.050 847.050 ;
        RECT 856.950 844.950 859.050 847.050 ;
        RECT 740.400 841.050 741.450 844.950 ;
        RECT 742.950 841.950 745.050 844.050 ;
        RECT 746.250 842.850 747.750 843.750 ;
        RECT 739.950 838.950 742.050 841.050 ;
        RECT 736.950 826.950 739.050 829.050 ;
        RECT 737.400 817.050 738.450 826.950 ;
        RECT 743.400 817.050 744.450 841.950 ;
        RECT 764.400 841.050 765.450 844.950 ;
        RECT 793.950 841.950 796.050 844.050 ;
        RECT 797.250 842.850 798.750 843.750 ;
        RECT 799.950 841.950 802.050 844.050 ;
        RECT 763.950 838.950 766.050 841.050 ;
        RECT 796.950 838.950 799.050 841.050 ;
        RECT 754.950 826.950 757.050 829.050 ;
        RECT 787.950 826.950 790.050 829.050 ;
        RECT 748.950 821.400 751.050 823.500 ;
        RECT 736.950 814.950 739.050 817.050 ;
        RECT 742.950 814.950 745.050 817.050 ;
        RECT 736.950 812.850 739.050 813.750 ;
        RECT 742.950 812.850 745.050 813.750 ;
        RECT 749.400 804.600 750.600 821.400 ;
        RECT 748.950 802.500 751.050 804.600 ;
        RECT 742.950 783.300 745.050 785.400 ;
        RECT 743.550 779.700 744.750 783.300 ;
        RECT 742.950 777.600 745.050 779.700 ;
        RECT 739.950 771.450 742.050 772.050 ;
        RECT 737.400 770.400 742.050 771.450 ;
        RECT 737.400 760.050 738.450 770.400 ;
        RECT 739.950 769.950 742.050 770.400 ;
        RECT 739.950 767.850 742.050 768.750 ;
        RECT 743.550 765.600 744.750 777.600 ;
        RECT 751.950 773.250 754.050 774.150 ;
        RECT 751.950 771.450 754.050 772.050 ;
        RECT 755.400 771.450 756.450 826.950 ;
        RECT 763.950 820.950 766.050 823.050 ;
        RECT 769.950 820.950 772.050 823.050 ;
        RECT 778.950 821.400 781.050 823.500 ;
        RECT 764.400 820.050 765.450 820.950 ;
        RECT 763.950 817.950 766.050 820.050 ;
        RECT 770.400 817.050 771.450 820.950 ;
        RECT 775.950 818.250 778.050 819.150 ;
        RECT 763.950 815.850 766.050 816.750 ;
        RECT 766.950 815.250 769.050 816.150 ;
        RECT 769.950 814.950 772.050 817.050 ;
        RECT 775.950 814.950 778.050 817.050 ;
        RECT 766.950 811.950 769.050 814.050 ;
        RECT 767.400 805.050 768.450 811.950 ;
        RECT 779.550 809.400 780.750 821.400 ;
        RECT 788.400 817.050 789.450 826.950 ;
        RECT 787.950 814.950 790.050 817.050 ;
        RECT 793.950 814.950 796.050 817.050 ;
        RECT 787.950 812.850 790.050 813.750 ;
        RECT 790.950 811.950 793.050 814.050 ;
        RECT 793.950 812.850 796.050 813.750 ;
        RECT 778.950 807.300 781.050 809.400 ;
        RECT 766.950 802.950 769.050 805.050 ;
        RECT 779.550 803.700 780.750 807.300 ;
        RECT 778.950 801.600 781.050 803.700 ;
        RECT 763.950 782.400 766.050 784.500 ;
        RECT 757.950 773.250 760.050 774.150 ;
        RECT 751.950 770.400 756.450 771.450 ;
        RECT 751.950 769.950 754.050 770.400 ;
        RECT 757.950 769.950 760.050 772.050 ;
        RECT 742.950 763.500 745.050 765.600 ;
        RECT 736.950 757.950 739.050 760.050 ;
        RECT 733.950 754.950 736.050 757.050 ;
        RECT 727.950 749.400 730.050 751.500 ;
        RECT 724.950 746.250 727.050 747.150 ;
        RECT 709.950 742.950 712.050 745.050 ;
        RECT 712.950 742.950 715.050 745.050 ;
        RECT 716.250 743.250 717.750 744.150 ;
        RECT 718.950 742.950 721.050 745.050 ;
        RECT 724.950 744.450 727.050 745.050 ;
        RECT 722.400 743.400 727.050 744.450 ;
        RECT 710.400 742.050 711.450 742.950 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 713.250 740.850 714.750 741.750 ;
        RECT 715.950 739.950 718.050 742.050 ;
        RECT 719.250 740.850 721.050 741.750 ;
        RECT 709.950 737.850 712.050 738.750 ;
        RECT 715.950 711.300 718.050 713.400 ;
        RECT 716.550 707.700 717.750 711.300 ;
        RECT 715.950 705.600 718.050 707.700 ;
        RECT 712.950 699.450 715.050 700.050 ;
        RECT 710.400 698.400 715.050 699.450 ;
        RECT 710.400 697.050 711.450 698.400 ;
        RECT 712.950 697.950 715.050 698.400 ;
        RECT 709.950 694.950 712.050 697.050 ;
        RECT 712.950 695.850 715.050 696.750 ;
        RECT 716.550 693.600 717.750 705.600 ;
        RECT 722.400 696.450 723.450 743.400 ;
        RECT 724.950 742.950 727.050 743.400 ;
        RECT 728.550 737.400 729.750 749.400 ;
        RECT 733.950 748.950 736.050 751.050 ;
        RECT 748.950 749.400 751.050 751.500 ;
        RECT 752.400 751.050 753.450 769.950 ;
        RECT 758.400 763.050 759.450 769.950 ;
        RECT 764.400 765.600 765.600 782.400 ;
        RECT 787.950 776.250 790.050 777.150 ;
        RECT 778.950 773.250 780.750 774.150 ;
        RECT 781.950 772.950 784.050 775.050 ;
        RECT 787.950 774.450 790.050 775.050 ;
        RECT 791.400 774.450 792.450 811.950 ;
        RECT 793.950 778.950 796.050 781.050 ;
        RECT 785.250 773.250 786.750 774.150 ;
        RECT 787.950 773.400 792.450 774.450 ;
        RECT 787.950 772.950 790.050 773.400 ;
        RECT 782.250 770.850 783.750 771.750 ;
        RECT 784.950 769.950 787.050 772.050 ;
        RECT 763.950 763.500 766.050 765.600 ;
        RECT 778.950 763.950 781.050 766.050 ;
        RECT 757.950 760.950 760.050 763.050 ;
        RECT 727.950 735.300 730.050 737.400 ;
        RECT 728.550 731.700 729.750 735.300 ;
        RECT 727.950 729.600 730.050 731.700 ;
        RECT 724.950 701.250 727.050 702.150 ;
        RECT 730.950 701.250 733.050 702.150 ;
        RECT 724.950 699.450 727.050 700.050 ;
        RECT 724.950 698.400 729.450 699.450 ;
        RECT 724.950 697.950 727.050 698.400 ;
        RECT 722.400 695.400 726.450 696.450 ;
        RECT 715.950 691.500 718.050 693.600 ;
        RECT 725.400 688.050 726.450 695.400 ;
        RECT 724.950 685.950 727.050 688.050 ;
        RECT 712.950 675.450 715.050 676.050 ;
        RECT 710.400 674.400 715.050 675.450 ;
        RECT 710.400 649.050 711.450 674.400 ;
        RECT 712.950 673.950 715.050 674.400 ;
        RECT 712.950 671.850 715.050 672.750 ;
        RECT 715.950 671.250 718.050 672.150 ;
        RECT 715.950 667.950 718.050 670.050 ;
        RECT 716.400 667.050 717.450 667.950 ;
        RECT 715.950 664.950 718.050 667.050 ;
        RECT 725.400 666.450 726.450 685.950 ;
        RECT 728.400 676.050 729.450 698.400 ;
        RECT 730.950 697.950 733.050 700.050 ;
        RECT 731.400 697.050 732.450 697.950 ;
        RECT 730.950 694.950 733.050 697.050 ;
        RECT 734.400 691.050 735.450 748.950 ;
        RECT 742.950 745.950 745.050 748.050 ;
        RECT 743.400 745.050 744.450 745.950 ;
        RECT 736.950 742.950 739.050 745.050 ;
        RECT 742.950 742.950 745.050 745.050 ;
        RECT 736.950 740.850 739.050 741.750 ;
        RECT 742.950 740.850 745.050 741.750 ;
        RECT 749.400 732.600 750.600 749.400 ;
        RECT 751.950 748.950 754.050 751.050 ;
        RECT 752.400 745.050 753.450 748.950 ;
        RECT 769.950 745.950 772.050 748.050 ;
        RECT 770.400 745.050 771.450 745.950 ;
        RECT 751.950 742.950 754.050 745.050 ;
        RECT 767.250 743.250 768.750 744.150 ;
        RECT 769.950 742.950 772.050 745.050 ;
        RECT 779.400 744.450 780.450 763.950 ;
        RECT 785.400 763.050 786.450 769.950 ;
        RECT 784.950 760.950 787.050 763.050 ;
        RECT 794.400 753.450 795.450 778.950 ;
        RECT 791.400 752.400 795.450 753.450 ;
        RECT 784.950 749.400 787.050 751.500 ;
        RECT 781.950 746.250 784.050 747.150 ;
        RECT 781.950 744.450 784.050 745.050 ;
        RECT 779.400 743.400 784.050 744.450 ;
        RECT 781.950 742.950 784.050 743.400 ;
        RECT 763.950 740.850 765.750 741.750 ;
        RECT 766.950 739.950 769.050 742.050 ;
        RECT 770.250 740.850 771.750 741.750 ;
        RECT 772.950 739.950 775.050 742.050 ;
        RECT 748.950 730.500 751.050 732.600 ;
        RECT 767.400 723.450 768.450 739.950 ;
        RECT 772.950 737.850 775.050 738.750 ;
        RECT 782.400 730.050 783.450 742.950 ;
        RECT 785.550 737.400 786.750 749.400 ;
        RECT 784.950 735.300 787.050 737.400 ;
        RECT 785.550 731.700 786.750 735.300 ;
        RECT 781.950 727.950 784.050 730.050 ;
        RECT 784.950 729.600 787.050 731.700 ;
        RECT 764.400 722.400 768.450 723.450 ;
        RECT 736.950 710.400 739.050 712.500 ;
        RECT 737.400 693.600 738.600 710.400 ;
        RECT 760.950 704.250 763.050 705.150 ;
        RECT 751.950 701.250 753.750 702.150 ;
        RECT 754.950 700.950 757.050 703.050 ;
        RECT 758.250 701.250 759.750 702.150 ;
        RECT 760.950 700.950 763.050 703.050 ;
        RECT 755.250 698.850 756.750 699.750 ;
        RECT 757.950 697.950 760.050 700.050 ;
        RECT 758.400 697.050 759.450 697.950 ;
        RECT 757.950 694.950 760.050 697.050 ;
        RECT 736.950 691.500 739.050 693.600 ;
        RECT 751.950 691.950 754.050 694.050 ;
        RECT 733.950 688.950 736.050 691.050 ;
        RECT 727.950 673.950 730.050 676.050 ;
        RECT 752.400 673.050 753.450 691.950 ;
        RECT 760.950 688.950 763.050 691.050 ;
        RECT 730.950 670.950 733.050 673.050 ;
        RECT 739.950 670.950 742.050 673.050 ;
        RECT 745.950 670.950 748.050 673.050 ;
        RECT 749.250 671.250 750.750 672.150 ;
        RECT 751.950 670.950 754.050 673.050 ;
        RECT 761.400 672.450 762.450 688.950 ;
        RECT 764.400 679.050 765.450 722.400 ;
        RECT 791.400 712.050 792.450 752.400 ;
        RECT 793.950 748.950 796.050 751.050 ;
        RECT 794.400 745.050 795.450 748.950 ;
        RECT 793.950 742.950 796.050 745.050 ;
        RECT 793.950 740.850 796.050 741.750 ;
        RECT 781.950 709.950 784.050 712.050 ;
        RECT 790.950 709.950 793.050 712.050 ;
        RECT 776.250 704.250 777.750 705.150 ;
        RECT 772.950 701.850 774.750 702.750 ;
        RECT 775.950 700.950 778.050 703.050 ;
        RECT 779.250 701.850 781.050 702.750 ;
        RECT 778.950 694.950 781.050 697.050 ;
        RECT 763.950 676.950 766.050 679.050 ;
        RECT 766.950 677.400 769.050 679.500 ;
        RECT 763.950 674.250 766.050 675.150 ;
        RECT 763.950 672.450 766.050 673.050 ;
        RECT 761.400 671.400 766.050 672.450 ;
        RECT 731.400 670.050 732.450 670.950 ;
        RECT 727.950 668.250 729.750 669.150 ;
        RECT 730.950 667.950 733.050 670.050 ;
        RECT 734.250 668.250 736.050 669.150 ;
        RECT 740.400 667.050 741.450 670.950 ;
        RECT 745.950 668.850 747.750 669.750 ;
        RECT 748.950 667.950 751.050 670.050 ;
        RECT 752.250 668.850 753.750 669.750 ;
        RECT 754.950 669.450 757.050 670.050 ;
        RECT 754.950 668.400 759.450 669.450 ;
        RECT 754.950 667.950 757.050 668.400 ;
        RECT 727.950 666.450 730.050 667.050 ;
        RECT 725.400 665.400 730.050 666.450 ;
        RECT 731.250 665.850 732.750 666.750 ;
        RECT 718.950 661.950 721.050 664.050 ;
        RECT 709.950 646.950 712.050 649.050 ;
        RECT 704.400 635.400 708.450 636.450 ;
        RECT 700.950 625.950 703.050 628.050 ;
        RECT 694.950 622.950 697.050 625.050 ;
        RECT 697.950 622.950 700.050 625.050 ;
        RECT 691.950 603.450 694.050 604.050 ;
        RECT 689.400 602.400 694.050 603.450 ;
        RECT 689.400 601.050 690.450 602.400 ;
        RECT 691.950 601.950 694.050 602.400 ;
        RECT 688.950 598.950 691.050 601.050 ;
        RECT 691.950 599.850 693.750 600.750 ;
        RECT 694.950 600.450 697.050 601.050 ;
        RECT 697.950 600.450 700.050 601.050 ;
        RECT 694.950 599.400 700.050 600.450 ;
        RECT 694.950 598.950 697.050 599.400 ;
        RECT 697.950 598.950 700.050 599.400 ;
        RECT 700.950 599.250 703.050 600.150 ;
        RECT 694.950 596.850 697.050 597.750 ;
        RECT 683.400 587.400 687.450 588.450 ;
        RECT 679.950 574.950 682.050 577.050 ;
        RECT 673.950 562.950 676.050 565.050 ;
        RECT 680.400 562.050 681.450 574.950 ;
        RECT 673.950 561.450 676.050 562.050 ;
        RECT 671.400 560.400 676.050 561.450 ;
        RECT 679.950 561.450 682.050 562.050 ;
        RECT 652.950 553.950 655.050 556.050 ;
        RECT 656.250 554.850 657.750 555.750 ;
        RECT 658.950 553.950 661.050 556.050 ;
        RECT 662.250 554.850 663.750 555.750 ;
        RECT 664.950 553.950 667.050 556.050 ;
        RECT 667.950 553.950 670.050 556.050 ;
        RECT 653.400 538.050 654.450 553.950 ;
        RECT 671.400 553.050 672.450 560.400 ;
        RECT 673.950 559.950 676.050 560.400 ;
        RECT 677.250 560.250 678.750 561.150 ;
        RECT 679.950 560.400 684.450 561.450 ;
        RECT 679.950 559.950 682.050 560.400 ;
        RECT 673.950 557.850 675.750 558.750 ;
        RECT 676.950 556.950 679.050 559.050 ;
        RECT 680.250 557.850 682.050 558.750 ;
        RECT 683.400 553.050 684.450 560.400 ;
        RECT 655.950 550.950 658.050 553.050 ;
        RECT 661.950 550.950 664.050 553.050 ;
        RECT 670.950 550.950 673.050 553.050 ;
        RECT 682.950 550.950 685.050 553.050 ;
        RECT 686.400 552.450 687.450 587.400 ;
        RECT 698.400 573.450 699.450 598.950 ;
        RECT 700.950 595.950 703.050 598.050 ;
        RECT 701.400 595.050 702.450 595.950 ;
        RECT 700.950 592.950 703.050 595.050 ;
        RECT 704.400 574.050 705.450 635.400 ;
        RECT 710.400 631.050 711.450 646.950 ;
        RECT 715.950 632.250 718.050 633.150 ;
        RECT 706.950 629.250 708.750 630.150 ;
        RECT 709.950 628.950 712.050 631.050 ;
        RECT 715.950 630.450 718.050 631.050 ;
        RECT 719.400 630.450 720.450 661.950 ;
        RECT 713.250 629.250 714.750 630.150 ;
        RECT 715.950 629.400 720.450 630.450 ;
        RECT 715.950 628.950 718.050 629.400 ;
        RECT 706.950 625.950 709.050 628.050 ;
        RECT 710.250 626.850 711.750 627.750 ;
        RECT 712.950 625.950 715.050 628.050 ;
        RECT 707.400 622.050 708.450 625.950 ;
        RECT 706.950 619.950 709.050 622.050 ;
        RECT 707.400 615.450 708.450 619.950 ;
        RECT 707.400 614.400 711.450 615.450 ;
        RECT 706.950 601.950 709.050 604.050 ;
        RECT 707.400 589.050 708.450 601.950 ;
        RECT 706.950 586.950 709.050 589.050 ;
        RECT 710.400 586.050 711.450 614.400 ;
        RECT 712.950 601.950 715.050 604.050 ;
        RECT 713.400 595.050 714.450 601.950 ;
        RECT 719.400 598.050 720.450 629.400 ;
        RECT 715.950 596.250 717.750 597.150 ;
        RECT 718.950 595.950 721.050 598.050 ;
        RECT 722.250 596.250 724.050 597.150 ;
        RECT 712.950 592.950 715.050 595.050 ;
        RECT 715.950 592.950 718.050 595.050 ;
        RECT 719.250 593.850 720.750 594.750 ;
        RECT 721.950 592.950 724.050 595.050 ;
        RECT 709.950 583.950 712.050 586.050 ;
        RECT 721.950 577.950 724.050 580.050 ;
        RECT 695.400 572.400 699.450 573.450 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 689.400 555.450 690.450 568.950 ;
        RECT 695.400 559.050 696.450 572.400 ;
        RECT 703.950 571.950 706.050 574.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 691.950 557.250 694.050 558.150 ;
        RECT 694.950 556.950 697.050 559.050 ;
        RECT 697.950 557.250 700.050 558.150 ;
        RECT 691.950 555.450 694.050 556.050 ;
        RECT 689.400 554.400 694.050 555.450 ;
        RECT 697.950 555.450 700.050 556.050 ;
        RECT 701.400 555.450 702.450 568.950 ;
        RECT 712.950 565.950 715.050 568.050 ;
        RECT 713.400 559.050 714.450 565.950 ;
        RECT 718.950 560.250 721.050 561.150 ;
        RECT 709.950 557.250 711.750 558.150 ;
        RECT 712.950 556.950 715.050 559.050 ;
        RECT 716.250 557.250 717.750 558.150 ;
        RECT 718.950 556.950 721.050 559.050 ;
        RECT 691.950 553.950 694.050 554.400 ;
        RECT 695.250 554.250 696.750 555.150 ;
        RECT 697.950 554.400 702.450 555.450 ;
        RECT 713.250 554.850 714.750 555.750 ;
        RECT 697.950 553.950 700.050 554.400 ;
        RECT 715.950 553.950 718.050 556.050 ;
        RECT 686.400 551.400 690.450 552.450 ;
        RECT 652.950 535.950 655.050 538.050 ;
        RECT 650.400 533.400 654.450 534.450 ;
        RECT 649.950 529.950 652.050 532.050 ;
        RECT 641.250 527.250 642.750 528.150 ;
        RECT 643.950 526.950 646.050 529.050 ;
        RECT 646.950 526.950 649.050 529.050 ;
        RECT 637.950 524.850 639.750 525.750 ;
        RECT 640.950 523.950 643.050 526.050 ;
        RECT 644.250 524.850 645.750 525.750 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 646.950 521.850 649.050 522.750 ;
        RECT 634.950 487.950 637.050 490.050 ;
        RECT 640.950 488.250 643.050 489.150 ;
        RECT 643.950 487.950 646.050 490.050 ;
        RECT 628.950 484.950 631.050 487.050 ;
        RECT 631.950 485.250 633.750 486.150 ;
        RECT 634.950 484.950 637.050 487.050 ;
        RECT 640.950 486.450 643.050 487.050 ;
        RECT 644.400 486.450 645.450 487.950 ;
        RECT 638.250 485.250 639.750 486.150 ;
        RECT 640.950 485.400 645.450 486.450 ;
        RECT 640.950 484.950 643.050 485.400 ;
        RECT 625.950 466.950 628.050 469.050 ;
        RECT 629.400 466.050 630.450 484.950 ;
        RECT 635.250 482.850 636.750 483.750 ;
        RECT 637.950 481.950 640.050 484.050 ;
        RECT 638.400 478.050 639.450 481.950 ;
        RECT 650.400 478.050 651.450 529.950 ;
        RECT 653.400 514.050 654.450 533.400 ;
        RECT 656.400 520.050 657.450 550.950 ;
        RECT 662.400 540.450 663.450 550.950 ;
        RECT 659.400 539.400 663.450 540.450 ;
        RECT 659.400 532.050 660.450 539.400 ;
        RECT 658.950 529.950 661.050 532.050 ;
        RECT 659.400 527.400 675.450 528.450 ;
        RECT 659.400 526.050 660.450 527.400 ;
        RECT 674.400 526.050 675.450 527.400 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 661.950 524.250 663.750 525.150 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 668.250 524.250 670.050 525.150 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 524.250 678.750 525.150 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 683.250 524.250 685.050 525.150 ;
        RECT 665.250 521.850 666.750 522.750 ;
        RECT 655.950 517.950 658.050 520.050 ;
        RECT 652.950 511.950 655.050 514.050 ;
        RECT 661.950 488.250 664.050 489.150 ;
        RECT 652.950 485.250 654.750 486.150 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 659.250 485.250 660.750 486.150 ;
        RECT 661.950 484.950 664.050 487.050 ;
        RECT 667.950 486.450 670.050 487.050 ;
        RECT 671.400 486.450 672.450 523.950 ;
        RECT 680.250 521.850 681.750 522.750 ;
        RECT 676.950 517.950 679.050 520.050 ;
        RECT 673.950 495.300 676.050 497.400 ;
        RECT 674.550 491.700 675.750 495.300 ;
        RECT 673.950 489.600 676.050 491.700 ;
        RECT 667.950 485.400 672.450 486.450 ;
        RECT 667.950 484.950 670.050 485.400 ;
        RECT 656.250 482.850 657.750 483.750 ;
        RECT 658.950 481.950 661.050 484.050 ;
        RECT 670.950 483.450 673.050 484.050 ;
        RECT 668.400 482.400 673.050 483.450 ;
        RECT 637.950 475.950 640.050 478.050 ;
        RECT 649.950 475.950 652.050 478.050 ;
        RECT 655.950 475.950 658.050 478.050 ;
        RECT 640.950 469.950 643.050 472.050 ;
        RECT 637.950 466.950 640.050 469.050 ;
        RECT 628.950 463.950 631.050 466.050 ;
        RECT 631.950 460.950 634.050 463.050 ;
        RECT 632.400 457.050 633.450 460.950 ;
        RECT 622.950 454.950 625.050 457.050 ;
        RECT 631.950 454.950 634.050 457.050 ;
        RECT 632.400 454.050 633.450 454.950 ;
        RECT 625.950 453.450 628.050 454.050 ;
        RECT 623.400 452.400 628.050 453.450 ;
        RECT 623.400 418.050 624.450 452.400 ;
        RECT 625.950 451.950 628.050 452.400 ;
        RECT 631.950 451.950 634.050 454.050 ;
        RECT 635.250 452.250 637.050 453.150 ;
        RECT 625.950 449.850 627.750 450.750 ;
        RECT 628.950 448.950 631.050 451.050 ;
        RECT 632.250 449.850 633.750 450.750 ;
        RECT 634.950 448.950 637.050 451.050 ;
        RECT 635.400 448.050 636.450 448.950 ;
        RECT 628.950 446.850 631.050 447.750 ;
        RECT 634.950 445.950 637.050 448.050 ;
        RECT 638.400 424.050 639.450 466.950 ;
        RECT 637.950 421.950 640.050 424.050 ;
        RECT 638.400 418.050 639.450 421.950 ;
        RECT 622.950 415.950 625.050 418.050 ;
        RECT 625.950 415.950 628.050 418.050 ;
        RECT 629.250 416.250 630.750 417.150 ;
        RECT 631.950 415.950 634.050 418.050 ;
        RECT 637.950 415.950 640.050 418.050 ;
        RECT 625.950 413.850 627.750 414.750 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 632.250 413.850 634.050 414.750 ;
        RECT 634.950 412.950 637.050 415.050 ;
        RECT 635.400 409.050 636.450 412.950 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 634.950 406.950 637.050 409.050 ;
        RECT 607.950 403.950 610.050 406.050 ;
        RECT 613.950 403.950 616.050 406.050 ;
        RECT 619.950 403.950 622.050 406.050 ;
        RECT 610.950 379.950 613.050 382.050 ;
        RECT 604.950 376.950 607.050 379.050 ;
        RECT 610.950 377.850 613.050 378.750 ;
        RECT 601.950 370.950 604.050 373.050 ;
        RECT 614.400 361.050 615.450 403.950 ;
        RECT 619.950 389.400 622.050 391.500 ;
        RECT 622.950 389.400 625.050 391.500 ;
        RECT 625.950 389.400 628.050 391.500 ;
        RECT 630.750 389.400 632.850 391.500 ;
        RECT 634.950 389.400 637.050 391.500 ;
        RECT 620.550 375.750 621.750 389.400 ;
        RECT 619.950 373.650 622.050 375.750 ;
        RECT 620.550 369.900 621.750 373.650 ;
        RECT 623.250 372.150 624.450 389.400 ;
        RECT 626.400 375.750 627.600 389.400 ;
        RECT 631.350 383.550 632.550 389.400 ;
        RECT 630.750 381.450 632.850 383.550 ;
        RECT 625.950 373.650 628.050 375.750 ;
        RECT 631.350 372.600 632.550 381.450 ;
        RECT 635.550 380.850 636.750 389.400 ;
        RECT 638.400 388.050 639.450 409.950 ;
        RECT 637.950 385.950 640.050 388.050 ;
        RECT 637.950 383.850 640.050 384.750 ;
        RECT 634.950 378.750 637.050 380.850 ;
        RECT 637.950 379.950 640.050 382.050 ;
        RECT 635.550 372.600 636.750 378.750 ;
        RECT 622.950 370.050 625.050 372.150 ;
        RECT 630.900 370.500 633.000 372.600 ;
        RECT 634.950 370.500 637.050 372.600 ;
        RECT 619.800 367.800 621.900 369.900 ;
        RECT 613.950 358.950 616.050 361.050 ;
        RECT 598.950 352.950 601.050 355.050 ;
        RECT 604.800 353.100 606.900 355.200 ;
        RECT 596.400 350.400 600.450 351.450 ;
        RECT 593.400 342.450 594.450 349.950 ;
        RECT 595.950 344.250 598.050 345.150 ;
        RECT 595.950 342.450 598.050 343.050 ;
        RECT 593.400 341.400 598.050 342.450 ;
        RECT 593.400 325.050 594.450 341.400 ;
        RECT 595.950 340.950 598.050 341.400 ;
        RECT 592.950 322.950 595.050 325.050 ;
        RECT 592.950 311.250 594.750 312.150 ;
        RECT 595.950 310.950 598.050 313.050 ;
        RECT 599.400 310.050 600.450 350.400 ;
        RECT 605.550 349.350 606.750 353.100 ;
        RECT 628.950 352.950 631.050 355.050 ;
        RECT 631.950 352.950 634.050 355.050 ;
        RECT 634.950 352.950 637.050 355.050 ;
        RECT 607.950 350.850 610.050 352.950 ;
        RECT 604.950 347.250 607.050 349.350 ;
        RECT 601.950 343.950 604.050 346.050 ;
        RECT 602.400 313.050 603.450 343.950 ;
        RECT 605.550 333.600 606.750 347.250 ;
        RECT 608.250 333.600 609.450 350.850 ;
        RECT 615.900 350.400 618.000 352.500 ;
        RECT 619.950 350.400 622.050 352.500 ;
        RECT 610.950 347.250 613.050 349.350 ;
        RECT 611.400 333.600 612.600 347.250 ;
        RECT 616.350 341.550 617.550 350.400 ;
        RECT 620.550 344.250 621.750 350.400 ;
        RECT 619.950 342.150 622.050 344.250 ;
        RECT 615.750 339.450 617.850 341.550 ;
        RECT 616.350 333.600 617.550 339.450 ;
        RECT 620.550 333.600 621.750 342.150 ;
        RECT 622.950 338.250 625.050 339.150 ;
        RECT 625.950 337.950 628.050 340.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 604.950 331.500 607.050 333.600 ;
        RECT 607.950 331.500 610.050 333.600 ;
        RECT 610.950 331.500 613.050 333.600 ;
        RECT 615.750 331.500 617.850 333.600 ;
        RECT 619.950 331.500 622.050 333.600 ;
        RECT 604.950 322.950 607.050 325.050 ;
        RECT 601.950 310.950 604.050 313.050 ;
        RECT 592.950 309.450 595.050 310.050 ;
        RECT 590.400 308.400 595.050 309.450 ;
        RECT 596.250 308.850 598.050 309.750 ;
        RECT 592.950 307.950 595.050 308.400 ;
        RECT 598.950 307.950 601.050 310.050 ;
        RECT 601.950 307.950 604.050 310.050 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 590.400 301.050 591.450 304.950 ;
        RECT 586.950 298.950 589.050 301.050 ;
        RECT 589.950 298.950 592.050 301.050 ;
        RECT 590.400 297.450 591.450 298.950 ;
        RECT 587.400 296.400 591.450 297.450 ;
        RECT 587.400 274.050 588.450 296.400 ;
        RECT 593.400 274.050 594.450 307.950 ;
        RECT 602.400 279.450 603.450 307.950 ;
        RECT 605.400 283.050 606.450 322.950 ;
        RECT 607.950 316.950 610.050 319.050 ;
        RECT 608.400 307.050 609.450 316.950 ;
        RECT 610.950 313.950 613.050 316.050 ;
        RECT 607.950 304.950 610.050 307.050 ;
        RECT 604.950 280.950 607.050 283.050 ;
        RECT 607.950 280.950 610.050 283.050 ;
        RECT 602.400 278.400 606.450 279.450 ;
        RECT 601.950 274.950 604.050 277.050 ;
        RECT 586.950 271.950 589.050 274.050 ;
        RECT 592.950 271.950 595.050 274.050 ;
        RECT 598.950 272.250 601.050 273.150 ;
        RECT 589.950 269.250 591.750 270.150 ;
        RECT 592.950 268.950 595.050 271.050 ;
        RECT 596.250 269.250 597.750 270.150 ;
        RECT 598.950 268.950 601.050 271.050 ;
        RECT 589.950 265.950 592.050 268.050 ;
        RECT 593.250 266.850 594.750 267.750 ;
        RECT 595.950 265.950 598.050 268.050 ;
        RECT 598.950 265.950 601.050 268.050 ;
        RECT 592.950 259.950 595.050 262.050 ;
        RECT 583.950 253.950 586.050 256.050 ;
        RECT 586.950 247.950 589.050 250.050 ;
        RECT 587.400 241.050 588.450 247.950 ;
        RECT 586.950 238.950 589.050 241.050 ;
        RECT 580.950 236.850 583.050 237.750 ;
        RECT 583.950 235.950 586.050 238.050 ;
        RECT 586.950 236.850 589.050 237.750 ;
        RECT 577.950 226.950 580.050 229.050 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 574.950 211.950 577.050 214.050 ;
        RECT 547.950 208.950 550.050 211.050 ;
        RECT 553.950 208.950 556.050 211.050 ;
        RECT 547.950 199.950 550.050 202.050 ;
        RECT 548.400 199.050 549.450 199.950 ;
        RECT 554.400 199.050 555.450 208.950 ;
        RECT 559.950 205.950 562.050 208.050 ;
        RECT 565.950 205.950 568.050 208.050 ;
        RECT 556.950 199.950 559.050 202.050 ;
        RECT 544.950 197.250 546.750 198.150 ;
        RECT 547.950 196.950 550.050 199.050 ;
        RECT 553.950 196.950 556.050 199.050 ;
        RECT 544.950 193.950 547.050 196.050 ;
        RECT 548.250 194.850 550.050 195.750 ;
        RECT 550.950 194.250 553.050 195.150 ;
        RECT 553.950 194.850 556.050 195.750 ;
        RECT 545.400 183.450 546.450 193.950 ;
        RECT 550.950 190.950 553.050 193.050 ;
        RECT 557.400 190.050 558.450 199.950 ;
        RECT 560.400 193.050 561.450 205.950 ;
        RECT 566.400 199.050 567.450 205.950 ;
        RECT 571.950 200.250 574.050 201.150 ;
        RECT 562.950 197.250 564.750 198.150 ;
        RECT 565.950 196.950 568.050 199.050 ;
        RECT 569.250 197.250 570.750 198.150 ;
        RECT 571.950 196.950 574.050 199.050 ;
        RECT 562.950 193.950 565.050 196.050 ;
        RECT 566.250 194.850 567.750 195.750 ;
        RECT 568.950 193.950 571.050 196.050 ;
        RECT 559.950 190.950 562.050 193.050 ;
        RECT 569.400 190.050 570.450 193.950 ;
        RECT 556.950 187.950 559.050 190.050 ;
        RECT 568.950 187.950 571.050 190.050 ;
        RECT 572.400 184.050 573.450 196.950 ;
        RECT 545.400 182.400 549.450 183.450 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 538.950 175.950 541.050 178.050 ;
        RECT 532.950 172.950 535.050 175.050 ;
        RECT 529.950 169.950 532.050 172.050 ;
        RECT 526.950 148.950 529.050 151.050 ;
        RECT 523.950 145.950 526.050 148.050 ;
        RECT 520.950 127.950 523.050 130.050 ;
        RECT 524.400 123.450 525.450 145.950 ;
        RECT 530.400 139.050 531.450 169.950 ;
        RECT 545.400 169.050 546.450 178.950 ;
        RECT 538.950 166.950 541.050 169.050 ;
        RECT 542.250 167.250 543.750 168.150 ;
        RECT 544.950 166.950 547.050 169.050 ;
        RECT 548.400 166.050 549.450 182.400 ;
        RECT 571.950 181.950 574.050 184.050 ;
        RECT 556.950 178.950 559.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 550.950 175.950 553.050 178.050 ;
        RECT 535.950 163.950 538.050 166.050 ;
        RECT 539.250 164.850 540.750 165.750 ;
        RECT 541.950 163.950 544.050 166.050 ;
        RECT 545.250 164.850 547.050 165.750 ;
        RECT 547.950 163.950 550.050 166.050 ;
        RECT 535.950 161.850 538.050 162.750 ;
        RECT 538.950 160.950 541.050 163.050 ;
        RECT 529.950 136.950 532.050 139.050 ;
        RECT 526.950 125.250 529.050 126.150 ;
        RECT 532.950 125.250 535.050 126.150 ;
        RECT 526.950 123.450 529.050 124.050 ;
        RECT 524.400 122.400 529.050 123.450 ;
        RECT 526.950 121.950 529.050 122.400 ;
        RECT 530.250 122.250 531.750 123.150 ;
        RECT 532.950 121.950 535.050 124.050 ;
        RECT 533.400 121.050 534.450 121.950 ;
        RECT 529.950 118.950 532.050 121.050 ;
        RECT 532.950 118.950 535.050 121.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 533.400 97.050 534.450 100.950 ;
        RECT 539.400 99.450 540.450 160.950 ;
        RECT 548.400 157.050 549.450 163.950 ;
        RECT 547.950 154.950 550.050 157.050 ;
        RECT 547.950 136.950 550.050 139.050 ;
        RECT 548.400 127.050 549.450 136.950 ;
        RECT 551.400 127.050 552.450 175.950 ;
        RECT 553.950 166.950 556.050 169.050 ;
        RECT 554.400 163.050 555.450 166.950 ;
        RECT 557.400 166.050 558.450 178.950 ;
        RECT 566.400 169.050 567.450 178.950 ;
        RECT 559.950 166.950 562.050 169.050 ;
        RECT 565.950 168.450 568.050 169.050 ;
        RECT 575.400 168.450 576.450 211.950 ;
        RECT 584.400 184.050 585.450 235.950 ;
        RECT 593.400 214.050 594.450 259.950 ;
        RECT 596.400 256.050 597.450 265.950 ;
        RECT 595.950 253.950 598.050 256.050 ;
        RECT 599.400 250.050 600.450 265.950 ;
        RECT 598.950 247.950 601.050 250.050 ;
        RECT 595.950 241.950 598.050 244.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 586.950 202.950 589.050 205.050 ;
        RECT 587.400 199.050 588.450 202.950 ;
        RECT 586.950 196.950 589.050 199.050 ;
        RECT 586.950 194.850 589.050 195.750 ;
        RECT 589.950 194.250 592.050 195.150 ;
        RECT 589.950 190.950 592.050 193.050 ;
        RECT 583.950 181.950 586.050 184.050 ;
        RECT 577.950 169.950 580.050 172.050 ;
        RECT 563.250 167.250 564.750 168.150 ;
        RECT 565.950 167.400 570.450 168.450 ;
        RECT 565.950 166.950 568.050 167.400 ;
        RECT 556.950 163.950 559.050 166.050 ;
        RECT 560.250 164.850 561.750 165.750 ;
        RECT 562.950 163.950 565.050 166.050 ;
        RECT 566.250 164.850 568.050 165.750 ;
        RECT 553.950 160.950 556.050 163.050 ;
        RECT 556.950 161.850 559.050 162.750 ;
        RECT 563.400 157.050 564.450 163.950 ;
        RECT 569.400 163.050 570.450 167.400 ;
        RECT 572.400 167.400 576.450 168.450 ;
        RECT 568.950 160.950 571.050 163.050 ;
        RECT 562.950 154.950 565.050 157.050 ;
        RECT 553.950 145.950 556.050 148.050 ;
        RECT 554.400 127.050 555.450 145.950 ;
        RECT 572.400 138.450 573.450 167.400 ;
        RECT 578.400 166.050 579.450 169.950 ;
        RECT 583.950 166.950 586.050 169.050 ;
        RECT 574.950 164.250 576.750 165.150 ;
        RECT 577.950 163.950 580.050 166.050 ;
        RECT 581.250 164.250 583.050 165.150 ;
        RECT 574.950 160.950 577.050 163.050 ;
        RECT 578.250 161.850 579.750 162.750 ;
        RECT 580.950 160.950 583.050 163.050 ;
        RECT 569.400 137.400 573.450 138.450 ;
        RECT 556.950 127.950 559.050 130.050 ;
        RECT 544.950 125.250 546.750 126.150 ;
        RECT 547.950 124.950 550.050 127.050 ;
        RECT 550.950 124.950 553.050 127.050 ;
        RECT 553.950 124.950 556.050 127.050 ;
        RECT 544.950 121.950 547.050 124.050 ;
        RECT 548.250 122.850 550.050 123.750 ;
        RECT 550.950 122.250 553.050 123.150 ;
        RECT 553.950 122.850 556.050 123.750 ;
        RECT 545.400 102.450 546.450 121.950 ;
        RECT 550.950 118.950 553.050 121.050 ;
        RECT 536.400 98.400 540.450 99.450 ;
        RECT 542.400 101.400 546.450 102.450 ;
        RECT 526.950 94.950 529.050 97.050 ;
        RECT 530.250 95.250 531.750 96.150 ;
        RECT 532.950 94.950 535.050 97.050 ;
        RECT 523.950 91.950 526.050 94.050 ;
        RECT 527.250 92.850 528.750 93.750 ;
        RECT 529.950 91.950 532.050 94.050 ;
        RECT 533.250 92.850 535.050 93.750 ;
        RECT 523.950 89.850 526.050 90.750 ;
        RECT 523.950 64.950 526.050 67.050 ;
        RECT 524.400 61.050 525.450 64.950 ;
        RECT 536.400 61.050 537.450 98.400 ;
        RECT 542.400 97.050 543.450 101.400 ;
        RECT 544.950 97.950 547.050 100.050 ;
        RECT 538.950 94.950 541.050 97.050 ;
        RECT 541.950 94.950 544.050 97.050 ;
        RECT 539.400 90.450 540.450 94.950 ;
        RECT 545.400 94.050 546.450 97.950 ;
        RECT 550.950 94.950 553.050 97.050 ;
        RECT 553.950 94.950 556.050 97.050 ;
        RECT 541.950 92.250 543.750 93.150 ;
        RECT 544.950 91.950 547.050 94.050 ;
        RECT 548.250 92.250 550.050 93.150 ;
        RECT 541.950 90.450 544.050 91.050 ;
        RECT 539.400 89.400 544.050 90.450 ;
        RECT 545.250 89.850 546.750 90.750 ;
        RECT 541.950 88.950 544.050 89.400 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 523.950 58.950 526.050 61.050 ;
        RECT 535.950 58.950 538.050 61.050 ;
        RECT 538.950 58.950 541.050 61.050 ;
        RECT 511.950 52.950 514.050 55.050 ;
        RECT 517.950 52.950 520.050 55.050 ;
        RECT 511.950 50.850 514.050 51.750 ;
        RECT 524.400 51.450 525.450 58.950 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 535.950 56.250 538.050 57.150 ;
        RECT 530.400 55.050 531.450 55.950 ;
        RECT 526.950 53.250 528.750 54.150 ;
        RECT 529.950 52.950 532.050 55.050 ;
        RECT 535.950 54.450 538.050 55.050 ;
        RECT 539.400 54.450 540.450 58.950 ;
        RECT 551.400 58.050 552.450 94.950 ;
        RECT 554.400 94.050 555.450 94.950 ;
        RECT 553.950 91.950 556.050 94.050 ;
        RECT 553.950 67.950 556.050 70.050 ;
        RECT 550.950 55.950 553.050 58.050 ;
        RECT 554.400 55.050 555.450 67.950 ;
        RECT 557.400 57.450 558.450 127.950 ;
        RECT 569.400 127.050 570.450 137.400 ;
        RECT 571.950 133.950 574.050 136.050 ;
        RECT 559.950 124.950 562.050 127.050 ;
        RECT 565.950 126.450 568.050 127.050 ;
        RECT 563.400 125.400 568.050 126.450 ;
        RECT 560.400 97.050 561.450 124.950 ;
        RECT 563.400 121.050 564.450 125.400 ;
        RECT 565.950 124.950 568.050 125.400 ;
        RECT 568.950 124.950 571.050 127.050 ;
        RECT 565.950 122.850 568.050 123.750 ;
        RECT 568.950 122.250 571.050 123.150 ;
        RECT 562.950 118.950 565.050 121.050 ;
        RECT 568.950 118.950 571.050 121.050 ;
        RECT 572.400 100.050 573.450 133.950 ;
        RECT 575.400 129.450 576.450 160.950 ;
        RECT 581.400 136.050 582.450 160.950 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 584.400 130.050 585.450 166.950 ;
        RECT 586.950 163.950 589.050 166.050 ;
        RECT 587.400 154.050 588.450 163.950 ;
        RECT 590.400 162.450 591.450 190.950 ;
        RECT 596.400 169.050 597.450 241.950 ;
        RECT 602.400 241.050 603.450 274.950 ;
        RECT 598.950 238.950 601.050 241.050 ;
        RECT 601.950 238.950 604.050 241.050 ;
        RECT 598.950 236.850 601.050 237.750 ;
        RECT 601.950 236.250 604.050 237.150 ;
        RECT 601.950 234.450 604.050 235.050 ;
        RECT 605.400 234.450 606.450 278.400 ;
        RECT 608.400 241.050 609.450 280.950 ;
        RECT 611.400 253.050 612.450 313.950 ;
        RECT 613.950 310.950 616.050 313.050 ;
        RECT 619.950 310.950 622.050 313.050 ;
        RECT 622.950 312.450 625.050 313.050 ;
        RECT 626.400 312.450 627.450 337.950 ;
        RECT 629.250 334.050 630.450 352.950 ;
        RECT 632.250 348.750 633.450 352.950 ;
        RECT 631.950 346.650 634.050 348.750 ;
        RECT 632.250 334.050 633.450 346.650 ;
        RECT 635.250 334.050 636.450 352.950 ;
        RECT 638.400 352.050 639.450 379.950 ;
        RECT 637.950 349.950 640.050 352.050 ;
        RECT 641.400 348.450 642.450 469.950 ;
        RECT 649.950 463.950 652.050 466.050 ;
        RECT 646.950 461.400 649.050 463.500 ;
        RECT 643.950 457.950 646.050 460.050 ;
        RECT 644.400 421.050 645.450 457.950 ;
        RECT 647.400 444.600 648.600 461.400 ;
        RECT 646.950 442.500 649.050 444.600 ;
        RECT 643.950 418.950 646.050 421.050 ;
        RECT 644.400 415.050 645.450 418.950 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 647.250 413.250 649.050 414.150 ;
        RECT 643.950 410.850 645.750 411.750 ;
        RECT 646.950 411.450 649.050 412.050 ;
        RECT 650.400 411.450 651.450 463.950 ;
        RECT 652.950 457.950 655.050 460.050 ;
        RECT 653.400 457.050 654.450 457.950 ;
        RECT 652.950 454.950 655.050 457.050 ;
        RECT 652.950 452.850 655.050 453.750 ;
        RECT 656.400 451.050 657.450 475.950 ;
        RECT 659.400 460.050 660.450 481.950 ;
        RECT 661.950 475.950 664.050 478.050 ;
        RECT 662.400 475.050 663.450 475.950 ;
        RECT 661.950 472.950 664.050 475.050 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 658.950 456.450 661.050 457.050 ;
        RECT 662.400 456.450 663.450 472.950 ;
        RECT 668.400 469.050 669.450 482.400 ;
        RECT 670.950 481.950 673.050 482.400 ;
        RECT 670.950 479.850 673.050 480.750 ;
        RECT 674.550 477.600 675.750 489.600 ;
        RECT 673.950 475.500 676.050 477.600 ;
        RECT 667.950 466.950 670.050 469.050 ;
        RECT 667.950 461.400 670.050 463.500 ;
        RECT 658.950 455.400 663.450 456.450 ;
        RECT 658.950 454.950 661.050 455.400 ;
        RECT 664.950 454.950 667.050 457.050 ;
        RECT 658.950 452.850 661.050 453.750 ;
        RECT 652.950 448.950 655.050 451.050 ;
        RECT 655.950 448.950 658.050 451.050 ;
        RECT 646.950 410.400 651.450 411.450 ;
        RECT 646.950 409.950 649.050 410.400 ;
        RECT 643.950 388.950 646.050 391.050 ;
        RECT 646.950 388.950 649.050 391.050 ;
        RECT 649.950 388.950 652.050 391.050 ;
        RECT 644.250 370.050 645.450 388.950 ;
        RECT 647.250 376.350 648.450 388.950 ;
        RECT 646.950 374.250 649.050 376.350 ;
        RECT 647.250 370.050 648.450 374.250 ;
        RECT 650.250 370.050 651.450 388.950 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 646.950 367.950 649.050 370.050 ;
        RECT 649.950 367.950 652.050 370.050 ;
        RECT 646.950 364.950 649.050 367.050 ;
        RECT 653.400 366.450 654.450 448.950 ;
        RECT 661.950 439.950 664.050 442.050 ;
        RECT 662.400 415.050 663.450 439.950 ;
        RECT 661.950 412.950 664.050 415.050 ;
        RECT 658.950 410.250 661.050 411.150 ;
        RECT 661.950 410.850 664.050 411.750 ;
        RECT 658.950 406.950 661.050 409.050 ;
        RECT 661.950 380.250 664.050 381.150 ;
        RECT 655.950 377.850 658.050 378.750 ;
        RECT 661.950 376.950 664.050 379.050 ;
        RECT 662.400 367.050 663.450 376.950 ;
        RECT 650.400 365.400 654.450 366.450 ;
        RECT 638.400 347.400 642.450 348.450 ;
        RECT 628.950 331.950 631.050 334.050 ;
        RECT 631.950 331.950 634.050 334.050 ;
        RECT 634.950 331.950 637.050 334.050 ;
        RECT 638.400 316.050 639.450 347.400 ;
        RECT 647.400 346.050 648.450 364.950 ;
        RECT 646.950 345.450 649.050 346.050 ;
        RECT 640.950 344.250 643.050 345.150 ;
        RECT 644.400 344.400 649.050 345.450 ;
        RECT 637.950 313.950 640.050 316.050 ;
        RECT 622.950 311.400 627.450 312.450 ;
        RECT 622.950 310.950 625.050 311.400 ;
        RECT 613.950 308.850 616.050 309.750 ;
        RECT 616.950 308.250 619.050 309.150 ;
        RECT 616.950 304.950 619.050 307.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 614.400 274.050 615.450 289.950 ;
        RECT 617.400 277.050 618.450 304.950 ;
        RECT 620.400 286.050 621.450 310.950 ;
        RECT 622.950 308.850 625.050 309.750 ;
        RECT 622.950 286.950 625.050 289.050 ;
        RECT 619.950 283.950 622.050 286.050 ;
        RECT 616.950 274.950 619.050 277.050 ;
        RECT 613.950 271.950 616.050 274.050 ;
        RECT 617.250 272.250 618.750 273.150 ;
        RECT 619.950 271.950 622.050 274.050 ;
        RECT 613.950 269.850 615.750 270.750 ;
        RECT 616.950 268.950 619.050 271.050 ;
        RECT 620.250 269.850 622.050 270.750 ;
        RECT 623.400 268.050 624.450 286.950 ;
        RECT 626.400 283.050 627.450 311.400 ;
        RECT 631.950 310.950 634.050 313.050 ;
        RECT 628.950 307.950 631.050 310.050 ;
        RECT 625.950 280.950 628.050 283.050 ;
        RECT 625.950 274.950 628.050 277.050 ;
        RECT 622.950 265.950 625.050 268.050 ;
        RECT 613.950 253.950 616.050 256.050 ;
        RECT 610.950 250.950 613.050 253.050 ;
        RECT 610.950 244.950 613.050 247.050 ;
        RECT 607.950 238.950 610.050 241.050 ;
        RECT 607.950 236.850 610.050 237.750 ;
        RECT 601.950 233.400 606.450 234.450 ;
        RECT 601.950 232.950 604.050 233.400 ;
        RECT 602.400 223.050 603.450 232.950 ;
        RECT 601.950 220.950 604.050 223.050 ;
        RECT 611.400 205.050 612.450 244.950 ;
        RECT 610.950 202.950 613.050 205.050 ;
        RECT 601.950 200.250 604.050 201.150 ;
        RECT 614.400 199.050 615.450 253.950 ;
        RECT 619.950 238.950 622.050 241.050 ;
        RECT 620.400 238.050 621.450 238.950 ;
        RECT 616.950 236.250 618.750 237.150 ;
        RECT 619.950 235.950 622.050 238.050 ;
        RECT 623.250 236.250 625.050 237.150 ;
        RECT 616.950 232.950 619.050 235.050 ;
        RECT 620.250 233.850 621.750 234.750 ;
        RECT 622.950 232.950 625.050 235.050 ;
        RECT 617.400 229.050 618.450 232.950 ;
        RECT 616.950 226.950 619.050 229.050 ;
        RECT 626.400 208.050 627.450 274.950 ;
        RECT 629.400 267.450 630.450 307.950 ;
        RECT 632.400 306.450 633.450 310.950 ;
        RECT 634.950 308.250 636.750 309.150 ;
        RECT 637.950 307.950 640.050 310.050 ;
        RECT 641.250 308.250 643.050 309.150 ;
        RECT 634.950 306.450 637.050 307.050 ;
        RECT 632.400 305.400 637.050 306.450 ;
        RECT 638.250 305.850 639.750 306.750 ;
        RECT 634.950 304.950 637.050 305.400 ;
        RECT 640.950 304.950 643.050 307.050 ;
        RECT 641.400 304.050 642.450 304.950 ;
        RECT 640.950 301.950 643.050 304.050 ;
        RECT 644.400 298.050 645.450 344.400 ;
        RECT 646.950 343.950 649.050 344.400 ;
        RECT 646.950 341.850 649.050 342.750 ;
        RECT 650.400 324.450 651.450 365.400 ;
        RECT 661.950 364.950 664.050 367.050 ;
        RECT 661.950 358.950 664.050 361.050 ;
        RECT 655.950 346.950 658.050 349.050 ;
        RECT 656.400 334.050 657.450 346.950 ;
        RECT 658.950 341.250 661.050 342.150 ;
        RECT 658.950 337.950 661.050 340.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 647.400 323.400 651.450 324.450 ;
        RECT 643.950 295.950 646.050 298.050 ;
        RECT 644.400 295.050 645.450 295.950 ;
        RECT 643.950 292.950 646.050 295.050 ;
        RECT 647.400 289.050 648.450 323.400 ;
        RECT 662.400 313.050 663.450 358.950 ;
        RECT 665.400 349.050 666.450 454.950 ;
        RECT 668.250 449.400 669.450 461.400 ;
        RECT 670.950 458.250 673.050 459.150 ;
        RECT 670.950 454.950 673.050 457.050 ;
        RECT 667.950 447.300 670.050 449.400 ;
        RECT 668.250 443.700 669.450 447.300 ;
        RECT 667.950 441.600 670.050 443.700 ;
        RECT 667.950 424.950 670.050 427.050 ;
        RECT 668.400 411.450 669.450 424.950 ;
        RECT 673.950 423.300 676.050 425.400 ;
        RECT 674.550 419.700 675.750 423.300 ;
        RECT 673.950 417.600 676.050 419.700 ;
        RECT 670.950 411.450 673.050 412.050 ;
        RECT 668.400 410.400 673.050 411.450 ;
        RECT 668.400 376.050 669.450 410.400 ;
        RECT 670.950 409.950 673.050 410.400 ;
        RECT 670.950 407.850 673.050 408.750 ;
        RECT 674.550 405.600 675.750 417.600 ;
        RECT 673.950 403.500 676.050 405.600 ;
        RECT 677.400 400.050 678.450 517.950 ;
        RECT 689.400 508.050 690.450 551.400 ;
        RECT 694.950 550.950 697.050 553.050 ;
        RECT 712.950 547.950 715.050 550.050 ;
        RECT 700.950 538.950 703.050 541.050 ;
        RECT 709.950 538.950 712.050 541.050 ;
        RECT 694.950 533.400 697.050 535.500 ;
        RECT 691.950 530.250 694.050 531.150 ;
        RECT 691.950 526.950 694.050 529.050 ;
        RECT 692.400 520.050 693.450 526.950 ;
        RECT 695.550 521.400 696.750 533.400 ;
        RECT 697.950 532.950 700.050 535.050 ;
        RECT 691.950 517.950 694.050 520.050 ;
        RECT 694.950 519.300 697.050 521.400 ;
        RECT 695.550 515.700 696.750 519.300 ;
        RECT 694.950 513.600 697.050 515.700 ;
        RECT 688.950 505.950 691.050 508.050 ;
        RECT 694.950 494.400 697.050 496.500 ;
        RECT 682.950 485.250 685.050 486.150 ;
        RECT 688.950 485.250 691.050 486.150 ;
        RECT 682.950 481.950 685.050 484.050 ;
        RECT 688.950 481.950 691.050 484.050 ;
        RECT 683.400 478.050 684.450 481.950 ;
        RECT 682.950 475.950 685.050 478.050 ;
        RECT 695.400 477.600 696.600 494.400 ;
        RECT 698.400 481.050 699.450 532.950 ;
        RECT 701.400 532.050 702.450 538.950 ;
        RECT 700.950 529.950 703.050 532.050 ;
        RECT 703.950 529.950 706.050 532.050 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 701.400 478.050 702.450 529.950 ;
        RECT 704.400 529.050 705.450 529.950 ;
        RECT 710.400 529.050 711.450 538.950 ;
        RECT 703.950 526.950 706.050 529.050 ;
        RECT 709.950 526.950 712.050 529.050 ;
        RECT 703.950 524.850 706.050 525.750 ;
        RECT 709.950 524.850 712.050 525.750 ;
        RECT 713.400 487.050 714.450 547.950 ;
        RECT 716.400 541.050 717.450 553.950 ;
        RECT 715.950 538.950 718.050 541.050 ;
        RECT 715.950 533.400 718.050 535.500 ;
        RECT 716.400 516.600 717.600 533.400 ;
        RECT 722.400 517.050 723.450 577.950 ;
        RECT 725.400 562.050 726.450 665.400 ;
        RECT 727.950 664.950 730.050 665.400 ;
        RECT 733.950 664.950 736.050 667.050 ;
        RECT 739.950 664.950 742.050 667.050 ;
        RECT 749.400 664.050 750.450 667.950 ;
        RECT 751.950 664.950 754.050 667.050 ;
        RECT 754.950 665.850 757.050 666.750 ;
        RECT 748.950 661.950 751.050 664.050 ;
        RECT 739.950 658.950 742.050 661.050 ;
        RECT 736.950 643.950 739.050 646.050 ;
        RECT 727.950 629.250 730.050 630.150 ;
        RECT 733.950 629.250 736.050 630.150 ;
        RECT 727.950 625.950 730.050 628.050 ;
        RECT 733.950 627.450 736.050 628.050 ;
        RECT 737.400 627.450 738.450 643.950 ;
        RECT 731.250 626.250 732.750 627.150 ;
        RECT 733.950 626.400 738.450 627.450 ;
        RECT 733.950 625.950 736.050 626.400 ;
        RECT 728.400 625.050 729.450 625.950 ;
        RECT 727.950 622.950 730.050 625.050 ;
        RECT 730.950 622.950 733.050 625.050 ;
        RECT 728.400 583.050 729.450 622.950 ;
        RECT 740.400 616.050 741.450 658.950 ;
        RECT 748.950 628.950 751.050 631.050 ;
        RECT 745.950 626.250 748.050 627.150 ;
        RECT 748.950 626.850 751.050 627.750 ;
        RECT 745.950 622.950 748.050 625.050 ;
        RECT 739.950 613.950 742.050 616.050 ;
        RECT 736.950 601.950 739.050 604.050 ;
        RECT 737.400 598.050 738.450 601.950 ;
        RECT 746.400 601.050 747.450 622.950 ;
        RECT 752.400 604.050 753.450 664.950 ;
        RECT 758.400 664.050 759.450 668.400 ;
        RECT 757.950 661.950 760.050 664.050 ;
        RECT 757.950 631.950 760.050 634.050 ;
        RECT 758.400 625.050 759.450 631.950 ;
        RECT 757.950 622.950 760.050 625.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 745.950 598.950 748.050 601.050 ;
        RECT 751.950 599.850 754.050 600.750 ;
        RECT 754.950 599.250 757.050 600.150 ;
        RECT 730.950 595.950 733.050 598.050 ;
        RECT 733.950 595.950 736.050 598.050 ;
        RECT 736.950 595.950 739.050 598.050 ;
        RECT 751.950 597.450 754.050 598.050 ;
        RECT 754.950 597.450 757.050 598.050 ;
        RECT 740.250 596.250 742.050 597.150 ;
        RECT 751.950 596.400 757.050 597.450 ;
        RECT 751.950 595.950 754.050 596.400 ;
        RECT 754.950 595.950 757.050 596.400 ;
        RECT 734.400 595.050 735.450 595.950 ;
        RECT 730.950 593.850 732.750 594.750 ;
        RECT 733.950 592.950 736.050 595.050 ;
        RECT 737.250 593.850 738.750 594.750 ;
        RECT 739.950 592.950 742.050 595.050 ;
        RECT 733.950 590.850 736.050 591.750 ;
        RECT 736.950 583.950 739.050 586.050 ;
        RECT 727.950 580.950 730.050 583.050 ;
        RECT 727.950 571.950 730.050 574.050 ;
        RECT 724.950 559.950 727.050 562.050 ;
        RECT 724.950 517.950 727.050 520.050 ;
        RECT 715.950 514.500 718.050 516.600 ;
        RECT 721.950 514.950 724.050 517.050 ;
        RECT 725.400 514.050 726.450 517.950 ;
        RECT 724.950 511.950 727.050 514.050 ;
        RECT 718.950 488.250 721.050 489.150 ;
        RECT 709.950 485.250 711.750 486.150 ;
        RECT 712.950 484.950 715.050 487.050 ;
        RECT 716.250 485.250 717.750 486.150 ;
        RECT 718.950 484.950 721.050 487.050 ;
        RECT 719.400 484.050 720.450 484.950 ;
        RECT 713.250 482.850 714.750 483.750 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 718.950 481.950 721.050 484.050 ;
        RECT 718.950 478.950 721.050 481.050 ;
        RECT 694.950 475.500 697.050 477.600 ;
        RECT 700.950 475.950 703.050 478.050 ;
        RECT 689.250 455.250 690.750 456.150 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 703.950 454.950 706.050 457.050 ;
        RECT 710.250 455.250 711.750 456.150 ;
        RECT 712.950 454.950 715.050 457.050 ;
        RECT 715.950 454.950 718.050 457.050 ;
        RECT 679.950 451.950 682.050 454.050 ;
        RECT 685.950 452.850 687.750 453.750 ;
        RECT 688.950 451.950 691.050 454.050 ;
        RECT 692.250 452.850 693.750 453.750 ;
        RECT 694.950 451.950 697.050 454.050 ;
        RECT 680.400 409.050 681.450 451.950 ;
        RECT 689.400 450.450 690.450 451.950 ;
        RECT 686.400 449.400 690.450 450.450 ;
        RECT 682.950 413.250 685.050 414.150 ;
        RECT 682.950 409.950 685.050 412.050 ;
        RECT 679.950 406.950 682.050 409.050 ;
        RECT 683.400 403.050 684.450 409.950 ;
        RECT 682.950 400.950 685.050 403.050 ;
        RECT 676.950 397.950 679.050 400.050 ;
        RECT 686.400 394.050 687.450 449.400 ;
        RECT 691.950 448.950 694.050 451.050 ;
        RECT 694.950 449.850 697.050 450.750 ;
        RECT 692.400 426.450 693.450 448.950 ;
        RECT 689.400 425.400 693.450 426.450 ;
        RECT 689.400 418.050 690.450 425.400 ;
        RECT 691.950 421.950 694.050 424.050 ;
        RECT 694.950 422.400 697.050 424.500 ;
        RECT 688.950 415.950 691.050 418.050 ;
        RECT 688.950 413.250 691.050 414.150 ;
        RECT 688.950 409.950 691.050 412.050 ;
        RECT 685.950 391.950 688.050 394.050 ;
        RECT 682.950 388.950 685.050 391.050 ;
        RECT 685.950 388.950 688.050 391.050 ;
        RECT 688.950 388.950 691.050 391.050 ;
        RECT 670.950 380.250 673.050 381.150 ;
        RECT 670.950 376.950 673.050 379.050 ;
        RECT 676.950 377.850 679.050 378.750 ;
        RECT 667.950 373.950 670.050 376.050 ;
        RECT 668.400 373.050 669.450 373.950 ;
        RECT 667.950 370.950 670.050 373.050 ;
        RECT 671.400 367.050 672.450 376.950 ;
        RECT 683.550 370.050 684.750 388.950 ;
        RECT 686.550 376.350 687.750 388.950 ;
        RECT 685.950 374.250 688.050 376.350 ;
        RECT 686.550 370.050 687.750 374.250 ;
        RECT 689.550 370.050 690.750 388.950 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 685.950 367.950 688.050 370.050 ;
        RECT 688.950 367.950 691.050 370.050 ;
        RECT 670.950 364.950 673.050 367.050 ;
        RECT 664.950 346.950 667.050 349.050 ;
        RECT 665.400 346.050 666.450 346.950 ;
        RECT 664.950 343.950 667.050 346.050 ;
        RECT 670.950 343.950 673.050 346.050 ;
        RECT 664.950 341.850 667.050 342.750 ;
        RECT 667.950 341.250 670.050 342.150 ;
        RECT 667.950 339.450 670.050 340.050 ;
        RECT 671.400 339.450 672.450 343.950 ;
        RECT 667.950 338.400 672.450 339.450 ;
        RECT 667.950 337.950 670.050 338.400 ;
        RECT 668.400 321.450 669.450 337.950 ;
        RECT 677.400 322.050 678.450 367.950 ;
        RECT 692.400 358.050 693.450 421.950 ;
        RECT 695.400 405.600 696.600 422.400 ;
        RECT 704.400 412.050 705.450 454.950 ;
        RECT 716.400 454.050 717.450 454.950 ;
        RECT 706.950 452.850 708.750 453.750 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 713.250 452.850 714.750 453.750 ;
        RECT 715.950 451.950 718.050 454.050 ;
        RECT 710.400 442.050 711.450 451.950 ;
        RECT 715.950 449.850 718.050 450.750 ;
        RECT 719.400 445.050 720.450 478.950 ;
        RECT 718.950 442.950 721.050 445.050 ;
        RECT 709.950 439.950 712.050 442.050 ;
        RECT 709.950 422.400 712.050 424.500 ;
        RECT 703.950 409.950 706.050 412.050 ;
        RECT 710.400 405.600 711.600 422.400 ;
        RECT 715.950 413.250 718.050 414.150 ;
        RECT 715.950 409.950 718.050 412.050 ;
        RECT 694.950 403.500 697.050 405.600 ;
        RECT 709.950 403.500 712.050 405.600 ;
        RECT 694.950 388.950 697.050 391.050 ;
        RECT 697.950 389.400 700.050 391.500 ;
        RECT 702.150 389.400 704.250 391.500 ;
        RECT 706.950 389.400 709.050 391.500 ;
        RECT 709.950 389.400 712.050 391.500 ;
        RECT 712.950 389.400 715.050 391.500 ;
        RECT 695.400 388.050 696.450 388.950 ;
        RECT 694.950 385.950 697.050 388.050 ;
        RECT 694.950 383.850 697.050 384.750 ;
        RECT 698.250 380.850 699.450 389.400 ;
        RECT 702.450 383.550 703.650 389.400 ;
        RECT 702.150 381.450 704.250 383.550 ;
        RECT 697.950 378.750 700.050 380.850 ;
        RECT 698.250 372.600 699.450 378.750 ;
        RECT 702.450 372.600 703.650 381.450 ;
        RECT 707.400 375.750 708.600 389.400 ;
        RECT 706.950 373.650 709.050 375.750 ;
        RECT 697.950 370.500 700.050 372.600 ;
        RECT 702.000 370.500 704.100 372.600 ;
        RECT 710.550 372.150 711.750 389.400 ;
        RECT 713.250 375.750 714.450 389.400 ;
        RECT 712.950 373.650 715.050 375.750 ;
        RECT 709.950 370.050 712.050 372.150 ;
        RECT 713.250 369.900 714.450 373.650 ;
        RECT 713.100 367.800 715.200 369.900 ;
        RECT 719.400 366.450 720.450 442.950 ;
        RECT 721.950 413.250 724.050 414.150 ;
        RECT 721.950 409.950 724.050 412.050 ;
        RECT 722.400 403.050 723.450 409.950 ;
        RECT 721.950 400.950 724.050 403.050 ;
        RECT 722.400 382.050 723.450 400.950 ;
        RECT 721.950 379.950 724.050 382.050 ;
        RECT 721.950 377.850 724.050 378.750 ;
        RECT 725.400 370.050 726.450 511.950 ;
        RECT 724.950 367.950 727.050 370.050 ;
        RECT 716.400 365.400 720.450 366.450 ;
        RECT 703.950 358.950 706.050 361.050 ;
        RECT 691.950 355.950 694.050 358.050 ;
        RECT 700.950 352.950 703.050 355.050 ;
        RECT 682.950 346.950 685.050 349.050 ;
        RECT 694.950 346.950 697.050 349.050 ;
        RECT 683.400 343.050 684.450 346.950 ;
        RECT 679.950 341.250 681.750 342.150 ;
        RECT 682.950 340.950 685.050 343.050 ;
        RECT 686.250 341.250 687.750 342.150 ;
        RECT 688.950 340.950 691.050 343.050 ;
        RECT 692.250 341.250 694.050 342.150 ;
        RECT 679.950 337.950 682.050 340.050 ;
        RECT 683.250 338.850 684.750 339.750 ;
        RECT 685.950 337.950 688.050 340.050 ;
        RECT 689.250 338.850 690.750 339.750 ;
        RECT 691.950 337.950 694.050 340.050 ;
        RECT 680.400 331.050 681.450 337.950 ;
        RECT 686.400 333.450 687.450 337.950 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 683.400 332.400 687.450 333.450 ;
        RECT 679.950 328.950 682.050 331.050 ;
        RECT 665.400 320.400 669.450 321.450 ;
        RECT 655.950 310.950 658.050 313.050 ;
        RECT 659.250 311.250 660.750 312.150 ;
        RECT 661.950 310.950 664.050 313.050 ;
        RECT 665.400 310.050 666.450 320.400 ;
        RECT 676.950 319.950 679.050 322.050 ;
        RECT 667.950 313.950 670.050 316.050 ;
        RECT 676.950 313.950 679.050 316.050 ;
        RECT 652.950 309.450 655.050 310.050 ;
        RECT 650.400 308.400 655.050 309.450 ;
        RECT 656.250 308.850 657.750 309.750 ;
        RECT 646.950 286.950 649.050 289.050 ;
        RECT 631.950 283.950 634.050 286.050 ;
        RECT 632.400 280.050 633.450 283.950 ;
        RECT 631.950 277.950 634.050 280.050 ;
        RECT 640.950 274.950 643.050 277.050 ;
        RECT 641.400 271.050 642.450 274.950 ;
        RECT 631.950 269.250 633.750 270.150 ;
        RECT 634.950 268.950 637.050 271.050 ;
        RECT 638.250 269.250 639.750 270.150 ;
        RECT 640.950 268.950 643.050 271.050 ;
        RECT 644.250 269.250 646.050 270.150 ;
        RECT 631.950 267.450 634.050 268.050 ;
        RECT 629.400 266.400 634.050 267.450 ;
        RECT 635.250 266.850 636.750 267.750 ;
        RECT 631.950 265.950 634.050 266.400 ;
        RECT 637.950 265.950 640.050 268.050 ;
        RECT 641.250 266.850 642.750 267.750 ;
        RECT 643.950 265.950 646.050 268.050 ;
        RECT 644.400 258.450 645.450 265.950 ;
        RECT 650.400 265.050 651.450 308.400 ;
        RECT 652.950 307.950 655.050 308.400 ;
        RECT 658.950 307.950 661.050 310.050 ;
        RECT 662.250 308.850 664.050 309.750 ;
        RECT 664.950 307.950 667.050 310.050 ;
        RECT 652.950 305.850 655.050 306.750 ;
        RECT 661.950 286.950 664.050 289.050 ;
        RECT 652.950 274.950 655.050 277.050 ;
        RECT 655.950 274.950 658.050 277.050 ;
        RECT 649.950 262.950 652.050 265.050 ;
        RECT 650.400 262.050 651.450 262.950 ;
        RECT 649.950 259.950 652.050 262.050 ;
        RECT 644.400 257.400 648.450 258.450 ;
        RECT 634.950 250.950 637.050 253.050 ;
        RECT 647.400 252.450 648.450 257.400 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 650.400 256.050 651.450 256.950 ;
        RECT 649.950 253.950 652.050 256.050 ;
        RECT 653.400 252.450 654.450 274.950 ;
        RECT 656.400 274.050 657.450 274.950 ;
        RECT 662.400 274.050 663.450 286.950 ;
        RECT 668.400 277.050 669.450 313.950 ;
        RECT 677.400 313.050 678.450 313.950 ;
        RECT 683.400 313.050 684.450 332.400 ;
        RECT 685.950 328.950 688.050 331.050 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 674.250 311.250 675.750 312.150 ;
        RECT 676.950 310.950 679.050 313.050 ;
        RECT 682.950 310.950 685.050 313.050 ;
        RECT 670.950 308.850 672.750 309.750 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 677.250 308.850 678.750 309.750 ;
        RECT 679.950 307.950 682.050 310.050 ;
        RECT 679.950 305.850 682.050 306.750 ;
        RECT 667.950 274.950 670.050 277.050 ;
        RECT 673.950 274.950 676.050 277.050 ;
        RECT 682.950 274.950 685.050 277.050 ;
        RECT 655.950 271.950 658.050 274.050 ;
        RECT 661.950 273.450 664.050 274.050 ;
        RECT 659.250 272.250 660.750 273.150 ;
        RECT 661.950 272.400 666.450 273.450 ;
        RECT 661.950 271.950 664.050 272.400 ;
        RECT 655.950 269.850 657.750 270.750 ;
        RECT 658.950 268.950 661.050 271.050 ;
        RECT 662.250 269.850 664.050 270.750 ;
        RECT 647.400 251.400 651.450 252.450 ;
        RECT 653.400 251.400 657.450 252.450 ;
        RECT 625.950 205.950 628.050 208.050 ;
        RECT 619.950 202.950 622.050 205.050 ;
        RECT 601.950 196.950 604.050 199.050 ;
        RECT 605.250 197.250 606.750 198.150 ;
        RECT 607.950 196.950 610.050 199.050 ;
        RECT 611.250 197.250 613.050 198.150 ;
        RECT 613.950 196.950 616.050 199.050 ;
        RECT 602.400 193.050 603.450 196.950 ;
        RECT 604.950 193.950 607.050 196.050 ;
        RECT 608.250 194.850 609.750 195.750 ;
        RECT 610.950 195.450 613.050 196.050 ;
        RECT 614.400 195.450 615.450 196.950 ;
        RECT 610.950 194.400 615.450 195.450 ;
        RECT 610.950 193.950 613.050 194.400 ;
        RECT 601.950 190.950 604.050 193.050 ;
        RECT 601.950 169.950 604.050 172.050 ;
        RECT 595.950 166.950 598.050 169.050 ;
        RECT 592.950 164.250 594.750 165.150 ;
        RECT 595.950 163.950 598.050 166.050 ;
        RECT 599.250 164.250 601.050 165.150 ;
        RECT 592.950 162.450 595.050 163.050 ;
        RECT 590.400 161.400 595.050 162.450 ;
        RECT 596.250 161.850 597.750 162.750 ;
        RECT 598.950 162.450 601.050 163.050 ;
        RECT 602.400 162.450 603.450 169.950 ;
        RECT 592.950 160.950 595.050 161.400 ;
        RECT 598.950 161.400 603.450 162.450 ;
        RECT 598.950 160.950 601.050 161.400 ;
        RECT 586.950 151.950 589.050 154.050 ;
        RECT 575.400 128.400 579.450 129.450 ;
        RECT 574.950 124.950 577.050 127.050 ;
        RECT 571.950 97.950 574.050 100.050 ;
        RECT 572.400 97.050 573.450 97.950 ;
        RECT 559.950 94.950 562.050 97.050 ;
        RECT 565.950 94.950 568.050 97.050 ;
        RECT 569.250 95.250 570.750 96.150 ;
        RECT 571.950 94.950 574.050 97.050 ;
        RECT 562.950 93.450 565.050 94.050 ;
        RECT 560.400 92.400 565.050 93.450 ;
        RECT 566.250 92.850 567.750 93.750 ;
        RECT 560.400 91.050 561.450 92.400 ;
        RECT 562.950 91.950 565.050 92.400 ;
        RECT 568.950 91.950 571.050 94.050 ;
        RECT 572.250 92.850 574.050 93.750 ;
        RECT 559.950 88.950 562.050 91.050 ;
        RECT 562.950 89.850 565.050 90.750 ;
        RECT 560.400 61.050 561.450 88.950 ;
        RECT 571.950 76.950 574.050 79.050 ;
        RECT 559.950 58.950 562.050 61.050 ;
        RECT 568.950 58.950 571.050 61.050 ;
        RECT 557.400 56.400 561.450 57.450 ;
        RECT 533.250 53.250 534.750 54.150 ;
        RECT 535.950 53.400 540.450 54.450 ;
        RECT 544.950 54.450 547.050 55.050 ;
        RECT 547.950 54.450 550.050 55.050 ;
        RECT 544.950 53.400 550.050 54.450 ;
        RECT 535.950 52.950 538.050 53.400 ;
        RECT 544.950 52.950 547.050 53.400 ;
        RECT 547.950 52.950 550.050 53.400 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 557.250 53.250 559.050 54.150 ;
        RECT 526.950 51.450 529.050 52.050 ;
        RECT 514.950 50.250 517.050 51.150 ;
        RECT 524.400 50.400 529.050 51.450 ;
        RECT 530.250 50.850 531.750 51.750 ;
        RECT 526.950 49.950 529.050 50.400 ;
        RECT 532.950 49.950 535.050 52.050 ;
        RECT 499.950 46.950 502.050 49.050 ;
        RECT 514.950 46.950 517.050 49.050 ;
        RECT 515.400 46.050 516.450 46.950 ;
        RECT 514.950 43.950 517.050 46.050 ;
        RECT 497.400 32.400 501.450 33.450 ;
        RECT 496.950 28.950 499.050 31.050 ;
        RECT 497.400 28.050 498.450 28.950 ;
        RECT 454.950 25.950 457.050 28.050 ;
        RECT 478.950 25.950 481.050 28.050 ;
        RECT 496.950 25.950 499.050 28.050 ;
        RECT 454.950 20.250 456.750 21.150 ;
        RECT 457.950 19.950 460.050 22.050 ;
        RECT 461.250 20.250 463.050 21.150 ;
        RECT 472.950 20.250 474.750 21.150 ;
        RECT 475.950 19.950 478.050 22.050 ;
        RECT 479.400 19.050 480.450 25.950 ;
        RECT 493.950 23.250 496.050 24.150 ;
        RECT 496.950 23.850 499.050 24.750 ;
        RECT 500.400 22.050 501.450 32.400 ;
        RECT 533.400 31.050 534.450 49.950 ;
        RECT 545.400 48.450 546.450 52.950 ;
        RECT 547.950 50.850 550.050 51.750 ;
        RECT 550.950 50.250 553.050 51.150 ;
        RECT 553.950 50.850 555.750 51.750 ;
        RECT 556.950 49.950 559.050 52.050 ;
        RECT 545.400 47.400 549.450 48.450 ;
        RECT 505.950 28.950 508.050 31.050 ;
        RECT 532.950 28.950 535.050 31.050 ;
        RECT 506.400 25.050 507.450 28.950 ;
        RECT 532.950 25.950 535.050 28.050 ;
        RECT 505.950 22.950 508.050 25.050 ;
        RECT 509.250 23.250 510.750 24.150 ;
        RECT 511.950 22.950 514.050 25.050 ;
        RECT 529.950 23.250 532.050 24.150 ;
        RECT 532.950 23.850 535.050 24.750 ;
        RECT 548.400 22.050 549.450 47.400 ;
        RECT 550.950 46.950 553.050 49.050 ;
        RECT 551.400 46.050 552.450 46.950 ;
        RECT 550.950 43.950 553.050 46.050 ;
        RECT 560.400 28.050 561.450 56.400 ;
        RECT 559.950 25.950 562.050 28.050 ;
        RECT 569.400 25.050 570.450 58.950 ;
        RECT 572.400 58.050 573.450 76.950 ;
        RECT 575.400 61.050 576.450 124.950 ;
        RECT 578.400 115.050 579.450 128.400 ;
        RECT 580.950 128.250 583.050 129.150 ;
        RECT 583.950 127.950 586.050 130.050 ;
        RECT 580.950 124.950 583.050 127.050 ;
        RECT 584.250 125.250 585.750 126.150 ;
        RECT 586.950 124.950 589.050 127.050 ;
        RECT 590.250 125.250 592.050 126.150 ;
        RECT 577.950 112.950 580.050 115.050 ;
        RECT 578.400 96.450 579.450 112.950 ;
        RECT 581.400 106.050 582.450 124.950 ;
        RECT 583.950 121.950 586.050 124.050 ;
        RECT 587.250 122.850 588.750 123.750 ;
        RECT 589.950 123.450 592.050 124.050 ;
        RECT 593.400 123.450 594.450 160.950 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 599.400 130.050 600.450 133.950 ;
        RECT 605.400 132.450 606.450 193.950 ;
        RECT 613.950 169.950 616.050 172.050 ;
        RECT 610.950 168.450 613.050 169.050 ;
        RECT 608.400 167.400 613.050 168.450 ;
        RECT 614.250 167.850 615.750 168.750 ;
        RECT 608.400 160.050 609.450 167.400 ;
        RECT 610.950 166.950 613.050 167.400 ;
        RECT 616.950 166.950 619.050 169.050 ;
        RECT 610.950 164.850 613.050 165.750 ;
        RECT 616.950 164.850 619.050 165.750 ;
        RECT 607.950 157.950 610.050 160.050 ;
        RECT 620.400 133.050 621.450 202.950 ;
        RECT 622.950 200.250 625.050 201.150 ;
        RECT 622.950 196.950 625.050 199.050 ;
        RECT 626.250 197.250 627.750 198.150 ;
        RECT 628.950 196.950 631.050 199.050 ;
        RECT 632.250 197.250 634.050 198.150 ;
        RECT 625.950 193.950 628.050 196.050 ;
        RECT 629.250 194.850 630.750 195.750 ;
        RECT 631.950 193.950 634.050 196.050 ;
        RECT 626.400 193.050 627.450 193.950 ;
        RECT 625.950 190.950 628.050 193.050 ;
        RECT 626.400 171.450 627.450 190.950 ;
        RECT 632.400 187.050 633.450 193.950 ;
        RECT 631.950 184.950 634.050 187.050 ;
        RECT 632.400 181.050 633.450 184.950 ;
        RECT 631.950 178.950 634.050 181.050 ;
        RECT 628.950 171.450 631.050 172.050 ;
        RECT 626.400 170.400 631.050 171.450 ;
        RECT 628.950 169.950 631.050 170.400 ;
        RECT 622.950 166.950 625.050 169.050 ;
        RECT 625.950 166.950 628.050 169.050 ;
        RECT 628.950 167.850 631.050 168.750 ;
        RECT 631.950 167.250 634.050 168.150 ;
        RECT 605.400 131.400 609.450 132.450 ;
        RECT 598.950 127.950 601.050 130.050 ;
        RECT 602.250 128.250 603.750 129.150 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 598.950 125.850 600.750 126.750 ;
        RECT 601.950 124.950 604.050 127.050 ;
        RECT 605.250 125.850 607.050 126.750 ;
        RECT 589.950 122.400 594.450 123.450 ;
        RECT 589.950 121.950 592.050 122.400 ;
        RECT 580.950 103.950 583.050 106.050 ;
        RECT 589.950 97.950 592.050 100.050 ;
        RECT 580.950 96.450 583.050 97.050 ;
        RECT 578.400 95.400 583.050 96.450 ;
        RECT 580.950 94.950 583.050 95.400 ;
        RECT 584.250 95.250 585.750 96.150 ;
        RECT 586.950 94.950 589.050 97.050 ;
        RECT 590.400 94.050 591.450 97.950 ;
        RECT 580.950 92.850 582.750 93.750 ;
        RECT 583.950 91.950 586.050 94.050 ;
        RECT 587.250 92.850 588.750 93.750 ;
        RECT 589.950 91.950 592.050 94.050 ;
        RECT 589.950 89.850 592.050 90.750 ;
        RECT 593.400 82.050 594.450 122.400 ;
        RECT 608.400 121.050 609.450 131.400 ;
        RECT 613.950 130.950 616.050 133.050 ;
        RECT 619.950 130.950 622.050 133.050 ;
        RECT 598.950 118.950 601.050 121.050 ;
        RECT 607.950 118.950 610.050 121.050 ;
        RECT 599.400 94.050 600.450 118.950 ;
        RECT 610.950 115.950 613.050 118.050 ;
        RECT 604.950 103.950 607.050 106.050 ;
        RECT 605.400 100.050 606.450 103.950 ;
        RECT 604.950 97.950 607.050 100.050 ;
        RECT 611.400 97.050 612.450 115.950 ;
        RECT 601.950 95.250 604.050 96.150 ;
        RECT 604.950 95.850 607.050 96.750 ;
        RECT 607.950 95.250 609.750 96.150 ;
        RECT 610.950 94.950 613.050 97.050 ;
        RECT 598.950 91.950 601.050 94.050 ;
        RECT 601.950 91.950 604.050 94.050 ;
        RECT 607.950 91.950 610.050 94.050 ;
        RECT 611.250 92.850 613.050 93.750 ;
        RECT 586.950 79.950 589.050 82.050 ;
        RECT 592.950 79.950 595.050 82.050 ;
        RECT 574.950 58.950 577.050 61.050 ;
        RECT 577.950 59.250 580.050 60.150 ;
        RECT 571.950 55.950 574.050 58.050 ;
        RECT 575.250 56.250 576.750 57.150 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 581.250 56.250 583.050 57.150 ;
        RECT 587.400 55.050 588.450 79.950 ;
        RECT 602.400 79.050 603.450 91.950 ;
        RECT 601.950 76.950 604.050 79.050 ;
        RECT 614.400 60.450 615.450 130.950 ;
        RECT 623.400 130.050 624.450 166.950 ;
        RECT 616.950 127.950 619.050 130.050 ;
        RECT 619.950 128.250 622.050 129.150 ;
        RECT 622.950 127.950 625.050 130.050 ;
        RECT 617.400 67.050 618.450 127.950 ;
        RECT 626.400 127.050 627.450 166.950 ;
        RECT 631.950 163.950 634.050 166.050 ;
        RECT 632.400 139.050 633.450 163.950 ;
        RECT 631.950 136.950 634.050 139.050 ;
        RECT 619.950 124.950 622.050 127.050 ;
        RECT 623.250 125.250 624.750 126.150 ;
        RECT 625.950 124.950 628.050 127.050 ;
        RECT 629.250 125.250 631.050 126.150 ;
        RECT 620.400 121.050 621.450 124.950 ;
        RECT 622.950 121.950 625.050 124.050 ;
        RECT 626.250 122.850 627.750 123.750 ;
        RECT 628.950 121.950 631.050 124.050 ;
        RECT 619.950 118.950 622.050 121.050 ;
        RECT 616.950 64.950 619.050 67.050 ;
        RECT 623.400 61.050 624.450 121.950 ;
        RECT 632.400 100.050 633.450 136.950 ;
        RECT 635.400 136.050 636.450 250.950 ;
        RECT 643.950 247.950 646.050 250.050 ;
        RECT 644.400 241.050 645.450 247.950 ;
        RECT 650.400 241.050 651.450 251.400 ;
        RECT 652.950 247.950 655.050 250.050 ;
        RECT 637.950 238.950 640.050 241.050 ;
        RECT 641.250 239.250 642.750 240.150 ;
        RECT 643.950 238.950 646.050 241.050 ;
        RECT 647.250 239.250 648.750 240.150 ;
        RECT 649.950 238.950 652.050 241.050 ;
        RECT 637.950 236.850 639.750 237.750 ;
        RECT 640.950 235.950 643.050 238.050 ;
        RECT 644.250 236.850 645.750 237.750 ;
        RECT 646.950 235.950 649.050 238.050 ;
        RECT 650.250 236.850 652.050 237.750 ;
        RECT 647.400 223.050 648.450 235.950 ;
        RECT 640.950 220.950 643.050 223.050 ;
        RECT 646.950 220.950 649.050 223.050 ;
        RECT 641.400 193.050 642.450 220.950 ;
        RECT 653.400 211.050 654.450 247.950 ;
        RECT 652.950 208.950 655.050 211.050 ;
        RECT 653.400 199.050 654.450 208.950 ;
        RECT 643.950 197.250 645.750 198.150 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 652.950 196.950 655.050 199.050 ;
        RECT 643.950 193.950 646.050 196.050 ;
        RECT 647.250 194.850 649.050 195.750 ;
        RECT 649.950 194.250 652.050 195.150 ;
        RECT 652.950 194.850 655.050 195.750 ;
        RECT 640.950 190.950 643.050 193.050 ;
        RECT 649.950 190.950 652.050 193.050 ;
        RECT 656.400 178.050 657.450 251.400 ;
        RECT 659.400 246.450 660.450 268.950 ;
        RECT 665.400 268.050 666.450 272.400 ;
        RECT 674.400 271.050 675.450 274.950 ;
        RECT 679.950 272.250 682.050 273.150 ;
        RECT 667.950 268.950 670.050 271.050 ;
        RECT 670.950 269.250 672.750 270.150 ;
        RECT 673.950 268.950 676.050 271.050 ;
        RECT 677.250 269.250 678.750 270.150 ;
        RECT 679.950 268.950 682.050 271.050 ;
        RECT 664.950 265.950 667.050 268.050 ;
        RECT 668.400 256.050 669.450 268.950 ;
        RECT 670.950 265.950 673.050 268.050 ;
        RECT 674.250 266.850 675.750 267.750 ;
        RECT 676.950 265.950 679.050 268.050 ;
        RECT 667.950 253.950 670.050 256.050 ;
        RECT 659.400 245.400 663.450 246.450 ;
        RECT 662.400 241.050 663.450 245.400 ;
        RECT 667.950 241.950 670.050 244.050 ;
        RECT 670.950 243.450 673.050 244.050 ;
        RECT 673.950 243.450 676.050 244.050 ;
        RECT 670.950 242.400 676.050 243.450 ;
        RECT 670.950 241.950 673.050 242.400 ;
        RECT 673.950 241.950 676.050 242.400 ;
        RECT 668.400 241.050 669.450 241.950 ;
        RECT 661.950 238.950 664.050 241.050 ;
        RECT 665.250 239.250 666.750 240.150 ;
        RECT 667.950 238.950 670.050 241.050 ;
        RECT 671.250 239.250 672.750 240.150 ;
        RECT 673.950 238.950 676.050 241.050 ;
        RECT 661.950 236.850 663.750 237.750 ;
        RECT 664.950 235.950 667.050 238.050 ;
        RECT 668.250 236.850 669.750 237.750 ;
        RECT 670.950 235.950 673.050 238.050 ;
        RECT 674.250 236.850 676.050 237.750 ;
        RECT 671.400 234.450 672.450 235.950 ;
        RECT 671.400 233.400 675.450 234.450 ;
        RECT 670.950 220.950 673.050 223.050 ;
        RECT 664.950 200.250 667.050 201.150 ;
        RECT 671.400 199.050 672.450 220.950 ;
        RECT 674.400 202.050 675.450 233.400 ;
        RECT 673.950 199.950 676.050 202.050 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 668.250 197.250 669.750 198.150 ;
        RECT 670.950 196.950 673.050 199.050 ;
        RECT 674.250 197.250 676.050 198.150 ;
        RECT 665.400 190.050 666.450 196.950 ;
        RECT 677.400 196.050 678.450 265.950 ;
        RECT 680.400 262.050 681.450 268.950 ;
        RECT 683.400 268.050 684.450 274.950 ;
        RECT 682.950 265.950 685.050 268.050 ;
        RECT 679.950 259.950 682.050 262.050 ;
        RECT 683.400 259.050 684.450 265.950 ;
        RECT 682.950 256.950 685.050 259.050 ;
        RECT 682.950 253.950 685.050 256.050 ;
        RECT 679.950 241.950 682.050 244.050 ;
        RECT 680.400 208.050 681.450 241.950 ;
        RECT 683.400 238.050 684.450 253.950 ;
        RECT 686.400 241.050 687.450 328.950 ;
        RECT 689.400 271.050 690.450 334.950 ;
        RECT 695.400 325.050 696.450 346.950 ;
        RECT 694.950 322.950 697.050 325.050 ;
        RECT 691.950 308.250 693.750 309.150 ;
        RECT 694.950 307.950 697.050 310.050 ;
        RECT 698.250 308.250 700.050 309.150 ;
        RECT 691.950 304.950 694.050 307.050 ;
        RECT 695.250 305.850 696.750 306.750 ;
        RECT 697.950 304.950 700.050 307.050 ;
        RECT 691.950 301.950 694.050 304.050 ;
        RECT 688.950 268.950 691.050 271.050 ;
        RECT 692.400 256.050 693.450 301.950 ;
        RECT 698.400 301.050 699.450 304.950 ;
        RECT 697.950 298.950 700.050 301.050 ;
        RECT 701.400 277.050 702.450 352.950 ;
        RECT 704.400 346.050 705.450 358.950 ;
        RECT 703.950 343.950 706.050 346.050 ;
        RECT 707.250 344.250 708.750 345.150 ;
        RECT 709.950 343.950 712.050 346.050 ;
        RECT 703.950 341.850 705.750 342.750 ;
        RECT 706.950 340.950 709.050 343.050 ;
        RECT 710.250 341.850 712.050 342.750 ;
        RECT 707.400 340.050 708.450 340.950 ;
        RECT 706.950 337.950 709.050 340.050 ;
        RECT 706.950 325.950 709.050 328.050 ;
        RECT 703.950 313.950 706.050 316.050 ;
        RECT 700.950 274.950 703.050 277.050 ;
        RECT 697.950 273.450 700.050 274.050 ;
        RECT 704.400 273.450 705.450 313.950 ;
        RECT 707.400 304.050 708.450 325.950 ;
        RECT 716.400 316.050 717.450 365.400 ;
        RECT 718.950 358.950 721.050 361.050 ;
        RECT 715.950 313.950 718.050 316.050 ;
        RECT 709.950 308.250 711.750 309.150 ;
        RECT 712.950 307.950 715.050 310.050 ;
        RECT 716.250 308.250 718.050 309.150 ;
        RECT 709.950 304.950 712.050 307.050 ;
        RECT 713.250 305.850 714.750 306.750 ;
        RECT 715.950 306.450 718.050 307.050 ;
        RECT 719.400 306.450 720.450 358.950 ;
        RECT 728.400 355.050 729.450 571.950 ;
        RECT 730.950 559.950 733.050 562.050 ;
        RECT 731.400 559.050 732.450 559.950 ;
        RECT 730.950 556.950 733.050 559.050 ;
        RECT 734.250 557.250 736.050 558.150 ;
        RECT 730.950 554.850 732.750 555.750 ;
        RECT 733.950 555.450 736.050 556.050 ;
        RECT 737.400 555.450 738.450 583.950 ;
        RECT 755.250 560.250 756.750 561.150 ;
        RECT 751.950 557.850 753.750 558.750 ;
        RECT 754.950 556.950 757.050 559.050 ;
        RECT 758.250 557.850 760.050 558.750 ;
        RECT 733.950 554.400 738.450 555.450 ;
        RECT 733.950 553.950 736.050 554.400 ;
        RECT 730.950 550.950 733.050 553.050 ;
        RECT 731.400 484.050 732.450 550.950 ;
        RECT 734.400 538.050 735.450 553.950 ;
        RECT 761.400 553.050 762.450 671.400 ;
        RECT 763.950 670.950 766.050 671.400 ;
        RECT 767.550 665.400 768.750 677.400 ;
        RECT 772.950 676.950 775.050 679.050 ;
        RECT 769.950 667.950 772.050 670.050 ;
        RECT 766.950 663.300 769.050 665.400 ;
        RECT 767.550 659.700 768.750 663.300 ;
        RECT 770.400 661.050 771.450 667.950 ;
        RECT 766.950 657.600 769.050 659.700 ;
        RECT 769.950 658.950 772.050 661.050 ;
        RECT 773.400 634.050 774.450 676.950 ;
        RECT 775.950 673.950 778.050 676.050 ;
        RECT 776.400 673.050 777.450 673.950 ;
        RECT 775.950 670.950 778.050 673.050 ;
        RECT 775.950 668.850 778.050 669.750 ;
        RECT 779.400 666.450 780.450 694.950 ;
        RECT 782.400 679.050 783.450 709.950 ;
        RECT 797.400 709.050 798.450 838.950 ;
        RECT 800.400 828.450 801.450 841.950 ;
        RECT 803.400 841.050 804.450 844.950 ;
        RECT 805.950 841.950 808.050 844.050 ;
        RECT 814.950 842.250 817.050 843.150 ;
        RECT 817.950 842.850 820.050 843.750 ;
        RECT 802.950 838.950 805.050 841.050 ;
        RECT 800.400 827.400 804.450 828.450 ;
        RECT 799.950 821.400 802.050 823.500 ;
        RECT 800.400 804.600 801.600 821.400 ;
        RECT 799.950 802.500 802.050 804.600 ;
        RECT 803.400 781.050 804.450 827.400 ;
        RECT 802.950 778.950 805.050 781.050 ;
        RECT 802.950 772.950 805.050 775.050 ;
        RECT 799.950 770.250 802.050 771.150 ;
        RECT 802.950 770.850 805.050 771.750 ;
        RECT 799.950 766.950 802.050 769.050 ;
        RECT 806.400 768.450 807.450 841.950 ;
        RECT 814.950 838.950 817.050 841.050 ;
        RECT 826.950 838.950 829.050 841.050 ;
        RECT 811.950 835.950 814.050 838.050 ;
        RECT 803.400 767.400 807.450 768.450 ;
        RECT 800.400 766.050 801.450 766.950 ;
        RECT 799.950 763.950 802.050 766.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 800.400 745.050 801.450 757.950 ;
        RECT 799.950 742.950 802.050 745.050 ;
        RECT 799.950 740.850 802.050 741.750 ;
        RECT 787.950 706.950 790.050 709.050 ;
        RECT 790.950 706.950 793.050 709.050 ;
        RECT 796.950 706.950 799.050 709.050 ;
        RECT 788.400 684.450 789.450 706.950 ;
        RECT 791.400 706.050 792.450 706.950 ;
        RECT 790.950 703.950 793.050 706.050 ;
        RECT 794.250 704.250 795.750 705.150 ;
        RECT 796.950 703.950 799.050 706.050 ;
        RECT 799.950 703.950 802.050 706.050 ;
        RECT 790.950 701.850 792.750 702.750 ;
        RECT 793.950 700.950 796.050 703.050 ;
        RECT 797.250 701.850 799.050 702.750 ;
        RECT 794.400 685.050 795.450 700.950 ;
        RECT 800.400 697.050 801.450 703.950 ;
        RECT 803.400 697.050 804.450 767.400 ;
        RECT 805.950 749.400 808.050 751.500 ;
        RECT 806.400 732.600 807.600 749.400 ;
        RECT 805.950 730.500 808.050 732.600 ;
        RECT 805.950 715.950 808.050 718.050 ;
        RECT 806.400 709.050 807.450 715.950 ;
        RECT 805.950 706.950 808.050 709.050 ;
        RECT 812.400 706.050 813.450 835.950 ;
        RECT 818.250 815.250 819.750 816.150 ;
        RECT 820.950 814.950 823.050 817.050 ;
        RECT 823.950 814.950 826.050 817.050 ;
        RECT 824.400 814.050 825.450 814.950 ;
        RECT 814.950 812.850 816.750 813.750 ;
        RECT 817.950 811.950 820.050 814.050 ;
        RECT 821.250 812.850 822.750 813.750 ;
        RECT 823.950 811.950 826.050 814.050 ;
        RECT 818.400 805.050 819.450 811.950 ;
        RECT 823.950 809.850 826.050 810.750 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 823.950 776.250 826.050 777.150 ;
        RECT 814.950 773.250 816.750 774.150 ;
        RECT 817.950 772.950 820.050 775.050 ;
        RECT 821.250 773.250 822.750 774.150 ;
        RECT 823.950 772.950 826.050 775.050 ;
        RECT 818.250 770.850 819.750 771.750 ;
        RECT 820.950 769.950 823.050 772.050 ;
        RECT 817.950 766.950 820.050 769.050 ;
        RECT 820.950 766.950 823.050 769.050 ;
        RECT 818.400 760.050 819.450 766.950 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 817.950 745.950 820.050 748.050 ;
        RECT 818.400 718.050 819.450 745.950 ;
        RECT 817.950 715.950 820.050 718.050 ;
        RECT 805.950 703.950 808.050 706.050 ;
        RECT 811.950 703.950 814.050 706.050 ;
        RECT 815.250 704.250 816.750 705.150 ;
        RECT 817.950 703.950 820.050 706.050 ;
        RECT 806.400 700.050 807.450 703.950 ;
        RECT 811.950 701.850 813.750 702.750 ;
        RECT 814.950 700.950 817.050 703.050 ;
        RECT 818.250 701.850 820.050 702.750 ;
        RECT 805.950 697.950 808.050 700.050 ;
        RECT 814.950 697.950 817.050 700.050 ;
        RECT 799.950 694.950 802.050 697.050 ;
        RECT 802.950 694.950 805.050 697.050 ;
        RECT 811.950 694.950 814.050 697.050 ;
        RECT 788.400 683.400 792.450 684.450 ;
        RECT 781.950 676.950 784.050 679.050 ;
        RECT 787.950 677.400 790.050 679.500 ;
        RECT 781.950 670.950 784.050 673.050 ;
        RECT 781.950 668.850 784.050 669.750 ;
        RECT 776.400 665.400 780.450 666.450 ;
        RECT 769.950 631.950 772.050 634.050 ;
        RECT 772.950 631.950 775.050 634.050 ;
        RECT 770.400 631.050 771.450 631.950 ;
        RECT 763.950 628.950 766.050 631.050 ;
        RECT 769.950 628.950 772.050 631.050 ;
        RECT 773.250 629.250 775.050 630.150 ;
        RECT 763.950 626.850 766.050 627.750 ;
        RECT 766.950 626.250 769.050 627.150 ;
        RECT 769.950 626.850 771.750 627.750 ;
        RECT 772.950 627.450 775.050 628.050 ;
        RECT 776.400 627.450 777.450 665.400 ;
        RECT 778.950 661.950 781.050 664.050 ;
        RECT 779.400 661.050 780.450 661.950 ;
        RECT 778.950 658.950 781.050 661.050 ;
        RECT 788.400 660.600 789.600 677.400 ;
        RECT 779.400 631.050 780.450 658.950 ;
        RECT 787.950 658.500 790.050 660.600 ;
        RECT 791.400 634.050 792.450 683.400 ;
        RECT 793.950 682.950 796.050 685.050 ;
        RECT 799.950 673.950 802.050 676.050 ;
        RECT 790.950 631.950 793.050 634.050 ;
        RECT 793.950 632.250 796.050 633.150 ;
        RECT 778.950 628.950 781.050 631.050 ;
        RECT 784.950 629.250 786.750 630.150 ;
        RECT 787.950 628.950 790.050 631.050 ;
        RECT 791.250 629.250 792.750 630.150 ;
        RECT 793.950 628.950 796.050 631.050 ;
        RECT 772.950 626.400 777.450 627.450 ;
        RECT 772.950 625.950 775.050 626.400 ;
        RECT 766.950 622.950 769.050 625.050 ;
        RECT 775.950 622.950 778.050 625.050 ;
        RECT 767.400 619.050 768.450 622.950 ;
        RECT 766.950 616.950 769.050 619.050 ;
        RECT 766.950 613.950 769.050 616.050 ;
        RECT 767.400 598.050 768.450 613.950 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 769.950 599.250 772.050 600.150 ;
        RECT 772.950 599.850 775.050 600.750 ;
        RECT 776.400 600.450 777.450 622.950 ;
        RECT 779.400 607.050 780.450 628.950 ;
        RECT 784.950 625.950 787.050 628.050 ;
        RECT 788.250 626.850 789.750 627.750 ;
        RECT 790.950 625.950 793.050 628.050 ;
        RECT 785.400 616.050 786.450 625.950 ;
        RECT 784.950 613.950 787.050 616.050 ;
        RECT 791.400 613.050 792.450 625.950 ;
        RECT 790.950 610.950 793.050 613.050 ;
        RECT 796.950 607.950 799.050 610.050 ;
        RECT 778.950 604.950 781.050 607.050 ;
        RECT 781.950 605.400 784.050 607.500 ;
        RECT 778.950 602.250 781.050 603.150 ;
        RECT 778.950 600.450 781.050 601.050 ;
        RECT 776.400 599.400 781.050 600.450 ;
        RECT 766.950 595.950 769.050 598.050 ;
        RECT 769.950 595.950 772.050 598.050 ;
        RECT 770.400 595.050 771.450 595.950 ;
        RECT 769.950 592.950 772.050 595.050 ;
        RECT 763.950 589.950 766.050 592.050 ;
        RECT 760.950 550.950 763.050 553.050 ;
        RECT 733.950 535.950 736.050 538.050 ;
        RECT 754.950 532.950 757.050 535.050 ;
        RECT 755.400 529.050 756.450 532.950 ;
        RECT 754.950 526.950 757.050 529.050 ;
        RECT 758.250 527.250 759.750 528.150 ;
        RECT 733.950 524.250 735.750 525.150 ;
        RECT 736.950 523.950 739.050 526.050 ;
        RECT 740.250 524.250 742.050 525.150 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 751.950 523.950 754.050 526.050 ;
        RECT 755.250 524.850 756.750 525.750 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 761.250 524.850 763.050 525.750 ;
        RECT 737.250 521.850 738.750 522.750 ;
        RECT 746.400 507.450 747.450 523.950 ;
        RECT 751.950 521.850 754.050 522.750 ;
        RECT 758.400 520.050 759.450 523.950 ;
        RECT 757.950 517.950 760.050 520.050 ;
        RECT 746.400 506.400 750.450 507.450 ;
        RECT 737.250 488.250 738.750 489.150 ;
        RECT 733.950 485.850 735.750 486.750 ;
        RECT 736.950 484.950 739.050 487.050 ;
        RECT 740.250 485.850 742.050 486.750 ;
        RECT 749.400 486.450 750.450 506.400 ;
        RECT 751.950 488.250 754.050 489.150 ;
        RECT 751.950 486.450 754.050 487.050 ;
        RECT 749.400 485.400 754.050 486.450 ;
        RECT 751.950 484.950 754.050 485.400 ;
        RECT 755.250 485.250 756.750 486.150 ;
        RECT 757.950 484.950 760.050 487.050 ;
        RECT 761.250 485.250 763.050 486.150 ;
        RECT 730.950 481.950 733.050 484.050 ;
        RECT 739.950 481.950 742.050 484.050 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 758.250 482.850 759.750 483.750 ;
        RECT 730.950 452.250 732.750 453.150 ;
        RECT 733.950 451.950 736.050 454.050 ;
        RECT 737.250 452.250 739.050 453.150 ;
        RECT 734.250 449.850 735.750 450.750 ;
        RECT 730.950 423.300 733.050 425.400 ;
        RECT 731.250 419.700 732.450 423.300 ;
        RECT 730.950 417.600 733.050 419.700 ;
        RECT 731.250 405.600 732.450 417.600 ;
        RECT 733.950 411.450 736.050 412.050 ;
        RECT 733.950 410.400 738.450 411.450 ;
        RECT 733.950 409.950 736.050 410.400 ;
        RECT 737.400 409.050 738.450 410.400 ;
        RECT 733.950 407.850 736.050 408.750 ;
        RECT 736.950 406.950 739.050 409.050 ;
        RECT 730.950 403.500 733.050 405.600 ;
        RECT 733.950 383.250 736.050 384.150 ;
        RECT 733.950 379.950 736.050 382.050 ;
        RECT 727.950 352.950 730.050 355.050 ;
        RECT 727.950 349.950 730.050 352.050 ;
        RECT 721.950 340.950 724.050 343.050 ;
        RECT 724.950 341.250 727.050 342.150 ;
        RECT 722.400 316.050 723.450 340.950 ;
        RECT 724.950 337.950 727.050 340.050 ;
        RECT 725.400 337.050 726.450 337.950 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 721.950 313.950 724.050 316.050 ;
        RECT 715.950 305.400 720.450 306.450 ;
        RECT 715.950 304.950 718.050 305.400 ;
        RECT 706.950 301.950 709.050 304.050 ;
        RECT 706.950 280.950 709.050 283.050 ;
        RECT 707.400 280.050 708.450 280.950 ;
        RECT 706.950 277.950 709.050 280.050 ;
        RECT 697.950 272.400 705.450 273.450 ;
        RECT 697.950 271.950 700.050 272.400 ;
        RECT 694.950 269.250 697.050 270.150 ;
        RECT 697.950 269.850 700.050 270.750 ;
        RECT 694.950 265.950 697.050 268.050 ;
        RECT 691.950 253.950 694.050 256.050 ;
        RECT 691.950 241.950 694.050 244.050 ;
        RECT 692.400 241.050 693.450 241.950 ;
        RECT 685.950 238.950 688.050 241.050 ;
        RECT 689.250 239.250 690.750 240.150 ;
        RECT 691.950 238.950 694.050 241.050 ;
        RECT 695.250 239.250 696.750 240.150 ;
        RECT 697.950 238.950 700.050 241.050 ;
        RECT 682.950 235.950 685.050 238.050 ;
        RECT 685.950 236.850 687.750 237.750 ;
        RECT 688.950 235.950 691.050 238.050 ;
        RECT 692.250 236.850 693.750 237.750 ;
        RECT 694.950 235.950 697.050 238.050 ;
        RECT 698.250 236.850 700.050 237.750 ;
        RECT 682.950 232.950 685.050 235.050 ;
        RECT 679.950 205.950 682.050 208.050 ;
        RECT 683.400 199.050 684.450 232.950 ;
        RECT 689.400 232.050 690.450 235.950 ;
        RECT 688.950 229.950 691.050 232.050 ;
        RECT 701.400 202.050 702.450 272.400 ;
        RECT 703.950 269.250 706.050 270.150 ;
        RECT 703.950 267.450 706.050 268.050 ;
        RECT 707.400 267.450 708.450 277.950 ;
        RECT 710.400 274.050 711.450 304.950 ;
        RECT 722.400 304.050 723.450 313.950 ;
        RECT 712.950 301.950 715.050 304.050 ;
        RECT 721.950 301.950 724.050 304.050 ;
        RECT 709.950 271.950 712.050 274.050 ;
        RECT 703.950 266.400 708.450 267.450 ;
        RECT 703.950 265.950 706.050 266.400 ;
        RECT 703.950 262.950 706.050 265.050 ;
        RECT 694.950 200.250 697.050 201.150 ;
        RECT 697.950 199.950 700.050 202.050 ;
        RECT 700.950 199.950 703.050 202.050 ;
        RECT 682.950 196.950 685.050 199.050 ;
        RECT 685.950 197.250 687.750 198.150 ;
        RECT 688.950 196.950 691.050 199.050 ;
        RECT 692.250 197.250 693.750 198.150 ;
        RECT 694.950 196.950 697.050 199.050 ;
        RECT 667.950 193.950 670.050 196.050 ;
        RECT 671.250 194.850 672.750 195.750 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 676.950 193.950 679.050 196.050 ;
        RECT 685.950 193.950 688.050 196.050 ;
        RECT 689.250 194.850 690.750 195.750 ;
        RECT 691.950 193.950 694.050 196.050 ;
        RECT 664.950 187.950 667.050 190.050 ;
        RECT 670.950 187.950 673.050 190.050 ;
        RECT 665.400 184.050 666.450 187.950 ;
        RECT 664.950 181.950 667.050 184.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 637.950 175.950 640.050 178.050 ;
        RECT 655.950 175.950 658.050 178.050 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 638.400 126.450 639.450 175.950 ;
        RECT 652.950 172.950 655.050 175.050 ;
        RECT 658.950 172.950 661.050 175.050 ;
        RECT 653.400 172.050 654.450 172.950 ;
        RECT 652.950 169.950 655.050 172.050 ;
        RECT 646.950 166.950 649.050 169.050 ;
        RECT 650.250 167.250 652.050 168.150 ;
        RECT 652.950 167.850 655.050 168.750 ;
        RECT 655.950 167.250 658.050 168.150 ;
        RECT 646.950 164.850 648.750 165.750 ;
        RECT 649.950 163.950 652.050 166.050 ;
        RECT 655.950 165.450 658.050 166.050 ;
        RECT 659.400 165.450 660.450 172.950 ;
        RECT 655.950 164.400 660.450 165.450 ;
        RECT 655.950 163.950 658.050 164.400 ;
        RECT 662.400 163.050 663.450 178.950 ;
        RECT 667.950 169.950 670.050 172.050 ;
        RECT 668.400 166.050 669.450 169.950 ;
        RECT 671.400 166.050 672.450 187.950 ;
        RECT 674.400 175.050 675.450 193.950 ;
        RECT 685.950 190.950 688.050 193.050 ;
        RECT 673.950 172.950 676.050 175.050 ;
        RECT 679.950 172.950 682.050 175.050 ;
        RECT 680.400 169.050 681.450 172.950 ;
        RECT 673.950 166.950 676.050 169.050 ;
        RECT 677.250 167.250 678.750 168.150 ;
        RECT 679.950 166.950 682.050 169.050 ;
        RECT 667.950 163.950 670.050 166.050 ;
        RECT 670.950 163.950 673.050 166.050 ;
        RECT 674.250 164.850 675.750 165.750 ;
        RECT 676.950 163.950 679.050 166.050 ;
        RECT 680.250 164.850 682.050 165.750 ;
        RECT 661.950 160.950 664.050 163.050 ;
        RECT 670.950 161.850 673.050 162.750 ;
        RECT 640.950 128.250 643.050 129.150 ;
        RECT 679.950 128.250 682.050 129.150 ;
        RECT 686.400 127.050 687.450 190.950 ;
        RECT 692.400 172.050 693.450 193.950 ;
        RECT 698.400 178.050 699.450 199.950 ;
        RECT 704.400 193.050 705.450 262.950 ;
        RECT 710.400 255.450 711.450 271.950 ;
        RECT 713.400 265.050 714.450 301.950 ;
        RECT 718.950 280.950 721.050 283.050 ;
        RECT 719.400 271.050 720.450 280.950 ;
        RECT 715.950 269.250 718.050 270.150 ;
        RECT 718.950 268.950 721.050 271.050 ;
        RECT 721.950 269.250 724.050 270.150 ;
        RECT 715.950 265.950 718.050 268.050 ;
        RECT 719.250 266.250 720.750 267.150 ;
        RECT 721.950 265.950 724.050 268.050 ;
        RECT 712.950 262.950 715.050 265.050 ;
        RECT 716.400 262.050 717.450 265.950 ;
        RECT 718.950 262.950 721.050 265.050 ;
        RECT 715.950 259.950 718.050 262.050 ;
        RECT 707.400 254.400 711.450 255.450 ;
        RECT 707.400 202.050 708.450 254.400 ;
        RECT 715.950 250.950 718.050 253.050 ;
        RECT 716.400 241.050 717.450 250.950 ;
        RECT 719.400 247.050 720.450 262.950 ;
        RECT 721.950 253.950 724.050 256.050 ;
        RECT 718.950 244.950 721.050 247.050 ;
        RECT 718.950 241.950 721.050 244.050 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 715.950 238.950 718.050 241.050 ;
        RECT 713.400 238.050 714.450 238.950 ;
        RECT 709.950 236.250 711.750 237.150 ;
        RECT 712.950 235.950 715.050 238.050 ;
        RECT 716.250 236.250 718.050 237.150 ;
        RECT 709.950 232.950 712.050 235.050 ;
        RECT 713.250 233.850 714.750 234.750 ;
        RECT 715.950 232.950 718.050 235.050 ;
        RECT 710.400 226.050 711.450 232.950 ;
        RECT 716.400 229.050 717.450 232.950 ;
        RECT 715.950 226.950 718.050 229.050 ;
        RECT 709.950 223.950 712.050 226.050 ;
        RECT 712.950 211.950 715.050 214.050 ;
        RECT 713.400 202.050 714.450 211.950 ;
        RECT 706.950 199.950 709.050 202.050 ;
        RECT 710.250 200.250 711.750 201.150 ;
        RECT 712.950 199.950 715.050 202.050 ;
        RECT 706.950 197.850 708.750 198.750 ;
        RECT 709.950 196.950 712.050 199.050 ;
        RECT 713.250 197.850 715.050 198.750 ;
        RECT 719.400 193.050 720.450 241.950 ;
        RECT 722.400 232.050 723.450 253.950 ;
        RECT 725.400 250.050 726.450 334.950 ;
        RECT 728.400 307.050 729.450 349.950 ;
        RECT 734.400 349.050 735.450 379.950 ;
        RECT 733.950 346.950 736.050 349.050 ;
        RECT 733.950 343.950 736.050 346.050 ;
        RECT 730.950 341.250 733.050 342.150 ;
        RECT 730.950 337.950 733.050 340.050 ;
        RECT 734.400 328.050 735.450 343.950 ;
        RECT 737.400 343.050 738.450 406.950 ;
        RECT 740.400 346.050 741.450 481.950 ;
        RECT 755.400 457.050 756.450 481.950 ;
        RECT 764.400 480.450 765.450 589.950 ;
        RECT 770.400 589.050 771.450 592.950 ;
        RECT 769.950 586.950 772.050 589.050 ;
        RECT 769.950 568.950 772.050 571.050 ;
        RECT 770.400 559.050 771.450 568.950 ;
        RECT 769.950 556.950 772.050 559.050 ;
        RECT 766.950 554.250 769.050 555.150 ;
        RECT 769.950 554.850 772.050 555.750 ;
        RECT 766.950 550.950 769.050 553.050 ;
        RECT 776.400 538.050 777.450 599.400 ;
        RECT 778.950 598.950 781.050 599.400 ;
        RECT 782.550 593.400 783.750 605.400 ;
        RECT 787.950 604.950 790.050 607.050 ;
        RECT 781.950 591.300 784.050 593.400 ;
        RECT 782.550 587.700 783.750 591.300 ;
        RECT 781.950 585.600 784.050 587.700 ;
        RECT 781.950 580.950 784.050 583.050 ;
        RECT 775.950 535.950 778.050 538.050 ;
        RECT 772.950 524.250 774.750 525.150 ;
        RECT 775.950 523.950 778.050 526.050 ;
        RECT 779.250 524.250 781.050 525.150 ;
        RECT 776.250 521.850 777.750 522.750 ;
        RECT 772.950 484.950 775.050 487.050 ;
        RECT 772.950 482.850 775.050 483.750 ;
        RECT 775.950 482.250 778.050 483.150 ;
        RECT 761.400 479.400 765.450 480.450 ;
        RECT 748.950 454.950 751.050 457.050 ;
        RECT 754.950 454.950 757.050 457.050 ;
        RECT 749.400 454.050 750.450 454.950 ;
        RECT 745.950 452.250 747.750 453.150 ;
        RECT 748.950 451.950 751.050 454.050 ;
        RECT 752.250 452.250 754.050 453.150 ;
        RECT 749.250 449.850 750.750 450.750 ;
        RECT 757.950 416.250 760.050 417.150 ;
        RECT 745.950 412.950 748.050 415.050 ;
        RECT 748.950 413.250 750.750 414.150 ;
        RECT 751.950 412.950 754.050 415.050 ;
        RECT 755.250 413.250 756.750 414.150 ;
        RECT 757.950 412.950 760.050 415.050 ;
        RECT 746.400 408.450 747.450 412.950 ;
        RECT 752.250 410.850 753.750 411.750 ;
        RECT 754.950 409.950 757.050 412.050 ;
        RECT 743.400 407.400 747.450 408.450 ;
        RECT 739.950 343.950 742.050 346.050 ;
        RECT 743.400 343.050 744.450 407.400 ;
        RECT 745.950 389.400 748.050 391.500 ;
        RECT 746.400 372.600 747.600 389.400 ;
        RECT 751.950 384.450 754.050 385.050 ;
        RECT 755.400 384.450 756.450 409.950 ;
        RECT 757.950 400.950 760.050 403.050 ;
        RECT 758.400 385.050 759.450 400.950 ;
        RECT 751.950 383.400 756.450 384.450 ;
        RECT 751.950 382.950 754.050 383.400 ;
        RECT 757.950 382.950 760.050 385.050 ;
        RECT 751.950 380.850 754.050 381.750 ;
        RECT 757.950 380.850 760.050 381.750 ;
        RECT 745.950 370.500 748.050 372.600 ;
        RECT 745.950 364.950 748.050 367.050 ;
        RECT 736.950 340.950 739.050 343.050 ;
        RECT 742.950 340.950 745.050 343.050 ;
        RECT 746.400 340.050 747.450 364.950 ;
        RECT 761.400 352.050 762.450 479.400 ;
        RECT 775.950 478.950 778.050 481.050 ;
        RECT 763.950 461.400 766.050 463.500 ;
        RECT 764.400 444.600 765.600 461.400 ;
        RECT 776.400 460.050 777.450 478.950 ;
        RECT 775.950 457.950 778.050 460.050 ;
        RECT 769.950 454.950 772.050 457.050 ;
        RECT 775.950 456.450 778.050 457.050 ;
        RECT 775.950 455.400 780.450 456.450 ;
        RECT 775.950 454.950 778.050 455.400 ;
        RECT 779.400 454.050 780.450 455.400 ;
        RECT 769.950 452.850 772.050 453.750 ;
        RECT 775.950 452.850 778.050 453.750 ;
        RECT 778.950 451.950 781.050 454.050 ;
        RECT 763.950 442.500 766.050 444.600 ;
        RECT 773.250 416.250 774.750 417.150 ;
        RECT 769.950 413.850 771.750 414.750 ;
        RECT 772.950 412.950 775.050 415.050 ;
        RECT 776.250 413.850 778.050 414.750 ;
        RECT 775.950 409.950 778.050 412.050 ;
        RECT 766.950 389.400 769.050 391.500 ;
        RECT 767.250 377.400 768.450 389.400 ;
        RECT 769.950 386.250 772.050 387.150 ;
        RECT 769.950 382.950 772.050 385.050 ;
        RECT 766.950 375.300 769.050 377.400 ;
        RECT 767.250 371.700 768.450 375.300 ;
        RECT 766.950 369.600 769.050 371.700 ;
        RECT 770.400 367.050 771.450 382.950 ;
        RECT 769.950 364.950 772.050 367.050 ;
        RECT 760.950 349.950 763.050 352.050 ;
        RECT 772.950 346.950 775.050 349.050 ;
        RECT 754.950 341.250 756.750 342.150 ;
        RECT 757.950 340.950 760.050 343.050 ;
        RECT 761.250 341.250 762.750 342.150 ;
        RECT 763.950 340.950 766.050 343.050 ;
        RECT 767.250 341.250 769.050 342.150 ;
        RECT 769.950 340.950 772.050 343.050 ;
        RECT 739.950 338.250 742.050 339.150 ;
        RECT 742.950 338.850 745.050 339.750 ;
        RECT 745.950 337.950 748.050 340.050 ;
        RECT 754.950 337.950 757.050 340.050 ;
        RECT 758.250 338.850 759.750 339.750 ;
        RECT 760.950 337.950 763.050 340.050 ;
        RECT 764.250 338.850 765.750 339.750 ;
        RECT 766.950 337.950 769.050 340.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 733.950 325.950 736.050 328.050 ;
        RECT 742.950 319.950 745.050 322.050 ;
        RECT 743.400 313.050 744.450 319.950 ;
        RECT 730.950 310.950 733.050 313.050 ;
        RECT 736.950 310.950 739.050 313.050 ;
        RECT 740.250 311.250 741.750 312.150 ;
        RECT 742.950 310.950 745.050 313.050 ;
        RECT 727.950 304.950 730.050 307.050 ;
        RECT 727.950 274.950 730.050 277.050 ;
        RECT 724.950 247.950 727.050 250.050 ;
        RECT 728.400 244.050 729.450 274.950 ;
        RECT 731.400 244.050 732.450 310.950 ;
        RECT 733.950 307.950 736.050 310.050 ;
        RECT 737.250 308.850 738.750 309.750 ;
        RECT 739.950 307.950 742.050 310.050 ;
        RECT 743.250 308.850 745.050 309.750 ;
        RECT 733.950 305.850 736.050 306.750 ;
        RECT 746.400 282.450 747.450 337.950 ;
        RECT 755.400 331.050 756.450 337.950 ;
        RECT 754.950 328.950 757.050 331.050 ;
        RECT 755.400 328.050 756.450 328.950 ;
        RECT 754.950 325.950 757.050 328.050 ;
        RECT 748.950 322.950 751.050 325.050 ;
        RECT 743.400 281.400 747.450 282.450 ;
        RECT 733.950 277.950 736.050 280.050 ;
        RECT 734.400 274.050 735.450 277.950 ;
        RECT 733.950 271.950 736.050 274.050 ;
        RECT 737.250 272.250 738.750 273.150 ;
        RECT 739.950 271.950 742.050 274.050 ;
        RECT 733.950 269.850 735.750 270.750 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 740.250 269.850 742.050 270.750 ;
        RECT 736.950 259.950 739.050 262.050 ;
        RECT 727.950 241.950 730.050 244.050 ;
        RECT 730.950 241.950 733.050 244.050 ;
        RECT 727.950 240.450 730.050 241.050 ;
        RECT 725.400 239.400 730.050 240.450 ;
        RECT 725.400 235.050 726.450 239.400 ;
        RECT 727.950 238.950 730.050 239.400 ;
        RECT 731.250 239.250 732.750 240.150 ;
        RECT 733.950 238.950 736.050 241.050 ;
        RECT 737.400 238.050 738.450 259.950 ;
        RECT 739.950 241.950 742.050 244.050 ;
        RECT 727.950 236.850 729.750 237.750 ;
        RECT 730.950 235.950 733.050 238.050 ;
        RECT 734.250 236.850 735.750 237.750 ;
        RECT 736.950 235.950 739.050 238.050 ;
        RECT 724.950 232.950 727.050 235.050 ;
        RECT 727.950 232.950 730.050 235.050 ;
        RECT 721.950 229.950 724.050 232.050 ;
        RECT 728.400 211.050 729.450 232.950 ;
        RECT 731.400 229.050 732.450 235.950 ;
        RECT 736.950 233.850 739.050 234.750 ;
        RECT 730.950 226.950 733.050 229.050 ;
        RECT 721.950 208.950 724.050 211.050 ;
        RECT 727.950 208.950 730.050 211.050 ;
        RECT 722.400 195.450 723.450 208.950 ;
        RECT 727.950 205.950 730.050 208.050 ;
        RECT 728.400 199.050 729.450 205.950 ;
        RECT 733.950 200.250 736.050 201.150 ;
        RECT 724.950 197.250 726.750 198.150 ;
        RECT 727.950 196.950 730.050 199.050 ;
        RECT 731.250 197.250 732.750 198.150 ;
        RECT 733.950 196.950 736.050 199.050 ;
        RECT 724.950 195.450 727.050 196.050 ;
        RECT 722.400 194.400 727.050 195.450 ;
        RECT 728.250 194.850 729.750 195.750 ;
        RECT 724.950 193.950 727.050 194.400 ;
        RECT 730.950 193.950 733.050 196.050 ;
        RECT 703.950 190.950 706.050 193.050 ;
        RECT 718.950 190.950 721.050 193.050 ;
        RECT 719.400 190.050 720.450 190.950 ;
        RECT 718.950 187.950 721.050 190.050 ;
        RECT 697.950 175.950 700.050 178.050 ;
        RECT 703.950 175.950 706.050 178.050 ;
        RECT 698.400 172.050 699.450 175.950 ;
        RECT 691.950 169.950 694.050 172.050 ;
        RECT 697.950 169.950 700.050 172.050 ;
        RECT 691.950 168.450 694.050 169.050 ;
        RECT 689.400 167.400 694.050 168.450 ;
        RECT 689.400 133.050 690.450 167.400 ;
        RECT 691.950 166.950 694.050 167.400 ;
        RECT 695.250 167.250 697.050 168.150 ;
        RECT 697.950 167.850 700.050 168.750 ;
        RECT 700.950 167.250 703.050 168.150 ;
        RECT 691.950 164.850 693.750 165.750 ;
        RECT 694.950 163.950 697.050 166.050 ;
        RECT 697.950 163.950 700.050 166.050 ;
        RECT 700.950 163.950 703.050 166.050 ;
        RECT 695.400 163.050 696.450 163.950 ;
        RECT 694.950 160.950 697.050 163.050 ;
        RECT 688.950 130.950 691.050 133.050 ;
        RECT 698.400 132.450 699.450 163.950 ;
        RECT 704.400 163.050 705.450 175.950 ;
        RECT 706.950 172.950 709.050 175.050 ;
        RECT 707.400 172.050 708.450 172.950 ;
        RECT 706.950 169.950 709.050 172.050 ;
        RECT 709.950 169.950 712.050 172.050 ;
        RECT 707.400 166.050 708.450 169.950 ;
        RECT 710.400 169.050 711.450 169.950 ;
        RECT 709.950 166.950 712.050 169.050 ;
        RECT 713.250 167.250 714.750 168.150 ;
        RECT 715.950 166.950 718.050 169.050 ;
        RECT 719.400 166.050 720.450 187.950 ;
        RECT 731.400 181.050 732.450 193.950 ;
        RECT 733.950 190.950 736.050 193.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 721.950 166.950 724.050 169.050 ;
        RECT 730.950 168.450 733.050 169.050 ;
        RECT 728.400 167.400 733.050 168.450 ;
        RECT 706.950 163.950 709.050 166.050 ;
        RECT 709.950 164.850 711.750 165.750 ;
        RECT 712.950 163.950 715.050 166.050 ;
        RECT 716.250 164.850 717.750 165.750 ;
        RECT 718.950 163.950 721.050 166.050 ;
        RECT 713.400 163.050 714.450 163.950 ;
        RECT 722.400 163.050 723.450 166.950 ;
        RECT 728.400 163.050 729.450 167.400 ;
        RECT 730.950 166.950 733.050 167.400 ;
        RECT 730.950 164.850 733.050 165.750 ;
        RECT 703.950 160.950 706.050 163.050 ;
        RECT 706.950 162.450 709.050 163.050 ;
        RECT 706.950 161.400 711.450 162.450 ;
        RECT 706.950 160.950 709.050 161.400 ;
        RECT 710.400 159.450 711.450 161.400 ;
        RECT 712.950 160.950 715.050 163.050 ;
        RECT 715.950 160.950 718.050 163.050 ;
        RECT 718.950 161.850 721.050 162.750 ;
        RECT 721.950 160.950 724.050 163.050 ;
        RECT 727.950 160.950 730.050 163.050 ;
        RECT 716.400 159.450 717.450 160.950 ;
        RECT 710.400 158.400 717.450 159.450 ;
        RECT 695.400 131.400 699.450 132.450 ;
        RECT 691.950 127.950 694.050 130.050 ;
        RECT 640.950 126.450 643.050 127.050 ;
        RECT 638.400 125.400 643.050 126.450 ;
        RECT 638.400 124.050 639.450 125.400 ;
        RECT 640.950 124.950 643.050 125.400 ;
        RECT 644.250 125.250 645.750 126.150 ;
        RECT 646.950 124.950 649.050 127.050 ;
        RECT 650.250 125.250 652.050 126.150 ;
        RECT 658.950 124.950 661.050 127.050 ;
        RECT 664.950 124.950 667.050 127.050 ;
        RECT 676.950 124.950 679.050 127.050 ;
        RECT 679.950 124.950 682.050 127.050 ;
        RECT 683.250 125.250 684.750 126.150 ;
        RECT 685.950 124.950 688.050 127.050 ;
        RECT 689.250 125.250 691.050 126.150 ;
        RECT 637.950 121.950 640.050 124.050 ;
        RECT 643.950 121.950 646.050 124.050 ;
        RECT 647.250 122.850 648.750 123.750 ;
        RECT 649.950 121.950 652.050 124.050 ;
        RECT 644.400 121.050 645.450 121.950 ;
        RECT 643.950 118.950 646.050 121.050 ;
        RECT 650.400 115.050 651.450 121.950 ;
        RECT 649.950 112.950 652.050 115.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 653.400 100.050 654.450 100.950 ;
        RECT 625.950 97.950 628.050 100.050 ;
        RECT 631.950 97.950 634.050 100.050 ;
        RECT 652.950 97.950 655.050 100.050 ;
        RECT 655.950 97.950 658.050 100.050 ;
        RECT 626.400 97.050 627.450 97.950 ;
        RECT 625.950 94.950 628.050 97.050 ;
        RECT 629.250 95.250 630.750 96.150 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 649.950 95.250 652.050 96.150 ;
        RECT 652.950 95.850 655.050 96.750 ;
        RECT 625.950 92.850 627.750 93.750 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 632.250 92.850 633.750 93.750 ;
        RECT 634.950 91.950 637.050 94.050 ;
        RECT 649.950 91.950 652.050 94.050 ;
        RECT 631.950 88.950 634.050 91.050 ;
        RECT 634.950 89.850 637.050 90.750 ;
        RECT 632.400 85.050 633.450 88.950 ;
        RECT 631.950 82.950 634.050 85.050 ;
        RECT 628.950 64.950 631.050 67.050 ;
        RECT 611.400 59.400 615.450 60.450 ;
        RECT 589.950 55.950 592.050 58.050 ;
        RECT 595.950 57.450 598.050 58.050 ;
        RECT 593.250 56.250 594.750 57.150 ;
        RECT 595.950 56.400 600.450 57.450 ;
        RECT 595.950 55.950 598.050 56.400 ;
        RECT 571.950 53.850 573.750 54.750 ;
        RECT 574.950 52.950 577.050 55.050 ;
        RECT 580.950 52.950 583.050 55.050 ;
        RECT 586.950 52.950 589.050 55.050 ;
        RECT 589.950 53.850 591.750 54.750 ;
        RECT 592.950 52.950 595.050 55.050 ;
        RECT 596.250 53.850 598.050 54.750 ;
        RECT 575.400 52.050 576.450 52.950 ;
        RECT 581.400 52.050 582.450 52.950 ;
        RECT 599.400 52.050 600.450 56.400 ;
        RECT 601.950 52.950 604.050 55.050 ;
        RECT 574.950 49.950 577.050 52.050 ;
        RECT 580.950 49.950 583.050 52.050 ;
        RECT 598.950 49.950 601.050 52.050 ;
        RECT 602.400 40.050 603.450 52.950 ;
        RECT 601.950 37.950 604.050 40.050 ;
        RECT 568.950 22.950 571.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 602.400 22.050 603.450 37.950 ;
        RECT 607.950 28.950 610.050 31.050 ;
        RECT 481.950 19.950 484.050 22.050 ;
        RECT 493.950 19.950 496.050 22.050 ;
        RECT 499.950 19.950 502.050 22.050 ;
        RECT 505.950 20.850 507.750 21.750 ;
        RECT 508.950 19.950 511.050 22.050 ;
        RECT 512.250 20.850 513.750 21.750 ;
        RECT 514.950 19.950 517.050 22.050 ;
        RECT 529.950 19.950 532.050 22.050 ;
        RECT 544.950 20.250 546.750 21.150 ;
        RECT 547.950 19.950 550.050 22.050 ;
        RECT 551.250 20.250 553.050 21.150 ;
        RECT 562.950 20.850 565.050 21.750 ;
        RECT 568.950 20.850 571.050 21.750 ;
        RECT 577.950 20.850 580.050 21.750 ;
        RECT 583.950 20.850 586.050 21.750 ;
        RECT 598.950 20.250 600.750 21.150 ;
        RECT 601.950 19.950 604.050 22.050 ;
        RECT 605.250 20.250 607.050 21.150 ;
        RECT 448.950 16.950 451.050 19.050 ;
        RECT 454.950 16.950 457.050 19.050 ;
        RECT 458.250 17.850 459.750 18.750 ;
        RECT 460.950 16.950 463.050 19.050 ;
        RECT 472.950 16.950 475.050 19.050 ;
        RECT 476.250 17.850 477.750 18.750 ;
        RECT 478.950 16.950 481.050 19.050 ;
        RECT 482.250 17.850 484.050 18.750 ;
        RECT 514.950 17.850 517.050 18.750 ;
        RECT 544.950 16.950 547.050 19.050 ;
        RECT 548.250 17.850 549.750 18.750 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 598.950 16.950 601.050 19.050 ;
        RECT 602.250 17.850 603.750 18.750 ;
        RECT 604.950 18.450 607.050 19.050 ;
        RECT 608.400 18.450 609.450 28.950 ;
        RECT 611.400 25.050 612.450 59.400 ;
        RECT 619.950 59.250 622.050 60.150 ;
        RECT 622.950 58.950 625.050 61.050 ;
        RECT 625.950 58.950 628.050 61.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 617.250 56.250 618.750 57.150 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 623.250 56.250 625.050 57.150 ;
        RECT 613.950 53.850 615.750 54.750 ;
        RECT 616.950 52.950 619.050 55.050 ;
        RECT 622.950 54.450 625.050 55.050 ;
        RECT 626.400 54.450 627.450 58.950 ;
        RECT 629.400 55.050 630.450 64.950 ;
        RECT 632.400 59.400 648.450 60.450 ;
        RECT 622.950 53.400 627.450 54.450 ;
        RECT 622.950 52.950 625.050 53.400 ;
        RECT 628.950 52.950 631.050 55.050 ;
        RECT 632.400 52.050 633.450 59.400 ;
        RECT 634.950 56.250 637.050 57.150 ;
        RECT 634.950 52.950 637.050 55.050 ;
        RECT 638.250 53.250 639.750 54.150 ;
        RECT 640.950 52.950 643.050 55.050 ;
        RECT 644.250 53.250 646.050 54.150 ;
        RECT 631.950 49.950 634.050 52.050 ;
        RECT 625.950 46.950 628.050 49.050 ;
        RECT 626.400 43.050 627.450 46.950 ;
        RECT 635.400 46.050 636.450 52.950 ;
        RECT 637.950 49.950 640.050 52.050 ;
        RECT 641.250 50.850 642.750 51.750 ;
        RECT 643.950 49.950 646.050 52.050 ;
        RECT 634.950 43.950 637.050 46.050 ;
        RECT 644.400 45.450 645.450 49.950 ;
        RECT 647.400 49.050 648.450 59.400 ;
        RECT 656.400 55.050 657.450 97.950 ;
        RECT 659.400 94.050 660.450 124.950 ;
        RECT 661.950 122.250 664.050 123.150 ;
        RECT 664.950 122.850 667.050 123.750 ;
        RECT 661.950 118.950 664.050 121.050 ;
        RECT 677.400 112.050 678.450 124.950 ;
        RECT 680.400 124.050 681.450 124.950 ;
        RECT 679.950 121.950 682.050 124.050 ;
        RECT 682.950 121.950 685.050 124.050 ;
        RECT 686.250 122.850 687.750 123.750 ;
        RECT 688.950 123.450 691.050 124.050 ;
        RECT 692.400 123.450 693.450 127.950 ;
        RECT 688.950 122.400 693.450 123.450 ;
        RECT 688.950 121.950 691.050 122.400 ;
        RECT 683.400 121.050 684.450 121.950 ;
        RECT 682.950 118.950 685.050 121.050 ;
        RECT 676.950 109.950 679.050 112.050 ;
        RECT 664.950 103.950 667.050 106.050 ;
        RECT 665.400 97.050 666.450 103.950 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 670.950 97.950 673.050 100.050 ;
        RECT 689.400 97.050 690.450 100.950 ;
        RECT 695.400 97.050 696.450 131.400 ;
        RECT 718.950 130.950 721.050 133.050 ;
        RECT 730.950 130.950 733.050 133.050 ;
        RECT 697.950 127.950 700.050 130.050 ;
        RECT 715.950 127.950 718.050 130.050 ;
        RECT 698.400 127.050 699.450 127.950 ;
        RECT 697.950 124.950 700.050 127.050 ;
        RECT 703.950 124.950 706.050 127.050 ;
        RECT 707.250 125.250 709.050 126.150 ;
        RECT 709.950 124.950 712.050 127.050 ;
        RECT 697.950 122.850 700.050 123.750 ;
        RECT 700.950 122.250 703.050 123.150 ;
        RECT 703.950 122.850 705.750 123.750 ;
        RECT 706.950 121.950 709.050 124.050 ;
        RECT 700.950 118.950 703.050 121.050 ;
        RECT 701.400 112.050 702.450 118.950 ;
        RECT 700.950 109.950 703.050 112.050 ;
        RECT 707.400 103.050 708.450 121.950 ;
        RECT 710.400 121.050 711.450 124.950 ;
        RECT 716.400 121.050 717.450 127.950 ;
        RECT 709.950 118.950 712.050 121.050 ;
        RECT 715.950 118.950 718.050 121.050 ;
        RECT 715.950 112.950 718.050 115.050 ;
        RECT 706.950 100.950 709.050 103.050 ;
        RECT 697.950 97.950 700.050 100.050 ;
        RECT 664.950 94.950 667.050 97.050 ;
        RECT 668.250 95.250 670.050 96.150 ;
        RECT 670.950 95.850 673.050 96.750 ;
        RECT 673.950 95.250 676.050 96.150 ;
        RECT 688.950 94.950 691.050 97.050 ;
        RECT 692.250 95.250 693.750 96.150 ;
        RECT 694.950 94.950 697.050 97.050 ;
        RECT 698.400 94.050 699.450 97.950 ;
        RECT 716.400 97.050 717.450 112.950 ;
        RECT 719.400 100.050 720.450 130.950 ;
        RECT 721.950 125.250 724.050 126.150 ;
        RECT 727.950 125.250 730.050 126.150 ;
        RECT 721.950 121.950 724.050 124.050 ;
        RECT 727.950 121.950 730.050 124.050 ;
        RECT 722.400 121.050 723.450 121.950 ;
        RECT 721.950 118.950 724.050 121.050 ;
        RECT 728.400 118.050 729.450 121.950 ;
        RECT 727.950 115.950 730.050 118.050 ;
        RECT 727.950 103.950 730.050 106.050 ;
        RECT 724.950 100.950 727.050 103.050 ;
        RECT 718.950 97.950 721.050 100.050 ;
        RECT 706.950 94.950 709.050 97.050 ;
        RECT 709.950 94.950 712.050 97.050 ;
        RECT 713.250 95.250 714.750 96.150 ;
        RECT 715.950 94.950 718.050 97.050 ;
        RECT 707.400 94.050 708.450 94.950 ;
        RECT 719.400 94.050 720.450 97.950 ;
        RECT 725.400 94.050 726.450 100.950 ;
        RECT 728.400 97.050 729.450 103.950 ;
        RECT 731.400 100.050 732.450 130.950 ;
        RECT 734.400 130.050 735.450 190.950 ;
        RECT 736.950 169.950 739.050 172.050 ;
        RECT 737.400 169.050 738.450 169.950 ;
        RECT 736.950 166.950 739.050 169.050 ;
        RECT 736.950 164.850 739.050 165.750 ;
        RECT 736.950 160.950 739.050 163.050 ;
        RECT 733.950 127.950 736.050 130.050 ;
        RECT 734.400 127.050 735.450 127.950 ;
        RECT 733.950 124.950 736.050 127.050 ;
        RECT 737.400 118.050 738.450 160.950 ;
        RECT 740.400 133.050 741.450 241.950 ;
        RECT 743.400 163.050 744.450 281.400 ;
        RECT 745.950 274.950 748.050 277.050 ;
        RECT 746.400 271.050 747.450 274.950 ;
        RECT 749.400 274.050 750.450 322.950 ;
        RECT 757.950 319.950 760.050 322.050 ;
        RECT 751.950 316.950 754.050 319.050 ;
        RECT 752.400 313.050 753.450 316.950 ;
        RECT 758.400 313.050 759.450 319.950 ;
        RECT 761.400 319.050 762.450 337.950 ;
        RECT 770.400 337.050 771.450 340.950 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 760.950 316.950 763.050 319.050 ;
        RECT 763.950 316.950 766.050 319.050 ;
        RECT 766.950 316.950 769.050 319.050 ;
        RECT 764.400 313.050 765.450 316.950 ;
        RECT 751.950 310.950 754.050 313.050 ;
        RECT 757.950 310.950 760.050 313.050 ;
        RECT 761.250 311.250 762.750 312.150 ;
        RECT 763.950 310.950 766.050 313.050 ;
        RECT 754.950 309.450 757.050 310.050 ;
        RECT 752.400 308.400 757.050 309.450 ;
        RECT 758.250 308.850 759.750 309.750 ;
        RECT 752.400 304.050 753.450 308.400 ;
        RECT 754.950 307.950 757.050 308.400 ;
        RECT 760.950 307.950 763.050 310.050 ;
        RECT 764.250 308.850 766.050 309.750 ;
        RECT 761.400 307.050 762.450 307.950 ;
        RECT 754.950 305.850 757.050 306.750 ;
        RECT 760.950 304.950 763.050 307.050 ;
        RECT 751.950 301.950 754.050 304.050 ;
        RECT 760.950 286.950 763.050 289.050 ;
        RECT 754.950 274.950 757.050 277.050 ;
        RECT 748.950 271.950 751.050 274.050 ;
        RECT 745.950 268.950 748.050 271.050 ;
        RECT 749.400 265.050 750.450 271.950 ;
        RECT 755.400 271.050 756.450 274.950 ;
        RECT 761.400 271.050 762.450 286.950 ;
        RECT 751.950 269.250 753.750 270.150 ;
        RECT 754.950 268.950 757.050 271.050 ;
        RECT 758.250 269.250 759.750 270.150 ;
        RECT 760.950 268.950 763.050 271.050 ;
        RECT 764.250 269.250 766.050 270.150 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 755.250 266.850 756.750 267.750 ;
        RECT 757.950 265.950 760.050 268.050 ;
        RECT 761.250 266.850 762.750 267.750 ;
        RECT 763.950 265.950 766.050 268.050 ;
        RECT 748.950 262.950 751.050 265.050 ;
        RECT 752.400 253.050 753.450 265.950 ;
        RECT 764.400 265.050 765.450 265.950 ;
        RECT 757.950 262.950 760.050 265.050 ;
        RECT 763.950 262.950 766.050 265.050 ;
        RECT 751.950 250.950 754.050 253.050 ;
        RECT 752.400 244.050 753.450 250.950 ;
        RECT 751.950 241.950 754.050 244.050 ;
        RECT 751.950 240.450 754.050 241.050 ;
        RECT 749.400 239.400 754.050 240.450 ;
        RECT 749.400 229.050 750.450 239.400 ;
        RECT 751.950 238.950 754.050 239.400 ;
        RECT 751.950 236.850 754.050 237.750 ;
        RECT 754.950 236.250 757.050 237.150 ;
        RECT 754.950 232.950 757.050 235.050 ;
        RECT 755.400 232.050 756.450 232.950 ;
        RECT 754.950 229.950 757.050 232.050 ;
        RECT 748.950 226.950 751.050 229.050 ;
        RECT 754.950 217.950 757.050 220.050 ;
        RECT 745.950 197.250 748.050 198.150 ;
        RECT 751.950 197.250 754.050 198.150 ;
        RECT 745.950 193.950 748.050 196.050 ;
        RECT 749.250 194.250 750.750 195.150 ;
        RECT 751.950 193.950 754.050 196.050 ;
        RECT 746.400 172.050 747.450 193.950 ;
        RECT 752.400 193.050 753.450 193.950 ;
        RECT 748.950 190.950 751.050 193.050 ;
        RECT 751.950 190.950 754.050 193.050 ;
        RECT 749.400 187.050 750.450 190.950 ;
        RECT 748.950 184.950 751.050 187.050 ;
        RECT 745.950 169.950 748.050 172.050 ;
        RECT 748.950 169.950 751.050 172.050 ;
        RECT 748.950 167.850 751.050 168.750 ;
        RECT 751.950 167.250 754.050 168.150 ;
        RECT 751.950 163.950 754.050 166.050 ;
        RECT 742.950 160.950 745.050 163.050 ;
        RECT 752.400 160.050 753.450 163.950 ;
        RECT 751.950 157.950 754.050 160.050 ;
        RECT 751.950 142.950 754.050 145.050 ;
        RECT 739.950 130.950 742.050 133.050 ;
        RECT 739.950 128.250 742.050 129.150 ;
        RECT 739.950 124.950 742.050 127.050 ;
        RECT 743.250 125.250 744.750 126.150 ;
        RECT 745.950 124.950 748.050 127.050 ;
        RECT 749.250 125.250 751.050 126.150 ;
        RECT 742.950 121.950 745.050 124.050 ;
        RECT 746.250 122.850 747.750 123.750 ;
        RECT 748.950 123.450 751.050 124.050 ;
        RECT 752.400 123.450 753.450 142.950 ;
        RECT 755.400 136.050 756.450 217.950 ;
        RECT 758.400 145.050 759.450 262.950 ;
        RECT 760.950 247.950 763.050 250.050 ;
        RECT 767.400 249.450 768.450 316.950 ;
        RECT 770.400 271.050 771.450 334.950 ;
        RECT 773.400 319.050 774.450 346.950 ;
        RECT 772.950 316.950 775.050 319.050 ;
        RECT 776.400 316.050 777.450 409.950 ;
        RECT 779.400 403.050 780.450 451.950 ;
        RECT 782.400 406.050 783.450 580.950 ;
        RECT 788.400 571.050 789.450 604.950 ;
        RECT 797.400 601.050 798.450 607.950 ;
        RECT 800.400 601.050 801.450 673.950 ;
        RECT 806.250 671.250 807.750 672.150 ;
        RECT 808.950 670.950 811.050 673.050 ;
        RECT 812.400 670.050 813.450 694.950 ;
        RECT 802.950 668.850 804.750 669.750 ;
        RECT 805.950 667.950 808.050 670.050 ;
        RECT 809.250 668.850 810.750 669.750 ;
        RECT 811.950 667.950 814.050 670.050 ;
        RECT 802.950 664.950 805.050 667.050 ;
        RECT 803.400 619.050 804.450 664.950 ;
        RECT 806.400 664.050 807.450 667.950 ;
        RECT 811.950 665.850 814.050 666.750 ;
        RECT 805.950 661.950 808.050 664.050 ;
        RECT 811.950 661.950 814.050 664.050 ;
        RECT 808.950 628.950 811.050 631.050 ;
        RECT 805.950 626.250 808.050 627.150 ;
        RECT 808.950 626.850 811.050 627.750 ;
        RECT 805.950 622.950 808.050 625.050 ;
        RECT 808.950 622.950 811.050 625.050 ;
        RECT 802.950 616.950 805.050 619.050 ;
        RECT 802.950 605.400 805.050 607.500 ;
        RECT 790.950 600.450 793.050 601.050 ;
        RECT 793.950 600.450 796.050 601.050 ;
        RECT 790.950 599.400 796.050 600.450 ;
        RECT 790.950 598.950 793.050 599.400 ;
        RECT 793.950 598.950 796.050 599.400 ;
        RECT 796.950 598.950 799.050 601.050 ;
        RECT 799.950 598.950 802.050 601.050 ;
        RECT 790.950 596.850 793.050 597.750 ;
        RECT 787.950 568.950 790.050 571.050 ;
        RECT 794.400 559.050 795.450 598.950 ;
        RECT 796.950 596.850 799.050 597.750 ;
        RECT 803.400 588.600 804.600 605.400 ;
        RECT 802.950 586.500 805.050 588.600 ;
        RECT 809.400 583.050 810.450 622.950 ;
        RECT 812.400 607.050 813.450 661.950 ;
        RECT 815.400 625.050 816.450 697.950 ;
        RECT 817.950 694.950 820.050 697.050 ;
        RECT 814.950 622.950 817.050 625.050 ;
        RECT 818.400 613.050 819.450 694.950 ;
        RECT 821.400 667.050 822.450 766.950 ;
        RECT 824.400 766.050 825.450 772.950 ;
        RECT 827.400 769.050 828.450 838.950 ;
        RECT 826.950 766.950 829.050 769.050 ;
        RECT 823.950 763.950 826.050 766.050 ;
        RECT 833.400 748.050 834.450 844.950 ;
        RECT 847.950 842.250 850.050 843.150 ;
        RECT 850.950 842.850 853.050 843.750 ;
        RECT 847.950 838.950 850.050 841.050 ;
        RECT 848.400 838.050 849.450 838.950 ;
        RECT 847.950 835.950 850.050 838.050 ;
        RECT 857.400 820.050 858.450 844.950 ;
        RECT 856.950 817.950 859.050 820.050 ;
        RECT 859.950 814.950 862.050 817.050 ;
        RECT 860.400 814.050 861.450 814.950 ;
        RECT 838.950 812.250 840.750 813.150 ;
        RECT 841.950 811.950 844.050 814.050 ;
        RECT 845.250 812.250 847.050 813.150 ;
        RECT 856.950 812.250 858.750 813.150 ;
        RECT 859.950 811.950 862.050 814.050 ;
        RECT 863.250 812.250 865.050 813.150 ;
        RECT 842.250 809.850 843.750 810.750 ;
        RECT 860.250 809.850 861.750 810.750 ;
        RECT 856.950 805.950 859.050 808.050 ;
        RECT 857.400 781.050 858.450 805.950 ;
        RECT 856.950 778.950 859.050 781.050 ;
        RECT 859.950 780.450 862.050 781.050 ;
        RECT 862.950 780.450 865.050 781.050 ;
        RECT 859.950 779.400 865.050 780.450 ;
        RECT 859.950 778.950 862.050 779.400 ;
        RECT 862.950 778.950 865.050 779.400 ;
        RECT 842.250 776.250 843.750 777.150 ;
        RECT 857.250 776.250 858.750 777.150 ;
        RECT 838.950 773.850 840.750 774.750 ;
        RECT 841.950 772.950 844.050 775.050 ;
        RECT 845.250 773.850 847.050 774.750 ;
        RECT 853.950 773.850 855.750 774.750 ;
        RECT 856.950 772.950 859.050 775.050 ;
        RECT 860.250 773.850 862.050 774.750 ;
        RECT 832.950 745.950 835.050 748.050 ;
        RECT 838.950 747.450 841.050 748.050 ;
        RECT 842.400 747.450 843.450 772.950 ;
        RECT 853.950 769.950 856.050 772.050 ;
        RECT 838.950 746.400 843.450 747.450 ;
        RECT 838.950 745.950 841.050 746.400 ;
        RECT 823.950 740.250 825.750 741.150 ;
        RECT 826.950 739.950 829.050 742.050 ;
        RECT 830.250 740.250 832.050 741.150 ;
        RECT 835.950 739.950 838.050 742.050 ;
        RECT 838.950 740.250 840.750 741.150 ;
        RECT 841.950 739.950 844.050 742.050 ;
        RECT 845.250 740.250 847.050 741.150 ;
        RECT 827.250 737.850 828.750 738.750 ;
        RECT 829.950 733.950 832.050 736.050 ;
        RECT 830.400 709.050 831.450 733.950 ;
        RECT 836.400 712.050 837.450 739.950 ;
        RECT 842.250 737.850 843.750 738.750 ;
        RECT 838.950 730.950 841.050 733.050 ;
        RECT 835.950 709.950 838.050 712.050 ;
        RECT 839.400 709.050 840.450 730.950 ;
        RECT 841.950 709.950 844.050 712.050 ;
        RECT 823.950 706.950 826.050 709.050 ;
        RECT 829.950 706.950 832.050 709.050 ;
        RECT 838.950 706.950 841.050 709.050 ;
        RECT 824.400 679.050 825.450 706.950 ;
        RECT 829.950 705.450 832.050 706.050 ;
        RECT 827.400 704.400 832.050 705.450 ;
        RECT 835.950 705.450 838.050 706.050 ;
        RECT 827.400 694.050 828.450 704.400 ;
        RECT 829.950 703.950 832.050 704.400 ;
        RECT 833.250 704.250 834.750 705.150 ;
        RECT 835.950 704.400 840.450 705.450 ;
        RECT 835.950 703.950 838.050 704.400 ;
        RECT 829.950 701.850 831.750 702.750 ;
        RECT 832.950 700.950 835.050 703.050 ;
        RECT 836.250 701.850 838.050 702.750 ;
        RECT 839.400 700.050 840.450 704.400 ;
        RECT 835.950 697.950 838.050 700.050 ;
        RECT 838.950 697.950 841.050 700.050 ;
        RECT 826.950 691.950 829.050 694.050 ;
        RECT 823.950 676.950 826.050 679.050 ;
        RECT 823.950 673.950 826.050 676.050 ;
        RECT 823.950 671.850 825.750 672.750 ;
        RECT 826.950 672.450 829.050 673.050 ;
        RECT 826.950 671.400 831.450 672.450 ;
        RECT 826.950 670.950 829.050 671.400 ;
        RECT 826.950 668.850 829.050 669.750 ;
        RECT 820.950 664.950 823.050 667.050 ;
        RECT 830.400 661.050 831.450 671.400 ;
        RECT 832.950 671.250 835.050 672.150 ;
        RECT 832.950 669.450 835.050 670.050 ;
        RECT 836.400 669.450 837.450 697.950 ;
        RECT 838.950 676.950 841.050 679.050 ;
        RECT 832.950 668.400 837.450 669.450 ;
        RECT 832.950 667.950 835.050 668.400 ;
        RECT 829.950 658.950 832.050 661.050 ;
        RECT 832.950 643.950 835.050 646.050 ;
        RECT 829.950 632.250 832.050 633.150 ;
        RECT 820.950 629.250 822.750 630.150 ;
        RECT 823.950 628.950 826.050 631.050 ;
        RECT 829.950 630.450 832.050 631.050 ;
        RECT 833.400 630.450 834.450 643.950 ;
        RECT 827.250 629.250 828.750 630.150 ;
        RECT 829.950 629.400 834.450 630.450 ;
        RECT 829.950 628.950 832.050 629.400 ;
        RECT 824.250 626.850 825.750 627.750 ;
        RECT 826.950 625.950 829.050 628.050 ;
        RECT 820.950 616.950 823.050 619.050 ;
        RECT 817.950 610.950 820.050 613.050 ;
        RECT 811.950 604.950 814.050 607.050 ;
        RECT 817.950 605.400 820.050 607.500 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 602.250 817.050 603.150 ;
        RECT 812.400 600.450 813.450 601.950 ;
        RECT 814.950 600.450 817.050 601.050 ;
        RECT 812.400 599.400 817.050 600.450 ;
        RECT 814.950 598.950 817.050 599.400 ;
        RECT 811.950 595.950 814.050 598.050 ;
        RECT 808.950 580.950 811.050 583.050 ;
        RECT 812.400 564.450 813.450 595.950 ;
        RECT 815.400 574.050 816.450 598.950 ;
        RECT 818.550 593.400 819.750 605.400 ;
        RECT 817.950 591.300 820.050 593.400 ;
        RECT 818.550 587.700 819.750 591.300 ;
        RECT 817.950 585.600 820.050 587.700 ;
        RECT 814.950 571.950 817.050 574.050 ;
        RECT 817.950 567.300 820.050 569.400 ;
        RECT 809.400 563.400 813.450 564.450 ;
        RECT 818.550 563.700 819.750 567.300 ;
        RECT 784.950 556.950 787.050 559.050 ;
        RECT 793.950 556.950 796.050 559.050 ;
        RECT 784.950 554.850 787.050 555.750 ;
        RECT 805.950 554.850 808.050 555.750 ;
        RECT 784.950 535.950 787.050 538.050 ;
        RECT 785.400 472.050 786.450 535.950 ;
        RECT 790.950 533.400 793.050 535.500 ;
        RECT 791.400 516.600 792.600 533.400 ;
        RECT 796.950 532.950 799.050 535.050 ;
        RECT 797.400 529.050 798.450 532.950 ;
        RECT 799.950 529.950 802.050 532.050 ;
        RECT 793.950 526.950 796.050 529.050 ;
        RECT 796.950 526.950 799.050 529.050 ;
        RECT 800.400 528.450 801.450 529.950 ;
        RECT 802.950 528.450 805.050 529.050 ;
        RECT 800.400 527.400 805.050 528.450 ;
        RECT 790.950 514.500 793.050 516.600 ;
        RECT 794.400 492.450 795.450 526.950 ;
        RECT 796.950 524.850 799.050 525.750 ;
        RECT 794.400 491.400 798.450 492.450 ;
        RECT 791.250 488.250 792.750 489.150 ;
        RECT 787.950 485.850 789.750 486.750 ;
        RECT 790.950 484.950 793.050 487.050 ;
        RECT 794.250 485.850 796.050 486.750 ;
        RECT 791.400 481.050 792.450 484.950 ;
        RECT 790.950 478.950 793.050 481.050 ;
        RECT 784.950 469.950 787.050 472.050 ;
        RECT 784.950 461.400 787.050 463.500 ;
        RECT 785.250 449.400 786.450 461.400 ;
        RECT 787.950 458.250 790.050 459.150 ;
        RECT 787.950 454.950 790.050 457.050 ;
        RECT 784.950 447.300 787.050 449.400 ;
        RECT 785.250 443.700 786.450 447.300 ;
        RECT 784.950 441.600 787.050 443.700 ;
        RECT 788.400 415.050 789.450 454.950 ;
        RECT 797.400 415.050 798.450 491.400 ;
        RECT 800.400 453.450 801.450 527.400 ;
        RECT 802.950 526.950 805.050 527.400 ;
        RECT 802.950 524.850 805.050 525.750 ;
        RECT 805.950 484.950 808.050 487.050 ;
        RECT 802.950 482.250 805.050 483.150 ;
        RECT 805.950 482.850 808.050 483.750 ;
        RECT 802.950 478.950 805.050 481.050 ;
        RECT 803.400 460.050 804.450 478.950 ;
        RECT 802.950 457.950 805.050 460.050 ;
        RECT 802.950 455.250 805.050 456.150 ;
        RECT 802.950 453.450 805.050 454.050 ;
        RECT 800.400 452.400 805.050 453.450 ;
        RECT 802.950 451.950 805.050 452.400 ;
        RECT 805.950 423.300 808.050 425.400 ;
        RECT 806.550 419.700 807.750 423.300 ;
        RECT 805.950 417.600 808.050 419.700 ;
        RECT 787.950 412.950 790.050 415.050 ;
        RECT 793.950 414.450 796.050 415.050 ;
        RECT 791.400 413.400 796.050 414.450 ;
        RECT 787.950 410.850 790.050 411.750 ;
        RECT 781.950 403.950 784.050 406.050 ;
        RECT 778.950 400.950 781.050 403.050 ;
        RECT 784.950 383.250 787.050 384.150 ;
        RECT 784.950 379.950 787.050 382.050 ;
        RECT 778.950 370.950 781.050 373.050 ;
        RECT 779.400 349.050 780.450 370.950 ;
        RECT 791.400 355.050 792.450 413.400 ;
        RECT 793.950 412.950 796.050 413.400 ;
        RECT 796.950 412.950 799.050 415.050 ;
        RECT 793.950 410.850 796.050 411.750 ;
        RECT 796.950 409.950 799.050 412.050 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 790.950 352.950 793.050 355.050 ;
        RECT 797.400 352.050 798.450 409.950 ;
        RECT 802.950 407.850 805.050 408.750 ;
        RECT 802.950 403.950 805.050 406.050 ;
        RECT 806.550 405.600 807.750 417.600 ;
        RECT 796.950 349.950 799.050 352.050 ;
        RECT 778.950 346.950 781.050 349.050 ;
        RECT 779.400 346.050 780.450 346.950 ;
        RECT 797.400 346.050 798.450 349.950 ;
        RECT 778.950 343.950 781.050 346.050 ;
        RECT 782.250 344.250 783.750 345.150 ;
        RECT 784.950 343.950 787.050 346.050 ;
        RECT 787.950 343.950 790.050 346.050 ;
        RECT 790.950 343.950 793.050 346.050 ;
        RECT 796.950 343.950 799.050 346.050 ;
        RECT 778.950 341.850 780.750 342.750 ;
        RECT 781.950 340.950 784.050 343.050 ;
        RECT 785.250 341.850 787.050 342.750 ;
        RECT 782.400 340.050 783.450 340.950 ;
        RECT 781.950 337.950 784.050 340.050 ;
        RECT 781.950 328.950 784.050 331.050 ;
        RECT 772.950 313.950 775.050 316.050 ;
        RECT 775.950 313.950 778.050 316.050 ;
        RECT 778.950 313.950 781.050 316.050 ;
        RECT 772.950 311.850 775.050 312.750 ;
        RECT 775.950 311.250 778.050 312.150 ;
        RECT 772.950 307.950 775.050 310.050 ;
        RECT 775.950 307.950 778.050 310.050 ;
        RECT 769.950 268.950 772.050 271.050 ;
        RECT 769.950 265.950 772.050 268.050 ;
        RECT 764.400 248.400 768.450 249.450 ;
        RECT 761.400 241.050 762.450 247.950 ;
        RECT 760.950 238.950 763.050 241.050 ;
        RECT 760.950 236.850 763.050 237.750 ;
        RECT 760.950 232.950 763.050 235.050 ;
        RECT 761.400 220.050 762.450 232.950 ;
        RECT 760.950 217.950 763.050 220.050 ;
        RECT 764.400 214.050 765.450 248.400 ;
        RECT 766.950 244.950 769.050 247.050 ;
        RECT 767.400 229.050 768.450 244.950 ;
        RECT 766.950 226.950 769.050 229.050 ;
        RECT 763.950 211.950 766.050 214.050 ;
        RECT 770.400 208.050 771.450 265.950 ;
        RECT 773.400 241.050 774.450 307.950 ;
        RECT 779.400 307.050 780.450 313.950 ;
        RECT 778.950 304.950 781.050 307.050 ;
        RECT 775.950 268.950 778.050 271.050 ;
        RECT 775.950 266.850 778.050 267.750 ;
        RECT 778.950 266.250 781.050 267.150 ;
        RECT 778.950 262.950 781.050 265.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 772.950 238.950 775.050 241.050 ;
        RECT 772.950 237.450 775.050 238.050 ;
        RECT 776.400 237.450 777.450 256.950 ;
        RECT 779.400 253.050 780.450 262.950 ;
        RECT 778.950 250.950 781.050 253.050 ;
        RECT 778.950 247.950 781.050 250.050 ;
        RECT 779.400 238.050 780.450 247.950 ;
        RECT 782.400 247.050 783.450 328.950 ;
        RECT 784.950 316.950 787.050 319.050 ;
        RECT 785.400 306.450 786.450 316.950 ;
        RECT 788.400 313.050 789.450 343.950 ;
        RECT 791.400 316.050 792.450 343.950 ;
        RECT 797.400 343.050 798.450 343.950 ;
        RECT 796.950 340.950 799.050 343.050 ;
        RECT 800.250 341.250 802.050 342.150 ;
        RECT 796.950 338.850 798.750 339.750 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 790.950 313.950 793.050 316.050 ;
        RECT 787.950 310.950 790.050 313.050 ;
        RECT 791.250 311.850 792.750 312.750 ;
        RECT 793.950 312.450 796.050 313.050 ;
        RECT 793.950 311.400 798.450 312.450 ;
        RECT 793.950 310.950 796.050 311.400 ;
        RECT 797.400 310.050 798.450 311.400 ;
        RECT 787.950 308.850 790.050 309.750 ;
        RECT 793.950 308.850 796.050 309.750 ;
        RECT 796.950 307.950 799.050 310.050 ;
        RECT 785.400 305.400 789.450 306.450 ;
        RECT 784.950 301.950 787.050 304.050 ;
        RECT 785.400 262.050 786.450 301.950 ;
        RECT 788.400 289.050 789.450 305.400 ;
        RECT 787.950 286.950 790.050 289.050 ;
        RECT 793.950 283.950 796.050 286.050 ;
        RECT 787.950 277.950 790.050 280.050 ;
        RECT 784.950 259.950 787.050 262.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 781.950 244.950 784.050 247.050 ;
        RECT 772.950 236.400 777.450 237.450 ;
        RECT 772.950 235.950 775.050 236.400 ;
        RECT 778.950 235.950 781.050 238.050 ;
        RECT 782.250 236.250 784.050 237.150 ;
        RECT 772.950 233.850 774.750 234.750 ;
        RECT 775.950 232.950 778.050 235.050 ;
        RECT 779.250 233.850 780.750 234.750 ;
        RECT 781.950 232.950 784.050 235.050 ;
        RECT 775.950 230.850 778.050 231.750 ;
        RECT 778.950 229.950 781.050 232.050 ;
        RECT 772.950 226.950 775.050 229.050 ;
        RECT 769.950 205.950 772.050 208.050 ;
        RECT 769.950 202.950 772.050 205.050 ;
        RECT 770.400 202.050 771.450 202.950 ;
        RECT 763.950 199.950 766.050 202.050 ;
        RECT 767.250 200.250 768.750 201.150 ;
        RECT 769.950 199.950 772.050 202.050 ;
        RECT 763.950 197.850 765.750 198.750 ;
        RECT 766.950 196.950 769.050 199.050 ;
        RECT 770.250 197.850 772.050 198.750 ;
        RECT 769.950 175.950 772.050 178.050 ;
        RECT 763.950 171.450 766.050 172.050 ;
        RECT 761.400 170.400 766.050 171.450 ;
        RECT 757.950 142.950 760.050 145.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 754.950 127.950 757.050 130.050 ;
        RECT 755.400 124.050 756.450 127.950 ;
        RECT 758.400 127.050 759.450 142.950 ;
        RECT 761.400 127.050 762.450 170.400 ;
        RECT 763.950 169.950 766.050 170.400 ;
        RECT 763.950 167.850 766.050 168.750 ;
        RECT 766.950 167.250 769.050 168.150 ;
        RECT 766.950 165.450 769.050 166.050 ;
        RECT 770.400 165.450 771.450 175.950 ;
        RECT 766.950 164.400 771.450 165.450 ;
        RECT 766.950 163.950 769.050 164.400 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 763.950 127.950 766.050 130.050 ;
        RECT 764.400 127.050 765.450 127.950 ;
        RECT 757.950 124.950 760.050 127.050 ;
        RECT 760.950 124.950 763.050 127.050 ;
        RECT 763.950 124.950 766.050 127.050 ;
        RECT 767.250 125.250 769.050 126.150 ;
        RECT 748.950 122.400 753.450 123.450 ;
        RECT 748.950 121.950 751.050 122.400 ;
        RECT 754.950 121.950 757.050 124.050 ;
        RECT 757.950 122.850 760.050 123.750 ;
        RECT 760.950 122.250 763.050 123.150 ;
        RECT 763.950 122.850 765.750 123.750 ;
        RECT 766.950 121.950 769.050 124.050 ;
        RECT 767.400 121.050 768.450 121.950 ;
        RECT 760.950 118.950 763.050 121.050 ;
        RECT 766.950 118.950 769.050 121.050 ;
        RECT 736.950 115.950 739.050 118.050 ;
        RECT 766.950 115.950 769.050 118.050 ;
        RECT 748.950 100.950 751.050 103.050 ;
        RECT 749.400 100.050 750.450 100.950 ;
        RECT 730.950 97.950 733.050 100.050 ;
        RECT 736.950 97.950 739.050 100.050 ;
        RECT 742.950 97.950 745.050 100.050 ;
        RECT 748.950 97.950 751.050 100.050 ;
        RECT 763.950 97.950 766.050 100.050 ;
        RECT 727.950 94.950 730.050 97.050 ;
        RECT 731.250 95.250 732.750 96.150 ;
        RECT 733.950 94.950 736.050 97.050 ;
        RECT 737.400 94.050 738.450 97.950 ;
        RECT 658.950 91.950 661.050 94.050 ;
        RECT 664.950 92.850 666.750 93.750 ;
        RECT 667.950 91.950 670.050 94.050 ;
        RECT 673.950 91.950 676.050 94.050 ;
        RECT 685.950 91.950 688.050 94.050 ;
        RECT 689.250 92.850 690.750 93.750 ;
        RECT 691.950 91.950 694.050 94.050 ;
        RECT 695.250 92.850 697.050 93.750 ;
        RECT 697.950 91.950 700.050 94.050 ;
        RECT 706.950 91.950 709.050 94.050 ;
        RECT 710.250 92.850 711.750 93.750 ;
        RECT 712.950 91.950 715.050 94.050 ;
        RECT 716.250 92.850 718.050 93.750 ;
        RECT 718.950 91.950 721.050 94.050 ;
        RECT 724.950 91.950 727.050 94.050 ;
        RECT 727.950 92.850 729.750 93.750 ;
        RECT 730.950 91.950 733.050 94.050 ;
        RECT 734.250 92.850 735.750 93.750 ;
        RECT 736.950 91.950 739.050 94.050 ;
        RECT 674.400 70.050 675.450 91.950 ;
        RECT 685.950 89.850 688.050 90.750 ;
        RECT 706.950 89.850 709.050 90.750 ;
        RECT 721.950 88.950 724.050 91.050 ;
        RECT 718.950 73.950 721.050 76.050 ;
        RECT 673.950 67.950 676.050 70.050 ;
        RECT 679.950 67.950 682.050 70.050 ;
        RECT 676.950 58.950 679.050 61.050 ;
        RECT 677.400 58.050 678.450 58.950 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 670.950 57.450 673.050 58.050 ;
        RECT 668.400 56.400 673.050 57.450 ;
        RECT 655.950 52.950 658.050 55.050 ;
        RECT 655.950 50.850 658.050 51.750 ;
        RECT 658.950 50.250 661.050 51.150 ;
        RECT 646.950 46.950 649.050 49.050 ;
        RECT 658.950 48.450 661.050 49.050 ;
        RECT 662.400 48.450 663.450 55.950 ;
        RECT 658.950 47.400 663.450 48.450 ;
        RECT 658.950 46.950 661.050 47.400 ;
        RECT 644.400 44.400 648.450 45.450 ;
        RECT 625.950 40.950 628.050 43.050 ;
        RECT 619.950 28.950 622.050 31.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 614.400 19.050 615.450 22.950 ;
        RECT 616.950 20.850 619.050 21.750 ;
        RECT 604.950 17.400 609.450 18.450 ;
        RECT 604.950 16.950 607.050 17.400 ;
        RECT 613.950 16.950 616.050 19.050 ;
        RECT 620.400 18.450 621.450 28.950 ;
        RECT 626.400 25.050 627.450 40.950 ;
        RECT 647.400 28.050 648.450 44.400 ;
        RECT 661.950 43.950 664.050 46.050 ;
        RECT 649.950 28.950 652.050 31.050 ;
        RECT 646.950 25.950 649.050 28.050 ;
        RECT 650.400 25.050 651.450 28.950 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 647.250 23.850 648.750 24.750 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 662.400 22.050 663.450 43.950 ;
        RECT 668.400 40.050 669.450 56.400 ;
        RECT 670.950 55.950 673.050 56.400 ;
        RECT 674.250 56.250 675.750 57.150 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 680.400 55.050 681.450 67.950 ;
        RECT 688.950 56.250 691.050 57.150 ;
        RECT 670.950 53.850 672.750 54.750 ;
        RECT 673.950 52.950 676.050 55.050 ;
        RECT 677.250 53.850 679.050 54.750 ;
        RECT 679.950 52.950 682.050 55.050 ;
        RECT 685.950 52.950 688.050 55.050 ;
        RECT 688.950 52.950 691.050 55.050 ;
        RECT 692.250 53.250 693.750 54.150 ;
        RECT 694.950 52.950 697.050 55.050 ;
        RECT 698.250 53.250 700.050 54.150 ;
        RECT 700.950 52.950 703.050 55.050 ;
        RECT 709.950 52.950 712.050 55.050 ;
        RECT 686.400 43.050 687.450 52.950 ;
        RECT 689.400 52.050 690.450 52.950 ;
        RECT 688.950 49.950 691.050 52.050 ;
        RECT 691.950 49.950 694.050 52.050 ;
        RECT 695.250 50.850 696.750 51.750 ;
        RECT 697.950 51.450 700.050 52.050 ;
        RECT 701.400 51.450 702.450 52.950 ;
        RECT 697.950 50.400 702.450 51.450 ;
        RECT 709.950 50.850 712.050 51.750 ;
        RECT 697.950 49.950 700.050 50.400 ;
        RECT 712.950 50.250 715.050 51.150 ;
        RECT 692.400 49.050 693.450 49.950 ;
        RECT 691.950 46.950 694.050 49.050 ;
        RECT 712.950 46.950 715.050 49.050 ;
        RECT 685.950 40.950 688.050 43.050 ;
        RECT 667.950 37.950 670.050 40.050 ;
        RECT 694.950 34.950 697.050 37.050 ;
        RECT 688.950 31.950 691.050 34.050 ;
        RECT 685.950 24.450 688.050 25.050 ;
        RECT 677.400 23.400 688.050 24.450 ;
        RECT 622.950 20.250 625.050 21.150 ;
        RECT 625.950 20.850 628.050 21.750 ;
        RECT 643.950 20.850 646.050 21.750 ;
        RECT 649.950 20.850 652.050 21.750 ;
        RECT 658.950 20.250 660.750 21.150 ;
        RECT 661.950 19.950 664.050 22.050 ;
        RECT 665.250 20.250 667.050 21.150 ;
        RECT 667.950 19.950 670.050 22.050 ;
        RECT 622.950 18.450 625.050 19.050 ;
        RECT 620.400 17.400 625.050 18.450 ;
        RECT 622.950 16.950 625.050 17.400 ;
        RECT 658.950 16.950 661.050 19.050 ;
        RECT 662.250 17.850 663.750 18.750 ;
        RECT 664.950 18.450 667.050 19.050 ;
        RECT 668.400 18.450 669.450 19.950 ;
        RECT 677.400 19.050 678.450 23.400 ;
        RECT 685.950 22.950 688.050 23.400 ;
        RECT 689.400 22.050 690.450 31.950 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 692.400 22.050 693.450 22.950 ;
        RECT 679.950 20.250 681.750 21.150 ;
        RECT 682.950 19.950 685.050 22.050 ;
        RECT 688.950 19.950 691.050 22.050 ;
        RECT 691.950 19.950 694.050 22.050 ;
        RECT 664.950 17.400 669.450 18.450 ;
        RECT 664.950 16.950 667.050 17.400 ;
        RECT 676.950 16.950 679.050 19.050 ;
        RECT 679.950 16.950 682.050 19.050 ;
        RECT 683.250 17.850 684.750 18.750 ;
        RECT 685.950 16.950 688.050 19.050 ;
        RECT 689.250 17.850 691.050 18.750 ;
        RECT 455.400 16.050 456.450 16.950 ;
        RECT 473.400 16.050 474.450 16.950 ;
        RECT 545.400 16.050 546.450 16.950 ;
        RECT 680.400 16.050 681.450 16.950 ;
        RECT 695.400 16.050 696.450 34.950 ;
        RECT 703.950 31.950 706.050 34.050 ;
        RECT 704.400 22.050 705.450 31.950 ;
        RECT 712.950 25.950 715.050 28.050 ;
        RECT 713.400 25.050 714.450 25.950 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 710.250 23.250 711.750 24.150 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 703.950 19.950 706.050 22.050 ;
        RECT 707.250 20.850 708.750 21.750 ;
        RECT 709.950 19.950 712.050 22.050 ;
        RECT 713.250 20.850 715.050 21.750 ;
        RECT 703.950 17.850 706.050 18.750 ;
        RECT 710.400 18.450 711.450 19.950 ;
        RECT 719.400 18.450 720.450 73.950 ;
        RECT 722.400 58.050 723.450 88.950 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 724.950 56.250 727.050 57.150 ;
        RECT 722.400 54.450 723.450 55.950 ;
        RECT 731.400 55.050 732.450 91.950 ;
        RECT 736.950 89.850 739.050 90.750 ;
        RECT 743.400 55.050 744.450 97.950 ;
        RECT 748.950 95.850 751.050 96.750 ;
        RECT 751.950 95.250 754.050 96.150 ;
        RECT 751.950 91.950 754.050 94.050 ;
        RECT 752.400 58.050 753.450 91.950 ;
        RECT 764.400 73.050 765.450 97.950 ;
        RECT 767.400 97.050 768.450 115.950 ;
        RECT 770.400 100.050 771.450 133.950 ;
        RECT 773.400 103.050 774.450 226.950 ;
        RECT 775.950 214.950 778.050 217.050 ;
        RECT 772.950 100.950 775.050 103.050 ;
        RECT 769.950 97.950 772.050 100.050 ;
        RECT 772.950 97.950 775.050 100.050 ;
        RECT 773.400 97.050 774.450 97.950 ;
        RECT 766.950 94.950 769.050 97.050 ;
        RECT 769.950 94.950 772.050 97.050 ;
        RECT 772.950 94.950 775.050 97.050 ;
        RECT 766.950 92.850 769.050 93.750 ;
        RECT 763.950 70.950 766.050 73.050 ;
        RECT 770.400 64.050 771.450 94.950 ;
        RECT 772.950 92.850 775.050 93.750 ;
        RECT 772.950 64.950 775.050 67.050 ;
        RECT 769.950 61.950 772.050 64.050 ;
        RECT 760.950 58.950 763.050 61.050 ;
        RECT 751.950 55.950 754.050 58.050 ;
        RECT 724.950 54.450 727.050 55.050 ;
        RECT 722.400 53.400 727.050 54.450 ;
        RECT 722.400 49.050 723.450 53.400 ;
        RECT 724.950 52.950 727.050 53.400 ;
        RECT 728.250 53.250 729.750 54.150 ;
        RECT 730.950 52.950 733.050 55.050 ;
        RECT 734.250 53.250 736.050 54.150 ;
        RECT 742.950 52.950 745.050 55.050 ;
        RECT 751.950 54.450 754.050 55.050 ;
        RECT 746.250 53.250 748.050 54.150 ;
        RECT 749.400 53.400 754.050 54.450 ;
        RECT 727.950 49.950 730.050 52.050 ;
        RECT 731.250 50.850 732.750 51.750 ;
        RECT 733.950 49.950 736.050 52.050 ;
        RECT 742.950 50.850 744.750 51.750 ;
        RECT 745.950 49.950 748.050 52.050 ;
        RECT 721.950 46.950 724.050 49.050 ;
        RECT 728.400 37.050 729.450 49.950 ;
        RECT 746.400 49.050 747.450 49.950 ;
        RECT 745.950 46.950 748.050 49.050 ;
        RECT 727.950 34.950 730.050 37.050 ;
        RECT 742.950 31.950 745.050 34.050 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 721.950 20.250 723.750 21.150 ;
        RECT 724.950 19.950 727.050 22.050 ;
        RECT 728.250 20.250 730.050 21.150 ;
        RECT 721.950 18.450 724.050 19.050 ;
        RECT 710.400 17.400 724.050 18.450 ;
        RECT 725.250 17.850 726.750 18.750 ;
        RECT 727.950 18.450 730.050 19.050 ;
        RECT 731.400 18.450 732.450 22.950 ;
        RECT 743.400 22.050 744.450 31.950 ;
        RECT 749.400 31.050 750.450 53.400 ;
        RECT 751.950 52.950 754.050 53.400 ;
        RECT 755.250 53.250 757.050 54.150 ;
        RECT 751.950 50.850 753.750 51.750 ;
        RECT 754.950 49.950 757.050 52.050 ;
        RECT 748.950 28.950 751.050 31.050 ;
        RECT 761.400 28.050 762.450 58.950 ;
        RECT 773.400 58.050 774.450 64.950 ;
        RECT 776.400 58.050 777.450 214.950 ;
        RECT 779.400 60.450 780.450 229.950 ;
        RECT 782.400 229.050 783.450 232.950 ;
        RECT 781.950 226.950 784.050 229.050 ;
        RECT 785.400 217.050 786.450 256.950 ;
        RECT 788.400 250.050 789.450 277.950 ;
        RECT 794.400 271.050 795.450 283.950 ;
        RECT 800.400 280.050 801.450 337.950 ;
        RECT 803.400 331.050 804.450 403.950 ;
        RECT 805.950 403.500 808.050 405.600 ;
        RECT 805.950 383.250 808.050 384.150 ;
        RECT 805.950 346.950 808.050 349.050 ;
        RECT 802.950 328.950 805.050 331.050 ;
        RECT 806.400 316.050 807.450 346.950 ;
        RECT 809.400 340.050 810.450 563.400 ;
        RECT 817.950 561.600 820.050 563.700 ;
        RECT 814.950 556.950 817.050 559.050 ;
        RECT 815.400 556.050 816.450 556.950 ;
        RECT 814.950 553.950 817.050 556.050 ;
        RECT 814.950 551.850 817.050 552.750 ;
        RECT 818.550 549.600 819.750 561.600 ;
        RECT 817.950 547.500 820.050 549.600 ;
        RECT 811.950 533.400 814.050 535.500 ;
        RECT 812.250 521.400 813.450 533.400 ;
        RECT 814.950 530.250 817.050 531.150 ;
        RECT 814.950 526.950 817.050 529.050 ;
        RECT 811.950 519.300 814.050 521.400 ;
        RECT 812.250 515.700 813.450 519.300 ;
        RECT 815.400 517.050 816.450 526.950 ;
        RECT 811.950 513.600 814.050 515.700 ;
        RECT 814.950 514.950 817.050 517.050 ;
        RECT 815.400 510.450 816.450 514.950 ;
        RECT 812.400 509.400 816.450 510.450 ;
        RECT 812.400 364.050 813.450 509.400 ;
        RECT 821.400 508.050 822.450 616.950 ;
        RECT 823.950 610.950 826.050 613.050 ;
        RECT 824.400 598.050 825.450 610.950 ;
        RECT 827.400 610.050 828.450 625.950 ;
        RECT 829.950 622.950 832.050 625.050 ;
        RECT 826.950 607.950 829.050 610.050 ;
        RECT 826.950 604.950 829.050 607.050 ;
        RECT 827.400 601.050 828.450 604.950 ;
        RECT 826.950 598.950 829.050 601.050 ;
        RECT 823.950 595.950 826.050 598.050 ;
        RECT 826.950 596.850 829.050 597.750 ;
        RECT 826.950 557.250 829.050 558.150 ;
        RECT 826.950 553.950 829.050 556.050 ;
        RECT 830.400 529.050 831.450 622.950 ;
        RECT 839.400 612.450 840.450 676.950 ;
        RECT 842.400 646.050 843.450 709.950 ;
        RECT 854.400 709.050 855.450 769.950 ;
        RECT 862.950 766.950 865.050 769.050 ;
        RECT 863.400 766.050 864.450 766.950 ;
        RECT 862.950 763.950 865.050 766.050 ;
        RECT 862.950 745.950 865.050 748.050 ;
        RECT 863.400 742.050 864.450 745.950 ;
        RECT 859.950 740.250 861.750 741.150 ;
        RECT 862.950 739.950 865.050 742.050 ;
        RECT 866.250 740.250 868.050 741.150 ;
        RECT 863.250 737.850 864.750 738.750 ;
        RECT 847.950 706.950 850.050 709.050 ;
        RECT 850.950 706.950 853.050 709.050 ;
        RECT 853.950 706.950 856.050 709.050 ;
        RECT 856.950 707.250 859.050 708.150 ;
        RECT 862.950 706.950 865.050 709.050 ;
        RECT 848.400 670.050 849.450 706.950 ;
        RECT 851.400 706.050 852.450 706.950 ;
        RECT 850.950 703.950 853.050 706.050 ;
        RECT 854.250 704.250 855.750 705.150 ;
        RECT 856.950 703.950 859.050 706.050 ;
        RECT 860.250 704.250 862.050 705.150 ;
        RECT 850.950 701.850 852.750 702.750 ;
        RECT 853.950 700.950 856.050 703.050 ;
        RECT 854.400 700.050 855.450 700.950 ;
        RECT 853.950 697.950 856.050 700.050 ;
        RECT 857.400 694.050 858.450 703.950 ;
        RECT 859.950 702.450 862.050 703.050 ;
        RECT 863.400 702.450 864.450 706.950 ;
        RECT 859.950 701.400 864.450 702.450 ;
        RECT 859.950 700.950 862.050 701.400 ;
        RECT 856.950 691.950 859.050 694.050 ;
        RECT 850.950 670.950 853.050 673.050 ;
        RECT 854.250 671.250 855.750 672.150 ;
        RECT 847.950 667.950 850.050 670.050 ;
        RECT 851.250 668.850 852.750 669.750 ;
        RECT 853.950 667.950 856.050 670.050 ;
        RECT 857.250 668.850 859.050 669.750 ;
        RECT 847.950 665.850 850.050 666.750 ;
        RECT 850.950 664.950 853.050 667.050 ;
        RECT 854.400 666.450 855.450 667.950 ;
        RECT 854.400 665.400 858.450 666.450 ;
        RECT 841.950 643.950 844.050 646.050 ;
        RECT 841.950 638.400 844.050 640.500 ;
        RECT 842.400 621.600 843.600 638.400 ;
        RECT 851.400 634.050 852.450 664.950 ;
        RECT 850.950 631.950 853.050 634.050 ;
        RECT 847.950 629.250 850.050 630.150 ;
        RECT 853.950 629.250 856.050 630.150 ;
        RECT 847.950 625.950 850.050 628.050 ;
        RECT 853.950 625.950 856.050 628.050 ;
        RECT 847.950 622.950 850.050 625.050 ;
        RECT 841.950 619.500 844.050 621.600 ;
        RECT 839.400 611.400 843.450 612.450 ;
        RECT 838.950 605.400 841.050 607.500 ;
        RECT 832.950 598.950 835.050 601.050 ;
        RECT 832.950 596.850 835.050 597.750 ;
        RECT 839.400 588.600 840.600 605.400 ;
        RECT 838.950 586.500 841.050 588.600 ;
        RECT 838.950 566.400 841.050 568.500 ;
        RECT 842.400 568.050 843.450 611.400 ;
        RECT 848.400 592.050 849.450 622.950 ;
        RECT 854.400 607.050 855.450 625.950 ;
        RECT 857.400 622.050 858.450 665.400 ;
        RECT 862.950 639.300 865.050 641.400 ;
        RECT 863.250 635.700 864.450 639.300 ;
        RECT 862.950 633.600 865.050 635.700 ;
        RECT 856.950 619.950 859.050 622.050 ;
        RECT 863.250 621.600 864.450 633.600 ;
        RECT 865.950 625.950 868.050 628.050 ;
        RECT 865.950 623.850 868.050 624.750 ;
        RECT 862.950 619.500 865.050 621.600 ;
        RECT 865.950 619.950 868.050 622.050 ;
        RECT 853.950 604.950 856.050 607.050 ;
        RECT 857.250 599.250 858.750 600.150 ;
        RECT 859.950 598.950 862.050 601.050 ;
        RECT 853.950 596.850 855.750 597.750 ;
        RECT 856.950 595.950 859.050 598.050 ;
        RECT 860.250 596.850 861.750 597.750 ;
        RECT 862.950 595.950 865.050 598.050 ;
        RECT 857.400 595.050 858.450 595.950 ;
        RECT 856.950 592.950 859.050 595.050 ;
        RECT 859.950 592.950 862.050 595.050 ;
        RECT 862.950 593.850 865.050 594.750 ;
        RECT 847.950 589.950 850.050 592.050 ;
        RECT 832.950 557.250 835.050 558.150 ;
        RECT 832.950 553.950 835.050 556.050 ;
        RECT 833.400 550.050 834.450 553.950 ;
        RECT 832.950 547.950 835.050 550.050 ;
        RECT 839.400 549.600 840.600 566.400 ;
        RECT 841.950 565.950 844.050 568.050 ;
        RECT 853.950 565.950 856.050 568.050 ;
        RECT 838.950 547.500 841.050 549.600 ;
        RECT 850.950 547.950 853.050 550.050 ;
        RECT 851.400 529.050 852.450 547.950 ;
        RECT 829.950 526.950 832.050 529.050 ;
        RECT 848.250 527.250 849.750 528.150 ;
        RECT 850.950 526.950 853.050 529.050 ;
        RECT 854.400 526.050 855.450 565.950 ;
        RECT 860.400 565.050 861.450 592.950 ;
        RECT 859.950 562.950 862.050 565.050 ;
        RECT 860.250 560.250 861.750 561.150 ;
        RECT 856.950 557.850 858.750 558.750 ;
        RECT 859.950 556.950 862.050 559.050 ;
        RECT 863.250 557.850 865.050 558.750 ;
        RECT 856.950 553.950 859.050 556.050 ;
        RECT 826.950 523.950 829.050 526.050 ;
        RECT 829.950 524.250 831.750 525.150 ;
        RECT 832.950 523.950 835.050 526.050 ;
        RECT 836.250 524.250 838.050 525.150 ;
        RECT 844.950 524.850 846.750 525.750 ;
        RECT 847.950 523.950 850.050 526.050 ;
        RECT 851.250 524.850 852.750 525.750 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 814.950 505.950 817.050 508.050 ;
        RECT 820.950 505.950 823.050 508.050 ;
        RECT 815.400 427.050 816.450 505.950 ;
        RECT 827.400 493.050 828.450 523.950 ;
        RECT 833.250 521.850 834.750 522.750 ;
        RECT 853.950 521.850 856.050 522.750 ;
        RECT 857.400 520.050 858.450 553.950 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 838.950 517.950 841.050 520.050 ;
        RECT 856.950 517.950 859.050 520.050 ;
        RECT 826.950 490.950 829.050 493.050 ;
        RECT 832.950 490.950 835.050 493.050 ;
        RECT 829.950 488.250 832.050 489.150 ;
        RECT 820.950 485.250 822.750 486.150 ;
        RECT 823.950 484.950 826.050 487.050 ;
        RECT 829.950 486.450 832.050 487.050 ;
        RECT 833.400 486.450 834.450 490.950 ;
        RECT 827.250 485.250 828.750 486.150 ;
        RECT 829.950 485.400 834.450 486.450 ;
        RECT 829.950 484.950 832.050 485.400 ;
        RECT 824.250 482.850 825.750 483.750 ;
        RECT 826.950 481.950 829.050 484.050 ;
        RECT 827.400 457.050 828.450 481.950 ;
        RECT 835.950 461.400 838.050 463.500 ;
        RECT 829.950 457.950 832.050 460.050 ;
        RECT 832.950 458.250 835.050 459.150 ;
        RECT 823.950 455.250 826.050 456.150 ;
        RECT 826.950 454.950 829.050 457.050 ;
        RECT 830.400 456.450 831.450 457.950 ;
        RECT 832.950 456.450 835.050 457.050 ;
        RECT 830.400 455.400 835.050 456.450 ;
        RECT 832.950 454.950 835.050 455.400 ;
        RECT 814.950 424.950 817.050 427.050 ;
        RECT 823.950 424.950 826.050 427.050 ;
        RECT 814.950 413.250 817.050 414.150 ;
        RECT 820.950 413.250 823.050 414.150 ;
        RECT 814.950 409.950 817.050 412.050 ;
        RECT 820.950 409.950 823.050 412.050 ;
        RECT 815.400 403.050 816.450 409.950 ;
        RECT 824.400 408.450 825.450 424.950 ;
        RECT 826.950 422.400 829.050 424.500 ;
        RECT 821.400 407.400 825.450 408.450 ;
        RECT 814.950 400.950 817.050 403.050 ;
        RECT 811.950 361.950 814.050 364.050 ;
        RECT 811.950 355.950 814.050 358.050 ;
        RECT 812.400 346.050 813.450 355.950 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 815.250 344.250 816.750 345.150 ;
        RECT 817.950 343.950 820.050 346.050 ;
        RECT 811.950 341.850 813.750 342.750 ;
        RECT 814.950 340.950 817.050 343.050 ;
        RECT 818.250 341.850 820.050 342.750 ;
        RECT 808.950 337.950 811.050 340.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 805.950 313.950 808.050 316.050 ;
        RECT 802.950 310.950 805.050 313.050 ;
        RECT 803.400 306.450 804.450 310.950 ;
        RECT 809.400 310.050 810.450 334.950 ;
        RECT 815.400 319.050 816.450 340.950 ;
        RECT 817.950 337.950 820.050 340.050 ;
        RECT 814.950 316.950 817.050 319.050 ;
        RECT 814.950 313.950 817.050 316.050 ;
        RECT 805.950 308.250 807.750 309.150 ;
        RECT 808.950 307.950 811.050 310.050 ;
        RECT 812.250 308.250 814.050 309.150 ;
        RECT 805.950 306.450 808.050 307.050 ;
        RECT 803.400 305.400 808.050 306.450 ;
        RECT 809.250 305.850 810.750 306.750 ;
        RECT 805.950 304.950 808.050 305.400 ;
        RECT 811.950 304.950 814.050 307.050 ;
        RECT 799.950 277.950 802.050 280.050 ;
        RECT 802.950 277.950 805.050 280.050 ;
        RECT 803.400 277.050 804.450 277.950 ;
        RECT 799.950 274.950 802.050 277.050 ;
        RECT 802.950 274.950 805.050 277.050 ;
        RECT 790.950 269.250 793.050 270.150 ;
        RECT 793.950 268.950 796.050 271.050 ;
        RECT 796.950 269.250 799.050 270.150 ;
        RECT 790.950 265.950 793.050 268.050 ;
        RECT 794.250 266.250 795.750 267.150 ;
        RECT 796.950 265.950 799.050 268.050 ;
        RECT 797.400 265.050 798.450 265.950 ;
        RECT 793.950 262.950 796.050 265.050 ;
        RECT 796.950 262.950 799.050 265.050 ;
        RECT 794.400 261.450 795.450 262.950 ;
        RECT 796.950 261.450 799.050 262.050 ;
        RECT 794.400 260.400 799.050 261.450 ;
        RECT 796.950 259.950 799.050 260.400 ;
        RECT 800.400 253.050 801.450 274.950 ;
        RECT 806.400 273.450 807.450 304.950 ;
        RECT 812.400 304.050 813.450 304.950 ;
        RECT 811.950 301.950 814.050 304.050 ;
        RECT 808.950 277.950 811.050 280.050 ;
        RECT 803.400 272.400 807.450 273.450 ;
        RECT 803.400 265.050 804.450 272.400 ;
        RECT 809.400 271.050 810.450 277.950 ;
        RECT 815.400 277.050 816.450 313.950 ;
        RECT 814.950 274.950 817.050 277.050 ;
        RECT 814.950 272.250 817.050 273.150 ;
        RECT 805.950 269.250 807.750 270.150 ;
        RECT 808.950 268.950 811.050 271.050 ;
        RECT 812.250 269.250 813.750 270.150 ;
        RECT 814.950 268.950 817.050 271.050 ;
        RECT 805.950 265.950 808.050 268.050 ;
        RECT 809.250 266.850 810.750 267.750 ;
        RECT 811.950 265.950 814.050 268.050 ;
        RECT 802.950 262.950 805.050 265.050 ;
        RECT 806.400 259.050 807.450 265.950 ;
        RECT 811.950 262.950 814.050 265.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 790.950 250.950 793.050 253.050 ;
        RECT 799.950 250.950 802.050 253.050 ;
        RECT 787.950 247.950 790.050 250.050 ;
        RECT 787.950 244.950 790.050 247.050 ;
        RECT 788.400 232.050 789.450 244.950 ;
        RECT 791.400 244.050 792.450 250.950 ;
        RECT 793.950 247.950 796.050 250.050 ;
        RECT 790.950 241.950 793.050 244.050 ;
        RECT 794.400 241.050 795.450 247.950 ;
        RECT 805.950 244.950 808.050 247.050 ;
        RECT 806.400 241.050 807.450 244.950 ;
        RECT 790.950 238.950 793.050 241.050 ;
        RECT 793.950 238.950 796.050 241.050 ;
        RECT 797.250 239.250 798.750 240.150 ;
        RECT 799.950 238.950 802.050 241.050 ;
        RECT 803.250 239.250 804.750 240.150 ;
        RECT 805.950 238.950 808.050 241.050 ;
        RECT 787.950 229.950 790.050 232.050 ;
        RECT 787.950 226.950 790.050 229.050 ;
        RECT 784.950 214.950 787.050 217.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 781.950 205.950 784.050 208.050 ;
        RECT 782.400 193.050 783.450 205.950 ;
        RECT 785.400 202.050 786.450 211.950 ;
        RECT 788.400 205.050 789.450 226.950 ;
        RECT 787.950 202.950 790.050 205.050 ;
        RECT 791.400 204.450 792.450 238.950 ;
        RECT 793.950 236.850 795.750 237.750 ;
        RECT 796.950 235.950 799.050 238.050 ;
        RECT 800.250 236.850 801.750 237.750 ;
        RECT 802.950 235.950 805.050 238.050 ;
        RECT 806.250 236.850 808.050 237.750 ;
        RECT 799.950 232.950 802.050 235.050 ;
        RECT 796.950 226.950 799.050 229.050 ;
        RECT 791.400 203.400 795.450 204.450 ;
        RECT 784.950 199.950 787.050 202.050 ;
        RECT 788.250 200.250 789.750 201.150 ;
        RECT 790.950 199.950 793.050 202.050 ;
        RECT 784.950 197.850 786.750 198.750 ;
        RECT 787.950 196.950 790.050 199.050 ;
        RECT 791.250 197.850 793.050 198.750 ;
        RECT 781.950 190.950 784.050 193.050 ;
        RECT 794.400 190.050 795.450 203.400 ;
        RECT 797.400 202.050 798.450 226.950 ;
        RECT 800.400 220.050 801.450 232.950 ;
        RECT 809.400 232.050 810.450 256.950 ;
        RECT 808.950 229.950 811.050 232.050 ;
        RECT 812.400 226.050 813.450 262.950 ;
        RECT 815.400 262.050 816.450 268.950 ;
        RECT 814.950 259.950 817.050 262.050 ;
        RECT 818.400 259.050 819.450 337.950 ;
        RECT 821.400 307.050 822.450 407.400 ;
        RECT 827.400 405.600 828.600 422.400 ;
        RECT 829.950 409.950 832.050 412.050 ;
        RECT 830.400 406.050 831.450 409.950 ;
        RECT 826.950 403.500 829.050 405.600 ;
        RECT 829.950 403.950 832.050 406.050 ;
        RECT 823.950 383.250 826.050 384.150 ;
        RECT 823.950 355.950 826.050 358.050 ;
        RECT 824.400 316.050 825.450 355.950 ;
        RECT 833.400 349.050 834.450 454.950 ;
        RECT 836.550 449.400 837.750 461.400 ;
        RECT 835.950 447.300 838.050 449.400 ;
        RECT 836.550 443.700 837.750 447.300 ;
        RECT 835.950 441.600 838.050 443.700 ;
        RECT 835.950 436.950 838.050 439.050 ;
        RECT 836.400 378.450 837.450 436.950 ;
        RECT 839.400 382.050 840.450 517.950 ;
        RECT 851.250 488.250 852.750 489.150 ;
        RECT 847.950 485.850 849.750 486.750 ;
        RECT 850.950 484.950 853.050 487.050 ;
        RECT 854.250 485.850 856.050 486.750 ;
        RECT 851.400 459.450 852.450 484.950 ;
        RECT 856.950 461.400 859.050 463.500 ;
        RECT 851.400 458.400 855.450 459.450 ;
        RECT 844.950 456.450 847.050 457.050 ;
        RECT 842.400 455.400 847.050 456.450 ;
        RECT 842.400 454.050 843.450 455.400 ;
        RECT 844.950 454.950 847.050 455.400 ;
        RECT 850.950 454.950 853.050 457.050 ;
        RECT 841.950 451.950 844.050 454.050 ;
        RECT 844.950 452.850 847.050 453.750 ;
        RECT 850.950 452.850 853.050 453.750 ;
        RECT 850.950 416.250 853.050 417.150 ;
        RECT 841.950 413.250 843.750 414.150 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 850.950 414.450 853.050 415.050 ;
        RECT 854.400 414.450 855.450 458.400 ;
        RECT 857.400 444.600 858.600 461.400 ;
        RECT 856.950 442.500 859.050 444.600 ;
        RECT 860.400 439.050 861.450 523.950 ;
        RECT 859.950 436.950 862.050 439.050 ;
        RECT 848.250 413.250 849.750 414.150 ;
        RECT 850.950 413.400 855.450 414.450 ;
        RECT 850.950 412.950 853.050 413.400 ;
        RECT 845.250 410.850 846.750 411.750 ;
        RECT 847.950 409.950 850.050 412.050 ;
        RECT 850.950 409.950 853.050 412.050 ;
        RECT 848.400 406.050 849.450 409.950 ;
        RECT 847.950 403.950 850.050 406.050 ;
        RECT 841.950 400.950 844.050 403.050 ;
        RECT 838.950 379.950 841.050 382.050 ;
        RECT 842.400 381.450 843.450 400.950 ;
        RECT 844.950 383.250 847.050 384.150 ;
        RECT 844.950 381.450 847.050 382.050 ;
        RECT 842.400 380.400 847.050 381.450 ;
        RECT 844.950 379.950 847.050 380.400 ;
        RECT 836.400 377.400 840.450 378.450 ;
        RECT 832.950 346.950 835.050 349.050 ;
        RECT 826.950 343.950 829.050 346.050 ;
        RECT 827.400 337.050 828.450 343.950 ;
        RECT 832.950 340.950 835.050 343.050 ;
        RECT 835.950 340.950 838.050 343.050 ;
        RECT 829.950 338.250 832.050 339.150 ;
        RECT 832.950 338.850 835.050 339.750 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 830.400 325.050 831.450 334.950 ;
        RECT 829.950 322.950 832.050 325.050 ;
        RECT 830.400 322.050 831.450 322.950 ;
        RECT 829.950 319.950 832.050 322.050 ;
        RECT 823.950 313.950 826.050 316.050 ;
        RECT 823.950 311.850 826.050 312.750 ;
        RECT 826.950 311.250 829.050 312.150 ;
        RECT 826.950 309.450 829.050 310.050 ;
        RECT 824.400 308.400 829.050 309.450 ;
        RECT 820.950 304.950 823.050 307.050 ;
        RECT 820.950 301.950 823.050 304.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 815.400 235.050 816.450 253.950 ;
        RECT 821.400 250.050 822.450 301.950 ;
        RECT 824.400 283.050 825.450 308.400 ;
        RECT 826.950 307.950 829.050 308.400 ;
        RECT 826.950 304.950 829.050 307.050 ;
        RECT 823.950 280.950 826.050 283.050 ;
        RECT 824.400 271.050 825.450 280.950 ;
        RECT 823.950 268.950 826.050 271.050 ;
        RECT 820.950 247.950 823.050 250.050 ;
        RECT 820.950 238.950 823.050 241.050 ;
        RECT 821.400 238.050 822.450 238.950 ;
        RECT 817.950 236.250 819.750 237.150 ;
        RECT 820.950 235.950 823.050 238.050 ;
        RECT 824.250 236.250 826.050 237.150 ;
        RECT 814.950 232.950 817.050 235.050 ;
        RECT 817.950 232.950 820.050 235.050 ;
        RECT 821.250 233.850 822.750 234.750 ;
        RECT 823.950 232.950 826.050 235.050 ;
        RECT 817.950 229.950 820.050 232.050 ;
        RECT 823.950 229.950 826.050 232.050 ;
        RECT 811.950 223.950 814.050 226.050 ;
        RECT 814.950 220.950 817.050 223.050 ;
        RECT 799.950 217.950 802.050 220.050 ;
        RECT 796.950 199.950 799.050 202.050 ;
        RECT 802.950 200.250 805.050 201.150 ;
        RECT 808.950 199.950 811.050 202.050 ;
        RECT 793.950 187.950 796.050 190.050 ;
        RECT 797.400 172.050 798.450 199.950 ;
        RECT 809.400 199.050 810.450 199.950 ;
        RECT 802.950 196.950 805.050 199.050 ;
        RECT 806.250 197.250 807.750 198.150 ;
        RECT 808.950 196.950 811.050 199.050 ;
        RECT 812.250 197.250 814.050 198.150 ;
        RECT 805.950 193.950 808.050 196.050 ;
        RECT 809.250 194.850 810.750 195.750 ;
        RECT 811.950 193.950 814.050 196.050 ;
        RECT 806.400 175.050 807.450 193.950 ;
        RECT 812.400 190.050 813.450 193.950 ;
        RECT 811.950 187.950 814.050 190.050 ;
        RECT 799.950 172.950 802.050 175.050 ;
        RECT 805.950 172.950 808.050 175.050 ;
        RECT 784.950 169.950 787.050 172.050 ;
        RECT 793.950 169.950 796.050 172.050 ;
        RECT 796.950 169.950 799.050 172.050 ;
        RECT 785.400 166.050 786.450 169.950 ;
        RECT 790.950 166.950 793.050 169.050 ;
        RECT 781.950 164.250 783.750 165.150 ;
        RECT 784.950 163.950 787.050 166.050 ;
        RECT 788.250 164.250 790.050 165.150 ;
        RECT 781.950 160.950 784.050 163.050 ;
        RECT 785.250 161.850 786.750 162.750 ;
        RECT 787.950 162.450 790.050 163.050 ;
        RECT 791.400 162.450 792.450 166.950 ;
        RECT 787.950 161.400 792.450 162.450 ;
        RECT 787.950 160.950 790.050 161.400 ;
        RECT 782.400 127.050 783.450 160.950 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 781.950 124.950 784.050 127.050 ;
        RECT 781.950 122.850 784.050 123.750 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 782.400 79.050 783.450 100.950 ;
        RECT 781.950 76.950 784.050 79.050 ;
        RECT 779.400 59.400 783.450 60.450 ;
        RECT 769.950 56.250 772.050 57.150 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 55.950 778.050 58.050 ;
        RECT 769.950 52.950 772.050 55.050 ;
        RECT 773.250 53.250 774.750 54.150 ;
        RECT 775.950 52.950 778.050 55.050 ;
        RECT 779.250 53.250 781.050 54.150 ;
        RECT 770.400 49.050 771.450 52.950 ;
        RECT 772.950 49.950 775.050 52.050 ;
        RECT 776.250 50.850 777.750 51.750 ;
        RECT 778.950 49.950 781.050 52.050 ;
        RECT 769.950 46.950 772.050 49.050 ;
        RECT 778.950 34.950 781.050 37.050 ;
        RECT 763.950 28.950 766.050 31.050 ;
        RECT 764.400 28.050 765.450 28.950 ;
        RECT 754.950 25.950 757.050 28.050 ;
        RECT 760.950 25.950 763.050 28.050 ;
        RECT 763.950 25.950 766.050 28.050 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 749.250 23.250 750.750 24.150 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 755.400 22.050 756.450 25.950 ;
        RECT 761.400 25.050 762.450 25.950 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 764.250 23.850 765.750 24.750 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 742.950 19.950 745.050 22.050 ;
        RECT 746.250 20.850 747.750 21.750 ;
        RECT 748.950 19.950 751.050 22.050 ;
        RECT 752.250 20.850 754.050 21.750 ;
        RECT 754.950 19.950 757.050 22.050 ;
        RECT 760.950 20.850 763.050 21.750 ;
        RECT 766.950 20.850 769.050 21.750 ;
        RECT 721.950 16.950 724.050 17.400 ;
        RECT 727.950 17.400 732.450 18.450 ;
        RECT 742.950 17.850 745.050 18.750 ;
        RECT 779.400 18.450 780.450 34.950 ;
        RECT 782.400 31.050 783.450 59.400 ;
        RECT 785.400 55.050 786.450 130.950 ;
        RECT 787.950 125.250 790.050 126.150 ;
        RECT 787.950 121.950 790.050 124.050 ;
        RECT 791.250 122.250 793.050 123.150 ;
        RECT 787.950 118.950 790.050 121.050 ;
        RECT 790.950 118.950 793.050 121.050 ;
        RECT 788.400 112.050 789.450 118.950 ;
        RECT 787.950 109.950 790.050 112.050 ;
        RECT 791.400 103.050 792.450 118.950 ;
        RECT 794.400 118.050 795.450 169.950 ;
        RECT 800.400 168.450 801.450 172.950 ;
        RECT 811.950 169.950 814.050 172.050 ;
        RECT 812.400 169.050 813.450 169.950 ;
        RECT 797.400 167.400 801.450 168.450 ;
        RECT 797.400 133.050 798.450 167.400 ;
        RECT 805.950 166.950 808.050 169.050 ;
        RECT 809.250 167.250 810.750 168.150 ;
        RECT 811.950 166.950 814.050 169.050 ;
        RECT 802.950 165.450 805.050 166.050 ;
        RECT 800.400 164.400 805.050 165.450 ;
        RECT 806.250 164.850 807.750 165.750 ;
        RECT 796.950 130.950 799.050 133.050 ;
        RECT 796.950 124.950 799.050 127.050 ;
        RECT 797.400 124.050 798.450 124.950 ;
        RECT 796.950 121.950 799.050 124.050 ;
        RECT 793.950 115.950 796.050 118.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 797.400 97.050 798.450 121.950 ;
        RECT 800.400 121.050 801.450 164.400 ;
        RECT 802.950 163.950 805.050 164.400 ;
        RECT 808.950 163.950 811.050 166.050 ;
        RECT 812.250 164.850 814.050 165.750 ;
        RECT 802.950 161.850 805.050 162.750 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 805.950 124.950 808.050 127.050 ;
        RECT 812.400 124.050 813.450 133.950 ;
        RECT 805.950 122.850 808.050 123.750 ;
        RECT 808.950 122.250 811.050 123.150 ;
        RECT 811.950 121.950 814.050 124.050 ;
        RECT 799.950 118.950 802.050 121.050 ;
        RECT 808.950 118.950 811.050 121.050 ;
        RECT 815.400 112.050 816.450 220.950 ;
        RECT 814.950 109.950 817.050 112.050 ;
        RECT 799.950 106.950 802.050 109.050 ;
        RECT 790.950 94.950 793.050 97.050 ;
        RECT 794.250 95.250 795.750 96.150 ;
        RECT 796.950 94.950 799.050 97.050 ;
        RECT 787.950 91.950 790.050 94.050 ;
        RECT 791.250 92.850 792.750 93.750 ;
        RECT 793.950 91.950 796.050 94.050 ;
        RECT 797.250 92.850 799.050 93.750 ;
        RECT 794.400 91.050 795.450 91.950 ;
        RECT 800.400 91.050 801.450 106.950 ;
        RECT 802.950 103.950 805.050 106.050 ;
        RECT 805.950 103.950 808.050 106.050 ;
        RECT 814.950 103.950 817.050 106.050 ;
        RECT 787.950 89.850 790.050 90.750 ;
        RECT 793.950 88.950 796.050 91.050 ;
        RECT 799.950 88.950 802.050 91.050 ;
        RECT 803.400 70.050 804.450 103.950 ;
        RECT 806.400 97.050 807.450 103.950 ;
        RECT 805.950 94.950 808.050 97.050 ;
        RECT 809.250 95.250 810.750 96.150 ;
        RECT 811.950 94.950 814.050 97.050 ;
        RECT 815.400 94.050 816.450 103.950 ;
        RECT 818.400 100.050 819.450 229.950 ;
        RECT 824.400 202.050 825.450 229.950 ;
        RECT 827.400 223.050 828.450 304.950 ;
        RECT 829.950 272.250 832.050 273.150 ;
        RECT 836.400 271.050 837.450 340.950 ;
        RECT 839.400 309.450 840.450 377.400 ;
        RECT 844.950 349.950 847.050 352.050 ;
        RECT 845.400 343.050 846.450 349.950 ;
        RECT 844.950 340.950 847.050 343.050 ;
        RECT 848.250 341.250 850.050 342.150 ;
        RECT 844.950 338.850 846.750 339.750 ;
        RECT 847.950 337.950 850.050 340.050 ;
        RECT 844.950 334.950 847.050 337.050 ;
        RECT 851.400 336.450 852.450 409.950 ;
        RECT 859.950 384.450 862.050 385.050 ;
        RECT 856.950 383.250 858.750 384.150 ;
        RECT 859.950 383.400 864.450 384.450 ;
        RECT 859.950 382.950 862.050 383.400 ;
        RECT 856.950 379.950 859.050 382.050 ;
        RECT 860.250 380.850 862.050 381.750 ;
        RECT 857.400 346.050 858.450 379.950 ;
        RECT 856.950 343.950 859.050 346.050 ;
        RECT 853.950 340.950 856.050 343.050 ;
        RECT 857.250 341.250 859.050 342.150 ;
        RECT 859.950 340.950 862.050 343.050 ;
        RECT 853.950 338.850 855.750 339.750 ;
        RECT 856.950 337.950 859.050 340.050 ;
        RECT 857.400 337.050 858.450 337.950 ;
        RECT 848.400 335.400 852.450 336.450 ;
        RECT 845.400 316.050 846.450 334.950 ;
        RECT 844.950 313.950 847.050 316.050 ;
        RECT 841.950 311.250 844.050 312.150 ;
        RECT 844.950 311.850 847.050 312.750 ;
        RECT 841.950 309.450 844.050 310.050 ;
        RECT 839.400 308.400 844.050 309.450 ;
        RECT 841.950 307.950 844.050 308.400 ;
        RECT 844.950 307.950 847.050 310.050 ;
        RECT 829.950 268.950 832.050 271.050 ;
        RECT 833.250 269.250 834.750 270.150 ;
        RECT 835.950 268.950 838.050 271.050 ;
        RECT 839.250 269.250 841.050 270.150 ;
        RECT 829.950 265.950 832.050 268.050 ;
        RECT 832.950 265.950 835.050 268.050 ;
        RECT 836.250 266.850 837.750 267.750 ;
        RECT 838.950 265.950 841.050 268.050 ;
        RECT 830.400 244.050 831.450 265.950 ;
        RECT 829.950 241.950 832.050 244.050 ;
        RECT 829.950 238.950 832.050 241.050 ;
        RECT 826.950 220.950 829.050 223.050 ;
        RECT 830.400 208.050 831.450 238.950 ;
        RECT 833.400 235.050 834.450 265.950 ;
        RECT 839.400 265.050 840.450 265.950 ;
        RECT 838.950 262.950 841.050 265.050 ;
        RECT 835.950 259.950 838.050 262.050 ;
        RECT 836.400 247.050 837.450 259.950 ;
        RECT 835.950 244.950 838.050 247.050 ;
        RECT 836.400 238.050 837.450 244.950 ;
        RECT 845.400 244.050 846.450 307.950 ;
        RECT 848.400 303.450 849.450 335.400 ;
        RECT 856.950 334.950 859.050 337.050 ;
        RECT 860.400 331.050 861.450 340.950 ;
        RECT 850.950 328.950 853.050 331.050 ;
        RECT 859.950 328.950 862.050 331.050 ;
        RECT 851.400 316.050 852.450 328.950 ;
        RECT 859.950 325.950 862.050 328.050 ;
        RECT 860.400 324.450 861.450 325.950 ;
        RECT 863.400 324.450 864.450 383.400 ;
        RECT 860.400 323.400 864.450 324.450 ;
        RECT 860.400 316.050 861.450 323.400 ;
        RECT 862.950 319.950 865.050 322.050 ;
        RECT 850.950 313.950 853.050 316.050 ;
        RECT 859.950 313.950 862.050 316.050 ;
        RECT 853.950 312.450 856.050 313.050 ;
        RECT 851.400 311.400 856.050 312.450 ;
        RECT 851.400 307.050 852.450 311.400 ;
        RECT 853.950 310.950 856.050 311.400 ;
        RECT 857.250 311.250 858.750 312.150 ;
        RECT 859.950 310.950 862.050 313.050 ;
        RECT 863.400 310.050 864.450 319.950 ;
        RECT 853.950 308.850 855.750 309.750 ;
        RECT 856.950 307.950 859.050 310.050 ;
        RECT 860.250 308.850 861.750 309.750 ;
        RECT 862.950 307.950 865.050 310.050 ;
        RECT 850.950 304.950 853.050 307.050 ;
        RECT 853.950 304.950 856.050 307.050 ;
        RECT 848.400 302.400 852.450 303.450 ;
        RECT 847.950 266.850 850.050 267.750 ;
        RECT 844.950 241.950 847.050 244.050 ;
        RECT 847.950 238.950 850.050 241.050 ;
        RECT 835.950 235.950 838.050 238.050 ;
        RECT 841.950 235.950 844.050 238.050 ;
        RECT 845.250 236.250 847.050 237.150 ;
        RECT 832.950 232.950 835.050 235.050 ;
        RECT 835.950 233.850 837.750 234.750 ;
        RECT 838.950 232.950 841.050 235.050 ;
        RECT 842.250 233.850 843.750 234.750 ;
        RECT 844.950 232.950 847.050 235.050 ;
        RECT 838.950 230.850 841.050 231.750 ;
        RECT 841.950 229.950 844.050 232.050 ;
        RECT 835.950 208.950 838.050 211.050 ;
        RECT 829.950 205.950 832.050 208.050 ;
        RECT 832.950 202.950 835.050 205.050 ;
        RECT 823.950 199.950 826.050 202.050 ;
        RECT 829.950 200.250 832.050 201.150 ;
        RECT 820.950 197.250 822.750 198.150 ;
        RECT 823.950 196.950 826.050 199.050 ;
        RECT 829.950 198.450 832.050 199.050 ;
        RECT 833.400 198.450 834.450 202.950 ;
        RECT 827.250 197.250 828.750 198.150 ;
        RECT 829.950 197.400 834.450 198.450 ;
        RECT 829.950 196.950 832.050 197.400 ;
        RECT 820.950 193.950 823.050 196.050 ;
        RECT 824.250 194.850 825.750 195.750 ;
        RECT 826.950 193.950 829.050 196.050 ;
        RECT 821.400 178.050 822.450 193.950 ;
        RECT 820.950 175.950 823.050 178.050 ;
        RECT 820.950 169.950 823.050 172.050 ;
        RECT 823.950 169.950 826.050 172.050 ;
        RECT 821.400 169.050 822.450 169.950 ;
        RECT 827.400 169.050 828.450 193.950 ;
        RECT 829.950 169.950 832.050 172.050 ;
        RECT 820.950 166.950 823.050 169.050 ;
        RECT 824.250 167.850 825.750 168.750 ;
        RECT 826.950 166.950 829.050 169.050 ;
        RECT 820.950 164.850 823.050 165.750 ;
        RECT 826.950 164.850 829.050 165.750 ;
        RECT 830.400 139.050 831.450 169.950 ;
        RECT 836.400 163.050 837.450 208.950 ;
        RECT 838.950 199.950 841.050 202.050 ;
        RECT 839.400 181.050 840.450 199.950 ;
        RECT 838.950 178.950 841.050 181.050 ;
        RECT 838.950 175.950 841.050 178.050 ;
        RECT 835.950 160.950 838.050 163.050 ;
        RECT 823.950 136.950 826.050 139.050 ;
        RECT 829.950 136.950 832.050 139.050 ;
        RECT 824.400 127.050 825.450 136.950 ;
        RECT 829.950 130.950 832.050 133.050 ;
        RECT 830.400 127.050 831.450 130.950 ;
        RECT 836.400 127.050 837.450 160.950 ;
        RECT 820.950 125.250 822.750 126.150 ;
        RECT 823.950 124.950 826.050 127.050 ;
        RECT 827.250 125.250 828.750 126.150 ;
        RECT 829.950 124.950 832.050 127.050 ;
        RECT 833.250 125.250 835.050 126.150 ;
        RECT 835.950 124.950 838.050 127.050 ;
        RECT 839.400 124.050 840.450 175.950 ;
        RECT 842.400 169.050 843.450 229.950 ;
        RECT 845.400 202.050 846.450 232.950 ;
        RECT 848.400 211.050 849.450 238.950 ;
        RECT 851.400 232.050 852.450 302.400 ;
        RECT 854.400 300.450 855.450 304.950 ;
        RECT 857.400 304.050 858.450 307.950 ;
        RECT 866.400 307.050 867.450 619.950 ;
        RECT 859.950 304.950 862.050 307.050 ;
        RECT 862.950 305.850 865.050 306.750 ;
        RECT 865.950 304.950 868.050 307.050 ;
        RECT 856.950 301.950 859.050 304.050 ;
        RECT 854.400 299.400 858.450 300.450 ;
        RECT 853.950 295.950 856.050 298.050 ;
        RECT 854.400 271.050 855.450 295.950 ;
        RECT 853.950 268.950 856.050 271.050 ;
        RECT 853.950 266.850 856.050 267.750 ;
        RECT 857.400 246.450 858.450 299.400 ;
        RECT 854.400 245.400 858.450 246.450 ;
        RECT 850.950 229.950 853.050 232.050 ;
        RECT 847.950 208.950 850.050 211.050 ;
        RECT 847.950 205.950 850.050 208.050 ;
        RECT 844.950 199.950 847.050 202.050 ;
        RECT 848.400 199.050 849.450 205.950 ;
        RECT 854.400 205.050 855.450 245.400 ;
        RECT 856.950 241.950 859.050 244.050 ;
        RECT 853.950 202.950 856.050 205.050 ;
        RECT 853.950 200.250 856.050 201.150 ;
        RECT 844.950 197.250 846.750 198.150 ;
        RECT 847.950 196.950 850.050 199.050 ;
        RECT 851.250 197.250 852.750 198.150 ;
        RECT 853.950 196.950 856.050 199.050 ;
        RECT 844.950 193.950 847.050 196.050 ;
        RECT 848.250 194.850 849.750 195.750 ;
        RECT 850.950 193.950 853.050 196.050 ;
        RECT 845.400 193.050 846.450 193.950 ;
        RECT 844.950 190.950 847.050 193.050 ;
        RECT 844.950 178.950 847.050 181.050 ;
        RECT 841.950 166.950 844.050 169.050 ;
        RECT 845.400 166.050 846.450 178.950 ;
        RECT 851.400 178.050 852.450 193.950 ;
        RECT 850.950 175.950 853.050 178.050 ;
        RECT 850.950 172.950 853.050 175.050 ;
        RECT 851.400 169.050 852.450 172.950 ;
        RECT 850.950 166.950 853.050 169.050 ;
        RECT 854.400 166.050 855.450 196.950 ;
        RECT 857.400 172.050 858.450 241.950 ;
        RECT 856.950 169.950 859.050 172.050 ;
        RECT 841.950 164.250 843.750 165.150 ;
        RECT 844.950 163.950 847.050 166.050 ;
        RECT 850.950 163.950 853.050 166.050 ;
        RECT 853.950 163.950 856.050 166.050 ;
        RECT 856.950 163.950 859.050 166.050 ;
        RECT 841.950 160.950 844.050 163.050 ;
        RECT 845.250 161.850 846.750 162.750 ;
        RECT 847.950 160.950 850.050 163.050 ;
        RECT 851.250 161.850 853.050 162.750 ;
        RECT 853.950 160.950 856.050 163.050 ;
        RECT 842.400 136.050 843.450 160.950 ;
        RECT 847.950 158.850 850.050 159.750 ;
        RECT 841.950 133.950 844.050 136.050 ;
        RECT 854.400 133.050 855.450 160.950 ;
        RECT 853.950 130.950 856.050 133.050 ;
        RECT 841.950 127.950 844.050 130.050 ;
        RECT 847.950 127.950 850.050 130.050 ;
        RECT 853.950 128.250 856.050 129.150 ;
        RECT 820.950 121.950 823.050 124.050 ;
        RECT 824.250 122.850 825.750 123.750 ;
        RECT 826.950 121.950 829.050 124.050 ;
        RECT 830.250 122.850 831.750 123.750 ;
        RECT 832.950 121.950 835.050 124.050 ;
        RECT 838.950 121.950 841.050 124.050 ;
        RECT 823.950 115.950 826.050 118.050 ;
        RECT 820.950 109.950 823.050 112.050 ;
        RECT 817.950 97.950 820.050 100.050 ;
        RECT 821.400 94.050 822.450 109.950 ;
        RECT 805.950 92.850 807.750 93.750 ;
        RECT 808.950 91.950 811.050 94.050 ;
        RECT 812.250 92.850 813.750 93.750 ;
        RECT 814.950 91.950 817.050 94.050 ;
        RECT 820.950 91.950 823.050 94.050 ;
        RECT 814.950 89.850 817.050 90.750 ;
        RECT 824.400 82.050 825.450 115.950 ;
        RECT 823.950 79.950 826.050 82.050 ;
        RECT 808.950 76.950 811.050 79.050 ;
        RECT 787.950 67.950 790.050 70.050 ;
        RECT 802.950 67.950 805.050 70.050 ;
        RECT 784.950 52.950 787.050 55.050 ;
        RECT 781.950 28.950 784.050 31.050 ;
        RECT 785.400 25.050 786.450 52.950 ;
        RECT 788.400 51.450 789.450 67.950 ;
        RECT 802.950 61.950 805.050 64.050 ;
        RECT 793.950 58.950 796.050 61.050 ;
        RECT 794.400 55.050 795.450 58.950 ;
        RECT 799.950 56.250 802.050 57.150 ;
        RECT 790.950 53.250 792.750 54.150 ;
        RECT 793.950 52.950 796.050 55.050 ;
        RECT 797.250 53.250 798.750 54.150 ;
        RECT 799.950 52.950 802.050 55.050 ;
        RECT 790.950 51.450 793.050 52.050 ;
        RECT 788.400 50.400 793.050 51.450 ;
        RECT 794.250 50.850 795.750 51.750 ;
        RECT 790.950 49.950 793.050 50.400 ;
        RECT 796.950 49.950 799.050 52.050 ;
        RECT 797.400 34.050 798.450 49.950 ;
        RECT 803.400 37.050 804.450 61.950 ;
        RECT 805.950 58.950 808.050 61.050 ;
        RECT 806.400 52.050 807.450 58.950 ;
        RECT 805.950 49.950 808.050 52.050 ;
        RECT 802.950 34.950 805.050 37.050 ;
        RECT 796.950 31.950 799.050 34.050 ;
        RECT 799.950 28.950 802.050 31.050 ;
        RECT 800.400 25.050 801.450 28.950 ;
        RECT 809.400 25.050 810.450 76.950 ;
        RECT 827.400 76.050 828.450 121.950 ;
        RECT 839.400 106.050 840.450 121.950 ;
        RECT 838.950 103.950 841.050 106.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 833.400 97.050 834.450 100.950 ;
        RECT 839.400 97.050 840.450 103.950 ;
        RECT 829.950 94.950 832.050 97.050 ;
        RECT 832.950 94.950 835.050 97.050 ;
        RECT 836.250 95.250 837.750 96.150 ;
        RECT 838.950 94.950 841.050 97.050 ;
        RECT 830.400 94.050 831.450 94.950 ;
        RECT 829.950 91.950 832.050 94.050 ;
        RECT 833.250 92.850 834.750 93.750 ;
        RECT 835.950 91.950 838.050 94.050 ;
        RECT 839.250 92.850 841.050 93.750 ;
        RECT 829.950 89.850 832.050 90.750 ;
        RECT 826.950 73.950 829.050 76.050 ;
        RECT 811.950 70.950 814.050 73.050 ;
        RECT 838.950 70.950 841.050 73.050 ;
        RECT 812.400 49.050 813.450 70.950 ;
        RECT 826.950 58.950 829.050 61.050 ;
        RECT 832.950 58.950 835.050 61.050 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 811.950 46.950 814.050 49.050 ;
        RECT 784.950 22.950 787.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 799.950 24.450 802.050 25.050 ;
        RECT 796.950 23.250 798.750 24.150 ;
        RECT 799.950 23.400 804.450 24.450 ;
        RECT 799.950 22.950 802.050 23.400 ;
        RECT 781.950 20.250 783.750 21.150 ;
        RECT 784.950 19.950 787.050 22.050 ;
        RECT 794.400 21.450 795.450 22.950 ;
        RECT 803.400 22.050 804.450 23.400 ;
        RECT 805.950 23.250 807.750 24.150 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 796.950 21.450 799.050 22.050 ;
        RECT 788.250 20.250 790.050 21.150 ;
        RECT 794.400 20.400 799.050 21.450 ;
        RECT 800.250 20.850 802.050 21.750 ;
        RECT 796.950 19.950 799.050 20.400 ;
        RECT 802.950 19.950 805.050 22.050 ;
        RECT 805.950 19.950 808.050 22.050 ;
        RECT 809.250 20.850 811.050 21.750 ;
        RECT 806.400 19.050 807.450 19.950 ;
        RECT 815.400 19.050 816.450 55.950 ;
        RECT 827.400 55.050 828.450 58.950 ;
        RECT 817.950 53.250 819.750 54.150 ;
        RECT 820.950 52.950 823.050 55.050 ;
        RECT 826.950 52.950 829.050 55.050 ;
        RECT 817.950 49.950 820.050 52.050 ;
        RECT 821.250 50.850 823.050 51.750 ;
        RECT 823.950 50.250 826.050 51.150 ;
        RECT 826.950 50.850 829.050 51.750 ;
        RECT 833.400 51.450 834.450 58.950 ;
        RECT 839.400 55.050 840.450 70.950 ;
        RECT 842.400 67.050 843.450 127.950 ;
        RECT 848.400 127.050 849.450 127.950 ;
        RECT 844.950 125.250 846.750 126.150 ;
        RECT 847.950 124.950 850.050 127.050 ;
        RECT 851.250 125.250 852.750 126.150 ;
        RECT 853.950 124.950 856.050 127.050 ;
        RECT 844.950 121.950 847.050 124.050 ;
        RECT 848.250 122.850 849.750 123.750 ;
        RECT 850.950 121.950 853.050 124.050 ;
        RECT 845.400 100.050 846.450 121.950 ;
        RECT 847.950 109.950 850.050 112.050 ;
        RECT 844.950 97.950 847.050 100.050 ;
        RECT 841.950 64.950 844.050 67.050 ;
        RECT 842.400 58.050 843.450 64.950 ;
        RECT 845.400 61.050 846.450 97.950 ;
        RECT 848.400 97.050 849.450 109.950 ;
        RECT 850.950 106.950 853.050 109.050 ;
        RECT 851.400 100.050 852.450 106.950 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 847.950 94.950 850.050 97.050 ;
        RECT 851.250 95.850 852.750 96.750 ;
        RECT 853.950 94.950 856.050 97.050 ;
        RECT 847.950 92.850 850.050 93.750 ;
        RECT 853.950 92.850 856.050 93.750 ;
        RECT 847.950 88.950 850.050 91.050 ;
        RECT 857.400 90.450 858.450 163.950 ;
        RECT 860.400 91.050 861.450 304.950 ;
        RECT 862.950 244.950 865.050 247.050 ;
        RECT 863.400 241.050 864.450 244.950 ;
        RECT 869.400 241.050 870.450 853.950 ;
        RECT 871.950 571.950 874.050 574.050 ;
        RECT 872.400 322.050 873.450 571.950 ;
        RECT 871.950 319.950 874.050 322.050 ;
        RECT 862.950 238.950 865.050 241.050 ;
        RECT 866.250 239.250 868.050 240.150 ;
        RECT 868.950 238.950 871.050 241.050 ;
        RECT 862.950 236.850 864.750 237.750 ;
        RECT 865.950 235.950 868.050 238.050 ;
        RECT 868.950 235.950 871.050 238.050 ;
        RECT 866.400 229.050 867.450 235.950 ;
        RECT 865.950 226.950 868.050 229.050 ;
        RECT 865.950 223.950 868.050 226.050 ;
        RECT 862.950 202.950 865.050 205.050 ;
        RECT 863.400 175.050 864.450 202.950 ;
        RECT 862.950 172.950 865.050 175.050 ;
        RECT 866.400 172.050 867.450 223.950 ;
        RECT 865.950 169.950 868.050 172.050 ;
        RECT 862.950 167.250 865.050 168.150 ;
        RECT 865.950 167.850 868.050 168.750 ;
        RECT 862.950 163.950 865.050 166.050 ;
        RECT 865.950 163.950 868.050 166.050 ;
        RECT 862.950 130.950 865.050 133.050 ;
        RECT 854.400 89.400 858.450 90.450 ;
        RECT 844.950 58.950 847.050 61.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 844.950 56.250 847.050 57.150 ;
        RECT 835.950 53.250 837.750 54.150 ;
        RECT 838.950 52.950 841.050 55.050 ;
        RECT 842.250 53.250 843.750 54.150 ;
        RECT 844.950 52.950 847.050 55.050 ;
        RECT 835.950 51.450 838.050 52.050 ;
        RECT 833.400 50.400 838.050 51.450 ;
        RECT 839.250 50.850 840.750 51.750 ;
        RECT 835.950 49.950 838.050 50.400 ;
        RECT 841.950 49.950 844.050 52.050 ;
        RECT 818.400 28.050 819.450 49.950 ;
        RECT 823.950 46.950 826.050 49.050 ;
        RECT 817.950 27.450 820.050 28.050 ;
        RECT 820.950 27.450 823.050 28.050 ;
        RECT 817.950 26.400 823.050 27.450 ;
        RECT 817.950 25.950 820.050 26.400 ;
        RECT 820.950 25.950 823.050 26.400 ;
        RECT 841.950 25.950 844.050 28.050 ;
        RECT 820.950 23.850 823.050 24.750 ;
        RECT 823.950 23.250 826.050 24.150 ;
        RECT 838.950 23.250 841.050 24.150 ;
        RECT 841.950 23.850 844.050 24.750 ;
        RECT 848.400 22.050 849.450 88.950 ;
        RECT 850.950 79.950 853.050 82.050 ;
        RECT 851.400 28.050 852.450 79.950 ;
        RECT 850.950 25.950 853.050 28.050 ;
        RECT 854.400 22.050 855.450 89.400 ;
        RECT 859.950 88.950 862.050 91.050 ;
        RECT 863.400 61.050 864.450 130.950 ;
        RECT 856.950 58.950 859.050 61.050 ;
        RECT 862.950 58.950 865.050 61.050 ;
        RECT 857.400 58.050 858.450 58.950 ;
        RECT 856.950 55.950 859.050 58.050 ;
        RECT 862.950 57.450 865.050 58.050 ;
        RECT 866.400 57.450 867.450 163.950 ;
        RECT 860.250 56.250 861.750 57.150 ;
        RECT 862.950 56.400 867.450 57.450 ;
        RECT 862.950 55.950 865.050 56.400 ;
        RECT 869.400 55.050 870.450 235.950 ;
        RECT 856.950 53.850 858.750 54.750 ;
        RECT 859.950 52.950 862.050 55.050 ;
        RECT 863.250 53.850 865.050 54.750 ;
        RECT 868.950 52.950 871.050 55.050 ;
        RECT 859.950 25.950 862.050 28.050 ;
        RECT 823.950 19.950 826.050 22.050 ;
        RECT 838.950 19.950 841.050 22.050 ;
        RECT 847.950 19.950 850.050 22.050 ;
        RECT 850.950 20.250 852.750 21.150 ;
        RECT 853.950 19.950 856.050 22.050 ;
        RECT 857.250 20.250 859.050 21.150 ;
        RECT 781.950 18.450 784.050 19.050 ;
        RECT 779.400 17.400 784.050 18.450 ;
        RECT 785.250 17.850 786.750 18.750 ;
        RECT 727.950 16.950 730.050 17.400 ;
        RECT 781.950 16.950 784.050 17.400 ;
        RECT 787.950 16.950 790.050 19.050 ;
        RECT 805.950 16.950 808.050 19.050 ;
        RECT 814.950 16.950 817.050 19.050 ;
        RECT 850.950 16.950 853.050 19.050 ;
        RECT 854.250 17.850 855.750 18.750 ;
        RECT 856.950 18.450 859.050 19.050 ;
        RECT 860.400 18.450 861.450 25.950 ;
        RECT 856.950 17.400 861.450 18.450 ;
        RECT 856.950 16.950 859.050 17.400 ;
        RECT 16.950 14.850 19.050 15.750 ;
        RECT 28.950 13.950 31.050 16.050 ;
        RECT 118.950 13.950 121.050 16.050 ;
        RECT 124.950 14.850 127.050 15.750 ;
        RECT 277.950 13.950 280.050 16.050 ;
        RECT 289.950 14.850 292.050 15.750 ;
        RECT 313.950 13.950 316.050 16.050 ;
        RECT 319.950 14.850 322.050 15.750 ;
        RECT 415.950 13.950 418.050 16.050 ;
        RECT 433.950 13.950 436.050 16.050 ;
        RECT 445.950 13.950 448.050 16.050 ;
        RECT 454.950 13.950 457.050 16.050 ;
        RECT 472.950 13.950 475.050 16.050 ;
        RECT 478.950 14.850 481.050 15.750 ;
        RECT 544.950 13.950 547.050 16.050 ;
        RECT 679.950 13.950 682.050 16.050 ;
        RECT 685.950 14.850 688.050 15.750 ;
        RECT 694.950 13.950 697.050 16.050 ;
      LAYER metal3 ;
        RECT 817.950 855.600 820.050 856.050 ;
        RECT 868.950 855.600 871.050 856.050 ;
        RECT 817.950 854.400 871.050 855.600 ;
        RECT 817.950 853.950 820.050 854.400 ;
        RECT 868.950 853.950 871.050 854.400 ;
        RECT 724.950 852.600 727.050 853.050 ;
        RECT 745.950 852.600 748.050 853.050 ;
        RECT 724.950 851.400 748.050 852.600 ;
        RECT 724.950 850.950 727.050 851.400 ;
        RECT 745.950 850.950 748.050 851.400 ;
        RECT 67.950 849.600 70.050 850.050 ;
        RECT 76.950 849.600 79.050 850.050 ;
        RECT 67.950 848.400 79.050 849.600 ;
        RECT 67.950 847.950 70.050 848.400 ;
        RECT 76.950 847.950 79.050 848.400 ;
        RECT 124.950 849.600 127.050 850.050 ;
        RECT 199.950 849.600 202.050 850.050 ;
        RECT 124.950 848.400 202.050 849.600 ;
        RECT 124.950 847.950 127.050 848.400 ;
        RECT 199.950 847.950 202.050 848.400 ;
        RECT 223.950 849.600 226.050 850.050 ;
        RECT 244.950 849.600 247.050 850.050 ;
        RECT 223.950 848.400 247.050 849.600 ;
        RECT 223.950 847.950 226.050 848.400 ;
        RECT 244.950 847.950 247.050 848.400 ;
        RECT 289.950 849.600 292.050 850.050 ;
        RECT 310.950 849.600 313.050 850.050 ;
        RECT 316.950 849.600 319.050 850.050 ;
        RECT 289.950 848.400 319.050 849.600 ;
        RECT 289.950 847.950 292.050 848.400 ;
        RECT 310.950 847.950 313.050 848.400 ;
        RECT 316.950 847.950 319.050 848.400 ;
        RECT 355.950 849.600 358.050 850.050 ;
        RECT 367.950 849.600 370.050 850.050 ;
        RECT 355.950 848.400 370.050 849.600 ;
        RECT 355.950 847.950 358.050 848.400 ;
        RECT 367.950 847.950 370.050 848.400 ;
        RECT 391.950 849.600 394.050 850.050 ;
        RECT 406.950 849.600 409.050 850.050 ;
        RECT 391.950 848.400 409.050 849.600 ;
        RECT 391.950 847.950 394.050 848.400 ;
        RECT 406.950 847.950 409.050 848.400 ;
        RECT 412.950 849.600 415.050 850.050 ;
        RECT 418.950 849.600 421.050 850.050 ;
        RECT 430.950 849.600 433.050 850.050 ;
        RECT 487.950 849.600 490.050 850.050 ;
        RECT 514.950 849.600 517.050 850.050 ;
        RECT 523.950 849.600 526.050 850.050 ;
        RECT 412.950 848.400 526.050 849.600 ;
        RECT 412.950 847.950 415.050 848.400 ;
        RECT 418.950 847.950 421.050 848.400 ;
        RECT 430.950 847.950 433.050 848.400 ;
        RECT 487.950 847.950 490.050 848.400 ;
        RECT 514.950 847.950 517.050 848.400 ;
        RECT 523.950 847.950 526.050 848.400 ;
        RECT 529.950 849.600 532.050 850.050 ;
        RECT 613.950 849.600 616.050 850.050 ;
        RECT 733.950 849.600 736.050 850.050 ;
        RECT 796.950 849.600 799.050 850.050 ;
        RECT 529.950 848.400 616.050 849.600 ;
        RECT 529.950 847.950 532.050 848.400 ;
        RECT 613.950 847.950 616.050 848.400 ;
        RECT 668.400 848.400 687.600 849.600 ;
        RECT 668.400 847.050 669.600 848.400 ;
        RECT 16.950 846.600 19.050 847.050 ;
        RECT 31.950 846.600 34.050 847.050 ;
        RECT 58.950 846.600 61.050 847.050 ;
        RECT 79.950 846.600 82.050 847.050 ;
        RECT 16.950 845.400 36.600 846.600 ;
        RECT 16.950 844.950 19.050 845.400 ;
        RECT 31.950 844.950 34.050 845.400 ;
        RECT 19.950 843.600 22.050 844.050 ;
        RECT 28.950 843.600 31.050 844.050 ;
        RECT 19.950 842.400 31.050 843.600 ;
        RECT 35.400 843.600 36.600 845.400 ;
        RECT 58.950 845.400 82.050 846.600 ;
        RECT 58.950 844.950 61.050 845.400 ;
        RECT 79.950 844.950 82.050 845.400 ;
        RECT 103.950 846.600 106.050 847.050 ;
        RECT 109.950 846.600 112.050 847.050 ;
        RECT 103.950 845.400 112.050 846.600 ;
        RECT 103.950 844.950 106.050 845.400 ;
        RECT 109.950 844.950 112.050 845.400 ;
        RECT 133.950 846.600 136.050 847.050 ;
        RECT 139.950 846.600 142.050 847.050 ;
        RECT 133.950 845.400 142.050 846.600 ;
        RECT 133.950 844.950 136.050 845.400 ;
        RECT 139.950 844.950 142.050 845.400 ;
        RECT 181.950 844.950 184.050 847.050 ;
        RECT 226.950 846.600 229.050 847.050 ;
        RECT 250.950 846.600 253.050 847.050 ;
        RECT 262.950 846.600 265.050 847.050 ;
        RECT 226.950 845.400 265.050 846.600 ;
        RECT 226.950 844.950 229.050 845.400 ;
        RECT 250.950 844.950 253.050 845.400 ;
        RECT 262.950 844.950 265.050 845.400 ;
        RECT 304.950 846.600 307.050 847.050 ;
        RECT 319.950 846.600 322.050 847.050 ;
        RECT 325.950 846.600 328.050 847.050 ;
        RECT 304.950 845.400 328.050 846.600 ;
        RECT 304.950 844.950 307.050 845.400 ;
        RECT 319.950 844.950 322.050 845.400 ;
        RECT 325.950 844.950 328.050 845.400 ;
        RECT 349.950 846.600 352.050 847.050 ;
        RECT 361.950 846.600 364.050 847.050 ;
        RECT 349.950 845.400 364.050 846.600 ;
        RECT 349.950 844.950 352.050 845.400 ;
        RECT 361.950 844.950 364.050 845.400 ;
        RECT 370.950 846.600 373.050 847.050 ;
        RECT 388.950 846.600 391.050 847.050 ;
        RECT 370.950 845.400 391.050 846.600 ;
        RECT 370.950 844.950 373.050 845.400 ;
        RECT 388.950 844.950 391.050 845.400 ;
        RECT 394.950 846.600 397.050 847.050 ;
        RECT 403.950 846.600 406.050 847.050 ;
        RECT 394.950 845.400 406.050 846.600 ;
        RECT 394.950 844.950 397.050 845.400 ;
        RECT 403.950 844.950 406.050 845.400 ;
        RECT 445.950 846.600 448.050 847.050 ;
        RECT 460.950 846.600 463.050 847.050 ;
        RECT 445.950 845.400 463.050 846.600 ;
        RECT 445.950 844.950 448.050 845.400 ;
        RECT 460.950 844.950 463.050 845.400 ;
        RECT 466.950 844.950 469.050 847.050 ;
        RECT 526.950 846.600 529.050 847.050 ;
        RECT 547.950 846.600 550.050 847.050 ;
        RECT 526.950 845.400 550.050 846.600 ;
        RECT 526.950 844.950 529.050 845.400 ;
        RECT 547.950 844.950 550.050 845.400 ;
        RECT 577.950 846.600 580.050 847.050 ;
        RECT 592.950 846.600 595.050 847.050 ;
        RECT 577.950 845.400 595.050 846.600 ;
        RECT 577.950 844.950 580.050 845.400 ;
        RECT 592.950 844.950 595.050 845.400 ;
        RECT 667.950 844.950 670.050 847.050 ;
        RECT 673.950 846.600 676.050 847.050 ;
        RECT 682.950 846.600 685.050 847.050 ;
        RECT 673.950 845.400 685.050 846.600 ;
        RECT 686.400 846.600 687.600 848.400 ;
        RECT 733.950 848.400 799.050 849.600 ;
        RECT 733.950 847.950 736.050 848.400 ;
        RECT 796.950 847.950 799.050 848.400 ;
        RECT 778.950 846.600 781.050 847.050 ;
        RECT 686.400 845.400 781.050 846.600 ;
        RECT 673.950 844.950 676.050 845.400 ;
        RECT 682.950 844.950 685.050 845.400 ;
        RECT 778.950 844.950 781.050 845.400 ;
        RECT 850.950 846.600 853.050 847.050 ;
        RECT 856.950 846.600 859.050 847.050 ;
        RECT 850.950 845.400 859.050 846.600 ;
        RECT 850.950 844.950 853.050 845.400 ;
        RECT 856.950 844.950 859.050 845.400 ;
        RECT 55.950 843.600 58.050 844.050 ;
        RECT 35.400 842.400 58.050 843.600 ;
        RECT 19.950 841.950 22.050 842.400 ;
        RECT 28.950 841.950 31.050 842.400 ;
        RECT 55.950 841.950 58.050 842.400 ;
        RECT 115.950 843.600 118.050 844.050 ;
        RECT 182.400 843.600 183.600 844.950 ;
        RECT 115.950 842.400 183.600 843.600 ;
        RECT 187.950 843.600 190.050 844.050 ;
        RECT 205.950 843.600 208.050 844.050 ;
        RECT 208.950 843.600 211.050 844.050 ;
        RECT 187.950 842.400 211.050 843.600 ;
        RECT 115.950 841.950 118.050 842.400 ;
        RECT 187.950 841.950 190.050 842.400 ;
        RECT 205.950 841.950 208.050 842.400 ;
        RECT 208.950 841.950 211.050 842.400 ;
        RECT 232.950 843.600 235.050 844.050 ;
        RECT 259.950 843.600 262.050 844.050 ;
        RECT 232.950 842.400 262.050 843.600 ;
        RECT 232.950 841.950 235.050 842.400 ;
        RECT 259.950 841.950 262.050 842.400 ;
        RECT 280.950 843.600 283.050 844.050 ;
        RECT 331.950 843.600 334.050 844.050 ;
        RECT 280.950 842.400 334.050 843.600 ;
        RECT 467.400 843.600 468.600 844.950 ;
        RECT 484.950 843.600 487.050 844.050 ;
        RECT 467.400 842.400 487.050 843.600 ;
        RECT 280.950 841.950 283.050 842.400 ;
        RECT 331.950 841.950 334.050 842.400 ;
        RECT 484.950 841.950 487.050 842.400 ;
        RECT 493.950 843.600 496.050 844.050 ;
        RECT 505.950 843.600 508.050 844.050 ;
        RECT 523.950 843.600 526.050 844.050 ;
        RECT 493.950 842.400 526.050 843.600 ;
        RECT 493.950 841.950 496.050 842.400 ;
        RECT 505.950 841.950 508.050 842.400 ;
        RECT 523.950 841.950 526.050 842.400 ;
        RECT 640.950 843.600 643.050 844.050 ;
        RECT 670.950 843.600 673.050 844.050 ;
        RECT 640.950 842.400 673.050 843.600 ;
        RECT 640.950 841.950 643.050 842.400 ;
        RECT 670.950 841.950 673.050 842.400 ;
        RECT 793.950 843.600 796.050 844.050 ;
        RECT 805.950 843.600 808.050 844.050 ;
        RECT 793.950 842.400 808.050 843.600 ;
        RECT 793.950 841.950 796.050 842.400 ;
        RECT 805.950 841.950 808.050 842.400 ;
        RECT 61.950 840.600 64.050 841.050 ;
        RECT 73.950 840.600 76.050 841.050 ;
        RECT 61.950 839.400 76.050 840.600 ;
        RECT 61.950 838.950 64.050 839.400 ;
        RECT 73.950 838.950 76.050 839.400 ;
        RECT 79.950 840.600 82.050 841.050 ;
        RECT 136.950 840.600 139.050 841.050 ;
        RECT 79.950 839.400 139.050 840.600 ;
        RECT 79.950 838.950 82.050 839.400 ;
        RECT 136.950 838.950 139.050 839.400 ;
        RECT 148.950 840.600 151.050 841.050 ;
        RECT 160.950 840.600 163.050 841.050 ;
        RECT 148.950 839.400 163.050 840.600 ;
        RECT 148.950 838.950 151.050 839.400 ;
        RECT 160.950 838.950 163.050 839.400 ;
        RECT 190.950 840.600 193.050 841.050 ;
        RECT 211.950 840.600 214.050 841.050 ;
        RECT 190.950 839.400 214.050 840.600 ;
        RECT 190.950 838.950 193.050 839.400 ;
        RECT 211.950 838.950 214.050 839.400 ;
        RECT 229.950 840.600 232.050 841.050 ;
        RECT 253.950 840.600 256.050 841.050 ;
        RECT 265.950 840.600 268.050 841.050 ;
        RECT 274.950 840.600 277.050 841.050 ;
        RECT 229.950 839.400 277.050 840.600 ;
        RECT 229.950 838.950 232.050 839.400 ;
        RECT 253.950 838.950 256.050 839.400 ;
        RECT 265.950 838.950 268.050 839.400 ;
        RECT 274.950 838.950 277.050 839.400 ;
        RECT 277.950 840.600 280.050 841.050 ;
        RECT 286.950 840.600 289.050 841.050 ;
        RECT 277.950 839.400 289.050 840.600 ;
        RECT 277.950 838.950 280.050 839.400 ;
        RECT 286.950 838.950 289.050 839.400 ;
        RECT 316.950 840.600 319.050 841.050 ;
        RECT 322.950 840.600 325.050 841.050 ;
        RECT 316.950 839.400 325.050 840.600 ;
        RECT 316.950 838.950 319.050 839.400 ;
        RECT 322.950 838.950 325.050 839.400 ;
        RECT 328.950 840.600 331.050 841.050 ;
        RECT 409.950 840.600 412.050 841.050 ;
        RECT 328.950 839.400 412.050 840.600 ;
        RECT 328.950 838.950 331.050 839.400 ;
        RECT 409.950 838.950 412.050 839.400 ;
        RECT 469.950 840.600 472.050 841.050 ;
        RECT 508.950 840.600 511.050 841.050 ;
        RECT 469.950 839.400 511.050 840.600 ;
        RECT 469.950 838.950 472.050 839.400 ;
        RECT 508.950 838.950 511.050 839.400 ;
        RECT 550.950 840.600 553.050 841.050 ;
        RECT 589.950 840.600 592.050 841.050 ;
        RECT 550.950 839.400 592.050 840.600 ;
        RECT 550.950 838.950 553.050 839.400 ;
        RECT 589.950 838.950 592.050 839.400 ;
        RECT 598.950 840.600 601.050 841.050 ;
        RECT 610.950 840.600 613.050 841.050 ;
        RECT 598.950 839.400 613.050 840.600 ;
        RECT 598.950 838.950 601.050 839.400 ;
        RECT 610.950 838.950 613.050 839.400 ;
        RECT 634.950 840.600 637.050 841.050 ;
        RECT 685.950 840.600 688.050 841.050 ;
        RECT 634.950 839.400 688.050 840.600 ;
        RECT 634.950 838.950 637.050 839.400 ;
        RECT 685.950 838.950 688.050 839.400 ;
        RECT 721.950 840.600 724.050 841.050 ;
        RECT 727.950 840.600 730.050 841.050 ;
        RECT 721.950 839.400 730.050 840.600 ;
        RECT 721.950 838.950 724.050 839.400 ;
        RECT 727.950 838.950 730.050 839.400 ;
        RECT 739.950 840.600 742.050 841.050 ;
        RECT 763.950 840.600 766.050 841.050 ;
        RECT 739.950 839.400 766.050 840.600 ;
        RECT 739.950 838.950 742.050 839.400 ;
        RECT 763.950 838.950 766.050 839.400 ;
        RECT 796.950 840.600 799.050 841.050 ;
        RECT 802.950 840.600 805.050 841.050 ;
        RECT 796.950 839.400 805.050 840.600 ;
        RECT 796.950 838.950 799.050 839.400 ;
        RECT 802.950 838.950 805.050 839.400 ;
        RECT 814.950 840.600 817.050 841.050 ;
        RECT 826.950 840.600 829.050 841.050 ;
        RECT 814.950 839.400 829.050 840.600 ;
        RECT 814.950 838.950 817.050 839.400 ;
        RECT 826.950 838.950 829.050 839.400 ;
        RECT 106.950 837.600 109.050 838.050 ;
        RECT 133.950 837.600 136.050 838.050 ;
        RECT 163.950 837.600 166.050 838.050 ;
        RECT 106.950 836.400 166.050 837.600 ;
        RECT 106.950 835.950 109.050 836.400 ;
        RECT 133.950 835.950 136.050 836.400 ;
        RECT 163.950 835.950 166.050 836.400 ;
        RECT 166.950 837.600 169.050 838.050 ;
        RECT 202.950 837.600 205.050 838.050 ;
        RECT 166.950 836.400 205.050 837.600 ;
        RECT 166.950 835.950 169.050 836.400 ;
        RECT 202.950 835.950 205.050 836.400 ;
        RECT 286.950 837.600 289.050 838.050 ;
        RECT 346.950 837.600 349.050 838.050 ;
        RECT 286.950 836.400 349.050 837.600 ;
        RECT 286.950 835.950 289.050 836.400 ;
        RECT 346.950 835.950 349.050 836.400 ;
        RECT 541.950 837.600 544.050 838.050 ;
        RECT 565.950 837.600 568.050 838.050 ;
        RECT 619.950 837.600 622.050 838.050 ;
        RECT 541.950 836.400 622.050 837.600 ;
        RECT 541.950 835.950 544.050 836.400 ;
        RECT 565.950 835.950 568.050 836.400 ;
        RECT 619.950 835.950 622.050 836.400 ;
        RECT 811.950 837.600 814.050 838.050 ;
        RECT 847.950 837.600 850.050 838.050 ;
        RECT 811.950 836.400 850.050 837.600 ;
        RECT 811.950 835.950 814.050 836.400 ;
        RECT 847.950 835.950 850.050 836.400 ;
        RECT 97.950 834.600 100.050 835.050 ;
        RECT 118.950 834.600 121.050 835.050 ;
        RECT 121.950 834.600 124.050 835.050 ;
        RECT 97.950 833.400 124.050 834.600 ;
        RECT 97.950 832.950 100.050 833.400 ;
        RECT 118.950 832.950 121.050 833.400 ;
        RECT 121.950 832.950 124.050 833.400 ;
        RECT 271.950 834.600 274.050 835.050 ;
        RECT 340.950 834.600 343.050 835.050 ;
        RECT 346.950 834.600 349.050 835.050 ;
        RECT 271.950 833.400 349.050 834.600 ;
        RECT 271.950 832.950 274.050 833.400 ;
        RECT 340.950 832.950 343.050 833.400 ;
        RECT 346.950 832.950 349.050 833.400 ;
        RECT 415.950 834.600 418.050 835.050 ;
        RECT 421.950 834.600 424.050 835.050 ;
        RECT 595.950 834.600 598.050 835.050 ;
        RECT 415.950 833.400 598.050 834.600 ;
        RECT 415.950 832.950 418.050 833.400 ;
        RECT 421.950 832.950 424.050 833.400 ;
        RECT 595.950 832.950 598.050 833.400 ;
        RECT 37.950 831.600 40.050 832.050 ;
        RECT 97.950 831.600 100.050 832.050 ;
        RECT 157.950 831.600 160.050 832.050 ;
        RECT 208.950 831.600 211.050 832.050 ;
        RECT 37.950 830.400 211.050 831.600 ;
        RECT 37.950 829.950 40.050 830.400 ;
        RECT 97.950 829.950 100.050 830.400 ;
        RECT 157.950 829.950 160.050 830.400 ;
        RECT 208.950 829.950 211.050 830.400 ;
        RECT 355.950 831.600 358.050 832.050 ;
        RECT 415.950 831.600 418.050 832.050 ;
        RECT 430.950 831.600 433.050 832.050 ;
        RECT 355.950 830.400 433.050 831.600 ;
        RECT 355.950 829.950 358.050 830.400 ;
        RECT 415.950 829.950 418.050 830.400 ;
        RECT 430.950 829.950 433.050 830.400 ;
        RECT 448.950 831.600 451.050 832.050 ;
        RECT 556.950 831.600 559.050 832.050 ;
        RECT 448.950 830.400 559.050 831.600 ;
        RECT 448.950 829.950 451.050 830.400 ;
        RECT 556.950 829.950 559.050 830.400 ;
        RECT 559.950 831.600 562.050 832.050 ;
        RECT 595.950 831.600 598.050 832.050 ;
        RECT 559.950 830.400 598.050 831.600 ;
        RECT 559.950 829.950 562.050 830.400 ;
        RECT 595.950 829.950 598.050 830.400 ;
        RECT 508.950 828.600 511.050 829.050 ;
        RECT 568.950 828.600 571.050 829.050 ;
        RECT 508.950 827.400 571.050 828.600 ;
        RECT 508.950 826.950 511.050 827.400 ;
        RECT 568.950 826.950 571.050 827.400 ;
        RECT 592.950 828.600 595.050 829.050 ;
        RECT 679.950 828.600 682.050 829.050 ;
        RECT 592.950 827.400 682.050 828.600 ;
        RECT 592.950 826.950 595.050 827.400 ;
        RECT 679.950 826.950 682.050 827.400 ;
        RECT 685.950 828.600 688.050 829.050 ;
        RECT 736.950 828.600 739.050 829.050 ;
        RECT 754.950 828.600 757.050 829.050 ;
        RECT 787.950 828.600 790.050 829.050 ;
        RECT 685.950 827.400 790.050 828.600 ;
        RECT 685.950 826.950 688.050 827.400 ;
        RECT 736.950 826.950 739.050 827.400 ;
        RECT 754.950 826.950 757.050 827.400 ;
        RECT 787.950 826.950 790.050 827.400 ;
        RECT 205.950 825.600 208.050 826.050 ;
        RECT 562.950 825.600 565.050 826.050 ;
        RECT 205.950 824.400 565.050 825.600 ;
        RECT 205.950 823.950 208.050 824.400 ;
        RECT 562.950 823.950 565.050 824.400 ;
        RECT 565.950 825.600 568.050 826.050 ;
        RECT 577.950 825.600 580.050 826.050 ;
        RECT 592.950 825.600 595.050 826.050 ;
        RECT 565.950 824.400 595.050 825.600 ;
        RECT 565.950 823.950 568.050 824.400 ;
        RECT 577.950 823.950 580.050 824.400 ;
        RECT 592.950 823.950 595.050 824.400 ;
        RECT 595.950 825.600 598.050 826.050 ;
        RECT 682.950 825.600 685.050 826.050 ;
        RECT 706.950 825.600 709.050 826.050 ;
        RECT 595.950 824.400 709.050 825.600 ;
        RECT 595.950 823.950 598.050 824.400 ;
        RECT 682.950 823.950 685.050 824.400 ;
        RECT 706.950 823.950 709.050 824.400 ;
        RECT 13.950 822.600 16.050 823.050 ;
        RECT 58.950 822.600 61.050 823.050 ;
        RECT 13.950 821.400 61.050 822.600 ;
        RECT 13.950 820.950 16.050 821.400 ;
        RECT 58.950 820.950 61.050 821.400 ;
        RECT 79.950 822.600 82.050 823.050 ;
        RECT 85.950 822.600 88.050 823.050 ;
        RECT 103.950 822.600 106.050 823.050 ;
        RECT 79.950 821.400 106.050 822.600 ;
        RECT 79.950 820.950 82.050 821.400 ;
        RECT 85.950 820.950 88.050 821.400 ;
        RECT 103.950 820.950 106.050 821.400 ;
        RECT 241.950 822.600 244.050 823.050 ;
        RECT 244.950 822.600 247.050 823.050 ;
        RECT 253.950 822.600 256.050 823.050 ;
        RECT 241.950 821.400 256.050 822.600 ;
        RECT 241.950 820.950 244.050 821.400 ;
        RECT 244.950 820.950 247.050 821.400 ;
        RECT 253.950 820.950 256.050 821.400 ;
        RECT 295.950 822.600 298.050 823.050 ;
        RECT 382.950 822.600 385.050 823.050 ;
        RECT 439.950 822.600 442.050 823.050 ;
        RECT 295.950 821.400 442.050 822.600 ;
        RECT 295.950 820.950 298.050 821.400 ;
        RECT 382.950 820.950 385.050 821.400 ;
        RECT 439.950 820.950 442.050 821.400 ;
        RECT 529.950 822.600 532.050 823.050 ;
        RECT 586.950 822.600 589.050 823.050 ;
        RECT 529.950 821.400 589.050 822.600 ;
        RECT 529.950 820.950 532.050 821.400 ;
        RECT 586.950 820.950 589.050 821.400 ;
        RECT 664.950 822.600 667.050 823.050 ;
        RECT 763.950 822.600 766.050 823.050 ;
        RECT 769.950 822.600 772.050 823.050 ;
        RECT 664.950 821.400 772.050 822.600 ;
        RECT 664.950 820.950 667.050 821.400 ;
        RECT 763.950 820.950 766.050 821.400 ;
        RECT 769.950 820.950 772.050 821.400 ;
        RECT 10.950 819.600 13.050 820.050 ;
        RECT 19.950 819.600 22.050 820.050 ;
        RECT 85.950 819.600 88.050 820.050 ;
        RECT 115.950 819.600 118.050 820.050 ;
        RECT 10.950 818.400 118.050 819.600 ;
        RECT 10.950 817.950 13.050 818.400 ;
        RECT 19.950 817.950 22.050 818.400 ;
        RECT 85.950 817.950 88.050 818.400 ;
        RECT 115.950 817.950 118.050 818.400 ;
        RECT 169.950 819.600 172.050 820.050 ;
        RECT 175.950 819.600 178.050 820.050 ;
        RECT 169.950 818.400 178.050 819.600 ;
        RECT 169.950 817.950 172.050 818.400 ;
        RECT 175.950 817.950 178.050 818.400 ;
        RECT 247.950 817.950 250.050 820.050 ;
        RECT 259.950 819.600 262.050 820.050 ;
        RECT 277.950 819.600 280.050 820.050 ;
        RECT 307.950 819.600 310.050 820.050 ;
        RECT 259.950 818.400 310.050 819.600 ;
        RECT 259.950 817.950 262.050 818.400 ;
        RECT 277.950 817.950 280.050 818.400 ;
        RECT 307.950 817.950 310.050 818.400 ;
        RECT 313.950 819.600 316.050 820.050 ;
        RECT 334.950 819.600 337.050 820.050 ;
        RECT 361.950 819.600 364.050 820.050 ;
        RECT 313.950 818.400 364.050 819.600 ;
        RECT 313.950 817.950 316.050 818.400 ;
        RECT 334.950 817.950 337.050 818.400 ;
        RECT 361.950 817.950 364.050 818.400 ;
        RECT 373.950 819.600 376.050 820.050 ;
        RECT 376.950 819.600 379.050 820.050 ;
        RECT 427.950 819.600 430.050 820.050 ;
        RECT 373.950 818.400 430.050 819.600 ;
        RECT 373.950 817.950 376.050 818.400 ;
        RECT 376.950 817.950 379.050 818.400 ;
        RECT 427.950 817.950 430.050 818.400 ;
        RECT 436.950 819.600 439.050 820.050 ;
        RECT 451.950 819.600 454.050 820.050 ;
        RECT 487.950 819.600 490.050 820.050 ;
        RECT 436.950 818.400 490.050 819.600 ;
        RECT 436.950 817.950 439.050 818.400 ;
        RECT 451.950 817.950 454.050 818.400 ;
        RECT 487.950 817.950 490.050 818.400 ;
        RECT 532.950 819.600 535.050 820.050 ;
        RECT 574.950 819.600 577.050 820.050 ;
        RECT 646.950 819.600 649.050 820.050 ;
        RECT 532.950 818.400 649.050 819.600 ;
        RECT 532.950 817.950 535.050 818.400 ;
        RECT 574.950 817.950 577.050 818.400 ;
        RECT 646.950 817.950 649.050 818.400 ;
        RECT 655.950 819.600 658.050 820.050 ;
        RECT 673.950 819.600 676.050 820.050 ;
        RECT 712.950 819.600 715.050 820.050 ;
        RECT 655.950 818.400 715.050 819.600 ;
        RECT 655.950 817.950 658.050 818.400 ;
        RECT 673.950 817.950 676.050 818.400 ;
        RECT 712.950 817.950 715.050 818.400 ;
        RECT 13.950 814.950 16.050 817.050 ;
        RECT 40.950 816.600 43.050 817.050 ;
        RECT 91.950 816.600 94.050 817.050 ;
        RECT 124.950 816.600 127.050 817.050 ;
        RECT 40.950 815.400 78.600 816.600 ;
        RECT 40.950 814.950 43.050 815.400 ;
        RECT 14.400 811.050 15.600 814.950 ;
        RECT 16.950 813.600 19.050 814.050 ;
        RECT 28.950 813.600 31.050 814.050 ;
        RECT 16.950 812.400 31.050 813.600 ;
        RECT 16.950 811.950 19.050 812.400 ;
        RECT 28.950 811.950 31.050 812.400 ;
        RECT 64.950 813.600 67.050 814.050 ;
        RECT 73.950 813.600 76.050 814.050 ;
        RECT 64.950 812.400 76.050 813.600 ;
        RECT 64.950 811.950 67.050 812.400 ;
        RECT 73.950 811.950 76.050 812.400 ;
        RECT 77.400 811.050 78.600 815.400 ;
        RECT 91.950 815.400 127.050 816.600 ;
        RECT 91.950 814.950 94.050 815.400 ;
        RECT 124.950 814.950 127.050 815.400 ;
        RECT 142.950 816.600 145.050 817.050 ;
        RECT 193.950 816.600 196.050 817.050 ;
        RECT 142.950 815.400 196.050 816.600 ;
        RECT 142.950 814.950 145.050 815.400 ;
        RECT 193.950 814.950 196.050 815.400 ;
        RECT 202.950 816.600 205.050 817.050 ;
        RECT 211.950 816.600 214.050 817.050 ;
        RECT 232.950 816.600 235.050 817.050 ;
        RECT 202.950 815.400 214.050 816.600 ;
        RECT 202.950 814.950 205.050 815.400 ;
        RECT 211.950 814.950 214.050 815.400 ;
        RECT 227.400 815.400 235.050 816.600 ;
        RECT 88.950 813.600 91.050 814.050 ;
        RECT 100.950 813.600 103.050 814.050 ;
        RECT 88.950 812.400 103.050 813.600 ;
        RECT 88.950 811.950 91.050 812.400 ;
        RECT 100.950 811.950 103.050 812.400 ;
        RECT 109.950 813.600 112.050 814.050 ;
        RECT 121.950 813.600 124.050 814.050 ;
        RECT 109.950 812.400 124.050 813.600 ;
        RECT 109.950 811.950 112.050 812.400 ;
        RECT 121.950 811.950 124.050 812.400 ;
        RECT 127.950 813.600 130.050 814.050 ;
        RECT 136.950 813.600 139.050 814.050 ;
        RECT 139.950 813.600 142.050 814.050 ;
        RECT 127.950 812.400 142.050 813.600 ;
        RECT 127.950 811.950 130.050 812.400 ;
        RECT 136.950 811.950 139.050 812.400 ;
        RECT 139.950 811.950 142.050 812.400 ;
        RECT 145.950 813.600 148.050 814.050 ;
        RECT 160.950 813.600 163.050 814.050 ;
        RECT 145.950 812.400 163.050 813.600 ;
        RECT 145.950 811.950 148.050 812.400 ;
        RECT 160.950 811.950 163.050 812.400 ;
        RECT 172.950 813.600 175.050 814.050 ;
        RECT 187.950 813.600 190.050 814.050 ;
        RECT 172.950 812.400 190.050 813.600 ;
        RECT 172.950 811.950 175.050 812.400 ;
        RECT 187.950 811.950 190.050 812.400 ;
        RECT 13.950 808.950 16.050 811.050 ;
        RECT 52.950 810.600 55.050 811.050 ;
        RECT 61.950 810.600 64.050 811.050 ;
        RECT 52.950 809.400 64.050 810.600 ;
        RECT 52.950 808.950 55.050 809.400 ;
        RECT 61.950 808.950 64.050 809.400 ;
        RECT 76.950 808.950 79.050 811.050 ;
        RECT 82.950 810.600 85.050 811.050 ;
        RECT 100.950 810.600 103.050 811.050 ;
        RECT 80.400 809.400 103.050 810.600 ;
        RECT 7.950 807.600 10.050 808.050 ;
        RECT 10.950 807.600 13.050 808.050 ;
        RECT 80.400 807.600 81.600 809.400 ;
        RECT 82.950 808.950 85.050 809.400 ;
        RECT 100.950 808.950 103.050 809.400 ;
        RECT 175.950 810.600 178.050 811.050 ;
        RECT 184.950 810.600 187.050 811.050 ;
        RECT 175.950 809.400 187.050 810.600 ;
        RECT 175.950 808.950 178.050 809.400 ;
        RECT 184.950 808.950 187.050 809.400 ;
        RECT 7.950 806.400 81.600 807.600 ;
        RECT 172.950 807.600 175.050 808.050 ;
        RECT 187.950 807.600 190.050 808.050 ;
        RECT 172.950 806.400 190.050 807.600 ;
        RECT 227.400 807.600 228.600 815.400 ;
        RECT 232.950 814.950 235.050 815.400 ;
        RECT 238.950 816.600 241.050 817.050 ;
        RECT 244.950 816.600 247.050 817.050 ;
        RECT 238.950 815.400 247.050 816.600 ;
        RECT 238.950 814.950 241.050 815.400 ;
        RECT 244.950 814.950 247.050 815.400 ;
        RECT 248.400 814.050 249.600 817.950 ;
        RECT 250.950 816.600 253.050 817.050 ;
        RECT 292.950 816.600 295.050 817.050 ;
        RECT 250.950 815.400 295.050 816.600 ;
        RECT 250.950 814.950 253.050 815.400 ;
        RECT 292.950 814.950 295.050 815.400 ;
        RECT 370.950 816.600 373.050 817.050 ;
        RECT 382.950 816.600 385.050 817.050 ;
        RECT 370.950 815.400 385.050 816.600 ;
        RECT 370.950 814.950 373.050 815.400 ;
        RECT 382.950 814.950 385.050 815.400 ;
        RECT 388.950 816.600 391.050 817.050 ;
        RECT 400.950 816.600 403.050 817.050 ;
        RECT 388.950 815.400 403.050 816.600 ;
        RECT 388.950 814.950 391.050 815.400 ;
        RECT 400.950 814.950 403.050 815.400 ;
        RECT 463.950 816.600 466.050 817.050 ;
        RECT 490.950 816.600 493.050 817.050 ;
        RECT 505.950 816.600 508.050 817.050 ;
        RECT 463.950 815.400 508.050 816.600 ;
        RECT 463.950 814.950 466.050 815.400 ;
        RECT 490.950 814.950 493.050 815.400 ;
        RECT 505.950 814.950 508.050 815.400 ;
        RECT 514.950 816.600 517.050 817.050 ;
        RECT 529.950 816.600 532.050 817.050 ;
        RECT 514.950 815.400 532.050 816.600 ;
        RECT 514.950 814.950 517.050 815.400 ;
        RECT 529.950 814.950 532.050 815.400 ;
        RECT 538.950 816.600 541.050 817.050 ;
        RECT 559.950 816.600 562.050 817.050 ;
        RECT 538.950 815.400 562.050 816.600 ;
        RECT 538.950 814.950 541.050 815.400 ;
        RECT 559.950 814.950 562.050 815.400 ;
        RECT 571.950 816.600 574.050 817.050 ;
        RECT 583.950 816.600 586.050 817.050 ;
        RECT 613.950 816.600 616.050 817.050 ;
        RECT 571.950 815.400 579.600 816.600 ;
        RECT 571.950 814.950 574.050 815.400 ;
        RECT 578.400 814.050 579.600 815.400 ;
        RECT 583.950 815.400 616.050 816.600 ;
        RECT 583.950 814.950 586.050 815.400 ;
        RECT 613.950 814.950 616.050 815.400 ;
        RECT 622.950 816.600 625.050 817.050 ;
        RECT 688.950 816.600 691.050 817.050 ;
        RECT 622.950 815.400 691.050 816.600 ;
        RECT 622.950 814.950 625.050 815.400 ;
        RECT 688.950 814.950 691.050 815.400 ;
        RECT 769.950 816.600 772.050 817.050 ;
        RECT 775.950 816.600 778.050 817.050 ;
        RECT 769.950 815.400 778.050 816.600 ;
        RECT 769.950 814.950 772.050 815.400 ;
        RECT 775.950 814.950 778.050 815.400 ;
        RECT 793.950 816.600 796.050 817.050 ;
        RECT 820.950 816.600 823.050 817.050 ;
        RECT 793.950 815.400 823.050 816.600 ;
        RECT 793.950 814.950 796.050 815.400 ;
        RECT 820.950 814.950 823.050 815.400 ;
        RECT 823.950 816.600 826.050 817.050 ;
        RECT 859.950 816.600 862.050 817.050 ;
        RECT 823.950 815.400 862.050 816.600 ;
        RECT 823.950 814.950 826.050 815.400 ;
        RECT 859.950 814.950 862.050 815.400 ;
        RECT 229.950 811.950 232.050 814.050 ;
        RECT 247.950 811.950 250.050 814.050 ;
        RECT 265.950 813.600 268.050 814.050 ;
        RECT 271.950 813.600 274.050 814.050 ;
        RECT 265.950 812.400 274.050 813.600 ;
        RECT 265.950 811.950 268.050 812.400 ;
        RECT 271.950 811.950 274.050 812.400 ;
        RECT 304.950 813.600 307.050 814.050 ;
        RECT 310.950 813.600 313.050 814.050 ;
        RECT 304.950 812.400 313.050 813.600 ;
        RECT 304.950 811.950 307.050 812.400 ;
        RECT 310.950 811.950 313.050 812.400 ;
        RECT 394.950 813.600 397.050 814.050 ;
        RECT 427.950 813.600 430.050 814.050 ;
        RECT 433.950 813.600 436.050 814.050 ;
        RECT 394.950 812.400 402.600 813.600 ;
        RECT 394.950 811.950 397.050 812.400 ;
        RECT 230.400 810.600 231.600 811.950 ;
        RECT 268.950 810.600 271.050 811.050 ;
        RECT 230.400 809.400 271.050 810.600 ;
        RECT 268.950 808.950 271.050 809.400 ;
        RECT 295.950 810.600 298.050 811.050 ;
        RECT 307.950 810.600 310.050 811.050 ;
        RECT 295.950 809.400 310.050 810.600 ;
        RECT 295.950 808.950 298.050 809.400 ;
        RECT 307.950 808.950 310.050 809.400 ;
        RECT 313.950 810.600 316.050 811.050 ;
        RECT 391.950 810.600 394.050 811.050 ;
        RECT 313.950 809.400 394.050 810.600 ;
        RECT 313.950 808.950 316.050 809.400 ;
        RECT 391.950 808.950 394.050 809.400 ;
        RECT 397.950 808.950 400.050 811.050 ;
        RECT 401.400 810.600 402.600 812.400 ;
        RECT 427.950 812.400 436.050 813.600 ;
        RECT 427.950 811.950 430.050 812.400 ;
        RECT 433.950 811.950 436.050 812.400 ;
        RECT 469.950 813.600 472.050 814.050 ;
        RECT 475.950 813.600 478.050 814.050 ;
        RECT 469.950 812.400 478.050 813.600 ;
        RECT 469.950 811.950 472.050 812.400 ;
        RECT 475.950 811.950 478.050 812.400 ;
        RECT 493.950 811.950 496.050 814.050 ;
        RECT 499.950 813.600 502.050 814.050 ;
        RECT 511.950 813.600 514.050 814.050 ;
        RECT 499.950 812.400 514.050 813.600 ;
        RECT 499.950 811.950 502.050 812.400 ;
        RECT 511.950 811.950 514.050 812.400 ;
        RECT 535.950 813.600 538.050 814.050 ;
        RECT 553.950 813.600 556.050 814.050 ;
        RECT 535.950 812.400 556.050 813.600 ;
        RECT 535.950 811.950 538.050 812.400 ;
        RECT 553.950 811.950 556.050 812.400 ;
        RECT 556.950 813.600 559.050 814.050 ;
        RECT 559.950 813.600 562.050 814.050 ;
        RECT 556.950 812.400 562.050 813.600 ;
        RECT 556.950 811.950 559.050 812.400 ;
        RECT 559.950 811.950 562.050 812.400 ;
        RECT 568.950 813.600 571.050 814.050 ;
        RECT 574.950 813.600 577.050 814.050 ;
        RECT 568.950 812.400 577.050 813.600 ;
        RECT 568.950 811.950 571.050 812.400 ;
        RECT 574.950 811.950 577.050 812.400 ;
        RECT 577.950 811.950 580.050 814.050 ;
        RECT 616.950 813.600 619.050 814.050 ;
        RECT 634.950 813.600 637.050 814.050 ;
        RECT 616.950 812.400 637.050 813.600 ;
        RECT 616.950 811.950 619.050 812.400 ;
        RECT 634.950 811.950 637.050 812.400 ;
        RECT 652.950 813.600 655.050 814.050 ;
        RECT 670.950 813.600 673.050 814.050 ;
        RECT 652.950 812.400 673.050 813.600 ;
        RECT 652.950 811.950 655.050 812.400 ;
        RECT 670.950 811.950 673.050 812.400 ;
        RECT 676.950 813.600 679.050 814.050 ;
        RECT 694.950 813.600 697.050 814.050 ;
        RECT 676.950 812.400 697.050 813.600 ;
        RECT 676.950 811.950 679.050 812.400 ;
        RECT 694.950 811.950 697.050 812.400 ;
        RECT 790.950 813.600 793.050 814.050 ;
        RECT 841.950 813.600 844.050 814.050 ;
        RECT 790.950 812.400 844.050 813.600 ;
        RECT 790.950 811.950 793.050 812.400 ;
        RECT 841.950 811.950 844.050 812.400 ;
        RECT 412.950 810.600 415.050 811.050 ;
        RECT 401.400 809.400 415.050 810.600 ;
        RECT 412.950 808.950 415.050 809.400 ;
        RECT 454.950 810.600 457.050 811.050 ;
        RECT 466.950 810.600 469.050 811.050 ;
        RECT 454.950 809.400 469.050 810.600 ;
        RECT 494.400 810.600 495.600 811.950 ;
        RECT 514.950 810.600 517.050 811.050 ;
        RECT 550.950 810.600 553.050 811.050 ;
        RECT 494.400 809.400 553.050 810.600 ;
        RECT 454.950 808.950 457.050 809.400 ;
        RECT 466.950 808.950 469.050 809.400 ;
        RECT 514.950 808.950 517.050 809.400 ;
        RECT 550.950 808.950 553.050 809.400 ;
        RECT 556.950 808.950 559.050 811.050 ;
        RECT 560.400 810.600 561.600 811.950 ;
        RECT 580.950 810.600 583.050 811.050 ;
        RECT 560.400 809.400 583.050 810.600 ;
        RECT 580.950 808.950 583.050 809.400 ;
        RECT 583.950 810.600 586.050 811.050 ;
        RECT 622.950 810.600 625.050 811.050 ;
        RECT 583.950 809.400 625.050 810.600 ;
        RECT 583.950 808.950 586.050 809.400 ;
        RECT 622.950 808.950 625.050 809.400 ;
        RECT 637.950 810.600 640.050 811.050 ;
        RECT 655.950 810.600 658.050 811.050 ;
        RECT 637.950 809.400 658.050 810.600 ;
        RECT 637.950 808.950 640.050 809.400 ;
        RECT 655.950 808.950 658.050 809.400 ;
        RECT 661.950 810.600 664.050 811.050 ;
        RECT 676.950 810.600 679.050 811.050 ;
        RECT 661.950 809.400 679.050 810.600 ;
        RECT 661.950 808.950 664.050 809.400 ;
        RECT 676.950 808.950 679.050 809.400 ;
        RECT 682.950 810.600 685.050 811.050 ;
        RECT 709.950 810.600 712.050 811.050 ;
        RECT 682.950 809.400 712.050 810.600 ;
        RECT 682.950 808.950 685.050 809.400 ;
        RECT 709.950 808.950 712.050 809.400 ;
        RECT 229.950 807.600 232.050 808.050 ;
        RECT 227.400 806.400 232.050 807.600 ;
        RECT 7.950 805.950 10.050 806.400 ;
        RECT 10.950 805.950 13.050 806.400 ;
        RECT 172.950 805.950 175.050 806.400 ;
        RECT 187.950 805.950 190.050 806.400 ;
        RECT 229.950 805.950 232.050 806.400 ;
        RECT 301.950 807.600 304.050 808.050 ;
        RECT 313.950 807.600 316.050 808.050 ;
        RECT 301.950 806.400 316.050 807.600 ;
        RECT 301.950 805.950 304.050 806.400 ;
        RECT 313.950 805.950 316.050 806.400 ;
        RECT 382.950 807.600 385.050 808.050 ;
        RECT 398.400 807.600 399.600 808.950 ;
        RECT 382.950 806.400 399.600 807.600 ;
        RECT 472.950 807.600 475.050 808.050 ;
        RECT 499.950 807.600 502.050 808.050 ;
        RECT 472.950 806.400 502.050 807.600 ;
        RECT 557.400 807.600 558.600 808.950 ;
        RECT 565.950 807.600 568.050 808.050 ;
        RECT 557.400 806.400 568.050 807.600 ;
        RECT 382.950 805.950 385.050 806.400 ;
        RECT 472.950 805.950 475.050 806.400 ;
        RECT 499.950 805.950 502.050 806.400 ;
        RECT 565.950 805.950 568.050 806.400 ;
        RECT 598.950 807.600 601.050 808.050 ;
        RECT 619.950 807.600 622.050 808.050 ;
        RECT 598.950 806.400 622.050 807.600 ;
        RECT 598.950 805.950 601.050 806.400 ;
        RECT 619.950 805.950 622.050 806.400 ;
        RECT 61.950 804.600 64.050 805.050 ;
        RECT 67.950 804.600 70.050 805.050 ;
        RECT 61.950 803.400 70.050 804.600 ;
        RECT 61.950 802.950 64.050 803.400 ;
        RECT 67.950 802.950 70.050 803.400 ;
        RECT 73.950 804.600 76.050 805.050 ;
        RECT 106.950 804.600 109.050 805.050 ;
        RECT 73.950 803.400 109.050 804.600 ;
        RECT 73.950 802.950 76.050 803.400 ;
        RECT 106.950 802.950 109.050 803.400 ;
        RECT 607.950 804.600 610.050 805.050 ;
        RECT 610.950 804.600 613.050 805.050 ;
        RECT 631.950 804.600 634.050 805.050 ;
        RECT 670.950 804.600 673.050 805.050 ;
        RECT 607.950 803.400 673.050 804.600 ;
        RECT 607.950 802.950 610.050 803.400 ;
        RECT 610.950 802.950 613.050 803.400 ;
        RECT 631.950 802.950 634.050 803.400 ;
        RECT 670.950 802.950 673.050 803.400 ;
        RECT 718.950 804.600 721.050 805.050 ;
        RECT 766.950 804.600 769.050 805.050 ;
        RECT 817.950 804.600 820.050 805.050 ;
        RECT 718.950 803.400 820.050 804.600 ;
        RECT 718.950 802.950 721.050 803.400 ;
        RECT 766.950 802.950 769.050 803.400 ;
        RECT 817.950 802.950 820.050 803.400 ;
        RECT 58.950 801.600 61.050 802.050 ;
        RECT 70.950 801.600 73.050 802.050 ;
        RECT 58.950 800.400 73.050 801.600 ;
        RECT 58.950 799.950 61.050 800.400 ;
        RECT 70.950 799.950 73.050 800.400 ;
        RECT 640.950 801.600 643.050 802.050 ;
        RECT 724.950 801.600 727.050 802.050 ;
        RECT 640.950 800.400 727.050 801.600 ;
        RECT 640.950 799.950 643.050 800.400 ;
        RECT 724.950 799.950 727.050 800.400 ;
        RECT 7.950 798.600 10.050 799.050 ;
        RECT 13.950 798.600 16.050 799.050 ;
        RECT 7.950 797.400 16.050 798.600 ;
        RECT 7.950 796.950 10.050 797.400 ;
        RECT 13.950 796.950 16.050 797.400 ;
        RECT 325.950 795.600 328.050 796.050 ;
        RECT 349.950 795.600 352.050 796.050 ;
        RECT 325.950 794.400 352.050 795.600 ;
        RECT 325.950 793.950 328.050 794.400 ;
        RECT 349.950 793.950 352.050 794.400 ;
        RECT 232.950 792.600 235.050 793.050 ;
        RECT 238.950 792.600 241.050 793.050 ;
        RECT 232.950 791.400 241.050 792.600 ;
        RECT 232.950 790.950 235.050 791.400 ;
        RECT 238.950 790.950 241.050 791.400 ;
        RECT 523.950 789.600 526.050 790.050 ;
        RECT 595.950 789.600 598.050 790.050 ;
        RECT 700.950 789.600 703.050 790.050 ;
        RECT 523.950 788.400 703.050 789.600 ;
        RECT 523.950 787.950 526.050 788.400 ;
        RECT 595.950 787.950 598.050 788.400 ;
        RECT 700.950 787.950 703.050 788.400 ;
        RECT 25.950 786.600 28.050 787.050 ;
        RECT 34.950 786.600 37.050 787.050 ;
        RECT 25.950 785.400 37.050 786.600 ;
        RECT 25.950 784.950 28.050 785.400 ;
        RECT 34.950 784.950 37.050 785.400 ;
        RECT 22.950 783.600 25.050 784.050 ;
        RECT 34.950 783.600 37.050 784.050 ;
        RECT 91.950 783.600 94.050 784.050 ;
        RECT 22.950 782.400 94.050 783.600 ;
        RECT 22.950 781.950 25.050 782.400 ;
        RECT 34.950 781.950 37.050 782.400 ;
        RECT 91.950 781.950 94.050 782.400 ;
        RECT 301.950 783.600 304.050 784.050 ;
        RECT 328.950 783.600 331.050 784.050 ;
        RECT 301.950 782.400 331.050 783.600 ;
        RECT 301.950 781.950 304.050 782.400 ;
        RECT 328.950 781.950 331.050 782.400 ;
        RECT 532.950 783.600 535.050 784.050 ;
        RECT 661.950 783.600 664.050 784.050 ;
        RECT 532.950 782.400 664.050 783.600 ;
        RECT 532.950 781.950 535.050 782.400 ;
        RECT 661.950 781.950 664.050 782.400 ;
        RECT 79.950 780.600 82.050 781.050 ;
        RECT 148.950 780.600 151.050 781.050 ;
        RECT 79.950 779.400 151.050 780.600 ;
        RECT 79.950 778.950 82.050 779.400 ;
        RECT 148.950 778.950 151.050 779.400 ;
        RECT 298.950 780.600 301.050 781.050 ;
        RECT 304.950 780.600 307.050 781.050 ;
        RECT 298.950 779.400 307.050 780.600 ;
        RECT 298.950 778.950 301.050 779.400 ;
        RECT 304.950 778.950 307.050 779.400 ;
        RECT 313.950 780.600 316.050 781.050 ;
        RECT 331.950 780.600 334.050 781.050 ;
        RECT 358.950 780.600 361.050 781.050 ;
        RECT 382.950 780.600 385.050 781.050 ;
        RECT 313.950 779.400 385.050 780.600 ;
        RECT 313.950 778.950 316.050 779.400 ;
        RECT 331.950 778.950 334.050 779.400 ;
        RECT 358.950 778.950 361.050 779.400 ;
        RECT 382.950 778.950 385.050 779.400 ;
        RECT 544.950 780.600 547.050 781.050 ;
        RECT 595.950 780.600 598.050 781.050 ;
        RECT 685.950 780.600 688.050 781.050 ;
        RECT 544.950 779.400 598.050 780.600 ;
        RECT 544.950 778.950 547.050 779.400 ;
        RECT 595.950 778.950 598.050 779.400 ;
        RECT 599.400 779.400 688.050 780.600 ;
        RECT 22.950 777.600 25.050 778.050 ;
        RECT 14.400 776.400 25.050 777.600 ;
        RECT 14.400 775.050 15.600 776.400 ;
        RECT 22.950 775.950 25.050 776.400 ;
        RECT 28.950 777.600 31.050 778.050 ;
        RECT 40.950 777.600 43.050 778.050 ;
        RECT 28.950 776.400 43.050 777.600 ;
        RECT 28.950 775.950 31.050 776.400 ;
        RECT 40.950 775.950 43.050 776.400 ;
        RECT 46.950 777.600 49.050 778.050 ;
        RECT 67.950 777.600 70.050 778.050 ;
        RECT 46.950 776.400 70.050 777.600 ;
        RECT 46.950 775.950 49.050 776.400 ;
        RECT 67.950 775.950 70.050 776.400 ;
        RECT 73.950 777.600 76.050 778.050 ;
        RECT 91.950 777.600 94.050 778.050 ;
        RECT 73.950 776.400 94.050 777.600 ;
        RECT 73.950 775.950 76.050 776.400 ;
        RECT 91.950 775.950 94.050 776.400 ;
        RECT 118.950 777.600 121.050 778.050 ;
        RECT 151.950 777.600 154.050 778.050 ;
        RECT 118.950 776.400 154.050 777.600 ;
        RECT 118.950 775.950 121.050 776.400 ;
        RECT 134.400 775.050 135.600 776.400 ;
        RECT 151.950 775.950 154.050 776.400 ;
        RECT 157.950 777.600 160.050 778.050 ;
        RECT 193.950 777.600 196.050 778.050 ;
        RECT 157.950 776.400 196.050 777.600 ;
        RECT 157.950 775.950 160.050 776.400 ;
        RECT 193.950 775.950 196.050 776.400 ;
        RECT 253.950 777.600 256.050 778.050 ;
        RECT 283.950 777.600 286.050 778.050 ;
        RECT 253.950 776.400 286.050 777.600 ;
        RECT 253.950 775.950 256.050 776.400 ;
        RECT 283.950 775.950 286.050 776.400 ;
        RECT 286.950 777.600 289.050 778.050 ;
        RECT 307.950 777.600 310.050 778.050 ;
        RECT 346.950 777.600 349.050 778.050 ;
        RECT 286.950 776.400 349.050 777.600 ;
        RECT 286.950 775.950 289.050 776.400 ;
        RECT 307.950 775.950 310.050 776.400 ;
        RECT 346.950 775.950 349.050 776.400 ;
        RECT 352.950 777.600 355.050 778.050 ;
        RECT 370.950 777.600 373.050 778.050 ;
        RECT 352.950 776.400 373.050 777.600 ;
        RECT 352.950 775.950 355.050 776.400 ;
        RECT 370.950 775.950 373.050 776.400 ;
        RECT 421.950 777.600 424.050 778.050 ;
        RECT 532.950 777.600 535.050 778.050 ;
        RECT 421.950 776.400 535.050 777.600 ;
        RECT 421.950 775.950 424.050 776.400 ;
        RECT 532.950 775.950 535.050 776.400 ;
        RECT 553.950 777.600 556.050 778.050 ;
        RECT 565.950 777.600 568.050 778.050 ;
        RECT 553.950 776.400 568.050 777.600 ;
        RECT 553.950 775.950 556.050 776.400 ;
        RECT 565.950 775.950 568.050 776.400 ;
        RECT 586.950 777.600 589.050 778.050 ;
        RECT 599.400 777.600 600.600 779.400 ;
        RECT 685.950 778.950 688.050 779.400 ;
        RECT 793.950 780.600 796.050 781.050 ;
        RECT 802.950 780.600 805.050 781.050 ;
        RECT 856.950 780.600 859.050 781.050 ;
        RECT 793.950 779.400 805.050 780.600 ;
        RECT 793.950 778.950 796.050 779.400 ;
        RECT 802.950 778.950 805.050 779.400 ;
        RECT 854.400 779.400 859.050 780.600 ;
        RECT 586.950 776.400 600.600 777.600 ;
        RECT 586.950 775.950 589.050 776.400 ;
        RECT 604.950 775.950 607.050 778.050 ;
        RECT 637.950 777.600 640.050 778.050 ;
        RECT 608.400 776.400 640.050 777.600 ;
        RECT 13.950 772.950 16.050 775.050 ;
        RECT 16.950 774.600 19.050 775.050 ;
        RECT 28.950 774.600 31.050 775.050 ;
        RECT 16.950 773.400 31.050 774.600 ;
        RECT 16.950 772.950 19.050 773.400 ;
        RECT 28.950 772.950 31.050 773.400 ;
        RECT 52.950 774.600 55.050 775.050 ;
        RECT 64.950 774.600 67.050 775.050 ;
        RECT 52.950 773.400 67.050 774.600 ;
        RECT 52.950 772.950 55.050 773.400 ;
        RECT 64.950 772.950 67.050 773.400 ;
        RECT 70.950 774.600 73.050 775.050 ;
        RECT 85.950 774.600 88.050 775.050 ;
        RECT 70.950 773.400 88.050 774.600 ;
        RECT 70.950 772.950 73.050 773.400 ;
        RECT 85.950 772.950 88.050 773.400 ;
        RECT 112.950 774.600 115.050 775.050 ;
        RECT 130.950 774.600 133.050 775.050 ;
        RECT 112.950 773.400 133.050 774.600 ;
        RECT 112.950 772.950 115.050 773.400 ;
        RECT 130.950 772.950 133.050 773.400 ;
        RECT 133.950 772.950 136.050 775.050 ;
        RECT 160.950 774.600 163.050 775.050 ;
        RECT 172.950 774.600 175.050 775.050 ;
        RECT 160.950 773.400 175.050 774.600 ;
        RECT 160.950 772.950 163.050 773.400 ;
        RECT 172.950 772.950 175.050 773.400 ;
        RECT 202.950 774.600 205.050 775.050 ;
        RECT 211.950 774.600 214.050 775.050 ;
        RECT 202.950 773.400 214.050 774.600 ;
        RECT 202.950 772.950 205.050 773.400 ;
        RECT 211.950 772.950 214.050 773.400 ;
        RECT 217.950 774.600 220.050 775.050 ;
        RECT 226.950 774.600 229.050 775.050 ;
        RECT 217.950 773.400 229.050 774.600 ;
        RECT 217.950 772.950 220.050 773.400 ;
        RECT 226.950 772.950 229.050 773.400 ;
        RECT 247.950 774.600 250.050 775.050 ;
        RECT 262.950 774.600 265.050 775.050 ;
        RECT 247.950 773.400 265.050 774.600 ;
        RECT 247.950 772.950 250.050 773.400 ;
        RECT 262.950 772.950 265.050 773.400 ;
        RECT 268.950 774.600 271.050 775.050 ;
        RECT 274.950 774.600 277.050 775.050 ;
        RECT 268.950 773.400 277.050 774.600 ;
        RECT 268.950 772.950 271.050 773.400 ;
        RECT 274.950 772.950 277.050 773.400 ;
        RECT 319.950 774.600 322.050 775.050 ;
        RECT 328.950 774.600 331.050 775.050 ;
        RECT 319.950 773.400 331.050 774.600 ;
        RECT 319.950 772.950 322.050 773.400 ;
        RECT 328.950 772.950 331.050 773.400 ;
        RECT 340.950 774.600 343.050 775.050 ;
        RECT 349.950 774.600 352.050 775.050 ;
        RECT 376.950 774.600 379.050 775.050 ;
        RECT 340.950 773.400 379.050 774.600 ;
        RECT 340.950 772.950 343.050 773.400 ;
        RECT 349.950 772.950 352.050 773.400 ;
        RECT 376.950 772.950 379.050 773.400 ;
        RECT 409.950 774.600 412.050 775.050 ;
        RECT 433.950 774.600 436.050 775.050 ;
        RECT 409.950 773.400 436.050 774.600 ;
        RECT 409.950 772.950 412.050 773.400 ;
        RECT 433.950 772.950 436.050 773.400 ;
        RECT 568.950 774.600 571.050 775.050 ;
        RECT 583.950 774.600 586.050 775.050 ;
        RECT 568.950 773.400 586.050 774.600 ;
        RECT 568.950 772.950 571.050 773.400 ;
        RECT 583.950 772.950 586.050 773.400 ;
        RECT 598.950 774.600 601.050 775.050 ;
        RECT 605.400 774.600 606.600 775.950 ;
        RECT 608.400 775.050 609.600 776.400 ;
        RECT 637.950 775.950 640.050 776.400 ;
        RECT 598.950 773.400 606.600 774.600 ;
        RECT 598.950 772.950 601.050 773.400 ;
        RECT 607.950 772.950 610.050 775.050 ;
        RECT 631.950 774.600 634.050 775.050 ;
        RECT 643.950 774.600 646.050 775.050 ;
        RECT 649.950 774.600 652.050 775.050 ;
        RECT 631.950 773.400 652.050 774.600 ;
        RECT 631.950 772.950 634.050 773.400 ;
        RECT 643.950 772.950 646.050 773.400 ;
        RECT 649.950 772.950 652.050 773.400 ;
        RECT 670.950 774.600 673.050 775.050 ;
        RECT 694.950 774.600 697.050 775.050 ;
        RECT 703.950 774.600 706.050 775.050 ;
        RECT 670.950 773.400 706.050 774.600 ;
        RECT 670.950 772.950 673.050 773.400 ;
        RECT 694.950 772.950 697.050 773.400 ;
        RECT 703.950 772.950 706.050 773.400 ;
        RECT 709.950 772.950 712.050 775.050 ;
        RECT 781.950 774.600 784.050 775.050 ;
        RECT 802.950 774.600 805.050 775.050 ;
        RECT 817.950 774.600 820.050 775.050 ;
        RECT 728.400 773.400 784.050 774.600 ;
        RECT 61.950 771.600 64.050 772.050 ;
        RECT 76.950 771.600 79.050 772.050 ;
        RECT 61.950 770.400 79.050 771.600 ;
        RECT 61.950 769.950 64.050 770.400 ;
        RECT 76.950 769.950 79.050 770.400 ;
        RECT 109.950 771.600 112.050 772.050 ;
        RECT 121.950 771.600 124.050 772.050 ;
        RECT 109.950 770.400 124.050 771.600 ;
        RECT 109.950 769.950 112.050 770.400 ;
        RECT 121.950 769.950 124.050 770.400 ;
        RECT 127.950 771.600 130.050 772.050 ;
        RECT 136.950 771.600 139.050 772.050 ;
        RECT 127.950 770.400 139.050 771.600 ;
        RECT 127.950 769.950 130.050 770.400 ;
        RECT 136.950 769.950 139.050 770.400 ;
        RECT 199.950 771.600 202.050 772.050 ;
        RECT 214.950 771.600 217.050 772.050 ;
        RECT 199.950 770.400 217.050 771.600 ;
        RECT 199.950 769.950 202.050 770.400 ;
        RECT 214.950 769.950 217.050 770.400 ;
        RECT 229.950 771.600 232.050 772.050 ;
        RECT 250.950 771.600 253.050 772.050 ;
        RECT 229.950 770.400 253.050 771.600 ;
        RECT 229.950 769.950 232.050 770.400 ;
        RECT 250.950 769.950 253.050 770.400 ;
        RECT 256.950 771.600 259.050 772.050 ;
        RECT 262.950 771.600 265.050 772.050 ;
        RECT 289.950 771.600 292.050 772.050 ;
        RECT 310.950 771.600 313.050 772.050 ;
        RECT 256.950 770.400 313.050 771.600 ;
        RECT 256.950 769.950 259.050 770.400 ;
        RECT 262.950 769.950 265.050 770.400 ;
        RECT 289.950 769.950 292.050 770.400 ;
        RECT 310.950 769.950 313.050 770.400 ;
        RECT 361.950 771.600 364.050 772.050 ;
        RECT 367.950 771.600 370.050 772.050 ;
        RECT 361.950 770.400 370.050 771.600 ;
        RECT 361.950 769.950 364.050 770.400 ;
        RECT 367.950 769.950 370.050 770.400 ;
        RECT 382.950 771.600 385.050 772.050 ;
        RECT 430.950 771.600 433.050 772.050 ;
        RECT 382.950 770.400 433.050 771.600 ;
        RECT 434.400 771.600 435.600 772.950 ;
        RECT 448.950 771.600 451.050 772.050 ;
        RECT 434.400 770.400 451.050 771.600 ;
        RECT 382.950 769.950 385.050 770.400 ;
        RECT 430.950 769.950 433.050 770.400 ;
        RECT 448.950 769.950 451.050 770.400 ;
        RECT 454.950 771.600 457.050 772.050 ;
        RECT 466.950 771.600 469.050 772.050 ;
        RECT 547.950 771.600 550.050 772.050 ;
        RECT 628.950 771.600 631.050 772.050 ;
        RECT 454.950 770.400 550.050 771.600 ;
        RECT 454.950 769.950 457.050 770.400 ;
        RECT 466.950 769.950 469.050 770.400 ;
        RECT 494.400 769.050 495.600 770.400 ;
        RECT 547.950 769.950 550.050 770.400 ;
        RECT 602.400 770.400 631.050 771.600 ;
        RECT 602.400 769.050 603.600 770.400 ;
        RECT 628.950 769.950 631.050 770.400 ;
        RECT 637.950 771.600 640.050 772.050 ;
        RECT 652.950 771.600 655.050 772.050 ;
        RECT 637.950 770.400 655.050 771.600 ;
        RECT 637.950 769.950 640.050 770.400 ;
        RECT 652.950 769.950 655.050 770.400 ;
        RECT 655.950 771.600 658.050 772.050 ;
        RECT 679.950 771.600 682.050 772.050 ;
        RECT 688.950 771.600 691.050 772.050 ;
        RECT 655.950 770.400 691.050 771.600 ;
        RECT 655.950 769.950 658.050 770.400 ;
        RECT 679.950 769.950 682.050 770.400 ;
        RECT 688.950 769.950 691.050 770.400 ;
        RECT 697.950 771.600 700.050 772.050 ;
        RECT 710.400 771.600 711.600 772.950 ;
        RECT 697.950 770.400 711.600 771.600 ;
        RECT 724.950 771.600 727.050 772.050 ;
        RECT 728.400 771.600 729.600 773.400 ;
        RECT 781.950 772.950 784.050 773.400 ;
        RECT 785.400 773.400 820.050 774.600 ;
        RECT 724.950 770.400 729.600 771.600 ;
        RECT 730.950 771.600 733.050 772.050 ;
        RECT 785.400 771.600 786.600 773.400 ;
        RECT 802.950 772.950 805.050 773.400 ;
        RECT 817.950 772.950 820.050 773.400 ;
        RECT 854.400 772.050 855.600 779.400 ;
        RECT 856.950 778.950 859.050 779.400 ;
        RECT 859.950 780.600 862.050 781.050 ;
        RECT 859.950 779.400 864.600 780.600 ;
        RECT 859.950 778.950 862.050 779.400 ;
        RECT 856.950 774.600 859.050 775.050 ;
        RECT 863.400 774.600 864.600 779.400 ;
        RECT 856.950 773.400 864.600 774.600 ;
        RECT 856.950 772.950 859.050 773.400 ;
        RECT 820.950 771.600 823.050 772.050 ;
        RECT 730.950 770.400 786.600 771.600 ;
        RECT 818.400 770.400 823.050 771.600 ;
        RECT 697.950 769.950 700.050 770.400 ;
        RECT 724.950 769.950 727.050 770.400 ;
        RECT 730.950 769.950 733.050 770.400 ;
        RECT 818.400 769.050 819.600 770.400 ;
        RECT 820.950 769.950 823.050 770.400 ;
        RECT 853.950 769.950 856.050 772.050 ;
        RECT 19.950 768.600 22.050 769.050 ;
        RECT 31.950 768.600 34.050 769.050 ;
        RECT 19.950 767.400 34.050 768.600 ;
        RECT 19.950 766.950 22.050 767.400 ;
        RECT 31.950 766.950 34.050 767.400 ;
        RECT 79.950 768.600 82.050 769.050 ;
        RECT 88.950 768.600 91.050 769.050 ;
        RECT 79.950 767.400 91.050 768.600 ;
        RECT 79.950 766.950 82.050 767.400 ;
        RECT 88.950 766.950 91.050 767.400 ;
        RECT 115.950 768.600 118.050 769.050 ;
        RECT 127.950 768.600 130.050 769.050 ;
        RECT 115.950 767.400 130.050 768.600 ;
        RECT 115.950 766.950 118.050 767.400 ;
        RECT 127.950 766.950 130.050 767.400 ;
        RECT 133.950 768.600 136.050 769.050 ;
        RECT 169.950 768.600 172.050 769.050 ;
        RECT 196.950 768.600 199.050 769.050 ;
        RECT 202.950 768.600 205.050 769.050 ;
        RECT 133.950 767.400 205.050 768.600 ;
        RECT 133.950 766.950 136.050 767.400 ;
        RECT 169.950 766.950 172.050 767.400 ;
        RECT 196.950 766.950 199.050 767.400 ;
        RECT 202.950 766.950 205.050 767.400 ;
        RECT 253.950 768.600 256.050 769.050 ;
        RECT 265.950 768.600 268.050 769.050 ;
        RECT 280.950 768.600 283.050 769.050 ;
        RECT 253.950 767.400 283.050 768.600 ;
        RECT 253.950 766.950 256.050 767.400 ;
        RECT 265.950 766.950 268.050 767.400 ;
        RECT 280.950 766.950 283.050 767.400 ;
        RECT 355.950 768.600 358.050 769.050 ;
        RECT 373.950 768.600 376.050 769.050 ;
        RECT 382.950 768.600 385.050 769.050 ;
        RECT 355.950 767.400 385.050 768.600 ;
        RECT 355.950 766.950 358.050 767.400 ;
        RECT 373.950 766.950 376.050 767.400 ;
        RECT 382.950 766.950 385.050 767.400 ;
        RECT 391.950 768.600 394.050 769.050 ;
        RECT 400.950 768.600 403.050 769.050 ;
        RECT 406.950 768.600 409.050 769.050 ;
        RECT 391.950 767.400 409.050 768.600 ;
        RECT 391.950 766.950 394.050 767.400 ;
        RECT 400.950 766.950 403.050 767.400 ;
        RECT 406.950 766.950 409.050 767.400 ;
        RECT 436.950 768.600 439.050 769.050 ;
        RECT 469.950 768.600 472.050 769.050 ;
        RECT 436.950 767.400 472.050 768.600 ;
        RECT 436.950 766.950 439.050 767.400 ;
        RECT 469.950 766.950 472.050 767.400 ;
        RECT 493.950 766.950 496.050 769.050 ;
        RECT 505.950 768.600 508.050 769.050 ;
        RECT 526.950 768.600 529.050 769.050 ;
        RECT 532.950 768.600 535.050 769.050 ;
        RECT 505.950 767.400 535.050 768.600 ;
        RECT 505.950 766.950 508.050 767.400 ;
        RECT 526.950 766.950 529.050 767.400 ;
        RECT 532.950 766.950 535.050 767.400 ;
        RECT 601.950 766.950 604.050 769.050 ;
        RECT 625.950 768.600 628.050 769.050 ;
        RECT 646.950 768.600 649.050 769.050 ;
        RECT 667.950 768.600 670.050 769.050 ;
        RECT 625.950 767.400 670.050 768.600 ;
        RECT 625.950 766.950 628.050 767.400 ;
        RECT 646.950 766.950 649.050 767.400 ;
        RECT 667.950 766.950 670.050 767.400 ;
        RECT 691.950 768.600 694.050 769.050 ;
        RECT 706.950 768.600 709.050 769.050 ;
        RECT 712.950 768.600 715.050 769.050 ;
        RECT 691.950 767.400 715.050 768.600 ;
        RECT 691.950 766.950 694.050 767.400 ;
        RECT 706.950 766.950 709.050 767.400 ;
        RECT 712.950 766.950 715.050 767.400 ;
        RECT 817.950 766.950 820.050 769.050 ;
        RECT 820.950 768.600 823.050 769.050 ;
        RECT 826.950 768.600 829.050 769.050 ;
        RECT 820.950 767.400 829.050 768.600 ;
        RECT 820.950 766.950 823.050 767.400 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 73.950 765.600 76.050 766.050 ;
        RECT 109.950 765.600 112.050 766.050 ;
        RECT 73.950 764.400 112.050 765.600 ;
        RECT 73.950 763.950 76.050 764.400 ;
        RECT 109.950 763.950 112.050 764.400 ;
        RECT 112.950 765.600 115.050 766.050 ;
        RECT 154.950 765.600 157.050 766.050 ;
        RECT 169.950 765.600 172.050 766.050 ;
        RECT 190.950 765.600 193.050 766.050 ;
        RECT 112.950 764.400 193.050 765.600 ;
        RECT 112.950 763.950 115.050 764.400 ;
        RECT 154.950 763.950 157.050 764.400 ;
        RECT 169.950 763.950 172.050 764.400 ;
        RECT 190.950 763.950 193.050 764.400 ;
        RECT 316.950 765.600 319.050 766.050 ;
        RECT 322.950 765.600 325.050 766.050 ;
        RECT 454.950 765.600 457.050 766.050 ;
        RECT 316.950 764.400 457.050 765.600 ;
        RECT 316.950 763.950 319.050 764.400 ;
        RECT 322.950 763.950 325.050 764.400 ;
        RECT 454.950 763.950 457.050 764.400 ;
        RECT 556.950 765.600 559.050 766.050 ;
        RECT 586.950 765.600 589.050 766.050 ;
        RECT 724.950 765.600 727.050 766.050 ;
        RECT 556.950 764.400 727.050 765.600 ;
        RECT 556.950 763.950 559.050 764.400 ;
        RECT 586.950 763.950 589.050 764.400 ;
        RECT 724.950 763.950 727.050 764.400 ;
        RECT 778.950 765.600 781.050 766.050 ;
        RECT 799.950 765.600 802.050 766.050 ;
        RECT 778.950 764.400 802.050 765.600 ;
        RECT 778.950 763.950 781.050 764.400 ;
        RECT 799.950 763.950 802.050 764.400 ;
        RECT 823.950 765.600 826.050 766.050 ;
        RECT 862.950 765.600 865.050 766.050 ;
        RECT 823.950 764.400 865.050 765.600 ;
        RECT 823.950 763.950 826.050 764.400 ;
        RECT 862.950 763.950 865.050 764.400 ;
        RECT 166.950 762.600 169.050 763.050 ;
        RECT 172.950 762.600 175.050 763.050 ;
        RECT 166.950 761.400 175.050 762.600 ;
        RECT 166.950 760.950 169.050 761.400 ;
        RECT 172.950 760.950 175.050 761.400 ;
        RECT 598.950 762.600 601.050 763.050 ;
        RECT 658.950 762.600 661.050 763.050 ;
        RECT 727.950 762.600 730.050 763.050 ;
        RECT 598.950 761.400 730.050 762.600 ;
        RECT 598.950 760.950 601.050 761.400 ;
        RECT 658.950 760.950 661.050 761.400 ;
        RECT 727.950 760.950 730.050 761.400 ;
        RECT 757.950 762.600 760.050 763.050 ;
        RECT 784.950 762.600 787.050 763.050 ;
        RECT 757.950 761.400 787.050 762.600 ;
        RECT 757.950 760.950 760.050 761.400 ;
        RECT 784.950 760.950 787.050 761.400 ;
        RECT 352.950 759.600 355.050 760.050 ;
        RECT 397.950 759.600 400.050 760.050 ;
        RECT 589.950 759.600 592.050 760.050 ;
        RECT 352.950 758.400 592.050 759.600 ;
        RECT 352.950 757.950 355.050 758.400 ;
        RECT 397.950 757.950 400.050 758.400 ;
        RECT 589.950 757.950 592.050 758.400 ;
        RECT 613.950 759.600 616.050 760.050 ;
        RECT 736.950 759.600 739.050 760.050 ;
        RECT 613.950 758.400 739.050 759.600 ;
        RECT 613.950 757.950 616.050 758.400 ;
        RECT 736.950 757.950 739.050 758.400 ;
        RECT 799.950 759.600 802.050 760.050 ;
        RECT 817.950 759.600 820.050 760.050 ;
        RECT 799.950 758.400 820.050 759.600 ;
        RECT 799.950 757.950 802.050 758.400 ;
        RECT 817.950 757.950 820.050 758.400 ;
        RECT 265.950 756.600 268.050 757.050 ;
        RECT 286.950 756.600 289.050 757.050 ;
        RECT 313.950 756.600 316.050 757.050 ;
        RECT 364.950 756.600 367.050 757.050 ;
        RECT 265.950 755.400 367.050 756.600 ;
        RECT 265.950 754.950 268.050 755.400 ;
        RECT 286.950 754.950 289.050 755.400 ;
        RECT 313.950 754.950 316.050 755.400 ;
        RECT 364.950 754.950 367.050 755.400 ;
        RECT 424.950 756.600 427.050 757.050 ;
        RECT 574.950 756.600 577.050 757.050 ;
        RECT 424.950 755.400 577.050 756.600 ;
        RECT 424.950 754.950 427.050 755.400 ;
        RECT 574.950 754.950 577.050 755.400 ;
        RECT 634.950 756.600 637.050 757.050 ;
        RECT 691.950 756.600 694.050 757.050 ;
        RECT 697.950 756.600 700.050 757.050 ;
        RECT 634.950 755.400 700.050 756.600 ;
        RECT 634.950 754.950 637.050 755.400 ;
        RECT 691.950 754.950 694.050 755.400 ;
        RECT 697.950 754.950 700.050 755.400 ;
        RECT 706.950 756.600 709.050 757.050 ;
        RECT 733.950 756.600 736.050 757.050 ;
        RECT 706.950 755.400 736.050 756.600 ;
        RECT 706.950 754.950 709.050 755.400 ;
        RECT 733.950 754.950 736.050 755.400 ;
        RECT 4.950 753.600 7.050 754.050 ;
        RECT 55.950 753.600 58.050 754.050 ;
        RECT 4.950 752.400 58.050 753.600 ;
        RECT 4.950 751.950 7.050 752.400 ;
        RECT 55.950 751.950 58.050 752.400 ;
        RECT 211.950 753.600 214.050 754.050 ;
        RECT 364.950 753.600 367.050 754.050 ;
        RECT 211.950 752.400 367.050 753.600 ;
        RECT 211.950 751.950 214.050 752.400 ;
        RECT 364.950 751.950 367.050 752.400 ;
        RECT 403.950 753.600 406.050 754.050 ;
        RECT 448.950 753.600 451.050 754.050 ;
        RECT 490.950 753.600 493.050 754.050 ;
        RECT 403.950 752.400 493.050 753.600 ;
        RECT 403.950 751.950 406.050 752.400 ;
        RECT 448.950 751.950 451.050 752.400 ;
        RECT 490.950 751.950 493.050 752.400 ;
        RECT 619.950 753.600 622.050 754.050 ;
        RECT 634.950 753.600 637.050 754.050 ;
        RECT 619.950 752.400 637.050 753.600 ;
        RECT 619.950 751.950 622.050 752.400 ;
        RECT 634.950 751.950 637.050 752.400 ;
        RECT 457.950 750.600 460.050 751.050 ;
        RECT 466.950 750.600 469.050 751.050 ;
        RECT 472.950 750.600 475.050 751.050 ;
        RECT 508.950 750.600 511.050 751.050 ;
        RECT 457.950 749.400 511.050 750.600 ;
        RECT 457.950 748.950 460.050 749.400 ;
        RECT 466.950 748.950 469.050 749.400 ;
        RECT 472.950 748.950 475.050 749.400 ;
        RECT 508.950 748.950 511.050 749.400 ;
        RECT 511.950 750.600 514.050 751.050 ;
        RECT 526.950 750.600 529.050 751.050 ;
        RECT 565.950 750.600 568.050 751.050 ;
        RECT 511.950 749.400 568.050 750.600 ;
        RECT 511.950 748.950 514.050 749.400 ;
        RECT 526.950 748.950 529.050 749.400 ;
        RECT 565.950 748.950 568.050 749.400 ;
        RECT 574.950 750.600 577.050 751.050 ;
        RECT 733.950 750.600 736.050 751.050 ;
        RECT 574.950 749.400 736.050 750.600 ;
        RECT 574.950 748.950 577.050 749.400 ;
        RECT 733.950 748.950 736.050 749.400 ;
        RECT 751.950 750.600 754.050 751.050 ;
        RECT 793.950 750.600 796.050 751.050 ;
        RECT 751.950 749.400 796.050 750.600 ;
        RECT 751.950 748.950 754.050 749.400 ;
        RECT 793.950 748.950 796.050 749.400 ;
        RECT 10.950 747.600 13.050 748.050 ;
        RECT 55.950 747.600 58.050 748.050 ;
        RECT 61.950 747.600 64.050 748.050 ;
        RECT 10.950 746.400 64.050 747.600 ;
        RECT 10.950 745.950 13.050 746.400 ;
        RECT 55.950 745.950 58.050 746.400 ;
        RECT 61.950 745.950 64.050 746.400 ;
        RECT 142.950 747.600 145.050 748.050 ;
        RECT 148.950 747.600 151.050 748.050 ;
        RECT 184.950 747.600 187.050 748.050 ;
        RECT 142.950 746.400 187.050 747.600 ;
        RECT 142.950 745.950 145.050 746.400 ;
        RECT 148.950 745.950 151.050 746.400 ;
        RECT 184.950 745.950 187.050 746.400 ;
        RECT 193.950 747.600 196.050 748.050 ;
        RECT 199.950 747.600 202.050 748.050 ;
        RECT 193.950 746.400 202.050 747.600 ;
        RECT 193.950 745.950 196.050 746.400 ;
        RECT 199.950 745.950 202.050 746.400 ;
        RECT 235.950 747.600 238.050 748.050 ;
        RECT 256.950 747.600 259.050 748.050 ;
        RECT 274.950 747.600 277.050 748.050 ;
        RECT 235.950 746.400 277.050 747.600 ;
        RECT 235.950 745.950 238.050 746.400 ;
        RECT 256.950 745.950 259.050 746.400 ;
        RECT 274.950 745.950 277.050 746.400 ;
        RECT 319.950 747.600 322.050 748.050 ;
        RECT 355.950 747.600 358.050 748.050 ;
        RECT 319.950 746.400 358.050 747.600 ;
        RECT 319.950 745.950 322.050 746.400 ;
        RECT 355.950 745.950 358.050 746.400 ;
        RECT 412.950 747.600 415.050 748.050 ;
        RECT 415.950 747.600 418.050 748.050 ;
        RECT 427.950 747.600 430.050 748.050 ;
        RECT 412.950 746.400 430.050 747.600 ;
        RECT 412.950 745.950 415.050 746.400 ;
        RECT 415.950 745.950 418.050 746.400 ;
        RECT 427.950 745.950 430.050 746.400 ;
        RECT 475.950 745.950 478.050 748.050 ;
        RECT 484.950 747.600 487.050 748.050 ;
        RECT 496.950 747.600 499.050 748.050 ;
        RECT 484.950 746.400 499.050 747.600 ;
        RECT 484.950 745.950 487.050 746.400 ;
        RECT 496.950 745.950 499.050 746.400 ;
        RECT 514.950 747.600 517.050 748.050 ;
        RECT 523.950 747.600 526.050 748.050 ;
        RECT 529.950 747.600 532.050 748.050 ;
        RECT 514.950 746.400 532.050 747.600 ;
        RECT 514.950 745.950 517.050 746.400 ;
        RECT 523.950 745.950 526.050 746.400 ;
        RECT 529.950 745.950 532.050 746.400 ;
        RECT 577.950 747.600 580.050 748.050 ;
        RECT 592.950 747.600 595.050 748.050 ;
        RECT 601.950 747.600 604.050 748.050 ;
        RECT 619.950 747.600 622.050 748.050 ;
        RECT 577.950 746.400 622.050 747.600 ;
        RECT 577.950 745.950 580.050 746.400 ;
        RECT 592.950 745.950 595.050 746.400 ;
        RECT 601.950 745.950 604.050 746.400 ;
        RECT 619.950 745.950 622.050 746.400 ;
        RECT 655.950 747.600 658.050 748.050 ;
        RECT 667.950 747.600 670.050 748.050 ;
        RECT 688.950 747.600 691.050 748.050 ;
        RECT 655.950 746.400 691.050 747.600 ;
        RECT 655.950 745.950 658.050 746.400 ;
        RECT 667.950 745.950 670.050 746.400 ;
        RECT 688.950 745.950 691.050 746.400 ;
        RECT 742.950 747.600 745.050 748.050 ;
        RECT 769.950 747.600 772.050 748.050 ;
        RECT 742.950 746.400 772.050 747.600 ;
        RECT 742.950 745.950 745.050 746.400 ;
        RECT 769.950 745.950 772.050 746.400 ;
        RECT 817.950 747.600 820.050 748.050 ;
        RECT 862.950 747.600 865.050 748.050 ;
        RECT 817.950 746.400 865.050 747.600 ;
        RECT 817.950 745.950 820.050 746.400 ;
        RECT 862.950 745.950 865.050 746.400 ;
        RECT 31.950 744.600 34.050 745.050 ;
        RECT 26.400 743.400 34.050 744.600 ;
        RECT 26.400 738.600 27.600 743.400 ;
        RECT 31.950 742.950 34.050 743.400 ;
        RECT 58.950 742.950 61.050 745.050 ;
        RECT 85.950 744.600 88.050 745.050 ;
        RECT 94.950 744.600 97.050 745.050 ;
        RECT 85.950 743.400 97.050 744.600 ;
        RECT 85.950 742.950 88.050 743.400 ;
        RECT 94.950 742.950 97.050 743.400 ;
        RECT 103.950 744.600 106.050 745.050 ;
        RECT 115.950 744.600 118.050 745.050 ;
        RECT 103.950 743.400 118.050 744.600 ;
        RECT 103.950 742.950 106.050 743.400 ;
        RECT 115.950 742.950 118.050 743.400 ;
        RECT 121.950 744.600 124.050 745.050 ;
        RECT 133.950 744.600 136.050 745.050 ;
        RECT 166.950 744.600 169.050 745.050 ;
        RECT 175.950 744.600 178.050 745.050 ;
        RECT 121.950 743.400 136.050 744.600 ;
        RECT 121.950 742.950 124.050 743.400 ;
        RECT 133.950 742.950 136.050 743.400 ;
        RECT 140.400 743.400 162.600 744.600 ;
        RECT 28.950 741.600 31.050 742.050 ;
        RECT 34.950 741.600 37.050 742.050 ;
        RECT 28.950 740.400 37.050 741.600 ;
        RECT 28.950 739.950 31.050 740.400 ;
        RECT 34.950 739.950 37.050 740.400 ;
        RECT 43.950 741.600 46.050 742.050 ;
        RECT 49.950 741.600 52.050 742.050 ;
        RECT 43.950 740.400 52.050 741.600 ;
        RECT 43.950 739.950 46.050 740.400 ;
        RECT 49.950 739.950 52.050 740.400 ;
        RECT 59.400 739.050 60.600 742.950 ;
        RECT 140.400 742.050 141.600 743.400 ;
        RECT 82.950 741.600 85.050 742.050 ;
        RECT 97.950 741.600 100.050 742.050 ;
        RECT 82.950 740.400 100.050 741.600 ;
        RECT 82.950 739.950 85.050 740.400 ;
        RECT 97.950 739.950 100.050 740.400 ;
        RECT 118.950 741.600 121.050 742.050 ;
        RECT 139.950 741.600 142.050 742.050 ;
        RECT 118.950 740.400 142.050 741.600 ;
        RECT 118.950 739.950 121.050 740.400 ;
        RECT 139.950 739.950 142.050 740.400 ;
        RECT 148.950 741.600 151.050 742.050 ;
        RECT 157.950 741.600 160.050 742.050 ;
        RECT 148.950 740.400 160.050 741.600 ;
        RECT 161.400 741.600 162.600 743.400 ;
        RECT 166.950 743.400 178.050 744.600 ;
        RECT 166.950 742.950 169.050 743.400 ;
        RECT 175.950 742.950 178.050 743.400 ;
        RECT 280.950 744.600 283.050 745.050 ;
        RECT 286.950 744.600 289.050 745.050 ;
        RECT 280.950 743.400 289.050 744.600 ;
        RECT 280.950 742.950 283.050 743.400 ;
        RECT 286.950 742.950 289.050 743.400 ;
        RECT 361.950 744.600 364.050 745.050 ;
        RECT 367.950 744.600 370.050 745.050 ;
        RECT 361.950 743.400 370.050 744.600 ;
        RECT 361.950 742.950 364.050 743.400 ;
        RECT 367.950 742.950 370.050 743.400 ;
        RECT 445.950 744.600 448.050 745.050 ;
        RECT 469.950 744.600 472.050 745.050 ;
        RECT 445.950 743.400 472.050 744.600 ;
        RECT 445.950 742.950 448.050 743.400 ;
        RECT 469.950 742.950 472.050 743.400 ;
        RECT 181.950 741.600 184.050 742.050 ;
        RECT 196.950 741.600 199.050 742.050 ;
        RECT 161.400 740.400 199.050 741.600 ;
        RECT 148.950 739.950 151.050 740.400 ;
        RECT 157.950 739.950 160.050 740.400 ;
        RECT 181.950 739.950 184.050 740.400 ;
        RECT 196.950 739.950 199.050 740.400 ;
        RECT 208.950 741.600 211.050 742.050 ;
        RECT 214.950 741.600 217.050 742.050 ;
        RECT 208.950 740.400 217.050 741.600 ;
        RECT 208.950 739.950 211.050 740.400 ;
        RECT 214.950 739.950 217.050 740.400 ;
        RECT 259.950 741.600 262.050 742.050 ;
        RECT 265.950 741.600 268.050 742.050 ;
        RECT 259.950 740.400 268.050 741.600 ;
        RECT 259.950 739.950 262.050 740.400 ;
        RECT 265.950 739.950 268.050 740.400 ;
        RECT 268.950 741.600 271.050 742.050 ;
        RECT 277.950 741.600 280.050 742.050 ;
        RECT 268.950 740.400 280.050 741.600 ;
        RECT 268.950 739.950 271.050 740.400 ;
        RECT 277.950 739.950 280.050 740.400 ;
        RECT 283.950 741.600 286.050 742.050 ;
        RECT 295.950 741.600 298.050 742.050 ;
        RECT 283.950 740.400 298.050 741.600 ;
        RECT 283.950 739.950 286.050 740.400 ;
        RECT 295.950 739.950 298.050 740.400 ;
        RECT 316.950 741.600 319.050 742.050 ;
        RECT 328.950 741.600 331.050 742.050 ;
        RECT 316.950 740.400 331.050 741.600 ;
        RECT 316.950 739.950 319.050 740.400 ;
        RECT 328.950 739.950 331.050 740.400 ;
        RECT 337.950 741.600 340.050 742.050 ;
        RECT 358.950 741.600 361.050 742.050 ;
        RECT 337.950 740.400 361.050 741.600 ;
        RECT 337.950 739.950 340.050 740.400 ;
        RECT 358.950 739.950 361.050 740.400 ;
        RECT 376.950 741.600 379.050 742.050 ;
        RECT 394.950 741.600 397.050 742.050 ;
        RECT 376.950 740.400 397.050 741.600 ;
        RECT 376.950 739.950 379.050 740.400 ;
        RECT 394.950 739.950 397.050 740.400 ;
        RECT 430.950 741.600 433.050 742.050 ;
        RECT 442.950 741.600 445.050 742.050 ;
        RECT 430.950 740.400 445.050 741.600 ;
        RECT 430.950 739.950 433.050 740.400 ;
        RECT 442.950 739.950 445.050 740.400 ;
        RECT 476.400 739.050 477.600 745.950 ;
        RECT 496.950 744.600 499.050 745.050 ;
        RECT 505.950 744.600 508.050 745.050 ;
        RECT 496.950 743.400 508.050 744.600 ;
        RECT 496.950 742.950 499.050 743.400 ;
        RECT 505.950 742.950 508.050 743.400 ;
        RECT 607.950 744.600 610.050 745.050 ;
        RECT 640.950 744.600 643.050 745.050 ;
        RECT 643.950 744.600 646.050 745.050 ;
        RECT 607.950 743.400 646.050 744.600 ;
        RECT 607.950 742.950 610.050 743.400 ;
        RECT 640.950 742.950 643.050 743.400 ;
        RECT 643.950 742.950 646.050 743.400 ;
        RECT 673.950 744.600 676.050 745.050 ;
        RECT 694.950 744.600 697.050 745.050 ;
        RECT 709.950 744.600 712.050 745.050 ;
        RECT 673.950 743.400 712.050 744.600 ;
        RECT 673.950 742.950 676.050 743.400 ;
        RECT 694.950 742.950 697.050 743.400 ;
        RECT 709.950 742.950 712.050 743.400 ;
        RECT 736.950 744.600 739.050 745.050 ;
        RECT 751.950 744.600 754.050 745.050 ;
        RECT 736.950 743.400 754.050 744.600 ;
        RECT 736.950 742.950 739.050 743.400 ;
        RECT 751.950 742.950 754.050 743.400 ;
        RECT 505.950 741.600 508.050 742.050 ;
        RECT 511.950 741.600 514.050 742.050 ;
        RECT 505.950 740.400 514.050 741.600 ;
        RECT 505.950 739.950 508.050 740.400 ;
        RECT 511.950 739.950 514.050 740.400 ;
        RECT 514.950 741.600 517.050 742.050 ;
        RECT 571.950 741.600 574.050 742.050 ;
        RECT 628.950 741.600 631.050 742.050 ;
        RECT 661.950 741.600 664.050 742.050 ;
        RECT 715.950 741.600 718.050 742.050 ;
        RECT 514.950 740.400 657.600 741.600 ;
        RECT 514.950 739.950 517.050 740.400 ;
        RECT 571.950 739.950 574.050 740.400 ;
        RECT 628.950 739.950 631.050 740.400 ;
        RECT 656.400 739.050 657.600 740.400 ;
        RECT 661.950 740.400 718.050 741.600 ;
        RECT 661.950 739.950 664.050 740.400 ;
        RECT 715.950 739.950 718.050 740.400 ;
        RECT 772.950 741.600 775.050 742.050 ;
        RECT 826.950 741.600 829.050 742.050 ;
        RECT 772.950 740.400 829.050 741.600 ;
        RECT 772.950 739.950 775.050 740.400 ;
        RECT 826.950 739.950 829.050 740.400 ;
        RECT 835.950 741.600 838.050 742.050 ;
        RECT 841.950 741.600 844.050 742.050 ;
        RECT 835.950 740.400 844.050 741.600 ;
        RECT 835.950 739.950 838.050 740.400 ;
        RECT 841.950 739.950 844.050 740.400 ;
        RECT 31.950 738.600 34.050 739.050 ;
        RECT 26.400 737.400 34.050 738.600 ;
        RECT 31.950 736.950 34.050 737.400 ;
        RECT 37.950 738.600 40.050 739.050 ;
        RECT 46.950 738.600 49.050 739.050 ;
        RECT 52.950 738.600 55.050 739.050 ;
        RECT 37.950 737.400 55.050 738.600 ;
        RECT 37.950 736.950 40.050 737.400 ;
        RECT 46.950 736.950 49.050 737.400 ;
        RECT 52.950 736.950 55.050 737.400 ;
        RECT 58.950 736.950 61.050 739.050 ;
        RECT 100.950 738.600 103.050 739.050 ;
        RECT 115.950 738.600 118.050 739.050 ;
        RECT 100.950 737.400 118.050 738.600 ;
        RECT 100.950 736.950 103.050 737.400 ;
        RECT 115.950 736.950 118.050 737.400 ;
        RECT 217.950 738.600 220.050 739.050 ;
        RECT 223.950 738.600 226.050 739.050 ;
        RECT 229.950 738.600 232.050 739.050 ;
        RECT 217.950 737.400 232.050 738.600 ;
        RECT 217.950 736.950 220.050 737.400 ;
        RECT 223.950 736.950 226.050 737.400 ;
        RECT 229.950 736.950 232.050 737.400 ;
        RECT 244.950 738.600 247.050 739.050 ;
        RECT 271.950 738.600 274.050 739.050 ;
        RECT 244.950 737.400 274.050 738.600 ;
        RECT 244.950 736.950 247.050 737.400 ;
        RECT 271.950 736.950 274.050 737.400 ;
        RECT 286.950 738.600 289.050 739.050 ;
        RECT 292.950 738.600 295.050 739.050 ;
        RECT 286.950 737.400 295.050 738.600 ;
        RECT 286.950 736.950 289.050 737.400 ;
        RECT 292.950 736.950 295.050 737.400 ;
        RECT 322.950 738.600 325.050 739.050 ;
        RECT 373.950 738.600 376.050 739.050 ;
        RECT 322.950 737.400 376.050 738.600 ;
        RECT 322.950 736.950 325.050 737.400 ;
        RECT 373.950 736.950 376.050 737.400 ;
        RECT 379.950 738.600 382.050 739.050 ;
        RECT 388.950 738.600 391.050 739.050 ;
        RECT 379.950 737.400 391.050 738.600 ;
        RECT 379.950 736.950 382.050 737.400 ;
        RECT 388.950 736.950 391.050 737.400 ;
        RECT 412.950 738.600 415.050 739.050 ;
        RECT 430.950 738.600 433.050 739.050 ;
        RECT 412.950 737.400 433.050 738.600 ;
        RECT 412.950 736.950 415.050 737.400 ;
        RECT 430.950 736.950 433.050 737.400 ;
        RECT 475.950 736.950 478.050 739.050 ;
        RECT 526.950 738.600 529.050 739.050 ;
        RECT 535.950 738.600 538.050 739.050 ;
        RECT 574.950 738.600 577.050 739.050 ;
        RECT 604.950 738.600 607.050 739.050 ;
        RECT 526.950 737.400 538.050 738.600 ;
        RECT 526.950 736.950 529.050 737.400 ;
        RECT 535.950 736.950 538.050 737.400 ;
        RECT 563.400 737.400 607.050 738.600 ;
        RECT 31.950 735.600 34.050 736.050 ;
        RECT 43.950 735.600 46.050 736.050 ;
        RECT 31.950 734.400 46.050 735.600 ;
        RECT 31.950 733.950 34.050 734.400 ;
        RECT 43.950 733.950 46.050 734.400 ;
        RECT 88.950 735.600 91.050 736.050 ;
        RECT 94.950 735.600 97.050 736.050 ;
        RECT 88.950 734.400 97.050 735.600 ;
        RECT 88.950 733.950 91.050 734.400 ;
        RECT 94.950 733.950 97.050 734.400 ;
        RECT 211.950 735.600 214.050 736.050 ;
        RECT 232.950 735.600 235.050 736.050 ;
        RECT 211.950 734.400 235.050 735.600 ;
        RECT 211.950 733.950 214.050 734.400 ;
        RECT 232.950 733.950 235.050 734.400 ;
        RECT 250.950 735.600 253.050 736.050 ;
        RECT 277.950 735.600 280.050 736.050 ;
        RECT 514.950 735.600 517.050 736.050 ;
        RECT 250.950 734.400 280.050 735.600 ;
        RECT 250.950 733.950 253.050 734.400 ;
        RECT 277.950 733.950 280.050 734.400 ;
        RECT 380.400 734.400 517.050 735.600 ;
        RECT 380.400 733.050 381.600 734.400 ;
        RECT 514.950 733.950 517.050 734.400 ;
        RECT 535.950 735.600 538.050 736.050 ;
        RECT 541.950 735.600 544.050 736.050 ;
        RECT 563.400 735.600 564.600 737.400 ;
        RECT 574.950 736.950 577.050 737.400 ;
        RECT 604.950 736.950 607.050 737.400 ;
        RECT 610.950 738.600 613.050 739.050 ;
        RECT 616.950 738.600 619.050 739.050 ;
        RECT 610.950 737.400 619.050 738.600 ;
        RECT 610.950 736.950 613.050 737.400 ;
        RECT 616.950 736.950 619.050 737.400 ;
        RECT 625.950 738.600 628.050 739.050 ;
        RECT 631.950 738.600 634.050 739.050 ;
        RECT 652.950 738.600 655.050 739.050 ;
        RECT 625.950 737.400 630.600 738.600 ;
        RECT 625.950 736.950 628.050 737.400 ;
        RECT 535.950 734.400 564.600 735.600 ;
        RECT 629.400 735.600 630.600 737.400 ;
        RECT 631.950 737.400 655.050 738.600 ;
        RECT 631.950 736.950 634.050 737.400 ;
        RECT 652.950 736.950 655.050 737.400 ;
        RECT 655.950 736.950 658.050 739.050 ;
        RECT 682.950 738.600 685.050 739.050 ;
        RECT 691.950 738.600 694.050 739.050 ;
        RECT 682.950 737.400 694.050 738.600 ;
        RECT 682.950 736.950 685.050 737.400 ;
        RECT 691.950 736.950 694.050 737.400 ;
        RECT 640.950 735.600 643.050 736.050 ;
        RECT 629.400 734.400 643.050 735.600 ;
        RECT 535.950 733.950 538.050 734.400 ;
        RECT 541.950 733.950 544.050 734.400 ;
        RECT 640.950 733.950 643.050 734.400 ;
        RECT 16.950 732.600 19.050 733.050 ;
        RECT 43.950 732.600 46.050 733.050 ;
        RECT 73.950 732.600 76.050 733.050 ;
        RECT 16.950 731.400 76.050 732.600 ;
        RECT 16.950 730.950 19.050 731.400 ;
        RECT 43.950 730.950 46.050 731.400 ;
        RECT 73.950 730.950 76.050 731.400 ;
        RECT 163.950 732.600 166.050 733.050 ;
        RECT 220.950 732.600 223.050 733.050 ;
        RECT 163.950 731.400 223.050 732.600 ;
        RECT 163.950 730.950 166.050 731.400 ;
        RECT 220.950 730.950 223.050 731.400 ;
        RECT 379.950 730.950 382.050 733.050 ;
        RECT 475.950 732.600 478.050 733.050 ;
        RECT 493.950 732.600 496.050 733.050 ;
        RECT 556.950 732.600 559.050 733.050 ;
        RECT 475.950 731.400 559.050 732.600 ;
        RECT 475.950 730.950 478.050 731.400 ;
        RECT 493.950 730.950 496.050 731.400 ;
        RECT 556.950 730.950 559.050 731.400 ;
        RECT 640.950 732.600 643.050 733.050 ;
        RECT 664.950 732.600 667.050 733.050 ;
        RECT 640.950 731.400 667.050 732.600 ;
        RECT 640.950 730.950 643.050 731.400 ;
        RECT 664.950 730.950 667.050 731.400 ;
        RECT 388.950 729.600 391.050 730.050 ;
        RECT 496.950 729.600 499.050 730.050 ;
        RECT 388.950 728.400 499.050 729.600 ;
        RECT 388.950 727.950 391.050 728.400 ;
        RECT 496.950 727.950 499.050 728.400 ;
        RECT 532.950 729.600 535.050 730.050 ;
        RECT 550.950 729.600 553.050 730.050 ;
        RECT 532.950 728.400 553.050 729.600 ;
        RECT 532.950 727.950 535.050 728.400 ;
        RECT 550.950 727.950 553.050 728.400 ;
        RECT 595.950 729.600 598.050 730.050 ;
        RECT 781.950 729.600 784.050 730.050 ;
        RECT 595.950 728.400 784.050 729.600 ;
        RECT 595.950 727.950 598.050 728.400 ;
        RECT 781.950 727.950 784.050 728.400 ;
        RECT 19.950 726.600 22.050 727.050 ;
        RECT 28.950 726.600 31.050 727.050 ;
        RECT 82.950 726.600 85.050 727.050 ;
        RECT 19.950 725.400 85.050 726.600 ;
        RECT 19.950 724.950 22.050 725.400 ;
        RECT 28.950 724.950 31.050 725.400 ;
        RECT 82.950 724.950 85.050 725.400 ;
        RECT 469.950 726.600 472.050 727.050 ;
        RECT 691.950 726.600 694.050 727.050 ;
        RECT 469.950 725.400 694.050 726.600 ;
        RECT 469.950 724.950 472.050 725.400 ;
        RECT 691.950 724.950 694.050 725.400 ;
        RECT 553.950 723.600 556.050 724.050 ;
        RECT 580.950 723.600 583.050 724.050 ;
        RECT 553.950 722.400 583.050 723.600 ;
        RECT 553.950 721.950 556.050 722.400 ;
        RECT 580.950 721.950 583.050 722.400 ;
        RECT 649.950 723.600 652.050 724.050 ;
        RECT 673.950 723.600 676.050 724.050 ;
        RECT 688.950 723.600 691.050 724.050 ;
        RECT 649.950 722.400 691.050 723.600 ;
        RECT 649.950 721.950 652.050 722.400 ;
        RECT 673.950 721.950 676.050 722.400 ;
        RECT 688.950 721.950 691.050 722.400 ;
        RECT 271.950 720.600 274.050 721.050 ;
        RECT 514.950 720.600 517.050 721.050 ;
        RECT 271.950 719.400 517.050 720.600 ;
        RECT 271.950 718.950 274.050 719.400 ;
        RECT 514.950 718.950 517.050 719.400 ;
        RECT 568.950 720.600 571.050 721.050 ;
        RECT 592.950 720.600 595.050 721.050 ;
        RECT 568.950 719.400 595.050 720.600 ;
        RECT 568.950 718.950 571.050 719.400 ;
        RECT 592.950 718.950 595.050 719.400 ;
        RECT 4.950 717.600 7.050 718.050 ;
        RECT 16.950 717.600 19.050 718.050 ;
        RECT 4.950 716.400 19.050 717.600 ;
        RECT 4.950 715.950 7.050 716.400 ;
        RECT 16.950 715.950 19.050 716.400 ;
        RECT 25.950 717.600 28.050 718.050 ;
        RECT 46.950 717.600 49.050 718.050 ;
        RECT 25.950 716.400 49.050 717.600 ;
        RECT 25.950 715.950 28.050 716.400 ;
        RECT 46.950 715.950 49.050 716.400 ;
        RECT 193.950 717.600 196.050 718.050 ;
        RECT 316.950 717.600 319.050 718.050 ;
        RECT 193.950 716.400 319.050 717.600 ;
        RECT 193.950 715.950 196.050 716.400 ;
        RECT 316.950 715.950 319.050 716.400 ;
        RECT 508.950 717.600 511.050 718.050 ;
        RECT 586.950 717.600 589.050 718.050 ;
        RECT 508.950 716.400 589.050 717.600 ;
        RECT 508.950 715.950 511.050 716.400 ;
        RECT 586.950 715.950 589.050 716.400 ;
        RECT 805.950 717.600 808.050 718.050 ;
        RECT 817.950 717.600 820.050 718.050 ;
        RECT 805.950 716.400 820.050 717.600 ;
        RECT 805.950 715.950 808.050 716.400 ;
        RECT 817.950 715.950 820.050 716.400 ;
        RECT 13.950 714.600 16.050 715.050 ;
        RECT 22.950 714.600 25.050 715.050 ;
        RECT 61.950 714.600 64.050 715.050 ;
        RECT 67.950 714.600 70.050 715.050 ;
        RECT 13.950 713.400 70.050 714.600 ;
        RECT 13.950 712.950 16.050 713.400 ;
        RECT 22.950 712.950 25.050 713.400 ;
        RECT 61.950 712.950 64.050 713.400 ;
        RECT 67.950 712.950 70.050 713.400 ;
        RECT 517.950 714.600 520.050 715.050 ;
        RECT 520.950 714.600 523.050 715.050 ;
        RECT 622.950 714.600 625.050 715.050 ;
        RECT 517.950 713.400 625.050 714.600 ;
        RECT 517.950 712.950 520.050 713.400 ;
        RECT 520.950 712.950 523.050 713.400 ;
        RECT 622.950 712.950 625.050 713.400 ;
        RECT 202.950 711.600 205.050 712.050 ;
        RECT 319.950 711.600 322.050 712.050 ;
        RECT 202.950 710.400 322.050 711.600 ;
        RECT 202.950 709.950 205.050 710.400 ;
        RECT 319.950 709.950 322.050 710.400 ;
        RECT 361.950 711.600 364.050 712.050 ;
        RECT 397.950 711.600 400.050 712.050 ;
        RECT 361.950 710.400 400.050 711.600 ;
        RECT 361.950 709.950 364.050 710.400 ;
        RECT 397.950 709.950 400.050 710.400 ;
        RECT 478.950 711.600 481.050 712.050 ;
        RECT 547.950 711.600 550.050 712.050 ;
        RECT 703.950 711.600 706.050 712.050 ;
        RECT 478.950 710.400 706.050 711.600 ;
        RECT 478.950 709.950 481.050 710.400 ;
        RECT 547.950 709.950 550.050 710.400 ;
        RECT 703.950 709.950 706.050 710.400 ;
        RECT 781.950 711.600 784.050 712.050 ;
        RECT 790.950 711.600 793.050 712.050 ;
        RECT 781.950 710.400 793.050 711.600 ;
        RECT 781.950 709.950 784.050 710.400 ;
        RECT 790.950 709.950 793.050 710.400 ;
        RECT 835.950 711.600 838.050 712.050 ;
        RECT 841.950 711.600 844.050 712.050 ;
        RECT 835.950 710.400 844.050 711.600 ;
        RECT 835.950 709.950 838.050 710.400 ;
        RECT 841.950 709.950 844.050 710.400 ;
        RECT 22.950 708.600 25.050 709.050 ;
        RECT 28.950 708.600 31.050 709.050 ;
        RECT 22.950 707.400 31.050 708.600 ;
        RECT 22.950 706.950 25.050 707.400 ;
        RECT 28.950 706.950 31.050 707.400 ;
        RECT 55.950 708.600 58.050 709.050 ;
        RECT 151.950 708.600 154.050 709.050 ;
        RECT 55.950 707.400 154.050 708.600 ;
        RECT 55.950 706.950 58.050 707.400 ;
        RECT 151.950 706.950 154.050 707.400 ;
        RECT 214.950 708.600 217.050 709.050 ;
        RECT 280.950 708.600 283.050 709.050 ;
        RECT 214.950 707.400 283.050 708.600 ;
        RECT 214.950 706.950 217.050 707.400 ;
        RECT 280.950 706.950 283.050 707.400 ;
        RECT 334.950 708.600 337.050 709.050 ;
        RECT 379.950 708.600 382.050 709.050 ;
        RECT 334.950 707.400 382.050 708.600 ;
        RECT 334.950 706.950 337.050 707.400 ;
        RECT 379.950 706.950 382.050 707.400 ;
        RECT 469.950 708.600 472.050 709.050 ;
        RECT 484.950 708.600 487.050 709.050 ;
        RECT 469.950 707.400 487.050 708.600 ;
        RECT 469.950 706.950 472.050 707.400 ;
        RECT 484.950 706.950 487.050 707.400 ;
        RECT 511.950 708.600 514.050 709.050 ;
        RECT 538.950 708.600 541.050 709.050 ;
        RECT 511.950 707.400 541.050 708.600 ;
        RECT 511.950 706.950 514.050 707.400 ;
        RECT 538.950 706.950 541.050 707.400 ;
        RECT 571.950 708.600 574.050 709.050 ;
        RECT 640.950 708.600 643.050 709.050 ;
        RECT 571.950 707.400 643.050 708.600 ;
        RECT 571.950 706.950 574.050 707.400 ;
        RECT 640.950 706.950 643.050 707.400 ;
        RECT 661.950 708.600 664.050 709.050 ;
        RECT 673.950 708.600 676.050 709.050 ;
        RECT 661.950 707.400 676.050 708.600 ;
        RECT 661.950 706.950 664.050 707.400 ;
        RECT 673.950 706.950 676.050 707.400 ;
        RECT 787.950 708.600 790.050 709.050 ;
        RECT 790.950 708.600 793.050 709.050 ;
        RECT 850.950 708.600 853.050 709.050 ;
        RECT 787.950 707.400 853.050 708.600 ;
        RECT 787.950 706.950 790.050 707.400 ;
        RECT 790.950 706.950 793.050 707.400 ;
        RECT 850.950 706.950 853.050 707.400 ;
        RECT 853.950 708.600 856.050 709.050 ;
        RECT 862.950 708.600 865.050 709.050 ;
        RECT 853.950 707.400 865.050 708.600 ;
        RECT 853.950 706.950 856.050 707.400 ;
        RECT 862.950 706.950 865.050 707.400 ;
        RECT 16.950 705.600 19.050 706.050 ;
        RECT 58.950 705.600 61.050 706.050 ;
        RECT 76.950 705.600 79.050 706.050 ;
        RECT 91.950 705.600 94.050 706.050 ;
        RECT 16.950 704.400 39.600 705.600 ;
        RECT 16.950 703.950 19.050 704.400 ;
        RECT 4.950 702.600 7.050 703.050 ;
        RECT 34.950 702.600 37.050 703.050 ;
        RECT 4.950 701.400 37.050 702.600 ;
        RECT 4.950 700.950 7.050 701.400 ;
        RECT 34.950 700.950 37.050 701.400 ;
        RECT 38.400 699.600 39.600 704.400 ;
        RECT 58.950 704.400 75.600 705.600 ;
        RECT 58.950 703.950 61.050 704.400 ;
        RECT 74.400 703.050 75.600 704.400 ;
        RECT 76.950 704.400 94.050 705.600 ;
        RECT 76.950 703.950 79.050 704.400 ;
        RECT 91.950 703.950 94.050 704.400 ;
        RECT 232.950 705.600 235.050 706.050 ;
        RECT 238.950 705.600 241.050 706.050 ;
        RECT 232.950 704.400 241.050 705.600 ;
        RECT 232.950 703.950 235.050 704.400 ;
        RECT 238.950 703.950 241.050 704.400 ;
        RECT 244.950 705.600 247.050 706.050 ;
        RECT 256.950 705.600 259.050 706.050 ;
        RECT 244.950 704.400 259.050 705.600 ;
        RECT 244.950 703.950 247.050 704.400 ;
        RECT 256.950 703.950 259.050 704.400 ;
        RECT 373.950 705.600 376.050 706.050 ;
        RECT 385.950 705.600 388.050 706.050 ;
        RECT 373.950 704.400 388.050 705.600 ;
        RECT 373.950 703.950 376.050 704.400 ;
        RECT 385.950 703.950 388.050 704.400 ;
        RECT 403.950 705.600 406.050 706.050 ;
        RECT 412.950 705.600 415.050 706.050 ;
        RECT 403.950 704.400 415.050 705.600 ;
        RECT 403.950 703.950 406.050 704.400 ;
        RECT 412.950 703.950 415.050 704.400 ;
        RECT 418.950 705.600 421.050 706.050 ;
        RECT 442.950 705.600 445.050 706.050 ;
        RECT 454.950 705.600 457.050 706.050 ;
        RECT 418.950 704.400 457.050 705.600 ;
        RECT 418.950 703.950 421.050 704.400 ;
        RECT 442.950 703.950 445.050 704.400 ;
        RECT 454.950 703.950 457.050 704.400 ;
        RECT 472.950 705.600 475.050 706.050 ;
        RECT 478.950 705.600 481.050 706.050 ;
        RECT 472.950 704.400 481.050 705.600 ;
        RECT 472.950 703.950 475.050 704.400 ;
        RECT 478.950 703.950 481.050 704.400 ;
        RECT 520.950 705.600 523.050 706.050 ;
        RECT 562.950 705.600 565.050 706.050 ;
        RECT 574.950 705.600 577.050 706.050 ;
        RECT 520.950 704.400 549.600 705.600 ;
        RECT 520.950 703.950 523.050 704.400 ;
        RECT 548.400 703.050 549.600 704.400 ;
        RECT 562.950 704.400 577.050 705.600 ;
        RECT 562.950 703.950 565.050 704.400 ;
        RECT 574.950 703.950 577.050 704.400 ;
        RECT 592.950 705.600 595.050 706.050 ;
        RECT 601.950 705.600 604.050 706.050 ;
        RECT 592.950 704.400 604.050 705.600 ;
        RECT 592.950 703.950 595.050 704.400 ;
        RECT 601.950 703.950 604.050 704.400 ;
        RECT 625.950 705.600 628.050 706.050 ;
        RECT 661.950 705.600 664.050 706.050 ;
        RECT 625.950 704.400 664.050 705.600 ;
        RECT 625.950 703.950 628.050 704.400 ;
        RECT 661.950 703.950 664.050 704.400 ;
        RECT 796.950 703.950 799.050 706.050 ;
        RECT 799.950 705.600 802.050 706.050 ;
        RECT 811.950 705.600 814.050 706.050 ;
        RECT 799.950 704.400 814.050 705.600 ;
        RECT 799.950 703.950 802.050 704.400 ;
        RECT 811.950 703.950 814.050 704.400 ;
        RECT 817.950 703.950 820.050 706.050 ;
        RECT 40.950 702.600 43.050 703.050 ;
        RECT 55.950 702.600 58.050 703.050 ;
        RECT 40.950 701.400 58.050 702.600 ;
        RECT 40.950 700.950 43.050 701.400 ;
        RECT 55.950 700.950 58.050 701.400 ;
        RECT 73.950 700.950 76.050 703.050 ;
        RECT 97.950 702.600 100.050 703.050 ;
        RECT 118.950 702.600 121.050 703.050 ;
        RECT 151.950 702.600 154.050 703.050 ;
        RECT 97.950 701.400 154.050 702.600 ;
        RECT 97.950 700.950 100.050 701.400 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 151.950 700.950 154.050 701.400 ;
        RECT 172.950 702.600 175.050 703.050 ;
        RECT 181.950 702.600 184.050 703.050 ;
        RECT 172.950 701.400 184.050 702.600 ;
        RECT 172.950 700.950 175.050 701.400 ;
        RECT 181.950 700.950 184.050 701.400 ;
        RECT 187.950 702.600 190.050 703.050 ;
        RECT 202.950 702.600 205.050 703.050 ;
        RECT 223.950 702.600 226.050 703.050 ;
        RECT 187.950 701.400 226.050 702.600 ;
        RECT 187.950 700.950 190.050 701.400 ;
        RECT 202.950 700.950 205.050 701.400 ;
        RECT 223.950 700.950 226.050 701.400 ;
        RECT 229.950 702.600 232.050 703.050 ;
        RECT 235.950 702.600 238.050 703.050 ;
        RECT 229.950 701.400 238.050 702.600 ;
        RECT 229.950 700.950 232.050 701.400 ;
        RECT 235.950 700.950 238.050 701.400 ;
        RECT 265.950 702.600 268.050 703.050 ;
        RECT 298.950 702.600 301.050 703.050 ;
        RECT 265.950 701.400 301.050 702.600 ;
        RECT 265.950 700.950 268.050 701.400 ;
        RECT 298.950 700.950 301.050 701.400 ;
        RECT 310.950 702.600 313.050 703.050 ;
        RECT 352.950 702.600 355.050 703.050 ;
        RECT 310.950 701.400 355.050 702.600 ;
        RECT 310.950 700.950 313.050 701.400 ;
        RECT 352.950 700.950 355.050 701.400 ;
        RECT 358.950 702.600 361.050 703.050 ;
        RECT 364.950 702.600 367.050 703.050 ;
        RECT 358.950 701.400 367.050 702.600 ;
        RECT 358.950 700.950 361.050 701.400 ;
        RECT 364.950 700.950 367.050 701.400 ;
        RECT 376.950 702.600 379.050 703.050 ;
        RECT 421.950 702.600 424.050 703.050 ;
        RECT 376.950 701.400 424.050 702.600 ;
        RECT 376.950 700.950 379.050 701.400 ;
        RECT 421.950 700.950 424.050 701.400 ;
        RECT 460.950 702.600 463.050 703.050 ;
        RECT 487.950 702.600 490.050 703.050 ;
        RECT 460.950 701.400 490.050 702.600 ;
        RECT 460.950 700.950 463.050 701.400 ;
        RECT 487.950 700.950 490.050 701.400 ;
        RECT 499.950 702.600 502.050 703.050 ;
        RECT 511.950 702.600 514.050 703.050 ;
        RECT 499.950 701.400 514.050 702.600 ;
        RECT 499.950 700.950 502.050 701.400 ;
        RECT 511.950 700.950 514.050 701.400 ;
        RECT 523.950 702.600 526.050 703.050 ;
        RECT 544.950 702.600 547.050 703.050 ;
        RECT 523.950 701.400 547.050 702.600 ;
        RECT 523.950 700.950 526.050 701.400 ;
        RECT 544.950 700.950 547.050 701.400 ;
        RECT 547.950 700.950 550.050 703.050 ;
        RECT 562.950 702.600 565.050 703.050 ;
        RECT 577.950 702.600 580.050 703.050 ;
        RECT 625.950 702.600 628.050 703.050 ;
        RECT 562.950 701.400 628.050 702.600 ;
        RECT 562.950 700.950 565.050 701.400 ;
        RECT 577.950 700.950 580.050 701.400 ;
        RECT 625.950 700.950 628.050 701.400 ;
        RECT 643.950 702.600 646.050 703.050 ;
        RECT 649.950 702.600 652.050 703.050 ;
        RECT 664.950 702.600 667.050 703.050 ;
        RECT 643.950 701.400 667.050 702.600 ;
        RECT 643.950 700.950 646.050 701.400 ;
        RECT 649.950 700.950 652.050 701.400 ;
        RECT 664.950 700.950 667.050 701.400 ;
        RECT 670.950 702.600 673.050 703.050 ;
        RECT 679.950 702.600 682.050 703.050 ;
        RECT 670.950 701.400 682.050 702.600 ;
        RECT 670.950 700.950 673.050 701.400 ;
        RECT 679.950 700.950 682.050 701.400 ;
        RECT 703.950 702.600 706.050 703.050 ;
        RECT 754.950 702.600 757.050 703.050 ;
        RECT 703.950 701.400 757.050 702.600 ;
        RECT 703.950 700.950 706.050 701.400 ;
        RECT 754.950 700.950 757.050 701.400 ;
        RECT 760.950 702.600 763.050 703.050 ;
        RECT 775.950 702.600 778.050 703.050 ;
        RECT 760.950 701.400 778.050 702.600 ;
        RECT 797.400 702.600 798.600 703.950 ;
        RECT 814.950 702.600 817.050 703.050 ;
        RECT 797.400 701.400 817.050 702.600 ;
        RECT 818.400 702.600 819.600 703.950 ;
        RECT 832.950 702.600 835.050 703.050 ;
        RECT 818.400 701.400 835.050 702.600 ;
        RECT 760.950 700.950 763.050 701.400 ;
        RECT 775.950 700.950 778.050 701.400 ;
        RECT 814.950 700.950 817.050 701.400 ;
        RECT 832.950 700.950 835.050 701.400 ;
        RECT 40.950 699.600 43.050 700.050 ;
        RECT 38.400 698.400 43.050 699.600 ;
        RECT 40.950 697.950 43.050 698.400 ;
        RECT 67.950 699.600 70.050 700.050 ;
        RECT 79.950 699.600 82.050 700.050 ;
        RECT 67.950 698.400 82.050 699.600 ;
        RECT 67.950 697.950 70.050 698.400 ;
        RECT 79.950 697.950 82.050 698.400 ;
        RECT 130.950 699.600 133.050 700.050 ;
        RECT 184.950 699.600 187.050 700.050 ;
        RECT 130.950 698.400 187.050 699.600 ;
        RECT 130.950 697.950 133.050 698.400 ;
        RECT 184.950 697.950 187.050 698.400 ;
        RECT 241.950 699.600 244.050 700.050 ;
        RECT 256.950 699.600 259.050 700.050 ;
        RECT 241.950 698.400 259.050 699.600 ;
        RECT 241.950 697.950 244.050 698.400 ;
        RECT 256.950 697.950 259.050 698.400 ;
        RECT 268.950 699.600 271.050 700.050 ;
        RECT 292.950 699.600 295.050 700.050 ;
        RECT 268.950 698.400 295.050 699.600 ;
        RECT 268.950 697.950 271.050 698.400 ;
        RECT 292.950 697.950 295.050 698.400 ;
        RECT 313.950 699.600 316.050 700.050 ;
        RECT 328.950 699.600 331.050 700.050 ;
        RECT 337.950 699.600 340.050 700.050 ;
        RECT 340.950 699.600 343.050 700.050 ;
        RECT 313.950 698.400 343.050 699.600 ;
        RECT 313.950 697.950 316.050 698.400 ;
        RECT 328.950 697.950 331.050 698.400 ;
        RECT 337.950 697.950 340.050 698.400 ;
        RECT 340.950 697.950 343.050 698.400 ;
        RECT 358.950 699.600 361.050 700.050 ;
        RECT 385.950 699.600 388.050 700.050 ;
        RECT 394.950 699.600 397.050 700.050 ;
        RECT 409.950 699.600 412.050 700.050 ;
        RECT 358.950 698.400 412.050 699.600 ;
        RECT 358.950 697.950 361.050 698.400 ;
        RECT 385.950 697.950 388.050 698.400 ;
        RECT 394.950 697.950 397.050 698.400 ;
        RECT 409.950 697.950 412.050 698.400 ;
        RECT 415.950 699.600 418.050 700.050 ;
        RECT 463.950 699.600 466.050 700.050 ;
        RECT 475.950 699.600 478.050 700.050 ;
        RECT 415.950 698.400 444.600 699.600 ;
        RECT 415.950 697.950 418.050 698.400 ;
        RECT 16.950 696.600 19.050 697.050 ;
        RECT 28.950 696.600 31.050 697.050 ;
        RECT 16.950 695.400 31.050 696.600 ;
        RECT 16.950 694.950 19.050 695.400 ;
        RECT 28.950 694.950 31.050 695.400 ;
        RECT 34.950 696.600 37.050 697.050 ;
        RECT 46.950 696.600 49.050 697.050 ;
        RECT 34.950 695.400 49.050 696.600 ;
        RECT 34.950 694.950 37.050 695.400 ;
        RECT 46.950 694.950 49.050 695.400 ;
        RECT 52.950 696.600 55.050 697.050 ;
        RECT 67.950 696.600 70.050 697.050 ;
        RECT 52.950 695.400 70.050 696.600 ;
        RECT 52.950 694.950 55.050 695.400 ;
        RECT 67.950 694.950 70.050 695.400 ;
        RECT 157.950 696.600 160.050 697.050 ;
        RECT 169.950 696.600 172.050 697.050 ;
        RECT 181.950 696.600 184.050 697.050 ;
        RECT 157.950 695.400 184.050 696.600 ;
        RECT 157.950 694.950 160.050 695.400 ;
        RECT 169.950 694.950 172.050 695.400 ;
        RECT 181.950 694.950 184.050 695.400 ;
        RECT 187.950 696.600 190.050 697.050 ;
        RECT 205.950 696.600 208.050 697.050 ;
        RECT 187.950 695.400 208.050 696.600 ;
        RECT 187.950 694.950 190.050 695.400 ;
        RECT 205.950 694.950 208.050 695.400 ;
        RECT 226.950 696.600 229.050 697.050 ;
        RECT 238.950 696.600 241.050 697.050 ;
        RECT 226.950 695.400 241.050 696.600 ;
        RECT 226.950 694.950 229.050 695.400 ;
        RECT 238.950 694.950 241.050 695.400 ;
        RECT 256.950 696.600 259.050 697.050 ;
        RECT 304.950 696.600 307.050 697.050 ;
        RECT 256.950 695.400 307.050 696.600 ;
        RECT 256.950 694.950 259.050 695.400 ;
        RECT 304.950 694.950 307.050 695.400 ;
        RECT 325.950 696.600 328.050 697.050 ;
        RECT 415.950 696.600 418.050 697.050 ;
        RECT 325.950 695.400 418.050 696.600 ;
        RECT 443.400 696.600 444.600 698.400 ;
        RECT 463.950 698.400 478.050 699.600 ;
        RECT 463.950 697.950 466.050 698.400 ;
        RECT 475.950 697.950 478.050 698.400 ;
        RECT 529.950 699.600 532.050 700.050 ;
        RECT 541.950 699.600 544.050 700.050 ;
        RECT 529.950 698.400 544.050 699.600 ;
        RECT 529.950 697.950 532.050 698.400 ;
        RECT 541.950 697.950 544.050 698.400 ;
        RECT 598.950 699.600 601.050 700.050 ;
        RECT 685.950 699.600 688.050 700.050 ;
        RECT 598.950 698.400 688.050 699.600 ;
        RECT 598.950 697.950 601.050 698.400 ;
        RECT 685.950 697.950 688.050 698.400 ;
        RECT 805.950 699.600 808.050 700.050 ;
        RECT 814.950 699.600 817.050 700.050 ;
        RECT 805.950 698.400 817.050 699.600 ;
        RECT 805.950 697.950 808.050 698.400 ;
        RECT 814.950 697.950 817.050 698.400 ;
        RECT 835.950 699.600 838.050 700.050 ;
        RECT 838.950 699.600 841.050 700.050 ;
        RECT 853.950 699.600 856.050 700.050 ;
        RECT 835.950 698.400 856.050 699.600 ;
        RECT 835.950 697.950 838.050 698.400 ;
        RECT 838.950 697.950 841.050 698.400 ;
        RECT 853.950 697.950 856.050 698.400 ;
        RECT 475.950 696.600 478.050 697.050 ;
        RECT 443.400 695.400 478.050 696.600 ;
        RECT 325.950 694.950 328.050 695.400 ;
        RECT 415.950 694.950 418.050 695.400 ;
        RECT 475.950 694.950 478.050 695.400 ;
        RECT 487.950 696.600 490.050 697.050 ;
        RECT 517.950 696.600 520.050 697.050 ;
        RECT 487.950 695.400 520.050 696.600 ;
        RECT 487.950 694.950 490.050 695.400 ;
        RECT 517.950 694.950 520.050 695.400 ;
        RECT 523.950 696.600 526.050 697.050 ;
        RECT 544.950 696.600 547.050 697.050 ;
        RECT 523.950 695.400 547.050 696.600 ;
        RECT 523.950 694.950 526.050 695.400 ;
        RECT 544.950 694.950 547.050 695.400 ;
        RECT 559.950 696.600 562.050 697.050 ;
        RECT 571.950 696.600 574.050 697.050 ;
        RECT 559.950 695.400 574.050 696.600 ;
        RECT 559.950 694.950 562.050 695.400 ;
        RECT 571.950 694.950 574.050 695.400 ;
        RECT 583.950 696.600 586.050 697.050 ;
        RECT 610.950 696.600 613.050 697.050 ;
        RECT 583.950 695.400 613.050 696.600 ;
        RECT 583.950 694.950 586.050 695.400 ;
        RECT 610.950 694.950 613.050 695.400 ;
        RECT 619.950 696.600 622.050 697.050 ;
        RECT 625.950 696.600 628.050 697.050 ;
        RECT 619.950 695.400 628.050 696.600 ;
        RECT 619.950 694.950 622.050 695.400 ;
        RECT 625.950 694.950 628.050 695.400 ;
        RECT 667.950 696.600 670.050 697.050 ;
        RECT 688.950 696.600 691.050 697.050 ;
        RECT 700.950 696.600 703.050 697.050 ;
        RECT 709.950 696.600 712.050 697.050 ;
        RECT 667.950 695.400 712.050 696.600 ;
        RECT 667.950 694.950 670.050 695.400 ;
        RECT 688.950 694.950 691.050 695.400 ;
        RECT 700.950 694.950 703.050 695.400 ;
        RECT 709.950 694.950 712.050 695.400 ;
        RECT 730.950 696.600 733.050 697.050 ;
        RECT 757.950 696.600 760.050 697.050 ;
        RECT 730.950 695.400 760.050 696.600 ;
        RECT 730.950 694.950 733.050 695.400 ;
        RECT 757.950 694.950 760.050 695.400 ;
        RECT 778.950 696.600 781.050 697.050 ;
        RECT 799.950 696.600 802.050 697.050 ;
        RECT 778.950 695.400 802.050 696.600 ;
        RECT 778.950 694.950 781.050 695.400 ;
        RECT 799.950 694.950 802.050 695.400 ;
        RECT 802.950 696.600 805.050 697.050 ;
        RECT 817.950 696.600 820.050 697.050 ;
        RECT 802.950 695.400 820.050 696.600 ;
        RECT 802.950 694.950 805.050 695.400 ;
        RECT 817.950 694.950 820.050 695.400 ;
        RECT 37.950 693.600 40.050 694.050 ;
        RECT 52.950 693.600 55.050 694.050 ;
        RECT 37.950 692.400 55.050 693.600 ;
        RECT 37.950 691.950 40.050 692.400 ;
        RECT 52.950 691.950 55.050 692.400 ;
        RECT 196.950 693.600 199.050 694.050 ;
        RECT 220.950 693.600 223.050 694.050 ;
        RECT 196.950 692.400 223.050 693.600 ;
        RECT 196.950 691.950 199.050 692.400 ;
        RECT 220.950 691.950 223.050 692.400 ;
        RECT 238.950 693.600 241.050 694.050 ;
        RECT 346.950 693.600 349.050 694.050 ;
        RECT 400.950 693.600 403.050 694.050 ;
        RECT 238.950 692.400 336.600 693.600 ;
        RECT 238.950 691.950 241.050 692.400 ;
        RECT 76.950 690.600 79.050 691.050 ;
        RECT 124.950 690.600 127.050 691.050 ;
        RECT 133.950 690.600 136.050 691.050 ;
        RECT 250.950 690.600 253.050 691.050 ;
        RECT 76.950 689.400 253.050 690.600 ;
        RECT 335.400 690.600 336.600 692.400 ;
        RECT 346.950 692.400 403.050 693.600 ;
        RECT 346.950 691.950 349.050 692.400 ;
        RECT 400.950 691.950 403.050 692.400 ;
        RECT 436.950 693.600 439.050 694.050 ;
        RECT 502.950 693.600 505.050 694.050 ;
        RECT 436.950 692.400 505.050 693.600 ;
        RECT 436.950 691.950 439.050 692.400 ;
        RECT 502.950 691.950 505.050 692.400 ;
        RECT 565.950 693.600 568.050 694.050 ;
        RECT 583.950 693.600 586.050 694.050 ;
        RECT 637.950 693.600 640.050 694.050 ;
        RECT 565.950 692.400 586.050 693.600 ;
        RECT 565.950 691.950 568.050 692.400 ;
        RECT 583.950 691.950 586.050 692.400 ;
        RECT 614.400 692.400 640.050 693.600 ;
        RECT 376.950 690.600 379.050 691.050 ;
        RECT 335.400 689.400 379.050 690.600 ;
        RECT 76.950 688.950 79.050 689.400 ;
        RECT 124.950 688.950 127.050 689.400 ;
        RECT 133.950 688.950 136.050 689.400 ;
        RECT 250.950 688.950 253.050 689.400 ;
        RECT 376.950 688.950 379.050 689.400 ;
        RECT 400.950 690.600 403.050 691.050 ;
        RECT 493.950 690.600 496.050 691.050 ;
        RECT 547.950 690.600 550.050 691.050 ;
        RECT 400.950 689.400 550.050 690.600 ;
        RECT 400.950 688.950 403.050 689.400 ;
        RECT 493.950 688.950 496.050 689.400 ;
        RECT 547.950 688.950 550.050 689.400 ;
        RECT 556.950 690.600 559.050 691.050 ;
        RECT 589.950 690.600 592.050 691.050 ;
        RECT 556.950 689.400 592.050 690.600 ;
        RECT 556.950 688.950 559.050 689.400 ;
        RECT 589.950 688.950 592.050 689.400 ;
        RECT 604.950 690.600 607.050 691.050 ;
        RECT 614.400 690.600 615.600 692.400 ;
        RECT 637.950 691.950 640.050 692.400 ;
        RECT 751.950 693.600 754.050 694.050 ;
        RECT 826.950 693.600 829.050 694.050 ;
        RECT 856.950 693.600 859.050 694.050 ;
        RECT 751.950 692.400 859.050 693.600 ;
        RECT 751.950 691.950 754.050 692.400 ;
        RECT 826.950 691.950 829.050 692.400 ;
        RECT 856.950 691.950 859.050 692.400 ;
        RECT 604.950 689.400 615.600 690.600 ;
        RECT 634.950 690.600 637.050 691.050 ;
        RECT 679.950 690.600 682.050 691.050 ;
        RECT 634.950 689.400 682.050 690.600 ;
        RECT 604.950 688.950 607.050 689.400 ;
        RECT 634.950 688.950 637.050 689.400 ;
        RECT 679.950 688.950 682.050 689.400 ;
        RECT 733.950 690.600 736.050 691.050 ;
        RECT 760.950 690.600 763.050 691.050 ;
        RECT 733.950 689.400 763.050 690.600 ;
        RECT 733.950 688.950 736.050 689.400 ;
        RECT 760.950 688.950 763.050 689.400 ;
        RECT 19.950 687.600 22.050 688.050 ;
        RECT 73.950 687.600 76.050 688.050 ;
        RECT 19.950 686.400 76.050 687.600 ;
        RECT 19.950 685.950 22.050 686.400 ;
        RECT 73.950 685.950 76.050 686.400 ;
        RECT 205.950 687.600 208.050 688.050 ;
        RECT 214.950 687.600 217.050 688.050 ;
        RECT 205.950 686.400 217.050 687.600 ;
        RECT 205.950 685.950 208.050 686.400 ;
        RECT 214.950 685.950 217.050 686.400 ;
        RECT 274.950 687.600 277.050 688.050 ;
        RECT 313.950 687.600 316.050 688.050 ;
        RECT 274.950 686.400 316.050 687.600 ;
        RECT 274.950 685.950 277.050 686.400 ;
        RECT 313.950 685.950 316.050 686.400 ;
        RECT 367.950 687.600 370.050 688.050 ;
        RECT 400.950 687.600 403.050 688.050 ;
        RECT 433.950 687.600 436.050 688.050 ;
        RECT 451.950 687.600 454.050 688.050 ;
        RECT 367.950 686.400 454.050 687.600 ;
        RECT 367.950 685.950 370.050 686.400 ;
        RECT 400.950 685.950 403.050 686.400 ;
        RECT 433.950 685.950 436.050 686.400 ;
        RECT 451.950 685.950 454.050 686.400 ;
        RECT 634.950 687.600 637.050 688.050 ;
        RECT 682.950 687.600 685.050 688.050 ;
        RECT 724.950 687.600 727.050 688.050 ;
        RECT 634.950 686.400 727.050 687.600 ;
        RECT 634.950 685.950 637.050 686.400 ;
        RECT 682.950 685.950 685.050 686.400 ;
        RECT 724.950 685.950 727.050 686.400 ;
        RECT 34.950 684.600 37.050 685.050 ;
        RECT 61.950 684.600 64.050 685.050 ;
        RECT 103.950 684.600 106.050 685.050 ;
        RECT 34.950 683.400 106.050 684.600 ;
        RECT 34.950 682.950 37.050 683.400 ;
        RECT 61.950 682.950 64.050 683.400 ;
        RECT 103.950 682.950 106.050 683.400 ;
        RECT 148.950 684.600 151.050 685.050 ;
        RECT 289.950 684.600 292.050 685.050 ;
        RECT 148.950 683.400 292.050 684.600 ;
        RECT 148.950 682.950 151.050 683.400 ;
        RECT 289.950 682.950 292.050 683.400 ;
        RECT 340.950 684.600 343.050 685.050 ;
        RECT 388.950 684.600 391.050 685.050 ;
        RECT 340.950 683.400 391.050 684.600 ;
        RECT 340.950 682.950 343.050 683.400 ;
        RECT 388.950 682.950 391.050 683.400 ;
        RECT 412.950 684.600 415.050 685.050 ;
        RECT 424.950 684.600 427.050 685.050 ;
        RECT 481.950 684.600 484.050 685.050 ;
        RECT 412.950 683.400 484.050 684.600 ;
        RECT 412.950 682.950 415.050 683.400 ;
        RECT 424.950 682.950 427.050 683.400 ;
        RECT 481.950 682.950 484.050 683.400 ;
        RECT 571.950 684.600 574.050 685.050 ;
        RECT 589.950 684.600 592.050 685.050 ;
        RECT 793.950 684.600 796.050 685.050 ;
        RECT 571.950 683.400 796.050 684.600 ;
        RECT 571.950 682.950 574.050 683.400 ;
        RECT 589.950 682.950 592.050 683.400 ;
        RECT 793.950 682.950 796.050 683.400 ;
        RECT 73.950 681.600 76.050 682.050 ;
        RECT 85.950 681.600 88.050 682.050 ;
        RECT 73.950 680.400 88.050 681.600 ;
        RECT 73.950 679.950 76.050 680.400 ;
        RECT 85.950 679.950 88.050 680.400 ;
        RECT 94.950 681.600 97.050 682.050 ;
        RECT 97.950 681.600 100.050 682.050 ;
        RECT 127.950 681.600 130.050 682.050 ;
        RECT 139.950 681.600 142.050 682.050 ;
        RECT 94.950 680.400 142.050 681.600 ;
        RECT 94.950 679.950 97.050 680.400 ;
        RECT 97.950 679.950 100.050 680.400 ;
        RECT 127.950 679.950 130.050 680.400 ;
        RECT 139.950 679.950 142.050 680.400 ;
        RECT 190.950 681.600 193.050 682.050 ;
        RECT 208.950 681.600 211.050 682.050 ;
        RECT 214.950 681.600 217.050 682.050 ;
        RECT 262.950 681.600 265.050 682.050 ;
        RECT 190.950 680.400 265.050 681.600 ;
        RECT 190.950 679.950 193.050 680.400 ;
        RECT 208.950 679.950 211.050 680.400 ;
        RECT 214.950 679.950 217.050 680.400 ;
        RECT 262.950 679.950 265.050 680.400 ;
        RECT 271.950 681.600 274.050 682.050 ;
        RECT 325.950 681.600 328.050 682.050 ;
        RECT 271.950 680.400 328.050 681.600 ;
        RECT 271.950 679.950 274.050 680.400 ;
        RECT 325.950 679.950 328.050 680.400 ;
        RECT 481.950 681.600 484.050 682.050 ;
        RECT 487.950 681.600 490.050 682.050 ;
        RECT 481.950 680.400 490.050 681.600 ;
        RECT 481.950 679.950 484.050 680.400 ;
        RECT 487.950 679.950 490.050 680.400 ;
        RECT 616.950 681.600 619.050 682.050 ;
        RECT 646.950 681.600 649.050 682.050 ;
        RECT 670.950 681.600 673.050 682.050 ;
        RECT 616.950 680.400 673.050 681.600 ;
        RECT 616.950 679.950 619.050 680.400 ;
        RECT 646.950 679.950 649.050 680.400 ;
        RECT 670.950 679.950 673.050 680.400 ;
        RECT 85.950 678.600 88.050 679.050 ;
        RECT 106.950 678.600 109.050 679.050 ;
        RECT 85.950 677.400 109.050 678.600 ;
        RECT 85.950 676.950 88.050 677.400 ;
        RECT 106.950 676.950 109.050 677.400 ;
        RECT 133.950 678.600 136.050 679.050 ;
        RECT 229.950 678.600 232.050 679.050 ;
        RECT 133.950 677.400 232.050 678.600 ;
        RECT 133.950 676.950 136.050 677.400 ;
        RECT 229.950 676.950 232.050 677.400 ;
        RECT 247.950 678.600 250.050 679.050 ;
        RECT 295.950 678.600 298.050 679.050 ;
        RECT 247.950 677.400 298.050 678.600 ;
        RECT 247.950 676.950 250.050 677.400 ;
        RECT 295.950 676.950 298.050 677.400 ;
        RECT 301.950 678.600 304.050 679.050 ;
        RECT 373.950 678.600 376.050 679.050 ;
        RECT 385.950 678.600 388.050 679.050 ;
        RECT 301.950 677.400 388.050 678.600 ;
        RECT 301.950 676.950 304.050 677.400 ;
        RECT 373.950 676.950 376.050 677.400 ;
        RECT 385.950 676.950 388.050 677.400 ;
        RECT 430.950 678.600 433.050 679.050 ;
        RECT 436.950 678.600 439.050 679.050 ;
        RECT 430.950 677.400 439.050 678.600 ;
        RECT 430.950 676.950 433.050 677.400 ;
        RECT 436.950 676.950 439.050 677.400 ;
        RECT 466.950 678.600 469.050 679.050 ;
        RECT 517.950 678.600 520.050 679.050 ;
        RECT 520.950 678.600 523.050 679.050 ;
        RECT 466.950 677.400 523.050 678.600 ;
        RECT 466.950 676.950 469.050 677.400 ;
        RECT 517.950 676.950 520.050 677.400 ;
        RECT 520.950 676.950 523.050 677.400 ;
        RECT 547.950 678.600 550.050 679.050 ;
        RECT 607.950 678.600 610.050 679.050 ;
        RECT 613.950 678.600 616.050 679.050 ;
        RECT 547.950 677.400 616.050 678.600 ;
        RECT 547.950 676.950 550.050 677.400 ;
        RECT 607.950 676.950 610.050 677.400 ;
        RECT 613.950 676.950 616.050 677.400 ;
        RECT 670.950 678.600 673.050 679.050 ;
        RECT 763.950 678.600 766.050 679.050 ;
        RECT 670.950 677.400 766.050 678.600 ;
        RECT 670.950 676.950 673.050 677.400 ;
        RECT 763.950 676.950 766.050 677.400 ;
        RECT 772.950 678.600 775.050 679.050 ;
        RECT 781.950 678.600 784.050 679.050 ;
        RECT 772.950 677.400 784.050 678.600 ;
        RECT 772.950 676.950 775.050 677.400 ;
        RECT 781.950 676.950 784.050 677.400 ;
        RECT 823.950 678.600 826.050 679.050 ;
        RECT 838.950 678.600 841.050 679.050 ;
        RECT 823.950 677.400 841.050 678.600 ;
        RECT 823.950 676.950 826.050 677.400 ;
        RECT 838.950 676.950 841.050 677.400 ;
        RECT 7.950 673.950 10.050 676.050 ;
        RECT 13.950 675.600 16.050 676.050 ;
        RECT 22.950 675.600 25.050 676.050 ;
        RECT 13.950 674.400 25.050 675.600 ;
        RECT 13.950 673.950 16.050 674.400 ;
        RECT 22.950 673.950 25.050 674.400 ;
        RECT 37.950 675.600 40.050 676.050 ;
        RECT 52.950 675.600 55.050 676.050 ;
        RECT 37.950 674.400 55.050 675.600 ;
        RECT 37.950 673.950 40.050 674.400 ;
        RECT 52.950 673.950 55.050 674.400 ;
        RECT 100.950 675.600 103.050 676.050 ;
        RECT 115.950 675.600 118.050 676.050 ;
        RECT 121.950 675.600 124.050 676.050 ;
        RECT 133.950 675.600 136.050 676.050 ;
        RECT 100.950 674.400 136.050 675.600 ;
        RECT 100.950 673.950 103.050 674.400 ;
        RECT 115.950 673.950 118.050 674.400 ;
        RECT 121.950 673.950 124.050 674.400 ;
        RECT 133.950 673.950 136.050 674.400 ;
        RECT 175.950 675.600 178.050 676.050 ;
        RECT 190.950 675.600 193.050 676.050 ;
        RECT 196.950 675.600 199.050 676.050 ;
        RECT 175.950 674.400 193.050 675.600 ;
        RECT 175.950 673.950 178.050 674.400 ;
        RECT 190.950 673.950 193.050 674.400 ;
        RECT 194.400 674.400 199.050 675.600 ;
        RECT 8.400 663.600 9.600 673.950 ;
        RECT 43.950 672.600 46.050 673.050 ;
        RECT 58.950 672.600 61.050 673.050 ;
        RECT 17.400 671.400 61.050 672.600 ;
        RECT 17.400 670.050 18.600 671.400 ;
        RECT 43.950 670.950 46.050 671.400 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 88.950 672.600 91.050 673.050 ;
        RECT 100.950 672.600 103.050 673.050 ;
        RECT 88.950 671.400 103.050 672.600 ;
        RECT 88.950 670.950 91.050 671.400 ;
        RECT 100.950 670.950 103.050 671.400 ;
        RECT 106.950 672.600 109.050 673.050 ;
        RECT 139.950 672.600 142.050 673.050 ;
        RECT 151.950 672.600 154.050 673.050 ;
        RECT 106.950 671.400 123.600 672.600 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 10.950 667.950 13.050 670.050 ;
        RECT 16.950 667.950 19.050 670.050 ;
        RECT 40.950 669.600 43.050 670.050 ;
        RECT 49.950 669.600 52.050 670.050 ;
        RECT 40.950 668.400 52.050 669.600 ;
        RECT 40.950 667.950 43.050 668.400 ;
        RECT 49.950 667.950 52.050 668.400 ;
        RECT 55.950 669.600 58.050 670.050 ;
        RECT 61.950 669.600 64.050 670.050 ;
        RECT 55.950 668.400 64.050 669.600 ;
        RECT 55.950 667.950 58.050 668.400 ;
        RECT 61.950 667.950 64.050 668.400 ;
        RECT 82.950 669.600 85.050 670.050 ;
        RECT 103.950 669.600 106.050 670.050 ;
        RECT 118.950 669.600 121.050 670.050 ;
        RECT 82.950 668.400 121.050 669.600 ;
        RECT 122.400 669.600 123.600 671.400 ;
        RECT 139.950 671.400 154.050 672.600 ;
        RECT 139.950 670.950 142.050 671.400 ;
        RECT 151.950 670.950 154.050 671.400 ;
        RECT 175.950 672.600 178.050 673.050 ;
        RECT 194.400 672.600 195.600 674.400 ;
        RECT 196.950 673.950 199.050 674.400 ;
        RECT 268.950 675.600 271.050 676.050 ;
        RECT 331.950 675.600 334.050 676.050 ;
        RECT 268.950 674.400 334.050 675.600 ;
        RECT 268.950 673.950 271.050 674.400 ;
        RECT 331.950 673.950 334.050 674.400 ;
        RECT 370.950 675.600 373.050 676.050 ;
        RECT 391.950 675.600 394.050 676.050 ;
        RECT 370.950 674.400 394.050 675.600 ;
        RECT 370.950 673.950 373.050 674.400 ;
        RECT 391.950 673.950 394.050 674.400 ;
        RECT 406.950 675.600 409.050 676.050 ;
        RECT 427.950 675.600 430.050 676.050 ;
        RECT 406.950 674.400 430.050 675.600 ;
        RECT 406.950 673.950 409.050 674.400 ;
        RECT 427.950 673.950 430.050 674.400 ;
        RECT 451.950 675.600 454.050 676.050 ;
        RECT 469.950 675.600 472.050 676.050 ;
        RECT 481.950 675.600 484.050 676.050 ;
        RECT 496.950 675.600 499.050 676.050 ;
        RECT 451.950 674.400 499.050 675.600 ;
        RECT 451.950 673.950 454.050 674.400 ;
        RECT 469.950 673.950 472.050 674.400 ;
        RECT 481.950 673.950 484.050 674.400 ;
        RECT 496.950 673.950 499.050 674.400 ;
        RECT 526.950 675.600 529.050 676.050 ;
        RECT 583.950 675.600 586.050 676.050 ;
        RECT 526.950 674.400 586.050 675.600 ;
        RECT 526.950 673.950 529.050 674.400 ;
        RECT 583.950 673.950 586.050 674.400 ;
        RECT 601.950 675.600 604.050 676.050 ;
        RECT 616.950 675.600 619.050 676.050 ;
        RECT 601.950 674.400 619.050 675.600 ;
        RECT 601.950 673.950 604.050 674.400 ;
        RECT 616.950 673.950 619.050 674.400 ;
        RECT 727.950 675.600 730.050 676.050 ;
        RECT 775.950 675.600 778.050 676.050 ;
        RECT 799.950 675.600 802.050 676.050 ;
        RECT 727.950 674.400 802.050 675.600 ;
        RECT 727.950 673.950 730.050 674.400 ;
        RECT 775.950 673.950 778.050 674.400 ;
        RECT 799.950 673.950 802.050 674.400 ;
        RECT 823.950 673.950 826.050 676.050 ;
        RECT 175.950 671.400 195.600 672.600 ;
        RECT 217.950 672.600 220.050 673.050 ;
        RECT 223.950 672.600 226.050 673.050 ;
        RECT 217.950 671.400 226.050 672.600 ;
        RECT 175.950 670.950 178.050 671.400 ;
        RECT 217.950 670.950 220.050 671.400 ;
        RECT 223.950 670.950 226.050 671.400 ;
        RECT 232.950 672.600 235.050 673.050 ;
        RECT 286.950 672.600 289.050 673.050 ;
        RECT 301.950 672.600 304.050 673.050 ;
        RECT 232.950 671.400 304.050 672.600 ;
        RECT 232.950 670.950 235.050 671.400 ;
        RECT 286.950 670.950 289.050 671.400 ;
        RECT 301.950 670.950 304.050 671.400 ;
        RECT 304.950 672.600 307.050 673.050 ;
        RECT 325.950 672.600 328.050 673.050 ;
        RECT 304.950 671.400 328.050 672.600 ;
        RECT 304.950 670.950 307.050 671.400 ;
        RECT 325.950 670.950 328.050 671.400 ;
        RECT 331.950 672.600 334.050 673.050 ;
        RECT 430.950 672.600 433.050 673.050 ;
        RECT 448.950 672.600 451.050 673.050 ;
        RECT 331.950 671.400 414.600 672.600 ;
        RECT 331.950 670.950 334.050 671.400 ;
        RECT 413.400 670.050 414.600 671.400 ;
        RECT 430.950 671.400 451.050 672.600 ;
        RECT 430.950 670.950 433.050 671.400 ;
        RECT 448.950 670.950 451.050 671.400 ;
        RECT 502.950 670.950 505.050 673.050 ;
        RECT 505.950 672.600 508.050 673.050 ;
        RECT 529.950 672.600 532.050 673.050 ;
        RECT 538.950 672.600 541.050 673.050 ;
        RECT 544.950 672.600 547.050 673.050 ;
        RECT 505.950 671.400 537.600 672.600 ;
        RECT 505.950 670.950 508.050 671.400 ;
        RECT 529.950 670.950 532.050 671.400 ;
        RECT 136.950 669.600 139.050 670.050 ;
        RECT 148.950 669.600 151.050 670.050 ;
        RECT 122.400 668.400 151.050 669.600 ;
        RECT 82.950 667.950 85.050 668.400 ;
        RECT 103.950 667.950 106.050 668.400 ;
        RECT 118.950 667.950 121.050 668.400 ;
        RECT 136.950 667.950 139.050 668.400 ;
        RECT 148.950 667.950 151.050 668.400 ;
        RECT 154.950 669.600 157.050 670.050 ;
        RECT 172.950 669.600 175.050 670.050 ;
        RECT 154.950 668.400 175.050 669.600 ;
        RECT 154.950 667.950 157.050 668.400 ;
        RECT 172.950 667.950 175.050 668.400 ;
        RECT 178.950 669.600 181.050 670.050 ;
        RECT 199.950 669.600 202.050 670.050 ;
        RECT 211.950 669.600 214.050 670.050 ;
        RECT 178.950 668.400 214.050 669.600 ;
        RECT 178.950 667.950 181.050 668.400 ;
        RECT 199.950 667.950 202.050 668.400 ;
        RECT 211.950 667.950 214.050 668.400 ;
        RECT 214.950 669.600 217.050 670.050 ;
        RECT 256.950 669.600 259.050 670.050 ;
        RECT 214.950 668.400 259.050 669.600 ;
        RECT 214.950 667.950 217.050 668.400 ;
        RECT 256.950 667.950 259.050 668.400 ;
        RECT 274.950 669.600 277.050 670.050 ;
        RECT 289.950 669.600 292.050 670.050 ;
        RECT 274.950 668.400 292.050 669.600 ;
        RECT 274.950 667.950 277.050 668.400 ;
        RECT 289.950 667.950 292.050 668.400 ;
        RECT 307.950 669.600 310.050 670.050 ;
        RECT 322.950 669.600 325.050 670.050 ;
        RECT 307.950 668.400 325.050 669.600 ;
        RECT 307.950 667.950 310.050 668.400 ;
        RECT 322.950 667.950 325.050 668.400 ;
        RECT 352.950 669.600 355.050 670.050 ;
        RECT 361.950 669.600 364.050 670.050 ;
        RECT 352.950 668.400 364.050 669.600 ;
        RECT 352.950 667.950 355.050 668.400 ;
        RECT 361.950 667.950 364.050 668.400 ;
        RECT 364.950 669.600 367.050 670.050 ;
        RECT 370.950 669.600 373.050 670.050 ;
        RECT 364.950 668.400 373.050 669.600 ;
        RECT 364.950 667.950 367.050 668.400 ;
        RECT 370.950 667.950 373.050 668.400 ;
        RECT 376.950 669.600 379.050 670.050 ;
        RECT 409.950 669.600 412.050 670.050 ;
        RECT 376.950 668.400 412.050 669.600 ;
        RECT 376.950 667.950 379.050 668.400 ;
        RECT 409.950 667.950 412.050 668.400 ;
        RECT 412.950 667.950 415.050 670.050 ;
        RECT 439.950 669.600 442.050 670.050 ;
        RECT 445.950 669.600 448.050 670.050 ;
        RECT 439.950 668.400 448.050 669.600 ;
        RECT 503.400 669.600 504.600 670.950 ;
        RECT 532.950 669.600 535.050 670.050 ;
        RECT 503.400 668.400 535.050 669.600 ;
        RECT 536.400 669.600 537.600 671.400 ;
        RECT 538.950 671.400 547.050 672.600 ;
        RECT 538.950 670.950 541.050 671.400 ;
        RECT 544.950 670.950 547.050 671.400 ;
        RECT 553.950 672.600 556.050 673.050 ;
        RECT 568.950 672.600 571.050 673.050 ;
        RECT 553.950 671.400 571.050 672.600 ;
        RECT 553.950 670.950 556.050 671.400 ;
        RECT 568.950 670.950 571.050 671.400 ;
        RECT 637.950 672.600 640.050 673.050 ;
        RECT 658.950 672.600 661.050 673.050 ;
        RECT 637.950 671.400 661.050 672.600 ;
        RECT 637.950 670.950 640.050 671.400 ;
        RECT 658.950 670.950 661.050 671.400 ;
        RECT 661.950 672.600 664.050 673.050 ;
        RECT 730.950 672.600 733.050 673.050 ;
        RECT 739.950 672.600 742.050 673.050 ;
        RECT 745.950 672.600 748.050 673.050 ;
        RECT 661.950 671.400 678.600 672.600 ;
        RECT 661.950 670.950 664.050 671.400 ;
        RECT 562.950 669.600 565.050 670.050 ;
        RECT 536.400 668.400 565.050 669.600 ;
        RECT 439.950 667.950 442.050 668.400 ;
        RECT 445.950 667.950 448.050 668.400 ;
        RECT 532.950 667.950 535.050 668.400 ;
        RECT 11.400 666.600 12.600 667.950 ;
        RECT 548.400 667.050 549.600 668.400 ;
        RECT 562.950 667.950 565.050 668.400 ;
        RECT 571.950 669.600 574.050 670.050 ;
        RECT 577.950 669.600 580.050 670.050 ;
        RECT 571.950 668.400 580.050 669.600 ;
        RECT 571.950 667.950 574.050 668.400 ;
        RECT 577.950 667.950 580.050 668.400 ;
        RECT 643.950 669.600 646.050 670.050 ;
        RECT 652.950 669.600 655.050 670.050 ;
        RECT 658.950 669.600 661.050 670.050 ;
        RECT 643.950 668.400 661.050 669.600 ;
        RECT 643.950 667.950 646.050 668.400 ;
        RECT 652.950 667.950 655.050 668.400 ;
        RECT 658.950 667.950 661.050 668.400 ;
        RECT 677.400 667.050 678.600 671.400 ;
        RECT 730.950 671.400 748.050 672.600 ;
        RECT 730.950 670.950 733.050 671.400 ;
        RECT 739.950 670.950 742.050 671.400 ;
        RECT 745.950 670.950 748.050 671.400 ;
        RECT 781.950 672.600 784.050 673.050 ;
        RECT 808.950 672.600 811.050 673.050 ;
        RECT 781.950 671.400 811.050 672.600 ;
        RECT 781.950 670.950 784.050 671.400 ;
        RECT 808.950 670.950 811.050 671.400 ;
        RECT 769.950 669.600 772.050 670.050 ;
        RECT 824.400 669.600 825.600 673.950 ;
        RECT 850.950 670.950 853.050 673.050 ;
        RECT 769.950 668.400 825.600 669.600 ;
        RECT 769.950 667.950 772.050 668.400 ;
        RECT 851.400 667.050 852.600 670.950 ;
        RECT 25.950 666.600 28.050 667.050 ;
        RECT 31.950 666.600 34.050 667.050 ;
        RECT 11.400 665.400 34.050 666.600 ;
        RECT 25.950 664.950 28.050 665.400 ;
        RECT 31.950 664.950 34.050 665.400 ;
        RECT 37.950 664.950 40.050 667.050 ;
        RECT 49.950 666.600 52.050 667.050 ;
        RECT 58.950 666.600 61.050 667.050 ;
        RECT 49.950 665.400 61.050 666.600 ;
        RECT 49.950 664.950 52.050 665.400 ;
        RECT 58.950 664.950 61.050 665.400 ;
        RECT 67.950 666.600 70.050 667.050 ;
        RECT 79.950 666.600 82.050 667.050 ;
        RECT 67.950 665.400 82.050 666.600 ;
        RECT 67.950 664.950 70.050 665.400 ;
        RECT 79.950 664.950 82.050 665.400 ;
        RECT 160.950 666.600 163.050 667.050 ;
        RECT 193.950 666.600 196.050 667.050 ;
        RECT 202.950 666.600 205.050 667.050 ;
        RECT 271.950 666.600 274.050 667.050 ;
        RECT 160.950 665.400 205.050 666.600 ;
        RECT 160.950 664.950 163.050 665.400 ;
        RECT 193.950 664.950 196.050 665.400 ;
        RECT 202.950 664.950 205.050 665.400 ;
        RECT 269.400 665.400 274.050 666.600 ;
        RECT 10.950 663.600 13.050 664.050 ;
        RECT 8.400 662.400 13.050 663.600 ;
        RECT 38.400 663.600 39.600 664.950 ;
        RECT 269.400 664.050 270.600 665.400 ;
        RECT 271.950 664.950 274.050 665.400 ;
        RECT 310.950 664.950 313.050 667.050 ;
        RECT 388.950 666.600 391.050 667.050 ;
        RECT 406.950 666.600 409.050 667.050 ;
        RECT 388.950 665.400 409.050 666.600 ;
        RECT 388.950 664.950 391.050 665.400 ;
        RECT 406.950 664.950 409.050 665.400 ;
        RECT 448.950 666.600 451.050 667.050 ;
        RECT 499.950 666.600 502.050 667.050 ;
        RECT 538.950 666.600 541.050 667.050 ;
        RECT 448.950 665.400 541.050 666.600 ;
        RECT 448.950 664.950 451.050 665.400 ;
        RECT 499.950 664.950 502.050 665.400 ;
        RECT 538.950 664.950 541.050 665.400 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 553.950 666.600 556.050 667.050 ;
        RECT 580.950 666.600 583.050 667.050 ;
        RECT 553.950 665.400 583.050 666.600 ;
        RECT 553.950 664.950 556.050 665.400 ;
        RECT 580.950 664.950 583.050 665.400 ;
        RECT 604.950 666.600 607.050 667.050 ;
        RECT 640.950 666.600 643.050 667.050 ;
        RECT 604.950 665.400 643.050 666.600 ;
        RECT 604.950 664.950 607.050 665.400 ;
        RECT 640.950 664.950 643.050 665.400 ;
        RECT 664.950 666.600 667.050 667.050 ;
        RECT 673.950 666.600 676.050 667.050 ;
        RECT 664.950 665.400 676.050 666.600 ;
        RECT 664.950 664.950 667.050 665.400 ;
        RECT 673.950 664.950 676.050 665.400 ;
        RECT 676.950 664.950 679.050 667.050 ;
        RECT 715.950 666.600 718.050 667.050 ;
        RECT 733.950 666.600 736.050 667.050 ;
        RECT 715.950 665.400 736.050 666.600 ;
        RECT 715.950 664.950 718.050 665.400 ;
        RECT 733.950 664.950 736.050 665.400 ;
        RECT 739.950 666.600 742.050 667.050 ;
        RECT 751.950 666.600 754.050 667.050 ;
        RECT 739.950 665.400 754.050 666.600 ;
        RECT 739.950 664.950 742.050 665.400 ;
        RECT 751.950 664.950 754.050 665.400 ;
        RECT 802.950 666.600 805.050 667.050 ;
        RECT 820.950 666.600 823.050 667.050 ;
        RECT 802.950 665.400 823.050 666.600 ;
        RECT 802.950 664.950 805.050 665.400 ;
        RECT 820.950 664.950 823.050 665.400 ;
        RECT 850.950 664.950 853.050 667.050 ;
        RECT 49.950 663.600 52.050 664.050 ;
        RECT 38.400 662.400 52.050 663.600 ;
        RECT 10.950 661.950 13.050 662.400 ;
        RECT 49.950 661.950 52.050 662.400 ;
        RECT 163.950 663.600 166.050 664.050 ;
        RECT 172.950 663.600 175.050 664.050 ;
        RECT 163.950 662.400 175.050 663.600 ;
        RECT 163.950 661.950 166.050 662.400 ;
        RECT 172.950 661.950 175.050 662.400 ;
        RECT 226.950 663.600 229.050 664.050 ;
        RECT 232.950 663.600 235.050 664.050 ;
        RECT 238.950 663.600 241.050 664.050 ;
        RECT 226.950 662.400 241.050 663.600 ;
        RECT 226.950 661.950 229.050 662.400 ;
        RECT 232.950 661.950 235.050 662.400 ;
        RECT 238.950 661.950 241.050 662.400 ;
        RECT 268.950 661.950 271.050 664.050 ;
        RECT 307.950 663.600 310.050 664.050 ;
        RECT 311.400 663.600 312.600 664.950 ;
        RECT 307.950 662.400 312.600 663.600 ;
        RECT 349.950 663.600 352.050 664.050 ;
        RECT 544.950 663.600 547.050 664.050 ;
        RECT 349.950 662.400 547.050 663.600 ;
        RECT 307.950 661.950 310.050 662.400 ;
        RECT 349.950 661.950 352.050 662.400 ;
        RECT 544.950 661.950 547.050 662.400 ;
        RECT 622.950 663.600 625.050 664.050 ;
        RECT 655.950 663.600 658.050 664.050 ;
        RECT 622.950 662.400 658.050 663.600 ;
        RECT 622.950 661.950 625.050 662.400 ;
        RECT 655.950 661.950 658.050 662.400 ;
        RECT 718.950 663.600 721.050 664.050 ;
        RECT 748.950 663.600 751.050 664.050 ;
        RECT 718.950 662.400 751.050 663.600 ;
        RECT 718.950 661.950 721.050 662.400 ;
        RECT 748.950 661.950 751.050 662.400 ;
        RECT 757.950 663.600 760.050 664.050 ;
        RECT 778.950 663.600 781.050 664.050 ;
        RECT 757.950 662.400 781.050 663.600 ;
        RECT 757.950 661.950 760.050 662.400 ;
        RECT 778.950 661.950 781.050 662.400 ;
        RECT 805.950 663.600 808.050 664.050 ;
        RECT 811.950 663.600 814.050 664.050 ;
        RECT 805.950 662.400 814.050 663.600 ;
        RECT 805.950 661.950 808.050 662.400 ;
        RECT 811.950 661.950 814.050 662.400 ;
        RECT 253.950 660.600 256.050 661.050 ;
        RECT 349.950 660.600 352.050 661.050 ;
        RECT 253.950 659.400 352.050 660.600 ;
        RECT 253.950 658.950 256.050 659.400 ;
        RECT 349.950 658.950 352.050 659.400 ;
        RECT 397.950 660.600 400.050 661.050 ;
        RECT 499.950 660.600 502.050 661.050 ;
        RECT 397.950 659.400 502.050 660.600 ;
        RECT 397.950 658.950 400.050 659.400 ;
        RECT 499.950 658.950 502.050 659.400 ;
        RECT 526.950 660.600 529.050 661.050 ;
        RECT 541.950 660.600 544.050 661.050 ;
        RECT 526.950 659.400 544.050 660.600 ;
        RECT 526.950 658.950 529.050 659.400 ;
        RECT 541.950 658.950 544.050 659.400 ;
        RECT 640.950 660.600 643.050 661.050 ;
        RECT 646.950 660.600 649.050 661.050 ;
        RECT 649.950 660.600 652.050 661.050 ;
        RECT 640.950 659.400 652.050 660.600 ;
        RECT 640.950 658.950 643.050 659.400 ;
        RECT 646.950 658.950 649.050 659.400 ;
        RECT 649.950 658.950 652.050 659.400 ;
        RECT 703.950 660.600 706.050 661.050 ;
        RECT 739.950 660.600 742.050 661.050 ;
        RECT 769.950 660.600 772.050 661.050 ;
        RECT 703.950 659.400 772.050 660.600 ;
        RECT 703.950 658.950 706.050 659.400 ;
        RECT 739.950 658.950 742.050 659.400 ;
        RECT 769.950 658.950 772.050 659.400 ;
        RECT 778.950 660.600 781.050 661.050 ;
        RECT 829.950 660.600 832.050 661.050 ;
        RECT 778.950 659.400 832.050 660.600 ;
        RECT 778.950 658.950 781.050 659.400 ;
        RECT 829.950 658.950 832.050 659.400 ;
        RECT 271.950 657.600 274.050 658.050 ;
        RECT 277.950 657.600 280.050 658.050 ;
        RECT 271.950 656.400 280.050 657.600 ;
        RECT 271.950 655.950 274.050 656.400 ;
        RECT 277.950 655.950 280.050 656.400 ;
        RECT 394.950 657.600 397.050 658.050 ;
        RECT 472.950 657.600 475.050 658.050 ;
        RECT 394.950 656.400 475.050 657.600 ;
        RECT 394.950 655.950 397.050 656.400 ;
        RECT 472.950 655.950 475.050 656.400 ;
        RECT 544.950 657.600 547.050 658.050 ;
        RECT 640.950 657.600 643.050 658.050 ;
        RECT 544.950 656.400 643.050 657.600 ;
        RECT 544.950 655.950 547.050 656.400 ;
        RECT 640.950 655.950 643.050 656.400 ;
        RECT 202.950 654.600 205.050 655.050 ;
        RECT 349.950 654.600 352.050 655.050 ;
        RECT 202.950 653.400 352.050 654.600 ;
        RECT 202.950 652.950 205.050 653.400 ;
        RECT 349.950 652.950 352.050 653.400 ;
        RECT 409.950 654.600 412.050 655.050 ;
        RECT 454.950 654.600 457.050 655.050 ;
        RECT 409.950 653.400 457.050 654.600 ;
        RECT 409.950 652.950 412.050 653.400 ;
        RECT 454.950 652.950 457.050 653.400 ;
        RECT 691.950 654.600 694.050 655.050 ;
        RECT 697.950 654.600 700.050 655.050 ;
        RECT 691.950 653.400 700.050 654.600 ;
        RECT 691.950 652.950 694.050 653.400 ;
        RECT 697.950 652.950 700.050 653.400 ;
        RECT 220.950 651.600 223.050 652.050 ;
        RECT 355.950 651.600 358.050 652.050 ;
        RECT 220.950 650.400 358.050 651.600 ;
        RECT 220.950 649.950 223.050 650.400 ;
        RECT 355.950 649.950 358.050 650.400 ;
        RECT 367.950 651.600 370.050 652.050 ;
        RECT 439.950 651.600 442.050 652.050 ;
        RECT 448.950 651.600 451.050 652.050 ;
        RECT 367.950 650.400 451.050 651.600 ;
        RECT 367.950 649.950 370.050 650.400 ;
        RECT 439.950 649.950 442.050 650.400 ;
        RECT 448.950 649.950 451.050 650.400 ;
        RECT 454.950 651.600 457.050 652.050 ;
        RECT 688.950 651.600 691.050 652.050 ;
        RECT 454.950 650.400 691.050 651.600 ;
        RECT 454.950 649.950 457.050 650.400 ;
        RECT 688.950 649.950 691.050 650.400 ;
        RECT 331.950 648.600 334.050 649.050 ;
        RECT 361.950 648.600 364.050 649.050 ;
        RECT 709.950 648.600 712.050 649.050 ;
        RECT 331.950 647.400 712.050 648.600 ;
        RECT 331.950 646.950 334.050 647.400 ;
        RECT 361.950 646.950 364.050 647.400 ;
        RECT 709.950 646.950 712.050 647.400 ;
        RECT 133.950 645.600 136.050 646.050 ;
        RECT 364.950 645.600 367.050 646.050 ;
        RECT 133.950 644.400 367.050 645.600 ;
        RECT 133.950 643.950 136.050 644.400 ;
        RECT 364.950 643.950 367.050 644.400 ;
        RECT 403.950 645.600 406.050 646.050 ;
        RECT 634.950 645.600 637.050 646.050 ;
        RECT 403.950 644.400 637.050 645.600 ;
        RECT 403.950 643.950 406.050 644.400 ;
        RECT 634.950 643.950 637.050 644.400 ;
        RECT 682.950 645.600 685.050 646.050 ;
        RECT 691.950 645.600 694.050 646.050 ;
        RECT 736.950 645.600 739.050 646.050 ;
        RECT 682.950 644.400 739.050 645.600 ;
        RECT 682.950 643.950 685.050 644.400 ;
        RECT 691.950 643.950 694.050 644.400 ;
        RECT 736.950 643.950 739.050 644.400 ;
        RECT 832.950 645.600 835.050 646.050 ;
        RECT 841.950 645.600 844.050 646.050 ;
        RECT 832.950 644.400 844.050 645.600 ;
        RECT 832.950 643.950 835.050 644.400 ;
        RECT 841.950 643.950 844.050 644.400 ;
        RECT 250.950 642.600 253.050 643.050 ;
        RECT 277.950 642.600 280.050 643.050 ;
        RECT 250.950 641.400 280.050 642.600 ;
        RECT 250.950 640.950 253.050 641.400 ;
        RECT 277.950 640.950 280.050 641.400 ;
        RECT 322.950 642.600 325.050 643.050 ;
        RECT 328.950 642.600 331.050 643.050 ;
        RECT 322.950 641.400 331.050 642.600 ;
        RECT 322.950 640.950 325.050 641.400 ;
        RECT 328.950 640.950 331.050 641.400 ;
        RECT 442.950 642.600 445.050 643.050 ;
        RECT 496.950 642.600 499.050 643.050 ;
        RECT 442.950 641.400 499.050 642.600 ;
        RECT 442.950 640.950 445.050 641.400 ;
        RECT 496.950 640.950 499.050 641.400 ;
        RECT 55.950 639.600 58.050 640.050 ;
        RECT 64.950 639.600 67.050 640.050 ;
        RECT 55.950 638.400 67.050 639.600 ;
        RECT 55.950 637.950 58.050 638.400 ;
        RECT 64.950 637.950 67.050 638.400 ;
        RECT 187.950 639.600 190.050 640.050 ;
        RECT 193.950 639.600 196.050 640.050 ;
        RECT 187.950 638.400 196.050 639.600 ;
        RECT 187.950 637.950 190.050 638.400 ;
        RECT 193.950 637.950 196.050 638.400 ;
        RECT 196.950 639.600 199.050 640.050 ;
        RECT 259.950 639.600 262.050 640.050 ;
        RECT 196.950 638.400 262.050 639.600 ;
        RECT 196.950 637.950 199.050 638.400 ;
        RECT 259.950 637.950 262.050 638.400 ;
        RECT 274.950 639.600 277.050 640.050 ;
        RECT 283.950 639.600 286.050 640.050 ;
        RECT 274.950 638.400 286.050 639.600 ;
        RECT 274.950 637.950 277.050 638.400 ;
        RECT 283.950 637.950 286.050 638.400 ;
        RECT 289.950 639.600 292.050 640.050 ;
        RECT 313.950 639.600 316.050 640.050 ;
        RECT 289.950 638.400 316.050 639.600 ;
        RECT 289.950 637.950 292.050 638.400 ;
        RECT 313.950 637.950 316.050 638.400 ;
        RECT 316.950 639.600 319.050 640.050 ;
        RECT 352.950 639.600 355.050 640.050 ;
        RECT 316.950 638.400 355.050 639.600 ;
        RECT 316.950 637.950 319.050 638.400 ;
        RECT 352.950 637.950 355.050 638.400 ;
        RECT 367.950 639.600 370.050 640.050 ;
        RECT 376.950 639.600 379.050 640.050 ;
        RECT 367.950 638.400 379.050 639.600 ;
        RECT 367.950 637.950 370.050 638.400 ;
        RECT 376.950 637.950 379.050 638.400 ;
        RECT 406.950 639.600 409.050 640.050 ;
        RECT 538.950 639.600 541.050 640.050 ;
        RECT 406.950 638.400 541.050 639.600 ;
        RECT 406.950 637.950 409.050 638.400 ;
        RECT 538.950 637.950 541.050 638.400 ;
        RECT 586.950 639.600 589.050 640.050 ;
        RECT 625.950 639.600 628.050 640.050 ;
        RECT 628.950 639.600 631.050 640.050 ;
        RECT 586.950 638.400 631.050 639.600 ;
        RECT 586.950 637.950 589.050 638.400 ;
        RECT 625.950 637.950 628.050 638.400 ;
        RECT 628.950 637.950 631.050 638.400 ;
        RECT 175.950 636.600 178.050 637.050 ;
        RECT 205.950 636.600 208.050 637.050 ;
        RECT 175.950 635.400 208.050 636.600 ;
        RECT 175.950 634.950 178.050 635.400 ;
        RECT 205.950 634.950 208.050 635.400 ;
        RECT 226.950 636.600 229.050 637.050 ;
        RECT 307.950 636.600 310.050 637.050 ;
        RECT 226.950 635.400 310.050 636.600 ;
        RECT 226.950 634.950 229.050 635.400 ;
        RECT 307.950 634.950 310.050 635.400 ;
        RECT 325.950 636.600 328.050 637.050 ;
        RECT 334.950 636.600 337.050 637.050 ;
        RECT 373.950 636.600 376.050 637.050 ;
        RECT 433.950 636.600 436.050 637.050 ;
        RECT 325.950 635.400 337.050 636.600 ;
        RECT 325.950 634.950 328.050 635.400 ;
        RECT 334.950 634.950 337.050 635.400 ;
        RECT 341.400 635.400 376.050 636.600 ;
        RECT 154.950 633.600 157.050 634.050 ;
        RECT 181.950 633.600 184.050 634.050 ;
        RECT 122.400 632.400 184.050 633.600 ;
        RECT 122.400 631.050 123.600 632.400 ;
        RECT 154.950 631.950 157.050 632.400 ;
        RECT 181.950 631.950 184.050 632.400 ;
        RECT 187.950 633.600 190.050 634.050 ;
        RECT 193.950 633.600 196.050 634.050 ;
        RECT 187.950 632.400 196.050 633.600 ;
        RECT 187.950 631.950 190.050 632.400 ;
        RECT 193.950 631.950 196.050 632.400 ;
        RECT 202.950 631.950 205.050 634.050 ;
        RECT 220.950 633.600 223.050 634.050 ;
        RECT 247.950 633.600 250.050 634.050 ;
        RECT 220.950 632.400 250.050 633.600 ;
        RECT 220.950 631.950 223.050 632.400 ;
        RECT 247.950 631.950 250.050 632.400 ;
        RECT 262.950 633.600 265.050 634.050 ;
        RECT 268.950 633.600 271.050 634.050 ;
        RECT 262.950 632.400 271.050 633.600 ;
        RECT 262.950 631.950 265.050 632.400 ;
        RECT 268.950 631.950 271.050 632.400 ;
        RECT 304.950 633.600 307.050 634.050 ;
        RECT 310.950 633.600 313.050 634.050 ;
        RECT 304.950 632.400 313.050 633.600 ;
        RECT 304.950 631.950 307.050 632.400 ;
        RECT 310.950 631.950 313.050 632.400 ;
        RECT 319.950 633.600 322.050 634.050 ;
        RECT 341.400 633.600 342.600 635.400 ;
        RECT 373.950 634.950 376.050 635.400 ;
        RECT 425.400 635.400 436.050 636.600 ;
        RECT 425.400 634.050 426.600 635.400 ;
        RECT 433.950 634.950 436.050 635.400 ;
        RECT 451.950 636.600 454.050 637.050 ;
        RECT 535.950 636.600 538.050 637.050 ;
        RECT 451.950 635.400 538.050 636.600 ;
        RECT 451.950 634.950 454.050 635.400 ;
        RECT 535.950 634.950 538.050 635.400 ;
        RECT 595.950 636.600 598.050 637.050 ;
        RECT 604.950 636.600 607.050 637.050 ;
        RECT 613.950 636.600 616.050 637.050 ;
        RECT 595.950 635.400 616.050 636.600 ;
        RECT 595.950 634.950 598.050 635.400 ;
        RECT 604.950 634.950 607.050 635.400 ;
        RECT 613.950 634.950 616.050 635.400 ;
        RECT 319.950 632.400 342.600 633.600 ;
        RECT 358.950 633.600 361.050 634.050 ;
        RECT 406.950 633.600 409.050 634.050 ;
        RECT 415.950 633.600 418.050 634.050 ;
        RECT 358.950 632.400 418.050 633.600 ;
        RECT 319.950 631.950 322.050 632.400 ;
        RECT 358.950 631.950 361.050 632.400 ;
        RECT 19.950 630.600 22.050 631.050 ;
        RECT 31.950 630.600 34.050 631.050 ;
        RECT 40.950 630.600 43.050 631.050 ;
        RECT 19.950 629.400 43.050 630.600 ;
        RECT 19.950 628.950 22.050 629.400 ;
        RECT 31.950 628.950 34.050 629.400 ;
        RECT 40.950 628.950 43.050 629.400 ;
        RECT 67.950 630.600 70.050 631.050 ;
        RECT 88.950 630.600 91.050 631.050 ;
        RECT 67.950 629.400 91.050 630.600 ;
        RECT 67.950 628.950 70.050 629.400 ;
        RECT 88.950 628.950 91.050 629.400 ;
        RECT 109.950 628.950 112.050 631.050 ;
        RECT 112.950 630.600 115.050 631.050 ;
        RECT 121.950 630.600 124.050 631.050 ;
        RECT 112.950 629.400 124.050 630.600 ;
        RECT 112.950 628.950 115.050 629.400 ;
        RECT 121.950 628.950 124.050 629.400 ;
        RECT 127.950 630.600 130.050 631.050 ;
        RECT 136.950 630.600 139.050 631.050 ;
        RECT 127.950 629.400 139.050 630.600 ;
        RECT 127.950 628.950 130.050 629.400 ;
        RECT 136.950 628.950 139.050 629.400 ;
        RECT 160.950 628.950 163.050 631.050 ;
        RECT 169.950 630.600 172.050 631.050 ;
        RECT 184.950 630.600 187.050 631.050 ;
        RECT 169.950 629.400 187.050 630.600 ;
        RECT 169.950 628.950 172.050 629.400 ;
        RECT 184.950 628.950 187.050 629.400 ;
        RECT 4.950 627.600 7.050 628.050 ;
        RECT 16.950 627.600 19.050 628.050 ;
        RECT 25.950 627.600 28.050 628.050 ;
        RECT 4.950 626.400 19.050 627.600 ;
        RECT 4.950 625.950 7.050 626.400 ;
        RECT 16.950 625.950 19.050 626.400 ;
        RECT 23.400 626.400 28.050 627.600 ;
        RECT 19.950 624.600 22.050 625.050 ;
        RECT 23.400 624.600 24.600 626.400 ;
        RECT 25.950 625.950 28.050 626.400 ;
        RECT 37.950 627.600 40.050 628.050 ;
        RECT 49.950 627.600 52.050 628.050 ;
        RECT 37.950 626.400 52.050 627.600 ;
        RECT 110.400 627.600 111.600 628.950 ;
        RECT 124.950 627.600 127.050 628.050 ;
        RECT 110.400 626.400 127.050 627.600 ;
        RECT 161.400 627.600 162.600 628.950 ;
        RECT 203.400 628.050 204.600 631.950 ;
        RECT 395.400 631.050 396.600 632.400 ;
        RECT 406.950 631.950 409.050 632.400 ;
        RECT 415.950 631.950 418.050 632.400 ;
        RECT 424.950 631.950 427.050 634.050 ;
        RECT 430.950 633.600 433.050 634.050 ;
        RECT 442.950 633.600 445.050 634.050 ;
        RECT 430.950 632.400 445.050 633.600 ;
        RECT 430.950 631.950 433.050 632.400 ;
        RECT 442.950 631.950 445.050 632.400 ;
        RECT 550.950 633.600 553.050 634.050 ;
        RECT 565.950 633.600 568.050 634.050 ;
        RECT 586.950 633.600 589.050 634.050 ;
        RECT 550.950 632.400 568.050 633.600 ;
        RECT 550.950 631.950 553.050 632.400 ;
        RECT 565.950 631.950 568.050 632.400 ;
        RECT 572.400 632.400 589.050 633.600 ;
        RECT 205.950 630.600 208.050 631.050 ;
        RECT 214.950 630.600 217.050 631.050 ;
        RECT 205.950 629.400 217.050 630.600 ;
        RECT 205.950 628.950 208.050 629.400 ;
        RECT 214.950 628.950 217.050 629.400 ;
        RECT 229.950 630.600 232.050 631.050 ;
        RECT 241.950 630.600 244.050 631.050 ;
        RECT 229.950 629.400 244.050 630.600 ;
        RECT 229.950 628.950 232.050 629.400 ;
        RECT 241.950 628.950 244.050 629.400 ;
        RECT 265.950 630.600 268.050 631.050 ;
        RECT 289.950 630.600 292.050 631.050 ;
        RECT 295.950 630.600 298.050 631.050 ;
        RECT 265.950 629.400 298.050 630.600 ;
        RECT 265.950 628.950 268.050 629.400 ;
        RECT 289.950 628.950 292.050 629.400 ;
        RECT 295.950 628.950 298.050 629.400 ;
        RECT 301.950 630.600 304.050 631.050 ;
        RECT 322.950 630.600 325.050 631.050 ;
        RECT 328.950 630.600 331.050 631.050 ;
        RECT 388.950 630.600 391.050 631.050 ;
        RECT 301.950 629.400 318.600 630.600 ;
        RECT 301.950 628.950 304.050 629.400 ;
        RECT 317.400 628.050 318.600 629.400 ;
        RECT 322.950 629.400 331.050 630.600 ;
        RECT 322.950 628.950 325.050 629.400 ;
        RECT 328.950 628.950 331.050 629.400 ;
        RECT 332.400 629.400 391.050 630.600 ;
        RECT 190.950 627.600 193.050 628.050 ;
        RECT 161.400 626.400 193.050 627.600 ;
        RECT 37.950 625.950 40.050 626.400 ;
        RECT 49.950 625.950 52.050 626.400 ;
        RECT 124.950 625.950 127.050 626.400 ;
        RECT 190.950 625.950 193.050 626.400 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 238.950 627.600 241.050 628.050 ;
        RECT 250.950 627.600 253.050 628.050 ;
        RECT 238.950 626.400 253.050 627.600 ;
        RECT 238.950 625.950 241.050 626.400 ;
        RECT 250.950 625.950 253.050 626.400 ;
        RECT 259.950 627.600 262.050 628.050 ;
        RECT 280.950 627.600 283.050 628.050 ;
        RECT 259.950 626.400 283.050 627.600 ;
        RECT 259.950 625.950 262.050 626.400 ;
        RECT 280.950 625.950 283.050 626.400 ;
        RECT 307.950 627.600 310.050 628.050 ;
        RECT 313.950 627.600 316.050 628.050 ;
        RECT 307.950 626.400 316.050 627.600 ;
        RECT 307.950 625.950 310.050 626.400 ;
        RECT 313.950 625.950 316.050 626.400 ;
        RECT 316.950 627.600 319.050 628.050 ;
        RECT 332.400 627.600 333.600 629.400 ;
        RECT 388.950 628.950 391.050 629.400 ;
        RECT 394.950 628.950 397.050 631.050 ;
        RECT 406.950 630.600 409.050 631.050 ;
        RECT 436.950 630.600 439.050 631.050 ;
        RECT 406.950 629.400 439.050 630.600 ;
        RECT 406.950 628.950 409.050 629.400 ;
        RECT 436.950 628.950 439.050 629.400 ;
        RECT 484.950 630.600 487.050 631.050 ;
        RECT 505.950 630.600 508.050 631.050 ;
        RECT 484.950 629.400 489.600 630.600 ;
        RECT 484.950 628.950 487.050 629.400 ;
        RECT 316.950 626.400 333.600 627.600 ;
        RECT 334.950 627.600 337.050 628.050 ;
        RECT 340.950 627.600 343.050 628.050 ;
        RECT 334.950 626.400 343.050 627.600 ;
        RECT 316.950 625.950 319.050 626.400 ;
        RECT 334.950 625.950 337.050 626.400 ;
        RECT 340.950 625.950 343.050 626.400 ;
        RECT 352.950 627.600 355.050 628.050 ;
        RECT 364.950 627.600 367.050 628.050 ;
        RECT 352.950 626.400 367.050 627.600 ;
        RECT 352.950 625.950 355.050 626.400 ;
        RECT 364.950 625.950 367.050 626.400 ;
        RECT 388.950 627.600 391.050 628.050 ;
        RECT 454.950 627.600 457.050 628.050 ;
        RECT 388.950 626.400 457.050 627.600 ;
        RECT 388.950 625.950 391.050 626.400 ;
        RECT 454.950 625.950 457.050 626.400 ;
        RECT 19.950 623.400 24.600 624.600 ;
        RECT 25.950 624.600 28.050 625.050 ;
        RECT 34.950 624.600 37.050 625.050 ;
        RECT 85.950 624.600 88.050 625.050 ;
        RECT 25.950 623.400 88.050 624.600 ;
        RECT 19.950 622.950 22.050 623.400 ;
        RECT 25.950 622.950 28.050 623.400 ;
        RECT 34.950 622.950 37.050 623.400 ;
        RECT 85.950 622.950 88.050 623.400 ;
        RECT 121.950 624.600 124.050 625.050 ;
        RECT 136.950 624.600 139.050 625.050 ;
        RECT 139.950 624.600 142.050 625.050 ;
        RECT 157.950 624.600 160.050 625.050 ;
        RECT 121.950 623.400 160.050 624.600 ;
        RECT 121.950 622.950 124.050 623.400 ;
        RECT 136.950 622.950 139.050 623.400 ;
        RECT 139.950 622.950 142.050 623.400 ;
        RECT 157.950 622.950 160.050 623.400 ;
        RECT 178.950 624.600 181.050 625.050 ;
        RECT 241.950 624.600 244.050 625.050 ;
        RECT 178.950 623.400 244.050 624.600 ;
        RECT 178.950 622.950 181.050 623.400 ;
        RECT 241.950 622.950 244.050 623.400 ;
        RECT 256.950 624.600 259.050 625.050 ;
        RECT 271.950 624.600 274.050 625.050 ;
        RECT 256.950 623.400 274.050 624.600 ;
        RECT 256.950 622.950 259.050 623.400 ;
        RECT 271.950 622.950 274.050 623.400 ;
        RECT 283.950 624.600 286.050 625.050 ;
        RECT 298.950 624.600 301.050 625.050 ;
        RECT 319.950 624.600 322.050 625.050 ;
        RECT 283.950 623.400 322.050 624.600 ;
        RECT 283.950 622.950 286.050 623.400 ;
        RECT 298.950 622.950 301.050 623.400 ;
        RECT 319.950 622.950 322.050 623.400 ;
        RECT 343.950 624.600 346.050 625.050 ;
        RECT 349.950 624.600 352.050 625.050 ;
        RECT 343.950 623.400 352.050 624.600 ;
        RECT 343.950 622.950 346.050 623.400 ;
        RECT 349.950 622.950 352.050 623.400 ;
        RECT 370.950 624.600 373.050 625.050 ;
        RECT 430.950 624.600 433.050 625.050 ;
        RECT 370.950 623.400 433.050 624.600 ;
        RECT 370.950 622.950 373.050 623.400 ;
        RECT 430.950 622.950 433.050 623.400 ;
        RECT 433.950 624.600 436.050 625.050 ;
        RECT 466.950 624.600 469.050 625.050 ;
        RECT 484.950 624.600 487.050 625.050 ;
        RECT 433.950 623.400 487.050 624.600 ;
        RECT 488.400 624.600 489.600 629.400 ;
        RECT 494.400 629.400 508.050 630.600 ;
        RECT 490.950 627.600 493.050 628.050 ;
        RECT 494.400 627.600 495.600 629.400 ;
        RECT 505.950 628.950 508.050 629.400 ;
        RECT 511.950 630.600 514.050 631.050 ;
        RECT 517.950 630.600 520.050 631.050 ;
        RECT 511.950 629.400 520.050 630.600 ;
        RECT 511.950 628.950 514.050 629.400 ;
        RECT 517.950 628.950 520.050 629.400 ;
        RECT 523.950 630.600 526.050 631.050 ;
        RECT 529.950 630.600 532.050 631.050 ;
        RECT 523.950 629.400 532.050 630.600 ;
        RECT 523.950 628.950 526.050 629.400 ;
        RECT 529.950 628.950 532.050 629.400 ;
        RECT 568.950 630.600 571.050 631.050 ;
        RECT 572.400 630.600 573.600 632.400 ;
        RECT 586.950 631.950 589.050 632.400 ;
        RECT 607.950 633.600 610.050 634.050 ;
        RECT 619.950 633.600 622.050 634.050 ;
        RECT 607.950 632.400 622.050 633.600 ;
        RECT 607.950 631.950 610.050 632.400 ;
        RECT 619.950 631.950 622.050 632.400 ;
        RECT 682.950 633.600 685.050 634.050 ;
        RECT 688.950 633.600 691.050 634.050 ;
        RECT 682.950 632.400 691.050 633.600 ;
        RECT 682.950 631.950 685.050 632.400 ;
        RECT 688.950 631.950 691.050 632.400 ;
        RECT 772.950 633.600 775.050 634.050 ;
        RECT 790.950 633.600 793.050 634.050 ;
        RECT 850.950 633.600 853.050 634.050 ;
        RECT 772.950 632.400 777.600 633.600 ;
        RECT 772.950 631.950 775.050 632.400 ;
        RECT 568.950 629.400 573.600 630.600 ;
        RECT 574.950 630.600 577.050 631.050 ;
        RECT 589.950 630.600 592.050 631.050 ;
        RECT 574.950 629.400 592.050 630.600 ;
        RECT 568.950 628.950 571.050 629.400 ;
        RECT 574.950 628.950 577.050 629.400 ;
        RECT 589.950 628.950 592.050 629.400 ;
        RECT 628.950 630.600 631.050 631.050 ;
        RECT 649.950 630.600 652.050 631.050 ;
        RECT 670.950 630.600 673.050 631.050 ;
        RECT 691.950 630.600 694.050 631.050 ;
        RECT 628.950 629.400 666.600 630.600 ;
        RECT 628.950 628.950 631.050 629.400 ;
        RECT 649.950 628.950 652.050 629.400 ;
        RECT 665.400 628.050 666.600 629.400 ;
        RECT 670.950 629.400 694.050 630.600 ;
        RECT 670.950 628.950 673.050 629.400 ;
        RECT 691.950 628.950 694.050 629.400 ;
        RECT 748.950 630.600 751.050 631.050 ;
        RECT 763.950 630.600 766.050 631.050 ;
        RECT 748.950 629.400 766.050 630.600 ;
        RECT 748.950 628.950 751.050 629.400 ;
        RECT 763.950 628.950 766.050 629.400 ;
        RECT 502.950 627.600 505.050 628.050 ;
        RECT 490.950 626.400 495.600 627.600 ;
        RECT 497.400 626.400 505.050 627.600 ;
        RECT 490.950 625.950 493.050 626.400 ;
        RECT 497.400 624.600 498.600 626.400 ;
        RECT 502.950 625.950 505.050 626.400 ;
        RECT 538.950 627.600 541.050 628.050 ;
        RECT 544.950 627.600 547.050 628.050 ;
        RECT 559.950 627.600 562.050 628.050 ;
        RECT 538.950 626.400 562.050 627.600 ;
        RECT 538.950 625.950 541.050 626.400 ;
        RECT 544.950 625.950 547.050 626.400 ;
        RECT 559.950 625.950 562.050 626.400 ;
        RECT 595.950 627.600 598.050 628.050 ;
        RECT 607.950 627.600 610.050 628.050 ;
        RECT 595.950 626.400 610.050 627.600 ;
        RECT 595.950 625.950 598.050 626.400 ;
        RECT 607.950 625.950 610.050 626.400 ;
        RECT 628.950 627.600 631.050 628.050 ;
        RECT 634.950 627.600 637.050 628.050 ;
        RECT 628.950 626.400 637.050 627.600 ;
        RECT 628.950 625.950 631.050 626.400 ;
        RECT 634.950 625.950 637.050 626.400 ;
        RECT 646.950 627.600 649.050 628.050 ;
        RECT 658.950 627.600 661.050 628.050 ;
        RECT 646.950 626.400 661.050 627.600 ;
        RECT 646.950 625.950 649.050 626.400 ;
        RECT 658.950 625.950 661.050 626.400 ;
        RECT 664.950 625.950 667.050 628.050 ;
        RECT 700.950 627.600 703.050 628.050 ;
        RECT 712.950 627.600 715.050 628.050 ;
        RECT 700.950 626.400 715.050 627.600 ;
        RECT 776.400 627.600 777.600 632.400 ;
        RECT 790.950 632.400 795.600 633.600 ;
        RECT 790.950 631.950 793.050 632.400 ;
        RECT 794.400 631.050 795.600 632.400 ;
        RECT 850.950 632.400 855.600 633.600 ;
        RECT 850.950 631.950 853.050 632.400 ;
        RECT 778.950 630.600 781.050 631.050 ;
        RECT 787.950 630.600 790.050 631.050 ;
        RECT 778.950 629.400 790.050 630.600 ;
        RECT 778.950 628.950 781.050 629.400 ;
        RECT 787.950 628.950 790.050 629.400 ;
        RECT 793.950 628.950 796.050 631.050 ;
        RECT 808.950 630.600 811.050 631.050 ;
        RECT 823.950 630.600 826.050 631.050 ;
        RECT 808.950 629.400 826.050 630.600 ;
        RECT 808.950 628.950 811.050 629.400 ;
        RECT 823.950 628.950 826.050 629.400 ;
        RECT 847.950 627.600 850.050 628.050 ;
        RECT 854.400 627.600 855.600 632.400 ;
        RECT 776.400 626.400 819.600 627.600 ;
        RECT 700.950 625.950 703.050 626.400 ;
        RECT 712.950 625.950 715.050 626.400 ;
        RECT 488.400 623.400 498.600 624.600 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 505.950 624.600 508.050 625.050 ;
        RECT 499.950 623.400 508.050 624.600 ;
        RECT 433.950 622.950 436.050 623.400 ;
        RECT 466.950 622.950 469.050 623.400 ;
        RECT 484.950 622.950 487.050 623.400 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 505.950 622.950 508.050 623.400 ;
        RECT 520.950 624.600 523.050 625.050 ;
        RECT 526.950 624.600 529.050 625.050 ;
        RECT 532.950 624.600 535.050 625.050 ;
        RECT 520.950 623.400 535.050 624.600 ;
        RECT 520.950 622.950 523.050 623.400 ;
        RECT 526.950 622.950 529.050 623.400 ;
        RECT 532.950 622.950 535.050 623.400 ;
        RECT 541.950 624.600 544.050 625.050 ;
        RECT 547.950 624.600 550.050 625.050 ;
        RECT 598.950 624.600 601.050 625.050 ;
        RECT 541.950 623.400 601.050 624.600 ;
        RECT 541.950 622.950 544.050 623.400 ;
        RECT 547.950 622.950 550.050 623.400 ;
        RECT 598.950 622.950 601.050 623.400 ;
        RECT 655.950 624.600 658.050 625.050 ;
        RECT 661.950 624.600 664.050 625.050 ;
        RECT 655.950 623.400 664.050 624.600 ;
        RECT 655.950 622.950 658.050 623.400 ;
        RECT 661.950 622.950 664.050 623.400 ;
        RECT 694.950 624.600 697.050 625.050 ;
        RECT 697.950 624.600 700.050 625.050 ;
        RECT 727.950 624.600 730.050 625.050 ;
        RECT 694.950 623.400 730.050 624.600 ;
        RECT 694.950 622.950 697.050 623.400 ;
        RECT 697.950 622.950 700.050 623.400 ;
        RECT 727.950 622.950 730.050 623.400 ;
        RECT 730.950 624.600 733.050 625.050 ;
        RECT 757.950 624.600 760.050 625.050 ;
        RECT 730.950 623.400 760.050 624.600 ;
        RECT 730.950 622.950 733.050 623.400 ;
        RECT 757.950 622.950 760.050 623.400 ;
        RECT 775.950 624.600 778.050 625.050 ;
        RECT 805.950 624.600 808.050 625.050 ;
        RECT 775.950 623.400 808.050 624.600 ;
        RECT 775.950 622.950 778.050 623.400 ;
        RECT 805.950 622.950 808.050 623.400 ;
        RECT 808.950 624.600 811.050 625.050 ;
        RECT 814.950 624.600 817.050 625.050 ;
        RECT 808.950 623.400 817.050 624.600 ;
        RECT 818.400 624.600 819.600 626.400 ;
        RECT 847.950 626.400 855.600 627.600 ;
        RECT 847.950 625.950 850.050 626.400 ;
        RECT 865.950 625.950 868.050 628.050 ;
        RECT 829.950 624.600 832.050 625.050 ;
        RECT 818.400 623.400 832.050 624.600 ;
        RECT 808.950 622.950 811.050 623.400 ;
        RECT 814.950 622.950 817.050 623.400 ;
        RECT 829.950 622.950 832.050 623.400 ;
        RECT 847.950 624.600 850.050 625.050 ;
        RECT 866.400 624.600 867.600 625.950 ;
        RECT 847.950 623.400 867.600 624.600 ;
        RECT 847.950 622.950 850.050 623.400 ;
        RECT 31.950 621.600 34.050 622.050 ;
        RECT 37.950 621.600 40.050 622.050 ;
        RECT 31.950 620.400 40.050 621.600 ;
        RECT 31.950 619.950 34.050 620.400 ;
        RECT 37.950 619.950 40.050 620.400 ;
        RECT 85.950 621.600 88.050 622.050 ;
        RECT 253.950 621.600 256.050 622.050 ;
        RECT 361.950 621.600 364.050 622.050 ;
        RECT 382.950 621.600 385.050 622.050 ;
        RECT 85.950 620.400 256.050 621.600 ;
        RECT 85.950 619.950 88.050 620.400 ;
        RECT 253.950 619.950 256.050 620.400 ;
        RECT 257.400 620.400 385.050 621.600 ;
        RECT 7.950 618.600 10.050 619.050 ;
        RECT 16.950 618.600 19.050 619.050 ;
        RECT 7.950 617.400 19.050 618.600 ;
        RECT 7.950 616.950 10.050 617.400 ;
        RECT 16.950 616.950 19.050 617.400 ;
        RECT 34.950 618.600 37.050 619.050 ;
        RECT 61.950 618.600 64.050 619.050 ;
        RECT 82.950 618.600 85.050 619.050 ;
        RECT 97.950 618.600 100.050 619.050 ;
        RECT 34.950 617.400 100.050 618.600 ;
        RECT 34.950 616.950 37.050 617.400 ;
        RECT 61.950 616.950 64.050 617.400 ;
        RECT 82.950 616.950 85.050 617.400 ;
        RECT 97.950 616.950 100.050 617.400 ;
        RECT 163.950 618.600 166.050 619.050 ;
        RECT 187.950 618.600 190.050 619.050 ;
        RECT 163.950 617.400 190.050 618.600 ;
        RECT 163.950 616.950 166.050 617.400 ;
        RECT 187.950 616.950 190.050 617.400 ;
        RECT 232.950 618.600 235.050 619.050 ;
        RECT 241.950 618.600 244.050 619.050 ;
        RECT 232.950 617.400 244.050 618.600 ;
        RECT 232.950 616.950 235.050 617.400 ;
        RECT 241.950 616.950 244.050 617.400 ;
        RECT 244.950 618.600 247.050 619.050 ;
        RECT 257.400 618.600 258.600 620.400 ;
        RECT 361.950 619.950 364.050 620.400 ;
        RECT 382.950 619.950 385.050 620.400 ;
        RECT 400.950 621.600 403.050 622.050 ;
        RECT 406.950 621.600 409.050 622.050 ;
        RECT 400.950 620.400 409.050 621.600 ;
        RECT 400.950 619.950 403.050 620.400 ;
        RECT 406.950 619.950 409.050 620.400 ;
        RECT 427.950 621.600 430.050 622.050 ;
        RECT 673.950 621.600 676.050 622.050 ;
        RECT 706.950 621.600 709.050 622.050 ;
        RECT 427.950 620.400 709.050 621.600 ;
        RECT 427.950 619.950 430.050 620.400 ;
        RECT 673.950 619.950 676.050 620.400 ;
        RECT 706.950 619.950 709.050 620.400 ;
        RECT 856.950 621.600 859.050 622.050 ;
        RECT 865.950 621.600 868.050 622.050 ;
        RECT 856.950 620.400 868.050 621.600 ;
        RECT 856.950 619.950 859.050 620.400 ;
        RECT 865.950 619.950 868.050 620.400 ;
        RECT 244.950 617.400 258.600 618.600 ;
        RECT 358.950 618.600 361.050 619.050 ;
        RECT 376.950 618.600 379.050 619.050 ;
        RECT 403.950 618.600 406.050 619.050 ;
        RECT 358.950 617.400 406.050 618.600 ;
        RECT 244.950 616.950 247.050 617.400 ;
        RECT 358.950 616.950 361.050 617.400 ;
        RECT 376.950 616.950 379.050 617.400 ;
        RECT 403.950 616.950 406.050 617.400 ;
        RECT 412.950 618.600 415.050 619.050 ;
        RECT 442.950 618.600 445.050 619.050 ;
        RECT 412.950 617.400 445.050 618.600 ;
        RECT 412.950 616.950 415.050 617.400 ;
        RECT 442.950 616.950 445.050 617.400 ;
        RECT 460.950 618.600 463.050 619.050 ;
        RECT 469.950 618.600 472.050 619.050 ;
        RECT 460.950 617.400 472.050 618.600 ;
        RECT 460.950 616.950 463.050 617.400 ;
        RECT 469.950 616.950 472.050 617.400 ;
        RECT 472.950 618.600 475.050 619.050 ;
        RECT 481.950 618.600 484.050 619.050 ;
        RECT 472.950 617.400 484.050 618.600 ;
        RECT 472.950 616.950 475.050 617.400 ;
        RECT 481.950 616.950 484.050 617.400 ;
        RECT 484.950 618.600 487.050 619.050 ;
        RECT 523.950 618.600 526.050 619.050 ;
        RECT 484.950 617.400 526.050 618.600 ;
        RECT 484.950 616.950 487.050 617.400 ;
        RECT 523.950 616.950 526.050 617.400 ;
        RECT 643.950 618.600 646.050 619.050 ;
        RECT 649.950 618.600 652.050 619.050 ;
        RECT 643.950 617.400 652.050 618.600 ;
        RECT 643.950 616.950 646.050 617.400 ;
        RECT 649.950 616.950 652.050 617.400 ;
        RECT 658.950 618.600 661.050 619.050 ;
        RECT 685.950 618.600 688.050 619.050 ;
        RECT 766.950 618.600 769.050 619.050 ;
        RECT 658.950 617.400 769.050 618.600 ;
        RECT 658.950 616.950 661.050 617.400 ;
        RECT 685.950 616.950 688.050 617.400 ;
        RECT 766.950 616.950 769.050 617.400 ;
        RECT 802.950 618.600 805.050 619.050 ;
        RECT 820.950 618.600 823.050 619.050 ;
        RECT 802.950 617.400 823.050 618.600 ;
        RECT 802.950 616.950 805.050 617.400 ;
        RECT 820.950 616.950 823.050 617.400 ;
        RECT 7.950 615.600 10.050 616.050 ;
        RECT 13.950 615.600 16.050 616.050 ;
        RECT 64.950 615.600 67.050 616.050 ;
        RECT 67.950 615.600 70.050 616.050 ;
        RECT 7.950 614.400 70.050 615.600 ;
        RECT 7.950 613.950 10.050 614.400 ;
        RECT 13.950 613.950 16.050 614.400 ;
        RECT 64.950 613.950 67.050 614.400 ;
        RECT 67.950 613.950 70.050 614.400 ;
        RECT 94.950 615.600 97.050 616.050 ;
        RECT 109.950 615.600 112.050 616.050 ;
        RECT 295.950 615.600 298.050 616.050 ;
        RECT 94.950 614.400 298.050 615.600 ;
        RECT 94.950 613.950 97.050 614.400 ;
        RECT 109.950 613.950 112.050 614.400 ;
        RECT 295.950 613.950 298.050 614.400 ;
        RECT 307.950 615.600 310.050 616.050 ;
        RECT 337.950 615.600 340.050 616.050 ;
        RECT 307.950 614.400 340.050 615.600 ;
        RECT 307.950 613.950 310.050 614.400 ;
        RECT 337.950 613.950 340.050 614.400 ;
        RECT 346.950 615.600 349.050 616.050 ;
        RECT 361.950 615.600 364.050 616.050 ;
        RECT 346.950 614.400 364.050 615.600 ;
        RECT 346.950 613.950 349.050 614.400 ;
        RECT 361.950 613.950 364.050 614.400 ;
        RECT 424.950 615.600 427.050 616.050 ;
        RECT 457.950 615.600 460.050 616.050 ;
        RECT 478.950 615.600 481.050 616.050 ;
        RECT 424.950 614.400 481.050 615.600 ;
        RECT 424.950 613.950 427.050 614.400 ;
        RECT 457.950 613.950 460.050 614.400 ;
        RECT 478.950 613.950 481.050 614.400 ;
        RECT 490.950 615.600 493.050 616.050 ;
        RECT 508.950 615.600 511.050 616.050 ;
        RECT 490.950 614.400 511.050 615.600 ;
        RECT 490.950 613.950 493.050 614.400 ;
        RECT 508.950 613.950 511.050 614.400 ;
        RECT 514.950 615.600 517.050 616.050 ;
        RECT 523.950 615.600 526.050 616.050 ;
        RECT 514.950 614.400 526.050 615.600 ;
        RECT 514.950 613.950 517.050 614.400 ;
        RECT 523.950 613.950 526.050 614.400 ;
        RECT 622.950 615.600 625.050 616.050 ;
        RECT 643.950 615.600 646.050 616.050 ;
        RECT 622.950 614.400 646.050 615.600 ;
        RECT 622.950 613.950 625.050 614.400 ;
        RECT 643.950 613.950 646.050 614.400 ;
        RECT 739.950 615.600 742.050 616.050 ;
        RECT 766.950 615.600 769.050 616.050 ;
        RECT 784.950 615.600 787.050 616.050 ;
        RECT 739.950 614.400 787.050 615.600 ;
        RECT 739.950 613.950 742.050 614.400 ;
        RECT 766.950 613.950 769.050 614.400 ;
        RECT 784.950 613.950 787.050 614.400 ;
        RECT 22.950 612.600 25.050 613.050 ;
        RECT 43.950 612.600 46.050 613.050 ;
        RECT 22.950 611.400 46.050 612.600 ;
        RECT 22.950 610.950 25.050 611.400 ;
        RECT 43.950 610.950 46.050 611.400 ;
        RECT 184.950 612.600 187.050 613.050 ;
        RECT 424.950 612.600 427.050 613.050 ;
        RECT 496.950 612.600 499.050 613.050 ;
        RECT 184.950 611.400 427.050 612.600 ;
        RECT 184.950 610.950 187.050 611.400 ;
        RECT 424.950 610.950 427.050 611.400 ;
        RECT 428.400 611.400 499.050 612.600 ;
        RECT 52.950 609.600 55.050 610.050 ;
        RECT 61.950 609.600 64.050 610.050 ;
        RECT 88.950 609.600 91.050 610.050 ;
        RECT 298.950 609.600 301.050 610.050 ;
        RECT 52.950 608.400 301.050 609.600 ;
        RECT 52.950 607.950 55.050 608.400 ;
        RECT 61.950 607.950 64.050 608.400 ;
        RECT 88.950 607.950 91.050 608.400 ;
        RECT 298.950 607.950 301.050 608.400 ;
        RECT 304.950 609.600 307.050 610.050 ;
        RECT 428.400 609.600 429.600 611.400 ;
        RECT 496.950 610.950 499.050 611.400 ;
        RECT 499.950 612.600 502.050 613.050 ;
        RECT 508.950 612.600 511.050 613.050 ;
        RECT 499.950 611.400 511.050 612.600 ;
        RECT 499.950 610.950 502.050 611.400 ;
        RECT 508.950 610.950 511.050 611.400 ;
        RECT 544.950 612.600 547.050 613.050 ;
        RECT 556.950 612.600 559.050 613.050 ;
        RECT 544.950 611.400 559.050 612.600 ;
        RECT 544.950 610.950 547.050 611.400 ;
        RECT 556.950 610.950 559.050 611.400 ;
        RECT 559.950 612.600 562.050 613.050 ;
        RECT 580.950 612.600 583.050 613.050 ;
        RECT 790.950 612.600 793.050 613.050 ;
        RECT 559.950 611.400 793.050 612.600 ;
        RECT 559.950 610.950 562.050 611.400 ;
        RECT 580.950 610.950 583.050 611.400 ;
        RECT 790.950 610.950 793.050 611.400 ;
        RECT 817.950 612.600 820.050 613.050 ;
        RECT 823.950 612.600 826.050 613.050 ;
        RECT 817.950 611.400 826.050 612.600 ;
        RECT 817.950 610.950 820.050 611.400 ;
        RECT 823.950 610.950 826.050 611.400 ;
        RECT 304.950 608.400 429.600 609.600 ;
        RECT 445.950 609.600 448.050 610.050 ;
        RECT 472.950 609.600 475.050 610.050 ;
        RECT 445.950 608.400 475.050 609.600 ;
        RECT 304.950 607.950 307.050 608.400 ;
        RECT 445.950 607.950 448.050 608.400 ;
        RECT 472.950 607.950 475.050 608.400 ;
        RECT 481.950 609.600 484.050 610.050 ;
        RECT 499.950 609.600 502.050 610.050 ;
        RECT 532.950 609.600 535.050 610.050 ;
        RECT 481.950 608.400 535.050 609.600 ;
        RECT 481.950 607.950 484.050 608.400 ;
        RECT 499.950 607.950 502.050 608.400 ;
        RECT 532.950 607.950 535.050 608.400 ;
        RECT 556.950 609.600 559.050 610.050 ;
        RECT 568.950 609.600 571.050 610.050 ;
        RECT 613.950 609.600 616.050 610.050 ;
        RECT 556.950 608.400 616.050 609.600 ;
        RECT 556.950 607.950 559.050 608.400 ;
        RECT 568.950 607.950 571.050 608.400 ;
        RECT 613.950 607.950 616.050 608.400 ;
        RECT 619.950 609.600 622.050 610.050 ;
        RECT 625.950 609.600 628.050 610.050 ;
        RECT 619.950 608.400 628.050 609.600 ;
        RECT 619.950 607.950 622.050 608.400 ;
        RECT 625.950 607.950 628.050 608.400 ;
        RECT 796.950 609.600 799.050 610.050 ;
        RECT 826.950 609.600 829.050 610.050 ;
        RECT 796.950 608.400 829.050 609.600 ;
        RECT 796.950 607.950 799.050 608.400 ;
        RECT 826.950 607.950 829.050 608.400 ;
        RECT 22.950 606.600 25.050 607.050 ;
        RECT 28.950 606.600 31.050 607.050 ;
        RECT 22.950 605.400 31.050 606.600 ;
        RECT 22.950 604.950 25.050 605.400 ;
        RECT 28.950 604.950 31.050 605.400 ;
        RECT 43.950 606.600 46.050 607.050 ;
        RECT 82.950 606.600 85.050 607.050 ;
        RECT 91.950 606.600 94.050 607.050 ;
        RECT 43.950 605.400 94.050 606.600 ;
        RECT 43.950 604.950 46.050 605.400 ;
        RECT 82.950 604.950 85.050 605.400 ;
        RECT 91.950 604.950 94.050 605.400 ;
        RECT 130.950 606.600 133.050 607.050 ;
        RECT 142.950 606.600 145.050 607.050 ;
        RECT 223.950 606.600 226.050 607.050 ;
        RECT 130.950 605.400 226.050 606.600 ;
        RECT 130.950 604.950 133.050 605.400 ;
        RECT 142.950 604.950 145.050 605.400 ;
        RECT 223.950 604.950 226.050 605.400 ;
        RECT 229.950 606.600 232.050 607.050 ;
        RECT 232.950 606.600 235.050 607.050 ;
        RECT 271.950 606.600 274.050 607.050 ;
        RECT 229.950 605.400 274.050 606.600 ;
        RECT 229.950 604.950 232.050 605.400 ;
        RECT 232.950 604.950 235.050 605.400 ;
        RECT 271.950 604.950 274.050 605.400 ;
        RECT 322.950 606.600 325.050 607.050 ;
        RECT 421.950 606.600 424.050 607.050 ;
        RECT 322.950 605.400 424.050 606.600 ;
        RECT 322.950 604.950 325.050 605.400 ;
        RECT 421.950 604.950 424.050 605.400 ;
        RECT 430.950 606.600 433.050 607.050 ;
        RECT 469.950 606.600 472.050 607.050 ;
        RECT 430.950 605.400 472.050 606.600 ;
        RECT 430.950 604.950 433.050 605.400 ;
        RECT 469.950 604.950 472.050 605.400 ;
        RECT 493.950 606.600 496.050 607.050 ;
        RECT 502.950 606.600 505.050 607.050 ;
        RECT 493.950 605.400 505.050 606.600 ;
        RECT 493.950 604.950 496.050 605.400 ;
        RECT 502.950 604.950 505.050 605.400 ;
        RECT 535.950 606.600 538.050 607.050 ;
        RECT 565.950 606.600 568.050 607.050 ;
        RECT 535.950 605.400 568.050 606.600 ;
        RECT 535.950 604.950 538.050 605.400 ;
        RECT 565.950 604.950 568.050 605.400 ;
        RECT 583.950 606.600 586.050 607.050 ;
        RECT 619.950 606.600 622.050 607.050 ;
        RECT 637.950 606.600 640.050 607.050 ;
        RECT 583.950 605.400 640.050 606.600 ;
        RECT 583.950 604.950 586.050 605.400 ;
        RECT 619.950 604.950 622.050 605.400 ;
        RECT 637.950 604.950 640.050 605.400 ;
        RECT 655.950 606.600 658.050 607.050 ;
        RECT 778.950 606.600 781.050 607.050 ;
        RECT 655.950 605.400 781.050 606.600 ;
        RECT 655.950 604.950 658.050 605.400 ;
        RECT 778.950 604.950 781.050 605.400 ;
        RECT 787.950 606.600 790.050 607.050 ;
        RECT 811.950 606.600 814.050 607.050 ;
        RECT 787.950 605.400 814.050 606.600 ;
        RECT 787.950 604.950 790.050 605.400 ;
        RECT 811.950 604.950 814.050 605.400 ;
        RECT 826.950 606.600 829.050 607.050 ;
        RECT 853.950 606.600 856.050 607.050 ;
        RECT 826.950 605.400 856.050 606.600 ;
        RECT 826.950 604.950 829.050 605.400 ;
        RECT 853.950 604.950 856.050 605.400 ;
        RECT 10.950 601.950 13.050 604.050 ;
        RECT 13.950 603.600 16.050 604.050 ;
        RECT 25.950 603.600 28.050 604.050 ;
        RECT 13.950 602.400 28.050 603.600 ;
        RECT 13.950 601.950 16.050 602.400 ;
        RECT 25.950 601.950 28.050 602.400 ;
        RECT 145.950 603.600 148.050 604.050 ;
        RECT 163.950 603.600 166.050 604.050 ;
        RECT 145.950 602.400 166.050 603.600 ;
        RECT 145.950 601.950 148.050 602.400 ;
        RECT 163.950 601.950 166.050 602.400 ;
        RECT 190.950 603.600 193.050 604.050 ;
        RECT 199.950 603.600 202.050 604.050 ;
        RECT 244.950 603.600 247.050 604.050 ;
        RECT 190.950 602.400 247.050 603.600 ;
        RECT 190.950 601.950 193.050 602.400 ;
        RECT 199.950 601.950 202.050 602.400 ;
        RECT 244.950 601.950 247.050 602.400 ;
        RECT 247.950 603.600 250.050 604.050 ;
        RECT 262.950 603.600 265.050 604.050 ;
        RECT 274.950 603.600 277.050 604.050 ;
        RECT 247.950 602.400 277.050 603.600 ;
        RECT 247.950 601.950 250.050 602.400 ;
        RECT 262.950 601.950 265.050 602.400 ;
        RECT 274.950 601.950 277.050 602.400 ;
        RECT 325.950 603.600 328.050 604.050 ;
        RECT 340.950 603.600 343.050 604.050 ;
        RECT 373.950 603.600 376.050 604.050 ;
        RECT 325.950 602.400 376.050 603.600 ;
        RECT 325.950 601.950 328.050 602.400 ;
        RECT 340.950 601.950 343.050 602.400 ;
        RECT 373.950 601.950 376.050 602.400 ;
        RECT 430.950 603.600 433.050 604.050 ;
        RECT 448.950 603.600 451.050 604.050 ;
        RECT 430.950 602.400 451.050 603.600 ;
        RECT 430.950 601.950 433.050 602.400 ;
        RECT 448.950 601.950 451.050 602.400 ;
        RECT 454.950 603.600 457.050 604.050 ;
        RECT 463.950 603.600 466.050 604.050 ;
        RECT 454.950 602.400 466.050 603.600 ;
        RECT 454.950 601.950 457.050 602.400 ;
        RECT 463.950 601.950 466.050 602.400 ;
        RECT 475.950 603.600 478.050 604.050 ;
        RECT 496.950 603.600 499.050 604.050 ;
        RECT 706.950 603.600 709.050 604.050 ;
        RECT 475.950 602.400 492.600 603.600 ;
        RECT 475.950 601.950 478.050 602.400 ;
        RECT 11.400 597.600 12.600 601.950 ;
        RECT 22.950 600.600 25.050 601.050 ;
        RECT 31.950 600.600 34.050 601.050 ;
        RECT 22.950 599.400 34.050 600.600 ;
        RECT 22.950 598.950 25.050 599.400 ;
        RECT 31.950 598.950 34.050 599.400 ;
        RECT 88.950 600.600 91.050 601.050 ;
        RECT 106.950 600.600 109.050 601.050 ;
        RECT 88.950 599.400 109.050 600.600 ;
        RECT 88.950 598.950 91.050 599.400 ;
        RECT 106.950 598.950 109.050 599.400 ;
        RECT 127.950 600.600 130.050 601.050 ;
        RECT 136.950 600.600 139.050 601.050 ;
        RECT 127.950 599.400 139.050 600.600 ;
        RECT 127.950 598.950 130.050 599.400 ;
        RECT 136.950 598.950 139.050 599.400 ;
        RECT 208.950 600.600 211.050 601.050 ;
        RECT 217.950 600.600 220.050 601.050 ;
        RECT 241.950 600.600 244.050 601.050 ;
        RECT 208.950 599.400 244.050 600.600 ;
        RECT 208.950 598.950 211.050 599.400 ;
        RECT 217.950 598.950 220.050 599.400 ;
        RECT 241.950 598.950 244.050 599.400 ;
        RECT 280.950 600.600 283.050 601.050 ;
        RECT 343.950 600.600 346.050 601.050 ;
        RECT 349.950 600.600 352.050 601.050 ;
        RECT 280.950 599.400 352.050 600.600 ;
        RECT 280.950 598.950 283.050 599.400 ;
        RECT 343.950 598.950 346.050 599.400 ;
        RECT 349.950 598.950 352.050 599.400 ;
        RECT 355.950 600.600 358.050 601.050 ;
        RECT 364.950 600.600 367.050 601.050 ;
        RECT 355.950 599.400 367.050 600.600 ;
        RECT 355.950 598.950 358.050 599.400 ;
        RECT 364.950 598.950 367.050 599.400 ;
        RECT 370.950 598.950 373.050 601.050 ;
        RECT 394.950 600.600 397.050 601.050 ;
        RECT 400.950 600.600 403.050 601.050 ;
        RECT 394.950 599.400 403.050 600.600 ;
        RECT 394.950 598.950 397.050 599.400 ;
        RECT 400.950 598.950 403.050 599.400 ;
        RECT 421.950 600.600 424.050 601.050 ;
        RECT 487.950 600.600 490.050 601.050 ;
        RECT 421.950 599.400 490.050 600.600 ;
        RECT 421.950 598.950 424.050 599.400 ;
        RECT 487.950 598.950 490.050 599.400 ;
        RECT 13.950 597.600 16.050 598.050 ;
        RECT 11.400 596.400 16.050 597.600 ;
        RECT 13.950 595.950 16.050 596.400 ;
        RECT 28.950 597.600 31.050 598.050 ;
        RECT 37.950 597.600 40.050 598.050 ;
        RECT 49.950 597.600 52.050 598.050 ;
        RECT 28.950 596.400 52.050 597.600 ;
        RECT 28.950 595.950 31.050 596.400 ;
        RECT 37.950 595.950 40.050 596.400 ;
        RECT 49.950 595.950 52.050 596.400 ;
        RECT 70.950 597.600 73.050 598.050 ;
        RECT 82.950 597.600 85.050 598.050 ;
        RECT 70.950 596.400 85.050 597.600 ;
        RECT 70.950 595.950 73.050 596.400 ;
        RECT 82.950 595.950 85.050 596.400 ;
        RECT 109.950 597.600 112.050 598.050 ;
        RECT 124.950 597.600 127.050 598.050 ;
        RECT 244.950 597.600 247.050 598.050 ;
        RECT 253.950 597.600 256.050 598.050 ;
        RECT 109.950 596.400 127.050 597.600 ;
        RECT 109.950 595.950 112.050 596.400 ;
        RECT 124.950 595.950 127.050 596.400 ;
        RECT 128.400 596.400 201.600 597.600 ;
        RECT 19.950 594.600 22.050 595.050 ;
        RECT 25.950 594.600 28.050 595.050 ;
        RECT 19.950 593.400 28.050 594.600 ;
        RECT 19.950 592.950 22.050 593.400 ;
        RECT 25.950 592.950 28.050 593.400 ;
        RECT 106.950 594.600 109.050 595.050 ;
        RECT 128.400 594.600 129.600 596.400 ;
        RECT 106.950 593.400 129.600 594.600 ;
        RECT 145.950 594.600 148.050 595.050 ;
        RECT 160.950 594.600 163.050 595.050 ;
        RECT 145.950 593.400 163.050 594.600 ;
        RECT 106.950 592.950 109.050 593.400 ;
        RECT 145.950 592.950 148.050 593.400 ;
        RECT 160.950 592.950 163.050 593.400 ;
        RECT 181.950 594.600 184.050 595.050 ;
        RECT 196.950 594.600 199.050 595.050 ;
        RECT 181.950 593.400 199.050 594.600 ;
        RECT 200.400 594.600 201.600 596.400 ;
        RECT 244.950 596.400 256.050 597.600 ;
        RECT 244.950 595.950 247.050 596.400 ;
        RECT 253.950 595.950 256.050 596.400 ;
        RECT 277.950 597.600 280.050 598.050 ;
        RECT 283.950 597.600 286.050 598.050 ;
        RECT 277.950 596.400 286.050 597.600 ;
        RECT 277.950 595.950 280.050 596.400 ;
        RECT 283.950 595.950 286.050 596.400 ;
        RECT 295.950 597.600 298.050 598.050 ;
        RECT 310.950 597.600 313.050 598.050 ;
        RECT 295.950 596.400 313.050 597.600 ;
        RECT 295.950 595.950 298.050 596.400 ;
        RECT 310.950 595.950 313.050 596.400 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 328.950 597.600 331.050 598.050 ;
        RECT 334.950 597.600 337.050 598.050 ;
        RECT 328.950 596.400 337.050 597.600 ;
        RECT 328.950 595.950 331.050 596.400 ;
        RECT 334.950 595.950 337.050 596.400 ;
        RECT 361.950 595.950 364.050 598.050 ;
        RECT 319.950 594.600 322.050 595.050 ;
        RECT 200.400 593.400 322.050 594.600 ;
        RECT 181.950 592.950 184.050 593.400 ;
        RECT 196.950 592.950 199.050 593.400 ;
        RECT 319.950 592.950 322.050 593.400 ;
        RECT 172.950 591.600 175.050 592.050 ;
        RECT 196.950 591.600 199.050 592.050 ;
        RECT 172.950 590.400 199.050 591.600 ;
        RECT 172.950 589.950 175.050 590.400 ;
        RECT 196.950 589.950 199.050 590.400 ;
        RECT 205.950 591.600 208.050 592.050 ;
        RECT 232.950 591.600 235.050 592.050 ;
        RECT 205.950 590.400 235.050 591.600 ;
        RECT 205.950 589.950 208.050 590.400 ;
        RECT 232.950 589.950 235.050 590.400 ;
        RECT 295.950 591.600 298.050 592.050 ;
        RECT 301.950 591.600 304.050 592.050 ;
        RECT 295.950 590.400 304.050 591.600 ;
        RECT 323.400 591.600 324.600 595.950 ;
        RECT 346.950 594.600 349.050 595.050 ;
        RECT 362.400 594.600 363.600 595.950 ;
        RECT 346.950 593.400 363.600 594.600 ;
        RECT 371.400 594.600 372.600 598.950 ;
        RECT 491.400 598.050 492.600 602.400 ;
        RECT 496.950 602.400 709.050 603.600 ;
        RECT 496.950 601.950 499.050 602.400 ;
        RECT 706.950 601.950 709.050 602.400 ;
        RECT 712.950 603.600 715.050 604.050 ;
        RECT 736.950 603.600 739.050 604.050 ;
        RECT 712.950 602.400 739.050 603.600 ;
        RECT 712.950 601.950 715.050 602.400 ;
        RECT 736.950 601.950 739.050 602.400 ;
        RECT 772.950 603.600 775.050 604.050 ;
        RECT 811.950 603.600 814.050 604.050 ;
        RECT 772.950 602.400 814.050 603.600 ;
        RECT 772.950 601.950 775.050 602.400 ;
        RECT 811.950 601.950 814.050 602.400 ;
        RECT 514.950 600.600 517.050 601.050 ;
        RECT 562.950 600.600 565.050 601.050 ;
        RECT 514.950 599.400 565.050 600.600 ;
        RECT 514.950 598.950 517.050 599.400 ;
        RECT 562.950 598.950 565.050 599.400 ;
        RECT 589.950 600.600 592.050 601.050 ;
        RECT 595.950 600.600 598.050 601.050 ;
        RECT 589.950 599.400 598.050 600.600 ;
        RECT 589.950 598.950 592.050 599.400 ;
        RECT 595.950 598.950 598.050 599.400 ;
        RECT 601.950 600.600 604.050 601.050 ;
        RECT 610.950 600.600 613.050 601.050 ;
        RECT 649.950 600.600 652.050 601.050 ;
        RECT 601.950 599.400 652.050 600.600 ;
        RECT 601.950 598.950 604.050 599.400 ;
        RECT 610.950 598.950 613.050 599.400 ;
        RECT 649.950 598.950 652.050 599.400 ;
        RECT 676.950 598.950 679.050 601.050 ;
        RECT 679.950 600.600 682.050 601.050 ;
        RECT 688.950 600.600 691.050 601.050 ;
        RECT 679.950 599.400 691.050 600.600 ;
        RECT 679.950 598.950 682.050 599.400 ;
        RECT 688.950 598.950 691.050 599.400 ;
        RECT 697.950 600.600 700.050 601.050 ;
        RECT 745.950 600.600 748.050 601.050 ;
        RECT 697.950 599.400 748.050 600.600 ;
        RECT 697.950 598.950 700.050 599.400 ;
        RECT 745.950 598.950 748.050 599.400 ;
        RECT 793.950 600.600 796.050 601.050 ;
        RECT 799.950 600.600 802.050 601.050 ;
        RECT 826.950 600.600 829.050 601.050 ;
        RECT 793.950 599.400 829.050 600.600 ;
        RECT 793.950 598.950 796.050 599.400 ;
        RECT 799.950 598.950 802.050 599.400 ;
        RECT 826.950 598.950 829.050 599.400 ;
        RECT 832.950 600.600 835.050 601.050 ;
        RECT 859.950 600.600 862.050 601.050 ;
        RECT 832.950 599.400 862.050 600.600 ;
        RECT 832.950 598.950 835.050 599.400 ;
        RECT 859.950 598.950 862.050 599.400 ;
        RECT 373.950 597.600 376.050 598.050 ;
        RECT 391.950 597.600 394.050 598.050 ;
        RECT 412.950 597.600 415.050 598.050 ;
        RECT 373.950 596.400 415.050 597.600 ;
        RECT 373.950 595.950 376.050 596.400 ;
        RECT 391.950 595.950 394.050 596.400 ;
        RECT 412.950 595.950 415.050 596.400 ;
        RECT 415.950 597.600 418.050 598.050 ;
        RECT 436.950 597.600 439.050 598.050 ;
        RECT 415.950 596.400 439.050 597.600 ;
        RECT 415.950 595.950 418.050 596.400 ;
        RECT 436.950 595.950 439.050 596.400 ;
        RECT 442.950 597.600 445.050 598.050 ;
        RECT 448.950 597.600 451.050 598.050 ;
        RECT 442.950 596.400 451.050 597.600 ;
        RECT 442.950 595.950 445.050 596.400 ;
        RECT 448.950 595.950 451.050 596.400 ;
        RECT 490.950 595.950 493.050 598.050 ;
        RECT 496.950 597.600 499.050 598.050 ;
        RECT 511.950 597.600 514.050 598.050 ;
        RECT 574.950 597.600 577.050 598.050 ;
        RECT 592.950 597.600 595.050 598.050 ;
        RECT 496.950 596.400 514.050 597.600 ;
        RECT 496.950 595.950 499.050 596.400 ;
        RECT 511.950 595.950 514.050 596.400 ;
        RECT 530.400 596.400 595.050 597.600 ;
        RECT 530.400 595.050 531.600 596.400 ;
        RECT 574.950 595.950 577.050 596.400 ;
        RECT 592.950 595.950 595.050 596.400 ;
        RECT 598.950 597.600 601.050 598.050 ;
        RECT 616.950 597.600 619.050 598.050 ;
        RECT 634.950 597.600 637.050 598.050 ;
        RECT 652.950 597.600 655.050 598.050 ;
        RECT 598.950 596.400 655.050 597.600 ;
        RECT 598.950 595.950 601.050 596.400 ;
        RECT 616.950 595.950 619.050 596.400 ;
        RECT 634.950 595.950 637.050 596.400 ;
        RECT 652.950 595.950 655.050 596.400 ;
        RECT 658.950 597.600 661.050 598.050 ;
        RECT 664.950 597.600 667.050 598.050 ;
        RECT 658.950 596.400 667.050 597.600 ;
        RECT 677.400 597.600 678.600 598.950 ;
        RECT 730.950 597.600 733.050 598.050 ;
        RECT 677.400 596.400 733.050 597.600 ;
        RECT 658.950 595.950 661.050 596.400 ;
        RECT 664.950 595.950 667.050 596.400 ;
        RECT 722.400 595.050 723.600 596.400 ;
        RECT 730.950 595.950 733.050 596.400 ;
        RECT 733.950 597.600 736.050 598.050 ;
        RECT 751.950 597.600 754.050 598.050 ;
        RECT 766.950 597.600 769.050 598.050 ;
        RECT 733.950 596.400 754.050 597.600 ;
        RECT 733.950 595.950 736.050 596.400 ;
        RECT 751.950 595.950 754.050 596.400 ;
        RECT 755.400 596.400 769.050 597.600 ;
        RECT 373.950 594.600 376.050 595.050 ;
        RECT 371.400 593.400 376.050 594.600 ;
        RECT 346.950 592.950 349.050 593.400 ;
        RECT 373.950 592.950 376.050 593.400 ;
        RECT 376.950 594.600 379.050 595.050 ;
        RECT 382.950 594.600 385.050 595.050 ;
        RECT 376.950 593.400 385.050 594.600 ;
        RECT 376.950 592.950 379.050 593.400 ;
        RECT 382.950 592.950 385.050 593.400 ;
        RECT 388.950 594.600 391.050 595.050 ;
        RECT 394.950 594.600 397.050 595.050 ;
        RECT 388.950 593.400 397.050 594.600 ;
        RECT 388.950 592.950 391.050 593.400 ;
        RECT 394.950 592.950 397.050 593.400 ;
        RECT 403.950 592.950 406.050 595.050 ;
        RECT 412.950 594.600 415.050 595.050 ;
        RECT 418.950 594.600 421.050 595.050 ;
        RECT 412.950 593.400 421.050 594.600 ;
        RECT 412.950 592.950 415.050 593.400 ;
        RECT 418.950 592.950 421.050 593.400 ;
        RECT 439.950 592.950 442.050 595.050 ;
        RECT 445.950 594.600 448.050 595.050 ;
        RECT 454.950 594.600 457.050 595.050 ;
        RECT 445.950 593.400 457.050 594.600 ;
        RECT 445.950 592.950 448.050 593.400 ;
        RECT 454.950 592.950 457.050 593.400 ;
        RECT 487.950 594.600 490.050 595.050 ;
        RECT 487.950 593.400 522.600 594.600 ;
        RECT 487.950 592.950 490.050 593.400 ;
        RECT 404.400 591.600 405.600 592.950 ;
        RECT 430.950 591.600 433.050 592.050 ;
        RECT 323.400 590.400 433.050 591.600 ;
        RECT 440.400 591.600 441.600 592.950 ;
        RECT 442.950 591.600 445.050 592.050 ;
        RECT 440.400 590.400 445.050 591.600 ;
        RECT 295.950 589.950 298.050 590.400 ;
        RECT 301.950 589.950 304.050 590.400 ;
        RECT 430.950 589.950 433.050 590.400 ;
        RECT 442.950 589.950 445.050 590.400 ;
        RECT 457.950 591.600 460.050 592.050 ;
        RECT 517.950 591.600 520.050 592.050 ;
        RECT 457.950 590.400 520.050 591.600 ;
        RECT 521.400 591.600 522.600 593.400 ;
        RECT 529.950 592.950 532.050 595.050 ;
        RECT 535.950 594.600 538.050 595.050 ;
        RECT 550.950 594.600 553.050 595.050 ;
        RECT 535.950 593.400 553.050 594.600 ;
        RECT 535.950 592.950 538.050 593.400 ;
        RECT 550.950 592.950 553.050 593.400 ;
        RECT 598.950 594.600 601.050 595.050 ;
        RECT 604.950 594.600 607.050 595.050 ;
        RECT 598.950 593.400 607.050 594.600 ;
        RECT 598.950 592.950 601.050 593.400 ;
        RECT 604.950 592.950 607.050 593.400 ;
        RECT 700.950 594.600 703.050 595.050 ;
        RECT 712.950 594.600 715.050 595.050 ;
        RECT 715.950 594.600 718.050 595.050 ;
        RECT 700.950 593.400 718.050 594.600 ;
        RECT 700.950 592.950 703.050 593.400 ;
        RECT 712.950 592.950 715.050 593.400 ;
        RECT 715.950 592.950 718.050 593.400 ;
        RECT 721.950 592.950 724.050 595.050 ;
        RECT 739.950 594.600 742.050 595.050 ;
        RECT 755.400 594.600 756.600 596.400 ;
        RECT 766.950 595.950 769.050 596.400 ;
        RECT 811.950 597.600 814.050 598.050 ;
        RECT 823.950 597.600 826.050 598.050 ;
        RECT 811.950 596.400 826.050 597.600 ;
        RECT 811.950 595.950 814.050 596.400 ;
        RECT 823.950 595.950 826.050 596.400 ;
        RECT 862.950 595.950 865.050 598.050 ;
        RECT 739.950 593.400 756.600 594.600 ;
        RECT 769.950 594.600 772.050 595.050 ;
        RECT 856.950 594.600 859.050 595.050 ;
        RECT 769.950 593.400 859.050 594.600 ;
        RECT 739.950 592.950 742.050 593.400 ;
        RECT 769.950 592.950 772.050 593.400 ;
        RECT 856.950 592.950 859.050 593.400 ;
        RECT 859.950 594.600 862.050 595.050 ;
        RECT 863.400 594.600 864.600 595.950 ;
        RECT 859.950 593.400 864.600 594.600 ;
        RECT 859.950 592.950 862.050 593.400 ;
        RECT 556.950 591.600 559.050 592.050 ;
        RECT 521.400 590.400 559.050 591.600 ;
        RECT 457.950 589.950 460.050 590.400 ;
        RECT 517.950 589.950 520.050 590.400 ;
        RECT 556.950 589.950 559.050 590.400 ;
        RECT 577.950 591.600 580.050 592.050 ;
        RECT 628.950 591.600 631.050 592.050 ;
        RECT 631.950 591.600 634.050 592.050 ;
        RECT 577.950 590.400 634.050 591.600 ;
        RECT 577.950 589.950 580.050 590.400 ;
        RECT 628.950 589.950 631.050 590.400 ;
        RECT 631.950 589.950 634.050 590.400 ;
        RECT 763.950 591.600 766.050 592.050 ;
        RECT 847.950 591.600 850.050 592.050 ;
        RECT 763.950 590.400 850.050 591.600 ;
        RECT 763.950 589.950 766.050 590.400 ;
        RECT 847.950 589.950 850.050 590.400 ;
        RECT 367.950 588.600 370.050 589.050 ;
        RECT 391.950 588.600 394.050 589.050 ;
        RECT 400.950 588.600 403.050 589.050 ;
        RECT 367.950 587.400 403.050 588.600 ;
        RECT 367.950 586.950 370.050 587.400 ;
        RECT 391.950 586.950 394.050 587.400 ;
        RECT 400.950 586.950 403.050 587.400 ;
        RECT 448.950 588.600 451.050 589.050 ;
        RECT 523.950 588.600 526.050 589.050 ;
        RECT 448.950 587.400 526.050 588.600 ;
        RECT 448.950 586.950 451.050 587.400 ;
        RECT 523.950 586.950 526.050 587.400 ;
        RECT 565.950 588.600 568.050 589.050 ;
        RECT 670.950 588.600 673.050 589.050 ;
        RECT 565.950 587.400 673.050 588.600 ;
        RECT 565.950 586.950 568.050 587.400 ;
        RECT 670.950 586.950 673.050 587.400 ;
        RECT 706.950 588.600 709.050 589.050 ;
        RECT 769.950 588.600 772.050 589.050 ;
        RECT 706.950 587.400 772.050 588.600 ;
        RECT 706.950 586.950 709.050 587.400 ;
        RECT 769.950 586.950 772.050 587.400 ;
        RECT 193.950 585.600 196.050 586.050 ;
        RECT 448.950 585.600 451.050 586.050 ;
        RECT 193.950 584.400 451.050 585.600 ;
        RECT 193.950 583.950 196.050 584.400 ;
        RECT 448.950 583.950 451.050 584.400 ;
        RECT 451.950 585.600 454.050 586.050 ;
        RECT 661.950 585.600 664.050 586.050 ;
        RECT 451.950 584.400 664.050 585.600 ;
        RECT 451.950 583.950 454.050 584.400 ;
        RECT 661.950 583.950 664.050 584.400 ;
        RECT 709.950 585.600 712.050 586.050 ;
        RECT 736.950 585.600 739.050 586.050 ;
        RECT 709.950 584.400 739.050 585.600 ;
        RECT 709.950 583.950 712.050 584.400 ;
        RECT 736.950 583.950 739.050 584.400 ;
        RECT 358.950 582.600 361.050 583.050 ;
        RECT 367.950 582.600 370.050 583.050 ;
        RECT 358.950 581.400 370.050 582.600 ;
        RECT 358.950 580.950 361.050 581.400 ;
        RECT 367.950 580.950 370.050 581.400 ;
        RECT 370.950 582.600 373.050 583.050 ;
        RECT 376.950 582.600 379.050 583.050 ;
        RECT 370.950 581.400 379.050 582.600 ;
        RECT 370.950 580.950 373.050 581.400 ;
        RECT 376.950 580.950 379.050 581.400 ;
        RECT 379.950 582.600 382.050 583.050 ;
        RECT 391.950 582.600 394.050 583.050 ;
        RECT 379.950 581.400 394.050 582.600 ;
        RECT 379.950 580.950 382.050 581.400 ;
        RECT 391.950 580.950 394.050 581.400 ;
        RECT 397.950 582.600 400.050 583.050 ;
        RECT 442.950 582.600 445.050 583.050 ;
        RECT 484.950 582.600 487.050 583.050 ;
        RECT 649.950 582.600 652.050 583.050 ;
        RECT 397.950 581.400 483.600 582.600 ;
        RECT 397.950 580.950 400.050 581.400 ;
        RECT 442.950 580.950 445.050 581.400 ;
        RECT 163.950 579.600 166.050 580.050 ;
        RECT 187.950 579.600 190.050 580.050 ;
        RECT 163.950 578.400 190.050 579.600 ;
        RECT 163.950 577.950 166.050 578.400 ;
        RECT 187.950 577.950 190.050 578.400 ;
        RECT 250.950 579.600 253.050 580.050 ;
        RECT 412.950 579.600 415.050 580.050 ;
        RECT 250.950 578.400 415.050 579.600 ;
        RECT 482.400 579.600 483.600 581.400 ;
        RECT 484.950 581.400 652.050 582.600 ;
        RECT 484.950 580.950 487.050 581.400 ;
        RECT 649.950 580.950 652.050 581.400 ;
        RECT 655.950 582.600 658.050 583.050 ;
        RECT 727.950 582.600 730.050 583.050 ;
        RECT 655.950 581.400 730.050 582.600 ;
        RECT 655.950 580.950 658.050 581.400 ;
        RECT 727.950 580.950 730.050 581.400 ;
        RECT 781.950 582.600 784.050 583.050 ;
        RECT 808.950 582.600 811.050 583.050 ;
        RECT 781.950 581.400 811.050 582.600 ;
        RECT 781.950 580.950 784.050 581.400 ;
        RECT 808.950 580.950 811.050 581.400 ;
        RECT 721.950 579.600 724.050 580.050 ;
        RECT 482.400 578.400 724.050 579.600 ;
        RECT 250.950 577.950 253.050 578.400 ;
        RECT 412.950 577.950 415.050 578.400 ;
        RECT 721.950 577.950 724.050 578.400 ;
        RECT 193.950 576.600 196.050 577.050 ;
        RECT 466.950 576.600 469.050 577.050 ;
        RECT 193.950 575.400 469.050 576.600 ;
        RECT 193.950 574.950 196.050 575.400 ;
        RECT 466.950 574.950 469.050 575.400 ;
        RECT 469.950 576.600 472.050 577.050 ;
        RECT 484.950 576.600 487.050 577.050 ;
        RECT 469.950 575.400 487.050 576.600 ;
        RECT 469.950 574.950 472.050 575.400 ;
        RECT 484.950 574.950 487.050 575.400 ;
        RECT 487.950 576.600 490.050 577.050 ;
        RECT 505.950 576.600 508.050 577.050 ;
        RECT 487.950 575.400 508.050 576.600 ;
        RECT 487.950 574.950 490.050 575.400 ;
        RECT 505.950 574.950 508.050 575.400 ;
        RECT 571.950 576.600 574.050 577.050 ;
        RECT 637.950 576.600 640.050 577.050 ;
        RECT 679.950 576.600 682.050 577.050 ;
        RECT 571.950 575.400 682.050 576.600 ;
        RECT 571.950 574.950 574.050 575.400 ;
        RECT 637.950 574.950 640.050 575.400 ;
        RECT 679.950 574.950 682.050 575.400 ;
        RECT 160.950 573.600 163.050 574.050 ;
        RECT 175.950 573.600 178.050 574.050 ;
        RECT 160.950 572.400 178.050 573.600 ;
        RECT 160.950 571.950 163.050 572.400 ;
        RECT 175.950 571.950 178.050 572.400 ;
        RECT 355.950 573.600 358.050 574.050 ;
        RECT 409.950 573.600 412.050 574.050 ;
        RECT 355.950 572.400 412.050 573.600 ;
        RECT 355.950 571.950 358.050 572.400 ;
        RECT 409.950 571.950 412.050 572.400 ;
        RECT 493.950 573.600 496.050 574.050 ;
        RECT 499.950 573.600 502.050 574.050 ;
        RECT 493.950 572.400 502.050 573.600 ;
        RECT 493.950 571.950 496.050 572.400 ;
        RECT 499.950 571.950 502.050 572.400 ;
        RECT 526.950 573.600 529.050 574.050 ;
        RECT 583.950 573.600 586.050 574.050 ;
        RECT 526.950 572.400 586.050 573.600 ;
        RECT 526.950 571.950 529.050 572.400 ;
        RECT 583.950 571.950 586.050 572.400 ;
        RECT 703.950 573.600 706.050 574.050 ;
        RECT 727.950 573.600 730.050 574.050 ;
        RECT 703.950 572.400 730.050 573.600 ;
        RECT 703.950 571.950 706.050 572.400 ;
        RECT 727.950 571.950 730.050 572.400 ;
        RECT 814.950 573.600 817.050 574.050 ;
        RECT 871.950 573.600 874.050 574.050 ;
        RECT 814.950 572.400 874.050 573.600 ;
        RECT 814.950 571.950 817.050 572.400 ;
        RECT 871.950 571.950 874.050 572.400 ;
        RECT 154.950 570.600 157.050 571.050 ;
        RECT 181.950 570.600 184.050 571.050 ;
        RECT 154.950 569.400 184.050 570.600 ;
        RECT 154.950 568.950 157.050 569.400 ;
        RECT 181.950 568.950 184.050 569.400 ;
        RECT 307.950 570.600 310.050 571.050 ;
        RECT 310.950 570.600 313.050 571.050 ;
        RECT 358.950 570.600 361.050 571.050 ;
        RECT 307.950 569.400 361.050 570.600 ;
        RECT 307.950 568.950 310.050 569.400 ;
        RECT 310.950 568.950 313.050 569.400 ;
        RECT 358.950 568.950 361.050 569.400 ;
        RECT 370.950 570.600 373.050 571.050 ;
        RECT 397.950 570.600 400.050 571.050 ;
        RECT 370.950 569.400 400.050 570.600 ;
        RECT 370.950 568.950 373.050 569.400 ;
        RECT 397.950 568.950 400.050 569.400 ;
        RECT 421.950 570.600 424.050 571.050 ;
        RECT 442.950 570.600 445.050 571.050 ;
        RECT 421.950 569.400 445.050 570.600 ;
        RECT 421.950 568.950 424.050 569.400 ;
        RECT 442.950 568.950 445.050 569.400 ;
        RECT 466.950 570.600 469.050 571.050 ;
        RECT 502.950 570.600 505.050 571.050 ;
        RECT 466.950 569.400 505.050 570.600 ;
        RECT 466.950 568.950 469.050 569.400 ;
        RECT 502.950 568.950 505.050 569.400 ;
        RECT 544.950 570.600 547.050 571.050 ;
        RECT 688.950 570.600 691.050 571.050 ;
        RECT 544.950 569.400 691.050 570.600 ;
        RECT 544.950 568.950 547.050 569.400 ;
        RECT 688.950 568.950 691.050 569.400 ;
        RECT 700.950 570.600 703.050 571.050 ;
        RECT 769.950 570.600 772.050 571.050 ;
        RECT 787.950 570.600 790.050 571.050 ;
        RECT 700.950 569.400 790.050 570.600 ;
        RECT 700.950 568.950 703.050 569.400 ;
        RECT 769.950 568.950 772.050 569.400 ;
        RECT 787.950 568.950 790.050 569.400 ;
        RECT 7.950 567.600 10.050 568.050 ;
        RECT 16.950 567.600 19.050 568.050 ;
        RECT 7.950 566.400 19.050 567.600 ;
        RECT 7.950 565.950 10.050 566.400 ;
        RECT 16.950 565.950 19.050 566.400 ;
        RECT 403.950 567.600 406.050 568.050 ;
        RECT 586.950 567.600 589.050 568.050 ;
        RECT 712.950 567.600 715.050 568.050 ;
        RECT 403.950 566.400 715.050 567.600 ;
        RECT 403.950 565.950 406.050 566.400 ;
        RECT 586.950 565.950 589.050 566.400 ;
        RECT 712.950 565.950 715.050 566.400 ;
        RECT 841.950 567.600 844.050 568.050 ;
        RECT 853.950 567.600 856.050 568.050 ;
        RECT 841.950 566.400 856.050 567.600 ;
        RECT 841.950 565.950 844.050 566.400 ;
        RECT 853.950 565.950 856.050 566.400 ;
        RECT 16.950 564.600 19.050 565.050 ;
        RECT 142.950 564.600 145.050 565.050 ;
        RECT 151.950 564.600 154.050 565.050 ;
        RECT 16.950 563.400 36.600 564.600 ;
        RECT 16.950 562.950 19.050 563.400 ;
        RECT 35.400 562.050 36.600 563.400 ;
        RECT 142.950 563.400 154.050 564.600 ;
        RECT 142.950 562.950 145.050 563.400 ;
        RECT 151.950 562.950 154.050 563.400 ;
        RECT 166.950 564.600 169.050 565.050 ;
        RECT 175.950 564.600 178.050 565.050 ;
        RECT 199.950 564.600 202.050 565.050 ;
        RECT 166.950 563.400 178.050 564.600 ;
        RECT 166.950 562.950 169.050 563.400 ;
        RECT 175.950 562.950 178.050 563.400 ;
        RECT 188.400 563.400 202.050 564.600 ;
        RECT 188.400 562.050 189.600 563.400 ;
        RECT 199.950 562.950 202.050 563.400 ;
        RECT 208.950 564.600 211.050 565.050 ;
        RECT 229.950 564.600 232.050 565.050 ;
        RECT 208.950 563.400 232.050 564.600 ;
        RECT 208.950 562.950 211.050 563.400 ;
        RECT 229.950 562.950 232.050 563.400 ;
        RECT 271.950 564.600 274.050 565.050 ;
        RECT 280.950 564.600 283.050 565.050 ;
        RECT 271.950 563.400 283.050 564.600 ;
        RECT 271.950 562.950 274.050 563.400 ;
        RECT 280.950 562.950 283.050 563.400 ;
        RECT 283.950 564.600 286.050 565.050 ;
        RECT 298.950 564.600 301.050 565.050 ;
        RECT 319.950 564.600 322.050 565.050 ;
        RECT 283.950 563.400 322.050 564.600 ;
        RECT 283.950 562.950 286.050 563.400 ;
        RECT 298.950 562.950 301.050 563.400 ;
        RECT 319.950 562.950 322.050 563.400 ;
        RECT 349.950 564.600 352.050 565.050 ;
        RECT 385.950 564.600 388.050 565.050 ;
        RECT 349.950 563.400 388.050 564.600 ;
        RECT 349.950 562.950 352.050 563.400 ;
        RECT 385.950 562.950 388.050 563.400 ;
        RECT 424.950 564.600 427.050 565.050 ;
        RECT 493.950 564.600 496.050 565.050 ;
        RECT 424.950 563.400 496.050 564.600 ;
        RECT 424.950 562.950 427.050 563.400 ;
        RECT 493.950 562.950 496.050 563.400 ;
        RECT 505.950 564.600 508.050 565.050 ;
        RECT 532.950 564.600 535.050 565.050 ;
        RECT 505.950 563.400 535.050 564.600 ;
        RECT 505.950 562.950 508.050 563.400 ;
        RECT 532.950 562.950 535.050 563.400 ;
        RECT 574.950 564.600 577.050 565.050 ;
        RECT 673.950 564.600 676.050 565.050 ;
        RECT 574.950 563.400 676.050 564.600 ;
        RECT 574.950 562.950 577.050 563.400 ;
        RECT 673.950 562.950 676.050 563.400 ;
        RECT 859.950 564.600 862.050 565.050 ;
        RECT 859.950 563.400 867.600 564.600 ;
        RECT 859.950 562.950 862.050 563.400 ;
        RECT 10.950 561.600 13.050 562.050 ;
        RECT 28.950 561.600 31.050 562.050 ;
        RECT 34.950 561.600 37.050 562.050 ;
        RECT 46.950 561.600 49.050 562.050 ;
        RECT 10.950 560.400 27.600 561.600 ;
        RECT 10.950 559.950 13.050 560.400 ;
        RECT 26.400 558.600 27.600 560.400 ;
        RECT 28.950 560.400 33.600 561.600 ;
        RECT 28.950 559.950 31.050 560.400 ;
        RECT 32.400 558.600 33.600 560.400 ;
        RECT 34.950 560.400 49.050 561.600 ;
        RECT 34.950 559.950 37.050 560.400 ;
        RECT 46.950 559.950 49.050 560.400 ;
        RECT 97.950 561.600 100.050 562.050 ;
        RECT 109.950 561.600 112.050 562.050 ;
        RECT 148.950 561.600 151.050 562.050 ;
        RECT 97.950 560.400 151.050 561.600 ;
        RECT 97.950 559.950 100.050 560.400 ;
        RECT 109.950 559.950 112.050 560.400 ;
        RECT 148.950 559.950 151.050 560.400 ;
        RECT 166.950 559.950 169.050 562.050 ;
        RECT 172.950 561.600 175.050 562.050 ;
        RECT 178.950 561.600 181.050 562.050 ;
        RECT 172.950 560.400 181.050 561.600 ;
        RECT 172.950 559.950 175.050 560.400 ;
        RECT 178.950 559.950 181.050 560.400 ;
        RECT 187.950 559.950 190.050 562.050 ;
        RECT 199.950 561.600 202.050 562.050 ;
        RECT 214.950 561.600 217.050 562.050 ;
        RECT 199.950 560.400 217.050 561.600 ;
        RECT 199.950 559.950 202.050 560.400 ;
        RECT 214.950 559.950 217.050 560.400 ;
        RECT 226.950 559.950 229.050 562.050 ;
        RECT 250.950 561.600 253.050 562.050 ;
        RECT 280.950 561.600 283.050 562.050 ;
        RECT 304.950 561.600 307.050 562.050 ;
        RECT 250.950 560.400 307.050 561.600 ;
        RECT 250.950 559.950 253.050 560.400 ;
        RECT 280.950 559.950 283.050 560.400 ;
        RECT 304.950 559.950 307.050 560.400 ;
        RECT 307.950 561.600 310.050 562.050 ;
        RECT 325.950 561.600 328.050 562.050 ;
        RECT 307.950 560.400 328.050 561.600 ;
        RECT 307.950 559.950 310.050 560.400 ;
        RECT 325.950 559.950 328.050 560.400 ;
        RECT 346.950 561.600 349.050 562.050 ;
        RECT 403.950 561.600 406.050 562.050 ;
        RECT 346.950 560.400 363.600 561.600 ;
        RECT 346.950 559.950 349.050 560.400 ;
        RECT 43.950 558.600 46.050 559.050 ;
        RECT 26.400 557.400 30.600 558.600 ;
        RECT 32.400 557.400 46.050 558.600 ;
        RECT 10.950 555.600 13.050 556.050 ;
        RECT 19.950 555.600 22.050 556.050 ;
        RECT 10.950 554.400 22.050 555.600 ;
        RECT 29.400 555.600 30.600 557.400 ;
        RECT 43.950 556.950 46.050 557.400 ;
        RECT 61.950 558.600 64.050 559.050 ;
        RECT 73.950 558.600 76.050 559.050 ;
        RECT 61.950 557.400 76.050 558.600 ;
        RECT 61.950 556.950 64.050 557.400 ;
        RECT 73.950 556.950 76.050 557.400 ;
        RECT 88.950 558.600 91.050 559.050 ;
        RECT 121.950 558.600 124.050 559.050 ;
        RECT 88.950 557.400 124.050 558.600 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 121.950 556.950 124.050 557.400 ;
        RECT 127.950 558.600 130.050 559.050 ;
        RECT 167.400 558.600 168.600 559.950 ;
        RECT 184.950 558.600 187.050 559.050 ;
        RECT 127.950 557.400 138.600 558.600 ;
        RECT 167.400 557.400 187.050 558.600 ;
        RECT 127.950 556.950 130.050 557.400 ;
        RECT 31.950 555.600 34.050 556.050 ;
        RECT 29.400 554.400 34.050 555.600 ;
        RECT 10.950 553.950 13.050 554.400 ;
        RECT 19.950 553.950 22.050 554.400 ;
        RECT 31.950 553.950 34.050 554.400 ;
        RECT 37.950 555.600 40.050 556.050 ;
        RECT 49.950 555.600 52.050 556.050 ;
        RECT 37.950 554.400 52.050 555.600 ;
        RECT 37.950 553.950 40.050 554.400 ;
        RECT 49.950 553.950 52.050 554.400 ;
        RECT 64.950 555.600 67.050 556.050 ;
        RECT 67.950 555.600 70.050 556.050 ;
        RECT 79.950 555.600 82.050 556.050 ;
        RECT 64.950 554.400 82.050 555.600 ;
        RECT 64.950 553.950 67.050 554.400 ;
        RECT 67.950 553.950 70.050 554.400 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 82.950 555.600 85.050 556.050 ;
        RECT 106.950 555.600 109.050 556.050 ;
        RECT 82.950 554.400 109.050 555.600 ;
        RECT 82.950 553.950 85.050 554.400 ;
        RECT 106.950 553.950 109.050 554.400 ;
        RECT 109.950 555.600 112.050 556.050 ;
        RECT 122.400 555.600 123.600 556.950 ;
        RECT 109.950 554.400 123.600 555.600 ;
        RECT 124.950 555.600 127.050 556.050 ;
        RECT 133.950 555.600 136.050 556.050 ;
        RECT 124.950 554.400 136.050 555.600 ;
        RECT 137.400 555.600 138.600 557.400 ;
        RECT 184.950 556.950 187.050 557.400 ;
        RECT 205.950 556.950 208.050 559.050 ;
        RECT 208.950 556.950 211.050 559.050 ;
        RECT 211.950 558.600 214.050 559.050 ;
        RECT 217.950 558.600 220.050 559.050 ;
        RECT 223.950 558.600 226.050 559.050 ;
        RECT 211.950 557.400 226.050 558.600 ;
        RECT 211.950 556.950 214.050 557.400 ;
        RECT 217.950 556.950 220.050 557.400 ;
        RECT 223.950 556.950 226.050 557.400 ;
        RECT 151.950 555.600 154.050 556.050 ;
        RECT 137.400 554.400 154.050 555.600 ;
        RECT 109.950 553.950 112.050 554.400 ;
        RECT 124.950 553.950 127.050 554.400 ;
        RECT 133.950 553.950 136.050 554.400 ;
        RECT 151.950 553.950 154.050 554.400 ;
        RECT 169.950 555.600 172.050 556.050 ;
        RECT 206.400 555.600 207.600 556.950 ;
        RECT 169.950 554.400 207.600 555.600 ;
        RECT 209.400 555.600 210.600 556.950 ;
        RECT 227.400 556.050 228.600 559.950 ;
        RECT 362.400 559.050 363.600 560.400 ;
        RECT 386.400 560.400 406.050 561.600 ;
        RECT 235.950 558.600 238.050 559.050 ;
        RECT 259.950 558.600 262.050 559.050 ;
        RECT 235.950 557.400 262.050 558.600 ;
        RECT 235.950 556.950 238.050 557.400 ;
        RECT 259.950 556.950 262.050 557.400 ;
        RECT 283.950 558.600 286.050 559.050 ;
        RECT 298.950 558.600 301.050 559.050 ;
        RECT 283.950 557.400 301.050 558.600 ;
        RECT 283.950 556.950 286.050 557.400 ;
        RECT 298.950 556.950 301.050 557.400 ;
        RECT 313.950 558.600 316.050 559.050 ;
        RECT 340.950 558.600 343.050 559.050 ;
        RECT 313.950 557.400 343.050 558.600 ;
        RECT 313.950 556.950 316.050 557.400 ;
        RECT 340.950 556.950 343.050 557.400 ;
        RECT 361.950 556.950 364.050 559.050 ;
        RECT 367.950 558.600 370.050 559.050 ;
        RECT 382.950 558.600 385.050 559.050 ;
        RECT 367.950 557.400 385.050 558.600 ;
        RECT 367.950 556.950 370.050 557.400 ;
        RECT 382.950 556.950 385.050 557.400 ;
        RECT 214.950 555.600 217.050 556.050 ;
        RECT 209.400 554.400 217.050 555.600 ;
        RECT 169.950 553.950 172.050 554.400 ;
        RECT 214.950 553.950 217.050 554.400 ;
        RECT 226.950 553.950 229.050 556.050 ;
        RECT 232.950 555.600 235.050 556.050 ;
        RECT 262.950 555.600 265.050 556.050 ;
        RECT 232.950 554.400 265.050 555.600 ;
        RECT 232.950 553.950 235.050 554.400 ;
        RECT 262.950 553.950 265.050 554.400 ;
        RECT 292.950 555.600 295.050 556.050 ;
        RECT 313.950 555.600 316.050 556.050 ;
        RECT 292.950 554.400 316.050 555.600 ;
        RECT 292.950 553.950 295.050 554.400 ;
        RECT 313.950 553.950 316.050 554.400 ;
        RECT 316.950 555.600 319.050 556.050 ;
        RECT 343.950 555.600 346.050 556.050 ;
        RECT 316.950 554.400 346.050 555.600 ;
        RECT 316.950 553.950 319.050 554.400 ;
        RECT 343.950 553.950 346.050 554.400 ;
        RECT 370.950 555.600 373.050 556.050 ;
        RECT 386.400 555.600 387.600 560.400 ;
        RECT 403.950 559.950 406.050 560.400 ;
        RECT 418.950 561.600 421.050 562.050 ;
        RECT 454.950 561.600 457.050 562.050 ;
        RECT 418.950 560.400 457.050 561.600 ;
        RECT 418.950 559.950 421.050 560.400 ;
        RECT 454.950 559.950 457.050 560.400 ;
        RECT 460.950 559.950 463.050 562.050 ;
        RECT 484.950 561.600 487.050 562.050 ;
        RECT 496.950 561.600 499.050 562.050 ;
        RECT 484.950 560.400 499.050 561.600 ;
        RECT 484.950 559.950 487.050 560.400 ;
        RECT 496.950 559.950 499.050 560.400 ;
        RECT 502.950 561.600 505.050 562.050 ;
        RECT 511.950 561.600 514.050 562.050 ;
        RECT 502.950 560.400 514.050 561.600 ;
        RECT 502.950 559.950 505.050 560.400 ;
        RECT 511.950 559.950 514.050 560.400 ;
        RECT 517.950 561.600 520.050 562.050 ;
        RECT 535.950 561.600 538.050 562.050 ;
        RECT 517.950 560.400 538.050 561.600 ;
        RECT 517.950 559.950 520.050 560.400 ;
        RECT 535.950 559.950 538.050 560.400 ;
        RECT 556.950 561.600 559.050 562.050 ;
        RECT 565.950 561.600 568.050 562.050 ;
        RECT 556.950 560.400 568.050 561.600 ;
        RECT 556.950 559.950 559.050 560.400 ;
        RECT 565.950 559.950 568.050 560.400 ;
        RECT 664.950 559.950 667.050 562.050 ;
        RECT 400.950 558.600 403.050 559.050 ;
        RECT 406.950 558.600 409.050 559.050 ;
        RECT 424.950 558.600 427.050 559.050 ;
        RECT 400.950 557.400 405.600 558.600 ;
        RECT 400.950 556.950 403.050 557.400 ;
        RECT 370.950 554.400 387.600 555.600 ;
        RECT 404.400 555.600 405.600 557.400 ;
        RECT 406.950 557.400 427.050 558.600 ;
        RECT 406.950 556.950 409.050 557.400 ;
        RECT 424.950 556.950 427.050 557.400 ;
        RECT 436.950 558.600 439.050 559.050 ;
        RECT 461.400 558.600 462.600 559.950 ;
        RECT 481.950 558.600 484.050 559.050 ;
        RECT 436.950 557.400 484.050 558.600 ;
        RECT 436.950 556.950 439.050 557.400 ;
        RECT 481.950 556.950 484.050 557.400 ;
        RECT 499.950 558.600 502.050 559.050 ;
        RECT 514.950 558.600 517.050 559.050 ;
        RECT 499.950 557.400 517.050 558.600 ;
        RECT 499.950 556.950 502.050 557.400 ;
        RECT 514.950 556.950 517.050 557.400 ;
        RECT 559.950 558.600 562.050 559.050 ;
        RECT 601.950 558.600 604.050 559.050 ;
        RECT 619.950 558.600 622.050 559.050 ;
        RECT 559.950 557.400 622.050 558.600 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 601.950 556.950 604.050 557.400 ;
        RECT 619.950 556.950 622.050 557.400 ;
        RECT 655.950 556.950 658.050 559.050 ;
        RECT 665.400 558.600 666.600 559.950 ;
        RECT 662.400 557.400 666.600 558.600 ;
        RECT 676.950 558.600 679.050 559.050 ;
        RECT 694.950 558.600 697.050 559.050 ;
        RECT 676.950 557.400 697.050 558.600 ;
        RECT 406.950 555.600 409.050 556.050 ;
        RECT 404.400 554.400 409.050 555.600 ;
        RECT 370.950 553.950 373.050 554.400 ;
        RECT 406.950 553.950 409.050 554.400 ;
        RECT 439.950 555.600 442.050 556.050 ;
        RECT 448.950 555.600 451.050 556.050 ;
        RECT 439.950 554.400 451.050 555.600 ;
        RECT 439.950 553.950 442.050 554.400 ;
        RECT 448.950 553.950 451.050 554.400 ;
        RECT 454.950 555.600 457.050 556.050 ;
        RECT 466.950 555.600 469.050 556.050 ;
        RECT 454.950 554.400 469.050 555.600 ;
        RECT 454.950 553.950 457.050 554.400 ;
        RECT 466.950 553.950 469.050 554.400 ;
        RECT 544.950 555.600 547.050 556.050 ;
        RECT 553.950 555.600 556.050 556.050 ;
        RECT 544.950 554.400 556.050 555.600 ;
        RECT 544.950 553.950 547.050 554.400 ;
        RECT 553.950 553.950 556.050 554.400 ;
        RECT 610.950 555.600 613.050 556.050 ;
        RECT 631.950 555.600 634.050 556.050 ;
        RECT 610.950 554.400 634.050 555.600 ;
        RECT 610.950 553.950 613.050 554.400 ;
        RECT 631.950 553.950 634.050 554.400 ;
        RECT 656.400 553.050 657.600 556.950 ;
        RECT 658.950 555.600 661.050 556.050 ;
        RECT 662.400 555.600 663.600 557.400 ;
        RECT 676.950 556.950 679.050 557.400 ;
        RECT 694.950 556.950 697.050 557.400 ;
        RECT 718.950 558.600 721.050 559.050 ;
        RECT 754.950 558.600 757.050 559.050 ;
        RECT 718.950 557.400 757.050 558.600 ;
        RECT 718.950 556.950 721.050 557.400 ;
        RECT 754.950 556.950 757.050 557.400 ;
        RECT 784.950 558.600 787.050 559.050 ;
        RECT 793.950 558.600 796.050 559.050 ;
        RECT 814.950 558.600 817.050 559.050 ;
        RECT 859.950 558.600 862.050 559.050 ;
        RECT 866.400 558.600 867.600 563.400 ;
        RECT 784.950 557.400 804.600 558.600 ;
        RECT 784.950 556.950 787.050 557.400 ;
        RECT 793.950 556.950 796.050 557.400 ;
        RECT 658.950 554.400 663.600 555.600 ;
        RECT 664.950 555.600 667.050 556.050 ;
        RECT 667.950 555.600 670.050 556.050 ;
        RECT 697.950 555.600 700.050 556.050 ;
        RECT 664.950 554.400 700.050 555.600 ;
        RECT 803.400 555.600 804.600 557.400 ;
        RECT 814.950 557.400 831.600 558.600 ;
        RECT 814.950 556.950 817.050 557.400 ;
        RECT 826.950 555.600 829.050 556.050 ;
        RECT 803.400 554.400 829.050 555.600 ;
        RECT 830.400 555.600 831.600 557.400 ;
        RECT 859.950 557.400 867.600 558.600 ;
        RECT 859.950 556.950 862.050 557.400 ;
        RECT 856.950 555.600 859.050 556.050 ;
        RECT 830.400 554.400 859.050 555.600 ;
        RECT 658.950 553.950 661.050 554.400 ;
        RECT 664.950 553.950 667.050 554.400 ;
        RECT 667.950 553.950 670.050 554.400 ;
        RECT 697.950 553.950 700.050 554.400 ;
        RECT 826.950 553.950 829.050 554.400 ;
        RECT 856.950 553.950 859.050 554.400 ;
        RECT 91.950 552.600 94.050 553.050 ;
        RECT 115.950 552.600 118.050 553.050 ;
        RECT 91.950 551.400 118.050 552.600 ;
        RECT 91.950 550.950 94.050 551.400 ;
        RECT 115.950 550.950 118.050 551.400 ;
        RECT 151.950 552.600 154.050 553.050 ;
        RECT 163.950 552.600 166.050 553.050 ;
        RECT 223.950 552.600 226.050 553.050 ;
        RECT 247.950 552.600 250.050 553.050 ;
        RECT 151.950 551.400 166.050 552.600 ;
        RECT 151.950 550.950 154.050 551.400 ;
        RECT 163.950 550.950 166.050 551.400 ;
        RECT 191.400 551.400 222.600 552.600 ;
        RECT 85.950 549.600 88.050 550.050 ;
        RECT 191.400 549.600 192.600 551.400 ;
        RECT 208.950 549.600 211.050 550.050 ;
        RECT 85.950 548.400 192.600 549.600 ;
        RECT 194.400 548.400 211.050 549.600 ;
        RECT 221.400 549.600 222.600 551.400 ;
        RECT 223.950 551.400 250.050 552.600 ;
        RECT 223.950 550.950 226.050 551.400 ;
        RECT 247.950 550.950 250.050 551.400 ;
        RECT 295.950 552.600 298.050 553.050 ;
        RECT 304.950 552.600 307.050 553.050 ;
        RECT 388.950 552.600 391.050 553.050 ;
        RECT 295.950 551.400 391.050 552.600 ;
        RECT 295.950 550.950 298.050 551.400 ;
        RECT 304.950 550.950 307.050 551.400 ;
        RECT 388.950 550.950 391.050 551.400 ;
        RECT 403.950 552.600 406.050 553.050 ;
        RECT 418.950 552.600 421.050 553.050 ;
        RECT 424.950 552.600 427.050 553.050 ;
        RECT 403.950 551.400 427.050 552.600 ;
        RECT 403.950 550.950 406.050 551.400 ;
        RECT 418.950 550.950 421.050 551.400 ;
        RECT 424.950 550.950 427.050 551.400 ;
        RECT 445.950 552.600 448.050 553.050 ;
        RECT 469.950 552.600 472.050 553.050 ;
        RECT 445.950 551.400 472.050 552.600 ;
        RECT 445.950 550.950 448.050 551.400 ;
        RECT 469.950 550.950 472.050 551.400 ;
        RECT 493.950 552.600 496.050 553.050 ;
        RECT 499.950 552.600 502.050 553.050 ;
        RECT 493.950 551.400 502.050 552.600 ;
        RECT 493.950 550.950 496.050 551.400 ;
        RECT 499.950 550.950 502.050 551.400 ;
        RECT 532.950 552.600 535.050 553.050 ;
        RECT 541.950 552.600 544.050 553.050 ;
        RECT 532.950 551.400 544.050 552.600 ;
        RECT 532.950 550.950 535.050 551.400 ;
        RECT 541.950 550.950 544.050 551.400 ;
        RECT 655.950 550.950 658.050 553.050 ;
        RECT 661.950 552.600 664.050 553.050 ;
        RECT 670.950 552.600 673.050 553.050 ;
        RECT 661.950 551.400 673.050 552.600 ;
        RECT 661.950 550.950 664.050 551.400 ;
        RECT 670.950 550.950 673.050 551.400 ;
        RECT 682.950 552.600 685.050 553.050 ;
        RECT 694.950 552.600 697.050 553.050 ;
        RECT 682.950 551.400 697.050 552.600 ;
        RECT 682.950 550.950 685.050 551.400 ;
        RECT 694.950 550.950 697.050 551.400 ;
        RECT 730.950 552.600 733.050 553.050 ;
        RECT 760.950 552.600 763.050 553.050 ;
        RECT 766.950 552.600 769.050 553.050 ;
        RECT 730.950 551.400 769.050 552.600 ;
        RECT 730.950 550.950 733.050 551.400 ;
        RECT 760.950 550.950 763.050 551.400 ;
        RECT 766.950 550.950 769.050 551.400 ;
        RECT 289.950 549.600 292.050 550.050 ;
        RECT 298.950 549.600 301.050 550.050 ;
        RECT 221.400 548.400 301.050 549.600 ;
        RECT 85.950 547.950 88.050 548.400 ;
        RECT 106.950 546.600 109.050 547.050 ;
        RECT 194.400 546.600 195.600 548.400 ;
        RECT 208.950 547.950 211.050 548.400 ;
        RECT 289.950 547.950 292.050 548.400 ;
        RECT 298.950 547.950 301.050 548.400 ;
        RECT 337.950 549.600 340.050 550.050 ;
        RECT 376.950 549.600 379.050 550.050 ;
        RECT 394.950 549.600 397.050 550.050 ;
        RECT 439.950 549.600 442.050 550.050 ;
        RECT 337.950 548.400 442.050 549.600 ;
        RECT 337.950 547.950 340.050 548.400 ;
        RECT 376.950 547.950 379.050 548.400 ;
        RECT 394.950 547.950 397.050 548.400 ;
        RECT 439.950 547.950 442.050 548.400 ;
        RECT 460.950 549.600 463.050 550.050 ;
        RECT 559.950 549.600 562.050 550.050 ;
        RECT 460.950 548.400 562.050 549.600 ;
        RECT 460.950 547.950 463.050 548.400 ;
        RECT 559.950 547.950 562.050 548.400 ;
        RECT 568.950 549.600 571.050 550.050 ;
        RECT 574.950 549.600 577.050 550.050 ;
        RECT 568.950 548.400 577.050 549.600 ;
        RECT 568.950 547.950 571.050 548.400 ;
        RECT 574.950 547.950 577.050 548.400 ;
        RECT 619.950 549.600 622.050 550.050 ;
        RECT 712.950 549.600 715.050 550.050 ;
        RECT 619.950 548.400 715.050 549.600 ;
        RECT 619.950 547.950 622.050 548.400 ;
        RECT 712.950 547.950 715.050 548.400 ;
        RECT 832.950 549.600 835.050 550.050 ;
        RECT 850.950 549.600 853.050 550.050 ;
        RECT 832.950 548.400 853.050 549.600 ;
        RECT 832.950 547.950 835.050 548.400 ;
        RECT 850.950 547.950 853.050 548.400 ;
        RECT 106.950 545.400 195.600 546.600 ;
        RECT 196.950 546.600 199.050 547.050 ;
        RECT 205.950 546.600 208.050 547.050 ;
        RECT 196.950 545.400 208.050 546.600 ;
        RECT 106.950 544.950 109.050 545.400 ;
        RECT 196.950 544.950 199.050 545.400 ;
        RECT 205.950 544.950 208.050 545.400 ;
        RECT 232.950 546.600 235.050 547.050 ;
        RECT 238.950 546.600 241.050 547.050 ;
        RECT 232.950 545.400 241.050 546.600 ;
        RECT 232.950 544.950 235.050 545.400 ;
        RECT 238.950 544.950 241.050 545.400 ;
        RECT 283.950 546.600 286.050 547.050 ;
        RECT 364.950 546.600 367.050 547.050 ;
        RECT 283.950 545.400 367.050 546.600 ;
        RECT 283.950 544.950 286.050 545.400 ;
        RECT 364.950 544.950 367.050 545.400 ;
        RECT 376.950 546.600 379.050 547.050 ;
        RECT 409.950 546.600 412.050 547.050 ;
        RECT 376.950 545.400 412.050 546.600 ;
        RECT 376.950 544.950 379.050 545.400 ;
        RECT 409.950 544.950 412.050 545.400 ;
        RECT 487.950 546.600 490.050 547.050 ;
        RECT 490.950 546.600 493.050 547.050 ;
        RECT 550.950 546.600 553.050 547.050 ;
        RECT 487.950 545.400 553.050 546.600 ;
        RECT 487.950 544.950 490.050 545.400 ;
        RECT 490.950 544.950 493.050 545.400 ;
        RECT 550.950 544.950 553.050 545.400 ;
        RECT 583.950 546.600 586.050 547.050 ;
        RECT 598.950 546.600 601.050 547.050 ;
        RECT 583.950 545.400 601.050 546.600 ;
        RECT 583.950 544.950 586.050 545.400 ;
        RECT 598.950 544.950 601.050 545.400 ;
        RECT 178.950 543.600 181.050 544.050 ;
        RECT 181.950 543.600 184.050 544.050 ;
        RECT 190.950 543.600 193.050 544.050 ;
        RECT 178.950 542.400 193.050 543.600 ;
        RECT 178.950 541.950 181.050 542.400 ;
        RECT 181.950 541.950 184.050 542.400 ;
        RECT 190.950 541.950 193.050 542.400 ;
        RECT 238.950 543.600 241.050 544.050 ;
        RECT 331.950 543.600 334.050 544.050 ;
        RECT 238.950 542.400 334.050 543.600 ;
        RECT 238.950 541.950 241.050 542.400 ;
        RECT 331.950 541.950 334.050 542.400 ;
        RECT 388.950 543.600 391.050 544.050 ;
        RECT 409.950 543.600 412.050 544.050 ;
        RECT 544.950 543.600 547.050 544.050 ;
        RECT 388.950 542.400 547.050 543.600 ;
        RECT 388.950 541.950 391.050 542.400 ;
        RECT 409.950 541.950 412.050 542.400 ;
        RECT 544.950 541.950 547.050 542.400 ;
        RECT 550.950 543.600 553.050 544.050 ;
        RECT 583.950 543.600 586.050 544.050 ;
        RECT 550.950 542.400 586.050 543.600 ;
        RECT 550.950 541.950 553.050 542.400 ;
        RECT 583.950 541.950 586.050 542.400 ;
        RECT 595.950 543.600 598.050 544.050 ;
        RECT 604.950 543.600 607.050 544.050 ;
        RECT 595.950 542.400 607.050 543.600 ;
        RECT 595.950 541.950 598.050 542.400 ;
        RECT 604.950 541.950 607.050 542.400 ;
        RECT 13.950 540.600 16.050 541.050 ;
        RECT 31.950 540.600 34.050 541.050 ;
        RECT 13.950 539.400 34.050 540.600 ;
        RECT 13.950 538.950 16.050 539.400 ;
        RECT 31.950 538.950 34.050 539.400 ;
        RECT 205.950 540.600 208.050 541.050 ;
        RECT 460.950 540.600 463.050 541.050 ;
        RECT 205.950 539.400 463.050 540.600 ;
        RECT 205.950 538.950 208.050 539.400 ;
        RECT 460.950 538.950 463.050 539.400 ;
        RECT 463.950 540.600 466.050 541.050 ;
        RECT 580.950 540.600 583.050 541.050 ;
        RECT 463.950 539.400 583.050 540.600 ;
        RECT 463.950 538.950 466.050 539.400 ;
        RECT 580.950 538.950 583.050 539.400 ;
        RECT 622.950 540.600 625.050 541.050 ;
        RECT 700.950 540.600 703.050 541.050 ;
        RECT 622.950 539.400 703.050 540.600 ;
        RECT 622.950 538.950 625.050 539.400 ;
        RECT 700.950 538.950 703.050 539.400 ;
        RECT 709.950 540.600 712.050 541.050 ;
        RECT 715.950 540.600 718.050 541.050 ;
        RECT 709.950 539.400 718.050 540.600 ;
        RECT 709.950 538.950 712.050 539.400 ;
        RECT 715.950 538.950 718.050 539.400 ;
        RECT 13.950 537.600 16.050 538.050 ;
        RECT 40.950 537.600 43.050 538.050 ;
        RECT 13.950 536.400 43.050 537.600 ;
        RECT 13.950 535.950 16.050 536.400 ;
        RECT 40.950 535.950 43.050 536.400 ;
        RECT 43.950 537.600 46.050 538.050 ;
        RECT 61.950 537.600 64.050 538.050 ;
        RECT 43.950 536.400 64.050 537.600 ;
        RECT 43.950 535.950 46.050 536.400 ;
        RECT 61.950 535.950 64.050 536.400 ;
        RECT 100.950 537.600 103.050 538.050 ;
        RECT 133.950 537.600 136.050 538.050 ;
        RECT 145.950 537.600 148.050 538.050 ;
        RECT 100.950 536.400 148.050 537.600 ;
        RECT 100.950 535.950 103.050 536.400 ;
        RECT 133.950 535.950 136.050 536.400 ;
        RECT 145.950 535.950 148.050 536.400 ;
        RECT 262.950 537.600 265.050 538.050 ;
        RECT 337.950 537.600 340.050 538.050 ;
        RECT 262.950 536.400 340.050 537.600 ;
        RECT 262.950 535.950 265.050 536.400 ;
        RECT 337.950 535.950 340.050 536.400 ;
        RECT 358.950 537.600 361.050 538.050 ;
        RECT 364.950 537.600 367.050 538.050 ;
        RECT 358.950 536.400 367.050 537.600 ;
        RECT 358.950 535.950 361.050 536.400 ;
        RECT 364.950 535.950 367.050 536.400 ;
        RECT 433.950 537.600 436.050 538.050 ;
        RECT 475.950 537.600 478.050 538.050 ;
        RECT 433.950 536.400 478.050 537.600 ;
        RECT 433.950 535.950 436.050 536.400 ;
        RECT 475.950 535.950 478.050 536.400 ;
        RECT 529.950 537.600 532.050 538.050 ;
        RECT 541.950 537.600 544.050 538.050 ;
        RECT 565.950 537.600 568.050 538.050 ;
        RECT 529.950 536.400 568.050 537.600 ;
        RECT 529.950 535.950 532.050 536.400 ;
        RECT 541.950 535.950 544.050 536.400 ;
        RECT 565.950 535.950 568.050 536.400 ;
        RECT 628.950 537.600 631.050 538.050 ;
        RECT 643.950 537.600 646.050 538.050 ;
        RECT 628.950 536.400 646.050 537.600 ;
        RECT 628.950 535.950 631.050 536.400 ;
        RECT 643.950 535.950 646.050 536.400 ;
        RECT 652.950 537.600 655.050 538.050 ;
        RECT 733.950 537.600 736.050 538.050 ;
        RECT 652.950 536.400 736.050 537.600 ;
        RECT 652.950 535.950 655.050 536.400 ;
        RECT 733.950 535.950 736.050 536.400 ;
        RECT 775.950 537.600 778.050 538.050 ;
        RECT 784.950 537.600 787.050 538.050 ;
        RECT 775.950 536.400 787.050 537.600 ;
        RECT 775.950 535.950 778.050 536.400 ;
        RECT 784.950 535.950 787.050 536.400 ;
        RECT 19.950 534.600 22.050 535.050 ;
        RECT 55.950 534.600 58.050 535.050 ;
        RECT 19.950 533.400 58.050 534.600 ;
        RECT 19.950 532.950 22.050 533.400 ;
        RECT 55.950 532.950 58.050 533.400 ;
        RECT 73.950 534.600 76.050 535.050 ;
        RECT 166.950 534.600 169.050 535.050 ;
        RECT 73.950 533.400 169.050 534.600 ;
        RECT 73.950 532.950 76.050 533.400 ;
        RECT 166.950 532.950 169.050 533.400 ;
        RECT 256.950 534.600 259.050 535.050 ;
        RECT 298.950 534.600 301.050 535.050 ;
        RECT 256.950 533.400 301.050 534.600 ;
        RECT 256.950 532.950 259.050 533.400 ;
        RECT 298.950 532.950 301.050 533.400 ;
        RECT 340.950 534.600 343.050 535.050 ;
        RECT 532.950 534.600 535.050 535.050 ;
        RECT 340.950 533.400 535.050 534.600 ;
        RECT 340.950 532.950 343.050 533.400 ;
        RECT 532.950 532.950 535.050 533.400 ;
        RECT 547.950 534.600 550.050 535.050 ;
        RECT 628.950 534.600 631.050 535.050 ;
        RECT 547.950 533.400 631.050 534.600 ;
        RECT 547.950 532.950 550.050 533.400 ;
        RECT 628.950 532.950 631.050 533.400 ;
        RECT 640.950 534.600 643.050 535.050 ;
        RECT 697.950 534.600 700.050 535.050 ;
        RECT 640.950 533.400 700.050 534.600 ;
        RECT 640.950 532.950 643.050 533.400 ;
        RECT 697.950 532.950 700.050 533.400 ;
        RECT 754.950 534.600 757.050 535.050 ;
        RECT 796.950 534.600 799.050 535.050 ;
        RECT 754.950 533.400 799.050 534.600 ;
        RECT 754.950 532.950 757.050 533.400 ;
        RECT 796.950 532.950 799.050 533.400 ;
        RECT 31.950 531.600 34.050 532.050 ;
        RECT 17.400 530.400 34.050 531.600 ;
        RECT 17.400 526.050 18.600 530.400 ;
        RECT 31.950 529.950 34.050 530.400 ;
        RECT 55.950 531.600 58.050 532.050 ;
        RECT 91.950 531.600 94.050 532.050 ;
        RECT 55.950 530.400 94.050 531.600 ;
        RECT 55.950 529.950 58.050 530.400 ;
        RECT 91.950 529.950 94.050 530.400 ;
        RECT 142.950 531.600 145.050 532.050 ;
        RECT 157.950 531.600 160.050 532.050 ;
        RECT 142.950 530.400 160.050 531.600 ;
        RECT 142.950 529.950 145.050 530.400 ;
        RECT 157.950 529.950 160.050 530.400 ;
        RECT 247.950 531.600 250.050 532.050 ;
        RECT 256.950 531.600 259.050 532.050 ;
        RECT 247.950 530.400 259.050 531.600 ;
        RECT 247.950 529.950 250.050 530.400 ;
        RECT 256.950 529.950 259.050 530.400 ;
        RECT 286.950 531.600 289.050 532.050 ;
        RECT 292.950 531.600 295.050 532.050 ;
        RECT 286.950 530.400 295.050 531.600 ;
        RECT 286.950 529.950 289.050 530.400 ;
        RECT 292.950 529.950 295.050 530.400 ;
        RECT 325.950 531.600 328.050 532.050 ;
        RECT 349.950 531.600 352.050 532.050 ;
        RECT 358.950 531.600 361.050 532.050 ;
        RECT 325.950 530.400 361.050 531.600 ;
        RECT 325.950 529.950 328.050 530.400 ;
        RECT 349.950 529.950 352.050 530.400 ;
        RECT 358.950 529.950 361.050 530.400 ;
        RECT 448.950 531.600 451.050 532.050 ;
        RECT 454.950 531.600 457.050 532.050 ;
        RECT 448.950 530.400 457.050 531.600 ;
        RECT 448.950 529.950 451.050 530.400 ;
        RECT 454.950 529.950 457.050 530.400 ;
        RECT 457.950 531.600 460.050 532.050 ;
        RECT 508.950 531.600 511.050 532.050 ;
        RECT 457.950 530.400 511.050 531.600 ;
        RECT 457.950 529.950 460.050 530.400 ;
        RECT 508.950 529.950 511.050 530.400 ;
        RECT 511.950 531.600 514.050 532.050 ;
        RECT 523.950 531.600 526.050 532.050 ;
        RECT 511.950 530.400 526.050 531.600 ;
        RECT 511.950 529.950 514.050 530.400 ;
        RECT 523.950 529.950 526.050 530.400 ;
        RECT 526.950 529.950 529.050 532.050 ;
        RECT 553.950 531.600 556.050 532.050 ;
        RECT 607.950 531.600 610.050 532.050 ;
        RECT 553.950 530.400 610.050 531.600 ;
        RECT 553.950 529.950 556.050 530.400 ;
        RECT 607.950 529.950 610.050 530.400 ;
        RECT 622.950 531.600 625.050 532.050 ;
        RECT 631.950 531.600 634.050 532.050 ;
        RECT 622.950 530.400 634.050 531.600 ;
        RECT 622.950 529.950 625.050 530.400 ;
        RECT 631.950 529.950 634.050 530.400 ;
        RECT 700.950 531.600 703.050 532.050 ;
        RECT 703.950 531.600 706.050 532.050 ;
        RECT 799.950 531.600 802.050 532.050 ;
        RECT 700.950 530.400 802.050 531.600 ;
        RECT 700.950 529.950 703.050 530.400 ;
        RECT 703.950 529.950 706.050 530.400 ;
        RECT 799.950 529.950 802.050 530.400 ;
        RECT 19.950 528.600 22.050 529.050 ;
        RECT 37.950 528.600 40.050 529.050 ;
        RECT 43.950 528.600 46.050 529.050 ;
        RECT 19.950 527.400 30.600 528.600 ;
        RECT 19.950 526.950 22.050 527.400 ;
        RECT 29.400 526.050 30.600 527.400 ;
        RECT 37.950 527.400 46.050 528.600 ;
        RECT 37.950 526.950 40.050 527.400 ;
        RECT 43.950 526.950 46.050 527.400 ;
        RECT 70.950 528.600 73.050 529.050 ;
        RECT 88.950 528.600 91.050 529.050 ;
        RECT 70.950 527.400 91.050 528.600 ;
        RECT 70.950 526.950 73.050 527.400 ;
        RECT 88.950 526.950 91.050 527.400 ;
        RECT 136.950 528.600 139.050 529.050 ;
        RECT 163.950 528.600 166.050 529.050 ;
        RECT 172.950 528.600 175.050 529.050 ;
        RECT 136.950 527.400 175.050 528.600 ;
        RECT 136.950 526.950 139.050 527.400 ;
        RECT 163.950 526.950 166.050 527.400 ;
        RECT 172.950 526.950 175.050 527.400 ;
        RECT 199.950 528.600 202.050 529.050 ;
        RECT 211.950 528.600 214.050 529.050 ;
        RECT 250.950 528.600 253.050 529.050 ;
        RECT 199.950 527.400 214.050 528.600 ;
        RECT 199.950 526.950 202.050 527.400 ;
        RECT 211.950 526.950 214.050 527.400 ;
        RECT 230.400 527.400 253.050 528.600 ;
        RECT 230.400 526.050 231.600 527.400 ;
        RECT 250.950 526.950 253.050 527.400 ;
        RECT 274.950 528.600 277.050 529.050 ;
        RECT 301.950 528.600 304.050 529.050 ;
        RECT 274.950 527.400 304.050 528.600 ;
        RECT 274.950 526.950 277.050 527.400 ;
        RECT 301.950 526.950 304.050 527.400 ;
        RECT 307.950 528.600 310.050 529.050 ;
        RECT 322.950 528.600 325.050 529.050 ;
        RECT 343.950 528.600 346.050 529.050 ;
        RECT 307.950 527.400 346.050 528.600 ;
        RECT 307.950 526.950 310.050 527.400 ;
        RECT 322.950 526.950 325.050 527.400 ;
        RECT 16.950 523.950 19.050 526.050 ;
        RECT 28.950 523.950 31.050 526.050 ;
        RECT 34.950 525.600 37.050 526.050 ;
        RECT 40.950 525.600 43.050 526.050 ;
        RECT 34.950 524.400 43.050 525.600 ;
        RECT 34.950 523.950 37.050 524.400 ;
        RECT 40.950 523.950 43.050 524.400 ;
        RECT 58.950 525.600 61.050 526.050 ;
        RECT 67.950 525.600 70.050 526.050 ;
        RECT 58.950 524.400 70.050 525.600 ;
        RECT 58.950 523.950 61.050 524.400 ;
        RECT 67.950 523.950 70.050 524.400 ;
        RECT 139.950 525.600 142.050 526.050 ;
        RECT 148.950 525.600 151.050 526.050 ;
        RECT 139.950 524.400 151.050 525.600 ;
        RECT 139.950 523.950 142.050 524.400 ;
        RECT 148.950 523.950 151.050 524.400 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 190.950 525.600 193.050 526.050 ;
        RECT 199.950 525.600 202.050 526.050 ;
        RECT 190.950 524.400 202.050 525.600 ;
        RECT 190.950 523.950 193.050 524.400 ;
        RECT 199.950 523.950 202.050 524.400 ;
        RECT 217.950 523.950 220.050 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 235.950 525.600 238.050 526.050 ;
        RECT 241.950 525.600 244.050 526.050 ;
        RECT 235.950 524.400 244.050 525.600 ;
        RECT 235.950 523.950 238.050 524.400 ;
        RECT 241.950 523.950 244.050 524.400 ;
        RECT 265.950 525.600 268.050 526.050 ;
        RECT 277.950 525.600 280.050 526.050 ;
        RECT 265.950 524.400 280.050 525.600 ;
        RECT 265.950 523.950 268.050 524.400 ;
        RECT 277.950 523.950 280.050 524.400 ;
        RECT 280.950 525.600 283.050 526.050 ;
        RECT 286.950 525.600 289.050 526.050 ;
        RECT 280.950 524.400 289.050 525.600 ;
        RECT 280.950 523.950 283.050 524.400 ;
        RECT 286.950 523.950 289.050 524.400 ;
        RECT 301.950 525.600 304.050 526.050 ;
        RECT 313.950 525.600 316.050 526.050 ;
        RECT 301.950 524.400 316.050 525.600 ;
        RECT 301.950 523.950 304.050 524.400 ;
        RECT 313.950 523.950 316.050 524.400 ;
        RECT 319.950 525.600 322.050 526.050 ;
        RECT 325.950 525.600 328.050 526.050 ;
        RECT 319.950 524.400 328.050 525.600 ;
        RECT 319.950 523.950 322.050 524.400 ;
        RECT 325.950 523.950 328.050 524.400 ;
        RECT 136.950 522.600 139.050 523.050 ;
        RECT 155.400 522.600 156.600 523.950 ;
        RECT 136.950 521.400 156.600 522.600 ;
        RECT 175.950 522.600 178.050 523.050 ;
        RECT 187.950 522.600 190.050 523.050 ;
        RECT 175.950 521.400 190.050 522.600 ;
        RECT 136.950 520.950 139.050 521.400 ;
        RECT 175.950 520.950 178.050 521.400 ;
        RECT 187.950 520.950 190.050 521.400 ;
        RECT 202.950 522.600 205.050 523.050 ;
        RECT 208.950 522.600 211.050 523.050 ;
        RECT 202.950 521.400 211.050 522.600 ;
        RECT 202.950 520.950 205.050 521.400 ;
        RECT 208.950 520.950 211.050 521.400 ;
        RECT 214.950 520.950 217.050 523.050 ;
        RECT 218.400 522.600 219.600 523.950 ;
        RECT 241.950 522.600 244.050 523.050 ;
        RECT 218.400 521.400 244.050 522.600 ;
        RECT 241.950 520.950 244.050 521.400 ;
        RECT 247.950 522.600 250.050 523.050 ;
        RECT 253.950 522.600 256.050 523.050 ;
        RECT 271.950 522.600 274.050 523.050 ;
        RECT 247.950 521.400 274.050 522.600 ;
        RECT 247.950 520.950 250.050 521.400 ;
        RECT 253.950 520.950 256.050 521.400 ;
        RECT 271.950 520.950 274.050 521.400 ;
        RECT 295.950 522.600 298.050 523.050 ;
        RECT 331.950 522.600 334.050 523.050 ;
        RECT 295.950 521.400 334.050 522.600 ;
        RECT 335.400 522.600 336.600 527.400 ;
        RECT 343.950 526.950 346.050 527.400 ;
        RECT 352.950 528.600 355.050 529.050 ;
        RECT 379.950 528.600 382.050 529.050 ;
        RECT 352.950 527.400 382.050 528.600 ;
        RECT 352.950 526.950 355.050 527.400 ;
        RECT 379.950 526.950 382.050 527.400 ;
        RECT 385.950 528.600 388.050 529.050 ;
        RECT 421.950 528.600 424.050 529.050 ;
        RECT 385.950 527.400 424.050 528.600 ;
        RECT 385.950 526.950 388.050 527.400 ;
        RECT 421.950 526.950 424.050 527.400 ;
        RECT 430.950 528.600 433.050 529.050 ;
        RECT 457.950 528.600 460.050 529.050 ;
        RECT 430.950 527.400 460.050 528.600 ;
        RECT 430.950 526.950 433.050 527.400 ;
        RECT 457.950 526.950 460.050 527.400 ;
        RECT 478.950 528.600 481.050 529.050 ;
        RECT 527.400 528.600 528.600 529.950 ;
        RECT 562.950 528.600 565.050 529.050 ;
        RECT 580.950 528.600 583.050 529.050 ;
        RECT 478.950 527.400 528.600 528.600 ;
        RECT 548.400 527.400 565.050 528.600 ;
        RECT 478.950 526.950 481.050 527.400 ;
        RECT 548.400 526.050 549.600 527.400 ;
        RECT 562.950 526.950 565.050 527.400 ;
        RECT 566.400 527.400 583.050 528.600 ;
        RECT 337.950 525.600 340.050 526.050 ;
        RECT 349.950 525.600 352.050 526.050 ;
        RECT 337.950 524.400 352.050 525.600 ;
        RECT 337.950 523.950 340.050 524.400 ;
        RECT 349.950 523.950 352.050 524.400 ;
        RECT 355.950 525.600 358.050 526.050 ;
        RECT 367.950 525.600 370.050 526.050 ;
        RECT 400.950 525.600 403.050 526.050 ;
        RECT 409.950 525.600 412.050 526.050 ;
        RECT 355.950 524.400 370.050 525.600 ;
        RECT 355.950 523.950 358.050 524.400 ;
        RECT 367.950 523.950 370.050 524.400 ;
        RECT 371.400 524.400 403.050 525.600 ;
        RECT 371.400 522.600 372.600 524.400 ;
        RECT 400.950 523.950 403.050 524.400 ;
        RECT 404.400 524.400 412.050 525.600 ;
        RECT 404.400 523.050 405.600 524.400 ;
        RECT 409.950 523.950 412.050 524.400 ;
        RECT 418.950 525.600 421.050 526.050 ;
        RECT 430.950 525.600 433.050 526.050 ;
        RECT 418.950 524.400 433.050 525.600 ;
        RECT 418.950 523.950 421.050 524.400 ;
        RECT 430.950 523.950 433.050 524.400 ;
        RECT 457.950 525.600 460.050 526.050 ;
        RECT 475.950 525.600 478.050 526.050 ;
        RECT 457.950 524.400 478.050 525.600 ;
        RECT 457.950 523.950 460.050 524.400 ;
        RECT 475.950 523.950 478.050 524.400 ;
        RECT 481.950 525.600 484.050 526.050 ;
        RECT 487.950 525.600 490.050 526.050 ;
        RECT 502.950 525.600 505.050 526.050 ;
        RECT 520.950 525.600 523.050 526.050 ;
        RECT 481.950 524.400 490.050 525.600 ;
        RECT 481.950 523.950 484.050 524.400 ;
        RECT 487.950 523.950 490.050 524.400 ;
        RECT 497.400 524.400 523.050 525.600 ;
        RECT 335.400 521.400 372.600 522.600 ;
        RECT 382.950 522.600 385.050 523.050 ;
        RECT 397.950 522.600 400.050 523.050 ;
        RECT 382.950 521.400 400.050 522.600 ;
        RECT 295.950 520.950 298.050 521.400 ;
        RECT 331.950 520.950 334.050 521.400 ;
        RECT 382.950 520.950 385.050 521.400 ;
        RECT 397.950 520.950 400.050 521.400 ;
        RECT 403.950 520.950 406.050 523.050 ;
        RECT 406.950 522.600 409.050 523.050 ;
        RECT 424.950 522.600 427.050 523.050 ;
        RECT 406.950 521.400 427.050 522.600 ;
        RECT 406.950 520.950 409.050 521.400 ;
        RECT 424.950 520.950 427.050 521.400 ;
        RECT 427.950 522.600 430.050 523.050 ;
        RECT 478.950 522.600 481.050 523.050 ;
        RECT 427.950 521.400 481.050 522.600 ;
        RECT 427.950 520.950 430.050 521.400 ;
        RECT 478.950 520.950 481.050 521.400 ;
        RECT 484.950 522.600 487.050 523.050 ;
        RECT 497.400 522.600 498.600 524.400 ;
        RECT 502.950 523.950 505.050 524.400 ;
        RECT 520.950 523.950 523.050 524.400 ;
        RECT 526.950 525.600 529.050 526.050 ;
        RECT 547.950 525.600 550.050 526.050 ;
        RECT 526.950 524.400 550.050 525.600 ;
        RECT 526.950 523.950 529.050 524.400 ;
        RECT 547.950 523.950 550.050 524.400 ;
        RECT 566.400 523.050 567.600 527.400 ;
        RECT 580.950 526.950 583.050 527.400 ;
        RECT 586.950 526.950 589.050 529.050 ;
        RECT 598.950 528.600 601.050 529.050 ;
        RECT 646.950 528.600 649.050 529.050 ;
        RECT 691.950 528.600 694.050 529.050 ;
        RECT 598.950 527.400 694.050 528.600 ;
        RECT 598.950 526.950 601.050 527.400 ;
        RECT 646.950 526.950 649.050 527.400 ;
        RECT 691.950 526.950 694.050 527.400 ;
        RECT 793.950 528.600 796.050 529.050 ;
        RECT 829.950 528.600 832.050 529.050 ;
        RECT 793.950 527.400 832.050 528.600 ;
        RECT 793.950 526.950 796.050 527.400 ;
        RECT 829.950 526.950 832.050 527.400 ;
        RECT 574.950 525.600 577.050 526.050 ;
        RECT 587.400 525.600 588.600 526.950 ;
        RECT 604.950 525.600 607.050 526.050 ;
        RECT 574.950 524.400 607.050 525.600 ;
        RECT 574.950 523.950 577.050 524.400 ;
        RECT 604.950 523.950 607.050 524.400 ;
        RECT 616.950 525.600 619.050 526.050 ;
        RECT 625.950 525.600 628.050 526.050 ;
        RECT 640.950 525.600 643.050 526.050 ;
        RECT 616.950 524.400 643.050 525.600 ;
        RECT 616.950 523.950 619.050 524.400 ;
        RECT 625.950 523.950 628.050 524.400 ;
        RECT 640.950 523.950 643.050 524.400 ;
        RECT 646.950 525.600 649.050 526.050 ;
        RECT 658.950 525.600 661.050 526.050 ;
        RECT 646.950 524.400 661.050 525.600 ;
        RECT 646.950 523.950 649.050 524.400 ;
        RECT 658.950 523.950 661.050 524.400 ;
        RECT 664.950 525.600 667.050 526.050 ;
        RECT 670.950 525.600 673.050 526.050 ;
        RECT 664.950 524.400 673.050 525.600 ;
        RECT 664.950 523.950 667.050 524.400 ;
        RECT 670.950 523.950 673.050 524.400 ;
        RECT 673.950 525.600 676.050 526.050 ;
        RECT 679.950 525.600 682.050 526.050 ;
        RECT 673.950 524.400 682.050 525.600 ;
        RECT 673.950 523.950 676.050 524.400 ;
        RECT 679.950 523.950 682.050 524.400 ;
        RECT 736.950 525.600 739.050 526.050 ;
        RECT 745.950 525.600 748.050 526.050 ;
        RECT 736.950 524.400 748.050 525.600 ;
        RECT 736.950 523.950 739.050 524.400 ;
        RECT 745.950 523.950 748.050 524.400 ;
        RECT 751.950 525.600 754.050 526.050 ;
        RECT 775.950 525.600 778.050 526.050 ;
        RECT 751.950 524.400 778.050 525.600 ;
        RECT 751.950 523.950 754.050 524.400 ;
        RECT 775.950 523.950 778.050 524.400 ;
        RECT 826.950 525.600 829.050 526.050 ;
        RECT 832.950 525.600 835.050 526.050 ;
        RECT 826.950 524.400 835.050 525.600 ;
        RECT 826.950 523.950 829.050 524.400 ;
        RECT 832.950 523.950 835.050 524.400 ;
        RECT 847.950 525.600 850.050 526.050 ;
        RECT 859.950 525.600 862.050 526.050 ;
        RECT 847.950 524.400 862.050 525.600 ;
        RECT 847.950 523.950 850.050 524.400 ;
        RECT 859.950 523.950 862.050 524.400 ;
        RECT 484.950 521.400 498.600 522.600 ;
        RECT 499.950 522.600 502.050 523.050 ;
        RECT 505.950 522.600 508.050 523.050 ;
        RECT 517.950 522.600 520.050 523.050 ;
        RECT 499.950 521.400 504.600 522.600 ;
        RECT 484.950 520.950 487.050 521.400 ;
        RECT 499.950 520.950 502.050 521.400 ;
        RECT 19.950 519.600 22.050 520.050 ;
        RECT 25.950 519.600 28.050 520.050 ;
        RECT 19.950 518.400 28.050 519.600 ;
        RECT 19.950 517.950 22.050 518.400 ;
        RECT 25.950 517.950 28.050 518.400 ;
        RECT 118.950 519.600 121.050 520.050 ;
        RECT 133.950 519.600 136.050 520.050 ;
        RECT 118.950 518.400 136.050 519.600 ;
        RECT 118.950 517.950 121.050 518.400 ;
        RECT 133.950 517.950 136.050 518.400 ;
        RECT 163.950 519.600 166.050 520.050 ;
        RECT 193.950 519.600 196.050 520.050 ;
        RECT 163.950 518.400 196.050 519.600 ;
        RECT 163.950 517.950 166.050 518.400 ;
        RECT 193.950 517.950 196.050 518.400 ;
        RECT 211.950 519.600 214.050 520.050 ;
        RECT 215.400 519.600 216.600 520.950 ;
        RECT 503.400 520.050 504.600 521.400 ;
        RECT 505.950 521.400 520.050 522.600 ;
        RECT 505.950 520.950 508.050 521.400 ;
        RECT 517.950 520.950 520.050 521.400 ;
        RECT 523.950 522.600 526.050 523.050 ;
        RECT 523.950 521.400 564.600 522.600 ;
        RECT 523.950 520.950 526.050 521.400 ;
        RECT 211.950 518.400 216.600 519.600 ;
        RECT 244.950 519.600 247.050 520.050 ;
        RECT 262.950 519.600 265.050 520.050 ;
        RECT 244.950 518.400 265.050 519.600 ;
        RECT 211.950 517.950 214.050 518.400 ;
        RECT 244.950 517.950 247.050 518.400 ;
        RECT 262.950 517.950 265.050 518.400 ;
        RECT 289.950 519.600 292.050 520.050 ;
        RECT 352.950 519.600 355.050 520.050 ;
        RECT 289.950 518.400 355.050 519.600 ;
        RECT 289.950 517.950 292.050 518.400 ;
        RECT 352.950 517.950 355.050 518.400 ;
        RECT 451.950 519.600 454.050 520.050 ;
        RECT 457.950 519.600 460.050 520.050 ;
        RECT 451.950 518.400 460.050 519.600 ;
        RECT 451.950 517.950 454.050 518.400 ;
        RECT 457.950 517.950 460.050 518.400 ;
        RECT 466.950 519.600 469.050 520.050 ;
        RECT 487.950 519.600 490.050 520.050 ;
        RECT 499.950 519.600 502.050 520.050 ;
        RECT 466.950 518.400 480.600 519.600 ;
        RECT 466.950 517.950 469.050 518.400 ;
        RECT 13.950 516.600 16.050 517.050 ;
        RECT 16.950 516.600 19.050 517.050 ;
        RECT 13.950 515.400 19.050 516.600 ;
        RECT 13.950 514.950 16.050 515.400 ;
        RECT 16.950 514.950 19.050 515.400 ;
        RECT 121.950 516.600 124.050 517.050 ;
        RECT 130.950 516.600 133.050 517.050 ;
        RECT 142.950 516.600 145.050 517.050 ;
        RECT 121.950 515.400 145.050 516.600 ;
        RECT 121.950 514.950 124.050 515.400 ;
        RECT 130.950 514.950 133.050 515.400 ;
        RECT 142.950 514.950 145.050 515.400 ;
        RECT 193.950 516.600 196.050 517.050 ;
        RECT 205.950 516.600 208.050 517.050 ;
        RECT 193.950 515.400 208.050 516.600 ;
        RECT 193.950 514.950 196.050 515.400 ;
        RECT 205.950 514.950 208.050 515.400 ;
        RECT 304.950 516.600 307.050 517.050 ;
        RECT 340.950 516.600 343.050 517.050 ;
        RECT 479.400 516.600 480.600 518.400 ;
        RECT 487.950 518.400 502.050 519.600 ;
        RECT 487.950 517.950 490.050 518.400 ;
        RECT 499.950 517.950 502.050 518.400 ;
        RECT 502.950 517.950 505.050 520.050 ;
        RECT 511.950 519.600 514.050 520.050 ;
        RECT 550.950 519.600 553.050 520.050 ;
        RECT 511.950 518.400 553.050 519.600 ;
        RECT 563.400 519.600 564.600 521.400 ;
        RECT 565.950 520.950 568.050 523.050 ;
        RECT 595.950 522.600 598.050 523.050 ;
        RECT 625.950 522.600 628.050 523.050 ;
        RECT 595.950 521.400 628.050 522.600 ;
        RECT 595.950 520.950 598.050 521.400 ;
        RECT 625.950 520.950 628.050 521.400 ;
        RECT 568.950 519.600 571.050 520.050 ;
        RECT 563.400 518.400 571.050 519.600 ;
        RECT 511.950 517.950 514.050 518.400 ;
        RECT 550.950 517.950 553.050 518.400 ;
        RECT 568.950 517.950 571.050 518.400 ;
        RECT 610.950 519.600 613.050 520.050 ;
        RECT 655.950 519.600 658.050 520.050 ;
        RECT 610.950 518.400 658.050 519.600 ;
        RECT 610.950 517.950 613.050 518.400 ;
        RECT 655.950 517.950 658.050 518.400 ;
        RECT 676.950 519.600 679.050 520.050 ;
        RECT 691.950 519.600 694.050 520.050 ;
        RECT 676.950 518.400 694.050 519.600 ;
        RECT 676.950 517.950 679.050 518.400 ;
        RECT 691.950 517.950 694.050 518.400 ;
        RECT 724.950 519.600 727.050 520.050 ;
        RECT 757.950 519.600 760.050 520.050 ;
        RECT 724.950 518.400 760.050 519.600 ;
        RECT 724.950 517.950 727.050 518.400 ;
        RECT 757.950 517.950 760.050 518.400 ;
        RECT 838.950 519.600 841.050 520.050 ;
        RECT 856.950 519.600 859.050 520.050 ;
        RECT 838.950 518.400 859.050 519.600 ;
        RECT 838.950 517.950 841.050 518.400 ;
        RECT 856.950 517.950 859.050 518.400 ;
        RECT 511.950 516.600 514.050 517.050 ;
        RECT 523.950 516.600 526.050 517.050 ;
        RECT 304.950 515.400 477.600 516.600 ;
        RECT 479.400 515.400 514.050 516.600 ;
        RECT 304.950 514.950 307.050 515.400 ;
        RECT 340.950 514.950 343.050 515.400 ;
        RECT 476.400 513.600 477.600 515.400 ;
        RECT 511.950 514.950 514.050 515.400 ;
        RECT 515.400 515.400 526.050 516.600 ;
        RECT 515.400 513.600 516.600 515.400 ;
        RECT 523.950 514.950 526.050 515.400 ;
        RECT 721.950 516.600 724.050 517.050 ;
        RECT 814.950 516.600 817.050 517.050 ;
        RECT 721.950 515.400 817.050 516.600 ;
        RECT 721.950 514.950 724.050 515.400 ;
        RECT 814.950 514.950 817.050 515.400 ;
        RECT 476.400 512.400 516.600 513.600 ;
        RECT 517.950 513.600 520.050 514.050 ;
        RECT 553.950 513.600 556.050 514.050 ;
        RECT 517.950 512.400 556.050 513.600 ;
        RECT 517.950 511.950 520.050 512.400 ;
        RECT 553.950 511.950 556.050 512.400 ;
        RECT 652.950 513.600 655.050 514.050 ;
        RECT 724.950 513.600 727.050 514.050 ;
        RECT 652.950 512.400 727.050 513.600 ;
        RECT 652.950 511.950 655.050 512.400 ;
        RECT 724.950 511.950 727.050 512.400 ;
        RECT 220.950 510.600 223.050 511.050 ;
        RECT 316.950 510.600 319.050 511.050 ;
        RECT 220.950 509.400 319.050 510.600 ;
        RECT 220.950 508.950 223.050 509.400 ;
        RECT 316.950 508.950 319.050 509.400 ;
        RECT 463.950 510.600 466.050 511.050 ;
        RECT 472.950 510.600 475.050 511.050 ;
        RECT 463.950 509.400 475.050 510.600 ;
        RECT 463.950 508.950 466.050 509.400 ;
        RECT 472.950 508.950 475.050 509.400 ;
        RECT 553.950 510.600 556.050 511.050 ;
        RECT 574.950 510.600 577.050 511.050 ;
        RECT 553.950 509.400 577.050 510.600 ;
        RECT 553.950 508.950 556.050 509.400 ;
        RECT 574.950 508.950 577.050 509.400 ;
        RECT 298.950 507.600 301.050 508.050 ;
        RECT 427.950 507.600 430.050 508.050 ;
        RECT 298.950 506.400 430.050 507.600 ;
        RECT 298.950 505.950 301.050 506.400 ;
        RECT 427.950 505.950 430.050 506.400 ;
        RECT 532.950 507.600 535.050 508.050 ;
        RECT 586.950 507.600 589.050 508.050 ;
        RECT 532.950 506.400 589.050 507.600 ;
        RECT 532.950 505.950 535.050 506.400 ;
        RECT 586.950 505.950 589.050 506.400 ;
        RECT 598.950 507.600 601.050 508.050 ;
        RECT 688.950 507.600 691.050 508.050 ;
        RECT 598.950 506.400 691.050 507.600 ;
        RECT 598.950 505.950 601.050 506.400 ;
        RECT 688.950 505.950 691.050 506.400 ;
        RECT 814.950 507.600 817.050 508.050 ;
        RECT 820.950 507.600 823.050 508.050 ;
        RECT 814.950 506.400 823.050 507.600 ;
        RECT 814.950 505.950 817.050 506.400 ;
        RECT 820.950 505.950 823.050 506.400 ;
        RECT 397.950 504.600 400.050 505.050 ;
        RECT 502.950 504.600 505.050 505.050 ;
        RECT 397.950 503.400 505.050 504.600 ;
        RECT 397.950 502.950 400.050 503.400 ;
        RECT 502.950 502.950 505.050 503.400 ;
        RECT 511.950 504.600 514.050 505.050 ;
        RECT 601.950 504.600 604.050 505.050 ;
        RECT 511.950 503.400 604.050 504.600 ;
        RECT 511.950 502.950 514.050 503.400 ;
        RECT 601.950 502.950 604.050 503.400 ;
        RECT 412.950 501.600 415.050 502.050 ;
        RECT 418.950 501.600 421.050 502.050 ;
        RECT 466.950 501.600 469.050 502.050 ;
        RECT 412.950 500.400 469.050 501.600 ;
        RECT 412.950 499.950 415.050 500.400 ;
        RECT 418.950 499.950 421.050 500.400 ;
        RECT 466.950 499.950 469.050 500.400 ;
        RECT 469.950 501.600 472.050 502.050 ;
        RECT 478.950 501.600 481.050 502.050 ;
        RECT 469.950 500.400 481.050 501.600 ;
        RECT 469.950 499.950 472.050 500.400 ;
        RECT 478.950 499.950 481.050 500.400 ;
        RECT 484.950 501.600 487.050 502.050 ;
        RECT 493.950 501.600 496.050 502.050 ;
        RECT 622.950 501.600 625.050 502.050 ;
        RECT 484.950 500.400 625.050 501.600 ;
        RECT 484.950 499.950 487.050 500.400 ;
        RECT 493.950 499.950 496.050 500.400 ;
        RECT 622.950 499.950 625.050 500.400 ;
        RECT 160.950 498.600 163.050 499.050 ;
        RECT 184.950 498.600 187.050 499.050 ;
        RECT 160.950 497.400 187.050 498.600 ;
        RECT 160.950 496.950 163.050 497.400 ;
        RECT 184.950 496.950 187.050 497.400 ;
        RECT 391.950 498.600 394.050 499.050 ;
        RECT 412.950 498.600 415.050 499.050 ;
        RECT 391.950 497.400 415.050 498.600 ;
        RECT 391.950 496.950 394.050 497.400 ;
        RECT 412.950 496.950 415.050 497.400 ;
        RECT 454.950 498.600 457.050 499.050 ;
        RECT 472.950 498.600 475.050 499.050 ;
        RECT 454.950 497.400 475.050 498.600 ;
        RECT 454.950 496.950 457.050 497.400 ;
        RECT 472.950 496.950 475.050 497.400 ;
        RECT 496.950 498.600 499.050 499.050 ;
        RECT 535.950 498.600 538.050 499.050 ;
        RECT 496.950 497.400 538.050 498.600 ;
        RECT 496.950 496.950 499.050 497.400 ;
        RECT 535.950 496.950 538.050 497.400 ;
        RECT 619.950 498.600 622.050 499.050 ;
        RECT 631.950 498.600 634.050 499.050 ;
        RECT 619.950 497.400 634.050 498.600 ;
        RECT 619.950 496.950 622.050 497.400 ;
        RECT 631.950 496.950 634.050 497.400 ;
        RECT 52.950 495.600 55.050 496.050 ;
        RECT 61.950 495.600 64.050 496.050 ;
        RECT 52.950 494.400 64.050 495.600 ;
        RECT 52.950 493.950 55.050 494.400 ;
        RECT 61.950 493.950 64.050 494.400 ;
        RECT 97.950 495.600 100.050 496.050 ;
        RECT 100.950 495.600 103.050 496.050 ;
        RECT 124.950 495.600 127.050 496.050 ;
        RECT 202.950 495.600 205.050 496.050 ;
        RECT 97.950 494.400 205.050 495.600 ;
        RECT 97.950 493.950 100.050 494.400 ;
        RECT 100.950 493.950 103.050 494.400 ;
        RECT 124.950 493.950 127.050 494.400 ;
        RECT 202.950 493.950 205.050 494.400 ;
        RECT 265.950 495.600 268.050 496.050 ;
        RECT 289.950 495.600 292.050 496.050 ;
        RECT 265.950 494.400 292.050 495.600 ;
        RECT 265.950 493.950 268.050 494.400 ;
        RECT 289.950 493.950 292.050 494.400 ;
        RECT 310.950 495.600 313.050 496.050 ;
        RECT 346.950 495.600 349.050 496.050 ;
        RECT 361.950 495.600 364.050 496.050 ;
        RECT 310.950 494.400 364.050 495.600 ;
        RECT 310.950 493.950 313.050 494.400 ;
        RECT 346.950 493.950 349.050 494.400 ;
        RECT 361.950 493.950 364.050 494.400 ;
        RECT 400.950 495.600 403.050 496.050 ;
        RECT 430.950 495.600 433.050 496.050 ;
        RECT 400.950 494.400 433.050 495.600 ;
        RECT 400.950 493.950 403.050 494.400 ;
        RECT 430.950 493.950 433.050 494.400 ;
        RECT 436.950 495.600 439.050 496.050 ;
        RECT 436.950 494.400 498.600 495.600 ;
        RECT 436.950 493.950 439.050 494.400 ;
        RECT 37.950 492.600 40.050 493.050 ;
        RECT 46.950 492.600 49.050 493.050 ;
        RECT 58.950 492.600 61.050 493.050 ;
        RECT 37.950 491.400 61.050 492.600 ;
        RECT 37.950 490.950 40.050 491.400 ;
        RECT 46.950 490.950 49.050 491.400 ;
        RECT 58.950 490.950 61.050 491.400 ;
        RECT 175.950 492.600 178.050 493.050 ;
        RECT 187.950 492.600 190.050 493.050 ;
        RECT 223.950 492.600 226.050 493.050 ;
        RECT 175.950 491.400 226.050 492.600 ;
        RECT 175.950 490.950 178.050 491.400 ;
        RECT 187.950 490.950 190.050 491.400 ;
        RECT 223.950 490.950 226.050 491.400 ;
        RECT 232.950 492.600 235.050 493.050 ;
        RECT 259.950 492.600 262.050 493.050 ;
        RECT 232.950 491.400 262.050 492.600 ;
        RECT 232.950 490.950 235.050 491.400 ;
        RECT 248.400 490.050 249.600 491.400 ;
        RECT 259.950 490.950 262.050 491.400 ;
        RECT 271.950 492.600 274.050 493.050 ;
        RECT 301.950 492.600 304.050 493.050 ;
        RECT 271.950 491.400 304.050 492.600 ;
        RECT 271.950 490.950 274.050 491.400 ;
        RECT 301.950 490.950 304.050 491.400 ;
        RECT 328.950 492.600 331.050 493.050 ;
        RECT 337.950 492.600 340.050 493.050 ;
        RECT 328.950 491.400 340.050 492.600 ;
        RECT 328.950 490.950 331.050 491.400 ;
        RECT 337.950 490.950 340.050 491.400 ;
        RECT 385.950 492.600 388.050 493.050 ;
        RECT 397.950 492.600 400.050 493.050 ;
        RECT 385.950 491.400 400.050 492.600 ;
        RECT 385.950 490.950 388.050 491.400 ;
        RECT 397.950 490.950 400.050 491.400 ;
        RECT 415.950 492.600 418.050 493.050 ;
        RECT 460.950 492.600 463.050 493.050 ;
        RECT 493.950 492.600 496.050 493.050 ;
        RECT 415.950 491.400 496.050 492.600 ;
        RECT 497.400 492.600 498.600 494.400 ;
        RECT 517.950 492.600 520.050 493.050 ;
        RECT 541.950 492.600 544.050 493.050 ;
        RECT 497.400 491.400 544.050 492.600 ;
        RECT 415.950 490.950 418.050 491.400 ;
        RECT 460.950 490.950 463.050 491.400 ;
        RECT 493.950 490.950 496.050 491.400 ;
        RECT 517.950 490.950 520.050 491.400 ;
        RECT 541.950 490.950 544.050 491.400 ;
        RECT 826.950 492.600 829.050 493.050 ;
        RECT 832.950 492.600 835.050 493.050 ;
        RECT 826.950 491.400 835.050 492.600 ;
        RECT 826.950 490.950 829.050 491.400 ;
        RECT 832.950 490.950 835.050 491.400 ;
        RECT 10.950 489.600 13.050 490.050 ;
        RECT 40.950 489.600 43.050 490.050 ;
        RECT 10.950 488.400 43.050 489.600 ;
        RECT 10.950 487.950 13.050 488.400 ;
        RECT 40.950 487.950 43.050 488.400 ;
        RECT 46.950 489.600 49.050 490.050 ;
        RECT 82.950 489.600 85.050 490.050 ;
        RECT 46.950 488.400 85.050 489.600 ;
        RECT 46.950 487.950 49.050 488.400 ;
        RECT 82.950 487.950 85.050 488.400 ;
        RECT 103.950 489.600 106.050 490.050 ;
        RECT 130.950 489.600 133.050 490.050 ;
        RECT 136.950 489.600 139.050 490.050 ;
        RECT 142.950 489.600 145.050 490.050 ;
        RECT 103.950 488.400 145.050 489.600 ;
        RECT 103.950 487.950 106.050 488.400 ;
        RECT 130.950 487.950 133.050 488.400 ;
        RECT 136.950 487.950 139.050 488.400 ;
        RECT 142.950 487.950 145.050 488.400 ;
        RECT 148.950 489.600 151.050 490.050 ;
        RECT 163.950 489.600 166.050 490.050 ;
        RECT 148.950 488.400 166.050 489.600 ;
        RECT 148.950 487.950 151.050 488.400 ;
        RECT 163.950 487.950 166.050 488.400 ;
        RECT 181.950 489.600 184.050 490.050 ;
        RECT 220.950 489.600 223.050 490.050 ;
        RECT 181.950 488.400 223.050 489.600 ;
        RECT 181.950 487.950 184.050 488.400 ;
        RECT 220.950 487.950 223.050 488.400 ;
        RECT 235.950 489.600 238.050 490.050 ;
        RECT 241.950 489.600 244.050 490.050 ;
        RECT 235.950 488.400 244.050 489.600 ;
        RECT 235.950 487.950 238.050 488.400 ;
        RECT 241.950 487.950 244.050 488.400 ;
        RECT 247.950 487.950 250.050 490.050 ;
        RECT 286.950 489.600 289.050 490.050 ;
        RECT 319.950 489.600 322.050 490.050 ;
        RECT 286.950 488.400 322.050 489.600 ;
        RECT 286.950 487.950 289.050 488.400 ;
        RECT 319.950 487.950 322.050 488.400 ;
        RECT 328.950 489.600 331.050 490.050 ;
        RECT 334.950 489.600 337.050 490.050 ;
        RECT 328.950 488.400 337.050 489.600 ;
        RECT 328.950 487.950 331.050 488.400 ;
        RECT 334.950 487.950 337.050 488.400 ;
        RECT 370.950 489.600 373.050 490.050 ;
        RECT 406.950 489.600 409.050 490.050 ;
        RECT 439.950 489.600 442.050 490.050 ;
        RECT 472.950 489.600 475.050 490.050 ;
        RECT 484.950 489.600 487.050 490.050 ;
        RECT 370.950 488.400 409.050 489.600 ;
        RECT 370.950 487.950 373.050 488.400 ;
        RECT 406.950 487.950 409.050 488.400 ;
        RECT 422.400 488.400 442.050 489.600 ;
        RECT 422.400 487.050 423.600 488.400 ;
        RECT 439.950 487.950 442.050 488.400 ;
        RECT 446.400 488.400 487.050 489.600 ;
        RECT 13.950 486.600 16.050 487.050 ;
        RECT 25.950 486.600 28.050 487.050 ;
        RECT 13.950 485.400 28.050 486.600 ;
        RECT 13.950 484.950 16.050 485.400 ;
        RECT 25.950 484.950 28.050 485.400 ;
        RECT 31.950 486.600 34.050 487.050 ;
        RECT 46.950 486.600 49.050 487.050 ;
        RECT 31.950 485.400 49.050 486.600 ;
        RECT 31.950 484.950 34.050 485.400 ;
        RECT 46.950 484.950 49.050 485.400 ;
        RECT 61.950 486.600 64.050 487.050 ;
        RECT 76.950 486.600 79.050 487.050 ;
        RECT 61.950 485.400 79.050 486.600 ;
        RECT 61.950 484.950 64.050 485.400 ;
        RECT 76.950 484.950 79.050 485.400 ;
        RECT 166.950 486.600 169.050 487.050 ;
        RECT 181.950 486.600 184.050 487.050 ;
        RECT 166.950 485.400 184.050 486.600 ;
        RECT 166.950 484.950 169.050 485.400 ;
        RECT 181.950 484.950 184.050 485.400 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 187.950 486.600 190.050 487.050 ;
        RECT 205.950 486.600 208.050 487.050 ;
        RECT 187.950 485.400 208.050 486.600 ;
        RECT 187.950 484.950 190.050 485.400 ;
        RECT 205.950 484.950 208.050 485.400 ;
        RECT 214.950 486.600 217.050 487.050 ;
        RECT 238.950 486.600 241.050 487.050 ;
        RECT 214.950 485.400 241.050 486.600 ;
        RECT 214.950 484.950 217.050 485.400 ;
        RECT 238.950 484.950 241.050 485.400 ;
        RECT 244.950 486.600 247.050 487.050 ;
        RECT 256.950 486.600 259.050 487.050 ;
        RECT 244.950 485.400 259.050 486.600 ;
        RECT 244.950 484.950 247.050 485.400 ;
        RECT 256.950 484.950 259.050 485.400 ;
        RECT 268.950 486.600 271.050 487.050 ;
        RECT 313.950 486.600 316.050 487.050 ;
        RECT 325.950 486.600 328.050 487.050 ;
        RECT 268.950 485.400 312.600 486.600 ;
        RECT 268.950 484.950 271.050 485.400 ;
        RECT 19.950 483.600 22.050 484.050 ;
        RECT 25.950 483.600 28.050 484.050 ;
        RECT 19.950 482.400 28.050 483.600 ;
        RECT 19.950 481.950 22.050 482.400 ;
        RECT 25.950 481.950 28.050 482.400 ;
        RECT 34.950 483.600 37.050 484.050 ;
        RECT 40.950 483.600 43.050 484.050 ;
        RECT 34.950 482.400 43.050 483.600 ;
        RECT 34.950 481.950 37.050 482.400 ;
        RECT 40.950 481.950 43.050 482.400 ;
        RECT 58.950 483.600 61.050 484.050 ;
        RECT 67.950 483.600 70.050 484.050 ;
        RECT 58.950 482.400 70.050 483.600 ;
        RECT 58.950 481.950 61.050 482.400 ;
        RECT 67.950 481.950 70.050 482.400 ;
        RECT 106.950 483.600 109.050 484.050 ;
        RECT 112.950 483.600 115.050 484.050 ;
        RECT 136.950 483.600 139.050 484.050 ;
        RECT 106.950 482.400 139.050 483.600 ;
        RECT 106.950 481.950 109.050 482.400 ;
        RECT 112.950 481.950 115.050 482.400 ;
        RECT 136.950 481.950 139.050 482.400 ;
        RECT 175.950 483.600 178.050 484.050 ;
        RECT 185.400 483.600 186.600 484.950 ;
        RECT 175.950 482.400 186.600 483.600 ;
        RECT 226.950 483.600 229.050 484.050 ;
        RECT 250.950 483.600 253.050 484.050 ;
        RECT 226.950 482.400 253.050 483.600 ;
        RECT 311.400 483.600 312.600 485.400 ;
        RECT 313.950 485.400 328.050 486.600 ;
        RECT 313.950 484.950 316.050 485.400 ;
        RECT 325.950 484.950 328.050 485.400 ;
        RECT 388.950 484.950 391.050 487.050 ;
        RECT 412.950 486.600 415.050 487.050 ;
        RECT 418.950 486.600 421.050 487.050 ;
        RECT 412.950 485.400 421.050 486.600 ;
        RECT 412.950 484.950 415.050 485.400 ;
        RECT 418.950 484.950 421.050 485.400 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 424.950 486.600 427.050 487.050 ;
        RECT 436.950 486.600 439.050 487.050 ;
        RECT 424.950 485.400 439.050 486.600 ;
        RECT 424.950 484.950 427.050 485.400 ;
        RECT 436.950 484.950 439.050 485.400 ;
        RECT 328.950 483.600 331.050 484.050 ;
        RECT 311.400 482.400 331.050 483.600 ;
        RECT 175.950 481.950 178.050 482.400 ;
        RECT 226.950 481.950 229.050 482.400 ;
        RECT 250.950 481.950 253.050 482.400 ;
        RECT 328.950 481.950 331.050 482.400 ;
        RECT 334.950 483.600 337.050 484.050 ;
        RECT 343.950 483.600 346.050 484.050 ;
        RECT 334.950 482.400 346.050 483.600 ;
        RECT 334.950 481.950 337.050 482.400 ;
        RECT 343.950 481.950 346.050 482.400 ;
        RECT 358.950 483.600 361.050 484.050 ;
        RECT 385.950 483.600 388.050 484.050 ;
        RECT 358.950 482.400 388.050 483.600 ;
        RECT 389.400 483.600 390.600 484.950 ;
        RECT 403.950 483.600 406.050 484.050 ;
        RECT 389.400 482.400 406.050 483.600 ;
        RECT 358.950 481.950 361.050 482.400 ;
        RECT 385.950 481.950 388.050 482.400 ;
        RECT 403.950 481.950 406.050 482.400 ;
        RECT 13.950 480.600 16.050 481.050 ;
        RECT 37.950 480.600 40.050 481.050 ;
        RECT 13.950 479.400 40.050 480.600 ;
        RECT 13.950 478.950 16.050 479.400 ;
        RECT 37.950 478.950 40.050 479.400 ;
        RECT 130.950 480.600 133.050 481.050 ;
        RECT 145.950 480.600 148.050 481.050 ;
        RECT 130.950 479.400 148.050 480.600 ;
        RECT 130.950 478.950 133.050 479.400 ;
        RECT 145.950 478.950 148.050 479.400 ;
        RECT 223.950 480.600 226.050 481.050 ;
        RECT 232.950 480.600 235.050 481.050 ;
        RECT 223.950 479.400 235.050 480.600 ;
        RECT 223.950 478.950 226.050 479.400 ;
        RECT 232.950 478.950 235.050 479.400 ;
        RECT 268.950 480.600 271.050 481.050 ;
        RECT 283.950 480.600 286.050 481.050 ;
        RECT 289.950 480.600 292.050 481.050 ;
        RECT 268.950 479.400 292.050 480.600 ;
        RECT 268.950 478.950 271.050 479.400 ;
        RECT 283.950 478.950 286.050 479.400 ;
        RECT 289.950 478.950 292.050 479.400 ;
        RECT 331.950 480.600 334.050 481.050 ;
        RECT 355.950 480.600 358.050 481.050 ;
        RECT 331.950 479.400 358.050 480.600 ;
        RECT 331.950 478.950 334.050 479.400 ;
        RECT 355.950 478.950 358.050 479.400 ;
        RECT 397.950 480.600 400.050 481.050 ;
        RECT 409.950 480.600 412.050 481.050 ;
        RECT 397.950 479.400 412.050 480.600 ;
        RECT 397.950 478.950 400.050 479.400 ;
        RECT 409.950 478.950 412.050 479.400 ;
        RECT 427.950 480.600 430.050 481.050 ;
        RECT 446.400 480.600 447.600 488.400 ;
        RECT 472.950 487.950 475.050 488.400 ;
        RECT 484.950 487.950 487.050 488.400 ;
        RECT 508.950 489.600 511.050 490.050 ;
        RECT 520.950 489.600 523.050 490.050 ;
        RECT 508.950 488.400 523.050 489.600 ;
        RECT 508.950 487.950 511.050 488.400 ;
        RECT 520.950 487.950 523.050 488.400 ;
        RECT 550.950 489.600 553.050 490.050 ;
        RECT 592.950 489.600 595.050 490.050 ;
        RECT 550.950 488.400 595.050 489.600 ;
        RECT 550.950 487.950 553.050 488.400 ;
        RECT 592.950 487.950 595.050 488.400 ;
        RECT 601.950 489.600 604.050 490.050 ;
        RECT 634.950 489.600 637.050 490.050 ;
        RECT 601.950 488.400 637.050 489.600 ;
        RECT 601.950 487.950 604.050 488.400 ;
        RECT 634.950 487.950 637.050 488.400 ;
        RECT 643.950 489.600 646.050 490.050 ;
        RECT 643.950 488.400 672.600 489.600 ;
        RECT 643.950 487.950 646.050 488.400 ;
        RECT 505.950 486.600 508.050 487.050 ;
        RECT 529.950 486.600 532.050 487.050 ;
        RECT 538.950 486.600 541.050 487.050 ;
        RECT 505.950 485.400 541.050 486.600 ;
        RECT 505.950 484.950 508.050 485.400 ;
        RECT 529.950 484.950 532.050 485.400 ;
        RECT 538.950 484.950 541.050 485.400 ;
        RECT 544.950 484.950 547.050 487.050 ;
        RECT 574.950 486.600 577.050 487.050 ;
        RECT 583.950 486.600 586.050 487.050 ;
        RECT 574.950 485.400 586.050 486.600 ;
        RECT 574.950 484.950 577.050 485.400 ;
        RECT 583.950 484.950 586.050 485.400 ;
        RECT 592.950 486.600 595.050 487.050 ;
        RECT 613.950 486.600 616.050 487.050 ;
        RECT 592.950 485.400 616.050 486.600 ;
        RECT 592.950 484.950 595.050 485.400 ;
        RECT 613.950 484.950 616.050 485.400 ;
        RECT 628.950 486.600 631.050 487.050 ;
        RECT 634.950 486.600 637.050 487.050 ;
        RECT 628.950 485.400 637.050 486.600 ;
        RECT 628.950 484.950 631.050 485.400 ;
        RECT 634.950 484.950 637.050 485.400 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 661.950 486.600 664.050 487.050 ;
        RECT 667.950 486.600 670.050 487.050 ;
        RECT 661.950 485.400 670.050 486.600 ;
        RECT 671.400 486.600 672.600 488.400 ;
        RECT 736.950 486.600 739.050 487.050 ;
        RECT 671.400 485.400 739.050 486.600 ;
        RECT 661.950 484.950 664.050 485.400 ;
        RECT 667.950 484.950 670.050 485.400 ;
        RECT 736.950 484.950 739.050 485.400 ;
        RECT 757.950 486.600 760.050 487.050 ;
        RECT 772.950 486.600 775.050 487.050 ;
        RECT 757.950 485.400 775.050 486.600 ;
        RECT 757.950 484.950 760.050 485.400 ;
        RECT 772.950 484.950 775.050 485.400 ;
        RECT 805.950 486.600 808.050 487.050 ;
        RECT 823.950 486.600 826.050 487.050 ;
        RECT 805.950 485.400 826.050 486.600 ;
        RECT 805.950 484.950 808.050 485.400 ;
        RECT 823.950 484.950 826.050 485.400 ;
        RECT 451.950 483.600 454.050 484.050 ;
        RECT 457.950 483.600 460.050 484.050 ;
        RECT 451.950 482.400 460.050 483.600 ;
        RECT 451.950 481.950 454.050 482.400 ;
        RECT 457.950 481.950 460.050 482.400 ;
        RECT 499.950 483.600 502.050 484.050 ;
        RECT 529.950 483.600 532.050 484.050 ;
        RECT 499.950 482.400 532.050 483.600 ;
        RECT 499.950 481.950 502.050 482.400 ;
        RECT 529.950 481.950 532.050 482.400 ;
        RECT 427.950 479.400 447.600 480.600 ;
        RECT 454.950 480.600 457.050 481.050 ;
        RECT 502.950 480.600 505.050 481.050 ;
        RECT 532.950 480.600 535.050 481.050 ;
        RECT 454.950 479.400 535.050 480.600 ;
        RECT 545.400 480.600 546.600 484.950 ;
        RECT 547.950 483.600 550.050 484.050 ;
        RECT 553.950 483.600 556.050 484.050 ;
        RECT 547.950 482.400 556.050 483.600 ;
        RECT 547.950 481.950 550.050 482.400 ;
        RECT 553.950 481.950 556.050 482.400 ;
        RECT 574.950 483.600 577.050 484.050 ;
        RECT 656.400 483.600 657.600 484.950 ;
        RECT 574.950 482.400 657.600 483.600 ;
        RECT 688.950 483.600 691.050 484.050 ;
        RECT 715.950 483.600 718.050 484.050 ;
        RECT 688.950 482.400 718.050 483.600 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 688.950 481.950 691.050 482.400 ;
        RECT 715.950 481.950 718.050 482.400 ;
        RECT 718.950 483.600 721.050 484.050 ;
        RECT 730.950 483.600 733.050 484.050 ;
        RECT 739.950 483.600 742.050 484.050 ;
        RECT 718.950 482.400 723.600 483.600 ;
        RECT 718.950 481.950 721.050 482.400 ;
        RECT 553.950 480.600 556.050 481.050 ;
        RECT 545.400 479.400 556.050 480.600 ;
        RECT 427.950 478.950 430.050 479.400 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 502.950 478.950 505.050 479.400 ;
        RECT 532.950 478.950 535.050 479.400 ;
        RECT 553.950 478.950 556.050 479.400 ;
        RECT 580.950 480.600 583.050 481.050 ;
        RECT 586.950 480.600 589.050 481.050 ;
        RECT 580.950 479.400 589.050 480.600 ;
        RECT 580.950 478.950 583.050 479.400 ;
        RECT 586.950 478.950 589.050 479.400 ;
        RECT 697.950 480.600 700.050 481.050 ;
        RECT 718.950 480.600 721.050 481.050 ;
        RECT 697.950 479.400 721.050 480.600 ;
        RECT 722.400 480.600 723.600 482.400 ;
        RECT 730.950 482.400 742.050 483.600 ;
        RECT 730.950 481.950 733.050 482.400 ;
        RECT 739.950 481.950 742.050 482.400 ;
        RECT 790.950 480.600 793.050 481.050 ;
        RECT 722.400 479.400 793.050 480.600 ;
        RECT 697.950 478.950 700.050 479.400 ;
        RECT 718.950 478.950 721.050 479.400 ;
        RECT 790.950 478.950 793.050 479.400 ;
        RECT 10.950 477.600 13.050 478.050 ;
        RECT 16.950 477.600 19.050 478.050 ;
        RECT 10.950 476.400 19.050 477.600 ;
        RECT 10.950 475.950 13.050 476.400 ;
        RECT 16.950 475.950 19.050 476.400 ;
        RECT 94.950 477.600 97.050 478.050 ;
        RECT 145.950 477.600 148.050 478.050 ;
        RECT 94.950 476.400 148.050 477.600 ;
        RECT 94.950 475.950 97.050 476.400 ;
        RECT 145.950 475.950 148.050 476.400 ;
        RECT 169.950 477.600 172.050 478.050 ;
        RECT 184.950 477.600 187.050 478.050 ;
        RECT 268.950 477.600 271.050 478.050 ;
        RECT 169.950 476.400 271.050 477.600 ;
        RECT 169.950 475.950 172.050 476.400 ;
        RECT 184.950 475.950 187.050 476.400 ;
        RECT 268.950 475.950 271.050 476.400 ;
        RECT 382.950 477.600 385.050 478.050 ;
        RECT 397.950 477.600 400.050 478.050 ;
        RECT 382.950 476.400 400.050 477.600 ;
        RECT 382.950 475.950 385.050 476.400 ;
        RECT 397.950 475.950 400.050 476.400 ;
        RECT 436.950 477.600 439.050 478.050 ;
        RECT 463.950 477.600 466.050 478.050 ;
        RECT 436.950 476.400 466.050 477.600 ;
        RECT 436.950 475.950 439.050 476.400 ;
        RECT 463.950 475.950 466.050 476.400 ;
        RECT 514.950 477.600 517.050 478.050 ;
        RECT 586.950 477.600 589.050 478.050 ;
        RECT 514.950 476.400 589.050 477.600 ;
        RECT 514.950 475.950 517.050 476.400 ;
        RECT 586.950 475.950 589.050 476.400 ;
        RECT 610.950 477.600 613.050 478.050 ;
        RECT 637.950 477.600 640.050 478.050 ;
        RECT 610.950 476.400 640.050 477.600 ;
        RECT 610.950 475.950 613.050 476.400 ;
        RECT 637.950 475.950 640.050 476.400 ;
        RECT 649.950 477.600 652.050 478.050 ;
        RECT 655.950 477.600 658.050 478.050 ;
        RECT 649.950 476.400 658.050 477.600 ;
        RECT 649.950 475.950 652.050 476.400 ;
        RECT 655.950 475.950 658.050 476.400 ;
        RECT 661.950 477.600 664.050 478.050 ;
        RECT 682.950 477.600 685.050 478.050 ;
        RECT 700.950 477.600 703.050 478.050 ;
        RECT 661.950 476.400 703.050 477.600 ;
        RECT 661.950 475.950 664.050 476.400 ;
        RECT 682.950 475.950 685.050 476.400 ;
        RECT 700.950 475.950 703.050 476.400 ;
        RECT 127.950 474.600 130.050 475.050 ;
        RECT 139.950 474.600 142.050 475.050 ;
        RECT 148.950 474.600 151.050 475.050 ;
        RECT 181.950 474.600 184.050 475.050 ;
        RECT 127.950 473.400 184.050 474.600 ;
        RECT 127.950 472.950 130.050 473.400 ;
        RECT 139.950 472.950 142.050 473.400 ;
        RECT 148.950 472.950 151.050 473.400 ;
        RECT 181.950 472.950 184.050 473.400 ;
        RECT 262.950 474.600 265.050 475.050 ;
        RECT 283.950 474.600 286.050 475.050 ;
        RECT 262.950 473.400 286.050 474.600 ;
        RECT 262.950 472.950 265.050 473.400 ;
        RECT 283.950 472.950 286.050 473.400 ;
        RECT 346.950 474.600 349.050 475.050 ;
        RECT 391.950 474.600 394.050 475.050 ;
        RECT 463.950 474.600 466.050 475.050 ;
        RECT 346.950 473.400 466.050 474.600 ;
        RECT 346.950 472.950 349.050 473.400 ;
        RECT 391.950 472.950 394.050 473.400 ;
        RECT 463.950 472.950 466.050 473.400 ;
        RECT 469.950 474.600 472.050 475.050 ;
        RECT 478.950 474.600 481.050 475.050 ;
        RECT 502.950 474.600 505.050 475.050 ;
        RECT 469.950 473.400 505.050 474.600 ;
        RECT 469.950 472.950 472.050 473.400 ;
        RECT 478.950 472.950 481.050 473.400 ;
        RECT 502.950 472.950 505.050 473.400 ;
        RECT 526.950 474.600 529.050 475.050 ;
        RECT 541.950 474.600 544.050 475.050 ;
        RECT 565.950 474.600 568.050 475.050 ;
        RECT 526.950 473.400 568.050 474.600 ;
        RECT 526.950 472.950 529.050 473.400 ;
        RECT 541.950 472.950 544.050 473.400 ;
        RECT 565.950 472.950 568.050 473.400 ;
        RECT 568.950 474.600 571.050 475.050 ;
        RECT 598.950 474.600 601.050 475.050 ;
        RECT 568.950 473.400 601.050 474.600 ;
        RECT 568.950 472.950 571.050 473.400 ;
        RECT 598.950 472.950 601.050 473.400 ;
        RECT 604.950 474.600 607.050 475.050 ;
        RECT 661.950 474.600 664.050 475.050 ;
        RECT 604.950 473.400 664.050 474.600 ;
        RECT 604.950 472.950 607.050 473.400 ;
        RECT 661.950 472.950 664.050 473.400 ;
        RECT 175.950 471.600 178.050 472.050 ;
        RECT 184.950 471.600 187.050 472.050 ;
        RECT 175.950 470.400 187.050 471.600 ;
        RECT 175.950 469.950 178.050 470.400 ;
        RECT 184.950 469.950 187.050 470.400 ;
        RECT 199.950 471.600 202.050 472.050 ;
        RECT 241.950 471.600 244.050 472.050 ;
        RECT 199.950 470.400 244.050 471.600 ;
        RECT 199.950 469.950 202.050 470.400 ;
        RECT 241.950 469.950 244.050 470.400 ;
        RECT 274.950 471.600 277.050 472.050 ;
        RECT 304.950 471.600 307.050 472.050 ;
        RECT 274.950 470.400 307.050 471.600 ;
        RECT 274.950 469.950 277.050 470.400 ;
        RECT 304.950 469.950 307.050 470.400 ;
        RECT 349.950 471.600 352.050 472.050 ;
        RECT 388.950 471.600 391.050 472.050 ;
        RECT 427.950 471.600 430.050 472.050 ;
        RECT 349.950 470.400 430.050 471.600 ;
        RECT 349.950 469.950 352.050 470.400 ;
        RECT 388.950 469.950 391.050 470.400 ;
        RECT 427.950 469.950 430.050 470.400 ;
        RECT 490.950 471.600 493.050 472.050 ;
        RECT 520.950 471.600 523.050 472.050 ;
        RECT 490.950 470.400 523.050 471.600 ;
        RECT 490.950 469.950 493.050 470.400 ;
        RECT 520.950 469.950 523.050 470.400 ;
        RECT 589.950 471.600 592.050 472.050 ;
        RECT 595.950 471.600 598.050 472.050 ;
        RECT 589.950 470.400 598.050 471.600 ;
        RECT 589.950 469.950 592.050 470.400 ;
        RECT 595.950 469.950 598.050 470.400 ;
        RECT 640.950 471.600 643.050 472.050 ;
        RECT 784.950 471.600 787.050 472.050 ;
        RECT 640.950 470.400 787.050 471.600 ;
        RECT 640.950 469.950 643.050 470.400 ;
        RECT 784.950 469.950 787.050 470.400 ;
        RECT 85.950 468.600 88.050 469.050 ;
        RECT 169.950 468.600 172.050 469.050 ;
        RECT 193.950 468.600 196.050 469.050 ;
        RECT 85.950 467.400 168.600 468.600 ;
        RECT 85.950 466.950 88.050 467.400 ;
        RECT 127.950 465.600 130.050 466.050 ;
        RECT 160.950 465.600 163.050 466.050 ;
        RECT 127.950 464.400 163.050 465.600 ;
        RECT 167.400 465.600 168.600 467.400 ;
        RECT 169.950 467.400 196.050 468.600 ;
        RECT 169.950 466.950 172.050 467.400 ;
        RECT 193.950 466.950 196.050 467.400 ;
        RECT 208.950 468.600 211.050 469.050 ;
        RECT 229.950 468.600 232.050 469.050 ;
        RECT 208.950 467.400 232.050 468.600 ;
        RECT 208.950 466.950 211.050 467.400 ;
        RECT 229.950 466.950 232.050 467.400 ;
        RECT 325.950 468.600 328.050 469.050 ;
        RECT 337.950 468.600 340.050 469.050 ;
        RECT 325.950 467.400 340.050 468.600 ;
        RECT 325.950 466.950 328.050 467.400 ;
        RECT 337.950 466.950 340.050 467.400 ;
        RECT 352.950 468.600 355.050 469.050 ;
        RECT 364.950 468.600 367.050 469.050 ;
        RECT 352.950 467.400 367.050 468.600 ;
        RECT 352.950 466.950 355.050 467.400 ;
        RECT 364.950 466.950 367.050 467.400 ;
        RECT 376.950 468.600 379.050 469.050 ;
        RECT 385.950 468.600 388.050 469.050 ;
        RECT 376.950 467.400 388.050 468.600 ;
        RECT 376.950 466.950 379.050 467.400 ;
        RECT 385.950 466.950 388.050 467.400 ;
        RECT 403.950 468.600 406.050 469.050 ;
        RECT 412.950 468.600 415.050 469.050 ;
        RECT 403.950 467.400 415.050 468.600 ;
        RECT 403.950 466.950 406.050 467.400 ;
        RECT 412.950 466.950 415.050 467.400 ;
        RECT 454.950 468.600 457.050 469.050 ;
        RECT 481.950 468.600 484.050 469.050 ;
        RECT 454.950 467.400 484.050 468.600 ;
        RECT 454.950 466.950 457.050 467.400 ;
        RECT 481.950 466.950 484.050 467.400 ;
        RECT 499.950 468.600 502.050 469.050 ;
        RECT 514.950 468.600 517.050 469.050 ;
        RECT 499.950 467.400 517.050 468.600 ;
        RECT 499.950 466.950 502.050 467.400 ;
        RECT 514.950 466.950 517.050 467.400 ;
        RECT 553.950 468.600 556.050 469.050 ;
        RECT 610.950 468.600 613.050 469.050 ;
        RECT 553.950 467.400 613.050 468.600 ;
        RECT 553.950 466.950 556.050 467.400 ;
        RECT 610.950 466.950 613.050 467.400 ;
        RECT 625.950 468.600 628.050 469.050 ;
        RECT 637.950 468.600 640.050 469.050 ;
        RECT 667.950 468.600 670.050 469.050 ;
        RECT 625.950 467.400 670.050 468.600 ;
        RECT 625.950 466.950 628.050 467.400 ;
        RECT 637.950 466.950 640.050 467.400 ;
        RECT 667.950 466.950 670.050 467.400 ;
        RECT 238.950 465.600 241.050 466.050 ;
        RECT 167.400 464.400 241.050 465.600 ;
        RECT 127.950 463.950 130.050 464.400 ;
        RECT 160.950 463.950 163.050 464.400 ;
        RECT 238.950 463.950 241.050 464.400 ;
        RECT 319.950 465.600 322.050 466.050 ;
        RECT 376.950 465.600 379.050 466.050 ;
        RECT 319.950 464.400 379.050 465.600 ;
        RECT 319.950 463.950 322.050 464.400 ;
        RECT 376.950 463.950 379.050 464.400 ;
        RECT 394.950 465.600 397.050 466.050 ;
        RECT 628.950 465.600 631.050 466.050 ;
        RECT 649.950 465.600 652.050 466.050 ;
        RECT 394.950 464.400 652.050 465.600 ;
        RECT 394.950 463.950 397.050 464.400 ;
        RECT 628.950 463.950 631.050 464.400 ;
        RECT 649.950 463.950 652.050 464.400 ;
        RECT 58.950 462.600 61.050 463.050 ;
        RECT 151.950 462.600 154.050 463.050 ;
        RECT 172.950 462.600 175.050 463.050 ;
        RECT 58.950 461.400 99.600 462.600 ;
        RECT 58.950 460.950 61.050 461.400 ;
        RECT 52.950 459.600 55.050 460.050 ;
        RECT 85.950 459.600 88.050 460.050 ;
        RECT 94.950 459.600 97.050 460.050 ;
        RECT 52.950 458.400 97.050 459.600 ;
        RECT 52.950 457.950 55.050 458.400 ;
        RECT 85.950 457.950 88.050 458.400 ;
        RECT 94.950 457.950 97.050 458.400 ;
        RECT 22.950 456.600 25.050 457.050 ;
        RECT 37.950 456.600 40.050 457.050 ;
        RECT 22.950 455.400 40.050 456.600 ;
        RECT 22.950 454.950 25.050 455.400 ;
        RECT 37.950 454.950 40.050 455.400 ;
        RECT 43.950 456.600 46.050 457.050 ;
        RECT 70.950 456.600 73.050 457.050 ;
        RECT 43.950 455.400 73.050 456.600 ;
        RECT 43.950 454.950 46.050 455.400 ;
        RECT 70.950 454.950 73.050 455.400 ;
        RECT 79.950 456.600 82.050 457.050 ;
        RECT 91.950 456.600 94.050 457.050 ;
        RECT 79.950 455.400 94.050 456.600 ;
        RECT 79.950 454.950 82.050 455.400 ;
        RECT 91.950 454.950 94.050 455.400 ;
        RECT 98.400 454.050 99.600 461.400 ;
        RECT 151.950 461.400 175.050 462.600 ;
        RECT 151.950 460.950 154.050 461.400 ;
        RECT 172.950 460.950 175.050 461.400 ;
        RECT 223.950 462.600 226.050 463.050 ;
        RECT 259.950 462.600 262.050 463.050 ;
        RECT 289.950 462.600 292.050 463.050 ;
        RECT 223.950 461.400 292.050 462.600 ;
        RECT 223.950 460.950 226.050 461.400 ;
        RECT 259.950 460.950 262.050 461.400 ;
        RECT 289.950 460.950 292.050 461.400 ;
        RECT 304.950 462.600 307.050 463.050 ;
        RECT 316.950 462.600 319.050 463.050 ;
        RECT 394.950 462.600 397.050 463.050 ;
        RECT 304.950 461.400 397.050 462.600 ;
        RECT 304.950 460.950 307.050 461.400 ;
        RECT 316.950 460.950 319.050 461.400 ;
        RECT 394.950 460.950 397.050 461.400 ;
        RECT 400.950 462.600 403.050 463.050 ;
        RECT 415.950 462.600 418.050 463.050 ;
        RECT 430.950 462.600 433.050 463.050 ;
        RECT 439.950 462.600 442.050 463.050 ;
        RECT 400.950 461.400 442.050 462.600 ;
        RECT 400.950 460.950 403.050 461.400 ;
        RECT 415.950 460.950 418.050 461.400 ;
        RECT 430.950 460.950 433.050 461.400 ;
        RECT 439.950 460.950 442.050 461.400 ;
        RECT 472.950 462.600 475.050 463.050 ;
        RECT 490.950 462.600 493.050 463.050 ;
        RECT 508.950 462.600 511.050 463.050 ;
        RECT 472.950 461.400 511.050 462.600 ;
        RECT 472.950 460.950 475.050 461.400 ;
        RECT 490.950 460.950 493.050 461.400 ;
        RECT 508.950 460.950 511.050 461.400 ;
        RECT 580.950 462.600 583.050 463.050 ;
        RECT 631.950 462.600 634.050 463.050 ;
        RECT 580.950 461.400 634.050 462.600 ;
        RECT 580.950 460.950 583.050 461.400 ;
        RECT 631.950 460.950 634.050 461.400 ;
        RECT 100.950 459.600 103.050 460.050 ;
        RECT 175.950 459.600 178.050 460.050 ;
        RECT 100.950 458.400 178.050 459.600 ;
        RECT 100.950 457.950 103.050 458.400 ;
        RECT 175.950 457.950 178.050 458.400 ;
        RECT 190.950 459.600 193.050 460.050 ;
        RECT 196.950 459.600 199.050 460.050 ;
        RECT 190.950 458.400 199.050 459.600 ;
        RECT 190.950 457.950 193.050 458.400 ;
        RECT 196.950 457.950 199.050 458.400 ;
        RECT 226.950 459.600 229.050 460.050 ;
        RECT 235.950 459.600 238.050 460.050 ;
        RECT 250.950 459.600 253.050 460.050 ;
        RECT 226.950 458.400 253.050 459.600 ;
        RECT 226.950 457.950 229.050 458.400 ;
        RECT 235.950 457.950 238.050 458.400 ;
        RECT 250.950 457.950 253.050 458.400 ;
        RECT 295.950 459.600 298.050 460.050 ;
        RECT 310.950 459.600 313.050 460.050 ;
        RECT 352.950 459.600 355.050 460.050 ;
        RECT 295.950 458.400 355.050 459.600 ;
        RECT 295.950 457.950 298.050 458.400 ;
        RECT 310.950 457.950 313.050 458.400 ;
        RECT 352.950 457.950 355.050 458.400 ;
        RECT 361.950 457.950 364.050 460.050 ;
        RECT 370.950 459.600 373.050 460.050 ;
        RECT 382.950 459.600 385.050 460.050 ;
        RECT 370.950 458.400 385.050 459.600 ;
        RECT 370.950 457.950 373.050 458.400 ;
        RECT 382.950 457.950 385.050 458.400 ;
        RECT 385.950 459.600 388.050 460.050 ;
        RECT 442.950 459.600 445.050 460.050 ;
        RECT 385.950 458.400 445.050 459.600 ;
        RECT 385.950 457.950 388.050 458.400 ;
        RECT 115.950 456.600 118.050 457.050 ;
        RECT 107.400 455.400 118.050 456.600 ;
        RECT 46.950 453.600 49.050 454.050 ;
        RECT 76.950 453.600 79.050 454.050 ;
        RECT 46.950 452.400 79.050 453.600 ;
        RECT 46.950 451.950 49.050 452.400 ;
        RECT 76.950 451.950 79.050 452.400 ;
        RECT 82.950 453.600 85.050 454.050 ;
        RECT 97.950 453.600 100.050 454.050 ;
        RECT 82.950 452.400 100.050 453.600 ;
        RECT 82.950 451.950 85.050 452.400 ;
        RECT 97.950 451.950 100.050 452.400 ;
        RECT 16.950 450.600 19.050 451.050 ;
        RECT 31.950 450.600 34.050 451.050 ;
        RECT 16.950 449.400 34.050 450.600 ;
        RECT 16.950 448.950 19.050 449.400 ;
        RECT 31.950 448.950 34.050 449.400 ;
        RECT 37.950 450.600 40.050 451.050 ;
        RECT 61.950 450.600 64.050 451.050 ;
        RECT 37.950 449.400 64.050 450.600 ;
        RECT 37.950 448.950 40.050 449.400 ;
        RECT 61.950 448.950 64.050 449.400 ;
        RECT 97.950 450.600 100.050 451.050 ;
        RECT 107.400 450.600 108.600 455.400 ;
        RECT 115.950 454.950 118.050 455.400 ;
        RECT 121.950 456.600 124.050 457.050 ;
        RECT 142.950 456.600 145.050 457.050 ;
        RECT 193.950 456.600 196.050 457.050 ;
        RECT 244.950 456.600 247.050 457.050 ;
        RECT 121.950 455.400 141.600 456.600 ;
        RECT 121.950 454.950 124.050 455.400 ;
        RECT 140.400 454.050 141.600 455.400 ;
        RECT 142.950 455.400 196.050 456.600 ;
        RECT 142.950 454.950 145.050 455.400 ;
        RECT 193.950 454.950 196.050 455.400 ;
        RECT 200.400 455.400 247.050 456.600 ;
        RECT 200.400 454.050 201.600 455.400 ;
        RECT 244.950 454.950 247.050 455.400 ;
        RECT 274.950 456.600 277.050 457.050 ;
        RECT 301.950 456.600 304.050 457.050 ;
        RECT 334.950 456.600 337.050 457.050 ;
        RECT 274.950 455.400 288.600 456.600 ;
        RECT 274.950 454.950 277.050 455.400 ;
        RECT 287.400 454.050 288.600 455.400 ;
        RECT 301.950 455.400 337.050 456.600 ;
        RECT 301.950 454.950 304.050 455.400 ;
        RECT 334.950 454.950 337.050 455.400 ;
        RECT 340.950 454.950 343.050 457.050 ;
        RECT 362.400 456.600 363.600 457.950 ;
        RECT 397.950 456.600 400.050 457.050 ;
        RECT 362.400 455.400 400.050 456.600 ;
        RECT 109.950 453.600 112.050 454.050 ;
        RECT 112.950 453.600 115.050 454.050 ;
        RECT 118.950 453.600 121.050 454.050 ;
        RECT 109.950 452.400 121.050 453.600 ;
        RECT 109.950 451.950 112.050 452.400 ;
        RECT 112.950 451.950 115.050 452.400 ;
        RECT 118.950 451.950 121.050 452.400 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 139.950 451.950 142.050 454.050 ;
        RECT 163.950 451.950 166.050 454.050 ;
        RECT 199.950 451.950 202.050 454.050 ;
        RECT 229.950 453.600 232.050 454.050 ;
        RECT 247.950 453.600 250.050 454.050 ;
        RECT 229.950 452.400 250.050 453.600 ;
        RECT 229.950 451.950 232.050 452.400 ;
        RECT 247.950 451.950 250.050 452.400 ;
        RECT 256.950 453.600 259.050 454.050 ;
        RECT 265.950 453.600 268.050 454.050 ;
        RECT 256.950 452.400 268.050 453.600 ;
        RECT 256.950 451.950 259.050 452.400 ;
        RECT 265.950 451.950 268.050 452.400 ;
        RECT 271.950 453.600 274.050 454.050 ;
        RECT 280.950 453.600 283.050 454.050 ;
        RECT 271.950 452.400 283.050 453.600 ;
        RECT 271.950 451.950 274.050 452.400 ;
        RECT 280.950 451.950 283.050 452.400 ;
        RECT 286.950 451.950 289.050 454.050 ;
        RECT 316.950 453.600 319.050 454.050 ;
        RECT 337.950 453.600 340.050 454.050 ;
        RECT 316.950 452.400 340.050 453.600 ;
        RECT 316.950 451.950 319.050 452.400 ;
        RECT 337.950 451.950 340.050 452.400 ;
        RECT 97.950 449.400 108.600 450.600 ;
        RECT 118.950 450.600 121.050 451.050 ;
        RECT 125.400 450.600 126.600 451.950 ;
        RECT 118.950 449.400 126.600 450.600 ;
        RECT 97.950 448.950 100.050 449.400 ;
        RECT 118.950 448.950 121.050 449.400 ;
        RECT 164.400 448.050 165.600 451.950 ;
        RECT 172.950 450.600 175.050 451.050 ;
        RECT 211.950 450.600 214.050 451.050 ;
        RECT 220.950 450.600 223.050 451.050 ;
        RECT 172.950 449.400 223.050 450.600 ;
        RECT 172.950 448.950 175.050 449.400 ;
        RECT 211.950 448.950 214.050 449.400 ;
        RECT 220.950 448.950 223.050 449.400 ;
        RECT 253.950 450.600 256.050 451.050 ;
        RECT 259.950 450.600 262.050 451.050 ;
        RECT 253.950 449.400 262.050 450.600 ;
        RECT 253.950 448.950 256.050 449.400 ;
        RECT 259.950 448.950 262.050 449.400 ;
        RECT 322.950 450.600 325.050 451.050 ;
        RECT 341.400 450.600 342.600 454.950 ;
        RECT 362.400 454.050 363.600 455.400 ;
        RECT 397.950 454.950 400.050 455.400 ;
        RECT 352.950 453.600 355.050 454.050 ;
        RECT 358.950 453.600 361.050 454.050 ;
        RECT 352.950 452.400 361.050 453.600 ;
        RECT 352.950 451.950 355.050 452.400 ;
        RECT 358.950 451.950 361.050 452.400 ;
        RECT 361.950 451.950 364.050 454.050 ;
        RECT 379.950 453.600 382.050 454.050 ;
        RECT 368.400 452.400 382.050 453.600 ;
        RECT 368.400 450.600 369.600 452.400 ;
        RECT 379.950 451.950 382.050 452.400 ;
        RECT 404.400 451.050 405.600 458.400 ;
        RECT 442.950 457.950 445.050 458.400 ;
        RECT 445.950 459.600 448.050 460.050 ;
        RECT 487.950 459.600 490.050 460.050 ;
        RECT 547.950 459.600 550.050 460.050 ;
        RECT 445.950 458.400 474.600 459.600 ;
        RECT 445.950 457.950 448.050 458.400 ;
        RECT 409.950 454.950 412.050 457.050 ;
        RECT 415.950 456.600 418.050 457.050 ;
        RECT 427.950 456.600 430.050 457.050 ;
        RECT 445.950 456.600 448.050 457.050 ;
        RECT 415.950 455.400 426.600 456.600 ;
        RECT 415.950 454.950 418.050 455.400 ;
        RECT 410.400 453.600 411.600 454.950 ;
        RECT 425.400 453.600 426.600 455.400 ;
        RECT 427.950 455.400 448.050 456.600 ;
        RECT 427.950 454.950 430.050 455.400 ;
        RECT 445.950 454.950 448.050 455.400 ;
        RECT 460.950 456.600 463.050 457.050 ;
        RECT 469.950 456.600 472.050 457.050 ;
        RECT 460.950 455.400 472.050 456.600 ;
        RECT 473.400 456.600 474.600 458.400 ;
        RECT 487.950 458.400 550.050 459.600 ;
        RECT 487.950 457.950 490.050 458.400 ;
        RECT 547.950 457.950 550.050 458.400 ;
        RECT 562.950 459.600 565.050 460.050 ;
        RECT 574.950 459.600 577.050 460.050 ;
        RECT 598.950 459.600 601.050 460.050 ;
        RECT 562.950 458.400 601.050 459.600 ;
        RECT 562.950 457.950 565.050 458.400 ;
        RECT 574.950 457.950 577.050 458.400 ;
        RECT 598.950 457.950 601.050 458.400 ;
        RECT 607.950 457.950 610.050 460.050 ;
        RECT 613.950 459.600 616.050 460.050 ;
        RECT 643.950 459.600 646.050 460.050 ;
        RECT 613.950 458.400 646.050 459.600 ;
        RECT 613.950 457.950 616.050 458.400 ;
        RECT 643.950 457.950 646.050 458.400 ;
        RECT 652.950 459.600 655.050 460.050 ;
        RECT 658.950 459.600 661.050 460.050 ;
        RECT 652.950 458.400 661.050 459.600 ;
        RECT 652.950 457.950 655.050 458.400 ;
        RECT 658.950 457.950 661.050 458.400 ;
        RECT 775.950 459.600 778.050 460.050 ;
        RECT 802.950 459.600 805.050 460.050 ;
        RECT 829.950 459.600 832.050 460.050 ;
        RECT 775.950 458.400 789.600 459.600 ;
        RECT 775.950 457.950 778.050 458.400 ;
        RECT 505.950 456.600 508.050 457.050 ;
        RECT 473.400 455.400 508.050 456.600 ;
        RECT 460.950 454.950 463.050 455.400 ;
        RECT 469.950 454.950 472.050 455.400 ;
        RECT 505.950 454.950 508.050 455.400 ;
        RECT 523.950 456.600 526.050 457.050 ;
        RECT 532.950 456.600 535.050 457.050 ;
        RECT 544.950 456.600 547.050 457.050 ;
        RECT 523.950 455.400 531.600 456.600 ;
        RECT 523.950 454.950 526.050 455.400 ;
        RECT 430.950 453.600 433.050 454.050 ;
        RECT 410.400 452.400 417.600 453.600 ;
        RECT 425.400 452.400 433.050 453.600 ;
        RECT 322.950 449.400 369.600 450.600 ;
        RECT 370.950 450.600 373.050 451.050 ;
        RECT 400.950 450.600 403.050 451.050 ;
        RECT 370.950 449.400 403.050 450.600 ;
        RECT 322.950 448.950 325.050 449.400 ;
        RECT 370.950 448.950 373.050 449.400 ;
        RECT 400.950 448.950 403.050 449.400 ;
        RECT 403.950 448.950 406.050 451.050 ;
        RECT 416.400 450.600 417.600 452.400 ;
        RECT 430.950 451.950 433.050 452.400 ;
        RECT 508.950 453.600 511.050 454.050 ;
        RECT 530.400 453.600 531.600 455.400 ;
        RECT 532.950 455.400 547.050 456.600 ;
        RECT 532.950 454.950 535.050 455.400 ;
        RECT 544.950 454.950 547.050 455.400 ;
        RECT 571.950 456.600 574.050 457.050 ;
        RECT 580.950 456.600 583.050 457.050 ;
        RECT 571.950 455.400 583.050 456.600 ;
        RECT 571.950 454.950 574.050 455.400 ;
        RECT 580.950 454.950 583.050 455.400 ;
        RECT 583.950 456.600 586.050 457.050 ;
        RECT 589.950 456.600 592.050 457.050 ;
        RECT 583.950 455.400 592.050 456.600 ;
        RECT 583.950 454.950 586.050 455.400 ;
        RECT 589.950 454.950 592.050 455.400 ;
        RECT 598.950 456.600 601.050 457.050 ;
        RECT 604.950 456.600 607.050 457.050 ;
        RECT 598.950 455.400 607.050 456.600 ;
        RECT 598.950 454.950 601.050 455.400 ;
        RECT 604.950 454.950 607.050 455.400 ;
        RECT 565.950 453.600 568.050 454.050 ;
        RECT 508.950 452.400 528.600 453.600 ;
        RECT 530.400 452.400 568.050 453.600 ;
        RECT 508.950 451.950 511.050 452.400 ;
        RECT 527.400 451.050 528.600 452.400 ;
        RECT 565.950 451.950 568.050 452.400 ;
        RECT 574.950 453.600 577.050 454.050 ;
        RECT 608.400 453.600 609.600 457.950 ;
        RECT 788.400 457.050 789.600 458.400 ;
        RECT 802.950 458.400 832.050 459.600 ;
        RECT 802.950 457.950 805.050 458.400 ;
        RECT 829.950 457.950 832.050 458.400 ;
        RECT 622.950 454.950 625.050 457.050 ;
        RECT 631.950 456.600 634.050 457.050 ;
        RECT 664.950 456.600 667.050 457.050 ;
        RECT 670.950 456.600 673.050 457.050 ;
        RECT 631.950 455.400 673.050 456.600 ;
        RECT 631.950 454.950 634.050 455.400 ;
        RECT 664.950 454.950 667.050 455.400 ;
        RECT 670.950 454.950 673.050 455.400 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 703.950 456.600 706.050 457.050 ;
        RECT 712.950 456.600 715.050 457.050 ;
        RECT 703.950 455.400 715.050 456.600 ;
        RECT 703.950 454.950 706.050 455.400 ;
        RECT 712.950 454.950 715.050 455.400 ;
        RECT 715.950 456.600 718.050 457.050 ;
        RECT 748.950 456.600 751.050 457.050 ;
        RECT 715.950 455.400 751.050 456.600 ;
        RECT 715.950 454.950 718.050 455.400 ;
        RECT 748.950 454.950 751.050 455.400 ;
        RECT 754.950 456.600 757.050 457.050 ;
        RECT 769.950 456.600 772.050 457.050 ;
        RECT 754.950 455.400 772.050 456.600 ;
        RECT 754.950 454.950 757.050 455.400 ;
        RECT 769.950 454.950 772.050 455.400 ;
        RECT 787.950 454.950 790.050 457.050 ;
        RECT 826.950 456.600 829.050 457.050 ;
        RECT 850.950 456.600 853.050 457.050 ;
        RECT 826.950 455.400 853.050 456.600 ;
        RECT 826.950 454.950 829.050 455.400 ;
        RECT 850.950 454.950 853.050 455.400 ;
        RECT 574.950 452.400 609.600 453.600 ;
        RECT 623.400 453.600 624.600 454.950 ;
        RECT 679.950 453.600 682.050 454.050 ;
        RECT 623.400 452.400 682.050 453.600 ;
        RECT 574.950 451.950 577.050 452.400 ;
        RECT 679.950 451.950 682.050 452.400 ;
        RECT 692.400 451.050 693.600 454.950 ;
        RECT 694.950 453.600 697.050 454.050 ;
        RECT 733.950 453.600 736.050 454.050 ;
        RECT 694.950 452.400 736.050 453.600 ;
        RECT 694.950 451.950 697.050 452.400 ;
        RECT 733.950 451.950 736.050 452.400 ;
        RECT 778.950 453.600 781.050 454.050 ;
        RECT 841.950 453.600 844.050 454.050 ;
        RECT 778.950 452.400 844.050 453.600 ;
        RECT 778.950 451.950 781.050 452.400 ;
        RECT 841.950 451.950 844.050 452.400 ;
        RECT 460.950 450.600 463.050 451.050 ;
        RECT 484.950 450.600 487.050 451.050 ;
        RECT 416.400 449.400 487.050 450.600 ;
        RECT 460.950 448.950 463.050 449.400 ;
        RECT 484.950 448.950 487.050 449.400 ;
        RECT 508.950 450.600 511.050 451.050 ;
        RECT 517.950 450.600 520.050 451.050 ;
        RECT 508.950 449.400 520.050 450.600 ;
        RECT 508.950 448.950 511.050 449.400 ;
        RECT 517.950 448.950 520.050 449.400 ;
        RECT 526.950 448.950 529.050 451.050 ;
        RECT 529.950 450.600 532.050 451.050 ;
        RECT 550.950 450.600 553.050 451.050 ;
        RECT 583.950 450.600 586.050 451.050 ;
        RECT 529.950 449.400 586.050 450.600 ;
        RECT 529.950 448.950 532.050 449.400 ;
        RECT 550.950 448.950 553.050 449.400 ;
        RECT 583.950 448.950 586.050 449.400 ;
        RECT 628.950 450.600 631.050 451.050 ;
        RECT 652.950 450.600 655.050 451.050 ;
        RECT 655.950 450.600 658.050 451.050 ;
        RECT 628.950 449.400 658.050 450.600 ;
        RECT 628.950 448.950 631.050 449.400 ;
        RECT 652.950 448.950 655.050 449.400 ;
        RECT 655.950 448.950 658.050 449.400 ;
        RECT 691.950 448.950 694.050 451.050 ;
        RECT 10.950 447.600 13.050 448.050 ;
        RECT 16.950 447.600 19.050 448.050 ;
        RECT 10.950 446.400 19.050 447.600 ;
        RECT 10.950 445.950 13.050 446.400 ;
        RECT 16.950 445.950 19.050 446.400 ;
        RECT 31.950 447.600 34.050 448.050 ;
        RECT 55.950 447.600 58.050 448.050 ;
        RECT 31.950 446.400 58.050 447.600 ;
        RECT 31.950 445.950 34.050 446.400 ;
        RECT 55.950 445.950 58.050 446.400 ;
        RECT 112.950 447.600 115.050 448.050 ;
        RECT 160.950 447.600 163.050 448.050 ;
        RECT 112.950 446.400 163.050 447.600 ;
        RECT 112.950 445.950 115.050 446.400 ;
        RECT 160.950 445.950 163.050 446.400 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 232.950 447.600 235.050 448.050 ;
        RECT 253.950 447.600 256.050 448.050 ;
        RECT 295.950 447.600 298.050 448.050 ;
        RECT 232.950 446.400 298.050 447.600 ;
        RECT 232.950 445.950 235.050 446.400 ;
        RECT 253.950 445.950 256.050 446.400 ;
        RECT 295.950 445.950 298.050 446.400 ;
        RECT 406.950 447.600 409.050 448.050 ;
        RECT 466.950 447.600 469.050 448.050 ;
        RECT 406.950 446.400 469.050 447.600 ;
        RECT 406.950 445.950 409.050 446.400 ;
        RECT 466.950 445.950 469.050 446.400 ;
        RECT 580.950 447.600 583.050 448.050 ;
        RECT 592.950 447.600 595.050 448.050 ;
        RECT 616.950 447.600 619.050 448.050 ;
        RECT 634.950 447.600 637.050 448.050 ;
        RECT 580.950 446.400 637.050 447.600 ;
        RECT 580.950 445.950 583.050 446.400 ;
        RECT 592.950 445.950 595.050 446.400 ;
        RECT 616.950 445.950 619.050 446.400 ;
        RECT 634.950 445.950 637.050 446.400 ;
        RECT 97.950 444.600 100.050 445.050 ;
        RECT 166.950 444.600 169.050 445.050 ;
        RECT 190.950 444.600 193.050 445.050 ;
        RECT 97.950 443.400 193.050 444.600 ;
        RECT 97.950 442.950 100.050 443.400 ;
        RECT 166.950 442.950 169.050 443.400 ;
        RECT 190.950 442.950 193.050 443.400 ;
        RECT 223.950 444.600 226.050 445.050 ;
        RECT 247.950 444.600 250.050 445.050 ;
        RECT 223.950 443.400 250.050 444.600 ;
        RECT 223.950 442.950 226.050 443.400 ;
        RECT 247.950 442.950 250.050 443.400 ;
        RECT 328.950 444.600 331.050 445.050 ;
        RECT 406.950 444.600 409.050 445.050 ;
        RECT 328.950 443.400 409.050 444.600 ;
        RECT 328.950 442.950 331.050 443.400 ;
        RECT 406.950 442.950 409.050 443.400 ;
        RECT 433.950 444.600 436.050 445.050 ;
        RECT 514.950 444.600 517.050 445.050 ;
        RECT 718.950 444.600 721.050 445.050 ;
        RECT 433.950 443.400 517.050 444.600 ;
        RECT 433.950 442.950 436.050 443.400 ;
        RECT 514.950 442.950 517.050 443.400 ;
        RECT 551.400 443.400 721.050 444.600 ;
        RECT 295.950 441.600 298.050 442.050 ;
        RECT 493.950 441.600 496.050 442.050 ;
        RECT 295.950 440.400 496.050 441.600 ;
        RECT 295.950 439.950 298.050 440.400 ;
        RECT 493.950 439.950 496.050 440.400 ;
        RECT 505.950 441.600 508.050 442.050 ;
        RECT 551.400 441.600 552.600 443.400 ;
        RECT 718.950 442.950 721.050 443.400 ;
        RECT 571.950 441.600 574.050 442.050 ;
        RECT 505.950 440.400 552.600 441.600 ;
        RECT 557.400 440.400 574.050 441.600 ;
        RECT 505.950 439.950 508.050 440.400 ;
        RECT 154.950 438.600 157.050 439.050 ;
        RECT 208.950 438.600 211.050 439.050 ;
        RECT 154.950 437.400 211.050 438.600 ;
        RECT 154.950 436.950 157.050 437.400 ;
        RECT 208.950 436.950 211.050 437.400 ;
        RECT 334.950 438.600 337.050 439.050 ;
        RECT 364.950 438.600 367.050 439.050 ;
        RECT 388.950 438.600 391.050 439.050 ;
        RECT 334.950 437.400 391.050 438.600 ;
        RECT 334.950 436.950 337.050 437.400 ;
        RECT 364.950 436.950 367.050 437.400 ;
        RECT 388.950 436.950 391.050 437.400 ;
        RECT 445.950 438.600 448.050 439.050 ;
        RECT 469.950 438.600 472.050 439.050 ;
        RECT 557.400 438.600 558.600 440.400 ;
        RECT 571.950 439.950 574.050 440.400 ;
        RECT 661.950 441.600 664.050 442.050 ;
        RECT 709.950 441.600 712.050 442.050 ;
        RECT 661.950 440.400 712.050 441.600 ;
        RECT 661.950 439.950 664.050 440.400 ;
        RECT 709.950 439.950 712.050 440.400 ;
        RECT 445.950 437.400 472.050 438.600 ;
        RECT 445.950 436.950 448.050 437.400 ;
        RECT 469.950 436.950 472.050 437.400 ;
        RECT 476.400 437.400 558.600 438.600 ;
        RECT 835.950 438.600 838.050 439.050 ;
        RECT 859.950 438.600 862.050 439.050 ;
        RECT 835.950 437.400 862.050 438.600 ;
        RECT 70.950 435.600 73.050 436.050 ;
        RECT 319.950 435.600 322.050 436.050 ;
        RECT 70.950 434.400 322.050 435.600 ;
        RECT 70.950 433.950 73.050 434.400 ;
        RECT 319.950 433.950 322.050 434.400 ;
        RECT 328.950 435.600 331.050 436.050 ;
        RECT 476.400 435.600 477.600 437.400 ;
        RECT 835.950 436.950 838.050 437.400 ;
        RECT 859.950 436.950 862.050 437.400 ;
        RECT 328.950 434.400 477.600 435.600 ;
        RECT 574.950 435.600 577.050 436.050 ;
        RECT 601.950 435.600 604.050 436.050 ;
        RECT 574.950 434.400 604.050 435.600 ;
        RECT 328.950 433.950 331.050 434.400 ;
        RECT 574.950 433.950 577.050 434.400 ;
        RECT 601.950 433.950 604.050 434.400 ;
        RECT 241.950 432.600 244.050 433.050 ;
        RECT 427.950 432.600 430.050 433.050 ;
        RECT 433.950 432.600 436.050 433.050 ;
        RECT 241.950 431.400 436.050 432.600 ;
        RECT 241.950 430.950 244.050 431.400 ;
        RECT 427.950 430.950 430.050 431.400 ;
        RECT 433.950 430.950 436.050 431.400 ;
        RECT 469.950 432.600 472.050 433.050 ;
        RECT 601.950 432.600 604.050 433.050 ;
        RECT 469.950 431.400 604.050 432.600 ;
        RECT 469.950 430.950 472.050 431.400 ;
        RECT 601.950 430.950 604.050 431.400 ;
        RECT 286.950 429.600 289.050 430.050 ;
        RECT 304.950 429.600 307.050 430.050 ;
        RECT 286.950 428.400 307.050 429.600 ;
        RECT 286.950 427.950 289.050 428.400 ;
        RECT 304.950 427.950 307.050 428.400 ;
        RECT 415.950 429.600 418.050 430.050 ;
        RECT 430.950 429.600 433.050 430.050 ;
        RECT 415.950 428.400 433.050 429.600 ;
        RECT 415.950 427.950 418.050 428.400 ;
        RECT 430.950 427.950 433.050 428.400 ;
        RECT 493.950 426.600 496.050 427.050 ;
        RECT 556.950 426.600 559.050 427.050 ;
        RECT 667.950 426.600 670.050 427.050 ;
        RECT 493.950 425.400 670.050 426.600 ;
        RECT 493.950 424.950 496.050 425.400 ;
        RECT 556.950 424.950 559.050 425.400 ;
        RECT 667.950 424.950 670.050 425.400 ;
        RECT 814.950 426.600 817.050 427.050 ;
        RECT 823.950 426.600 826.050 427.050 ;
        RECT 814.950 425.400 826.050 426.600 ;
        RECT 814.950 424.950 817.050 425.400 ;
        RECT 823.950 424.950 826.050 425.400 ;
        RECT 73.950 423.600 76.050 424.050 ;
        RECT 127.950 423.600 130.050 424.050 ;
        RECT 73.950 422.400 130.050 423.600 ;
        RECT 73.950 421.950 76.050 422.400 ;
        RECT 127.950 421.950 130.050 422.400 ;
        RECT 193.950 423.600 196.050 424.050 ;
        RECT 307.950 423.600 310.050 424.050 ;
        RECT 193.950 422.400 310.050 423.600 ;
        RECT 193.950 421.950 196.050 422.400 ;
        RECT 307.950 421.950 310.050 422.400 ;
        RECT 316.950 423.600 319.050 424.050 ;
        RECT 325.950 423.600 328.050 424.050 ;
        RECT 316.950 422.400 328.050 423.600 ;
        RECT 316.950 421.950 319.050 422.400 ;
        RECT 325.950 421.950 328.050 422.400 ;
        RECT 385.950 423.600 388.050 424.050 ;
        RECT 454.950 423.600 457.050 424.050 ;
        RECT 385.950 422.400 457.050 423.600 ;
        RECT 385.950 421.950 388.050 422.400 ;
        RECT 454.950 421.950 457.050 422.400 ;
        RECT 466.950 423.600 469.050 424.050 ;
        RECT 577.950 423.600 580.050 424.050 ;
        RECT 580.950 423.600 583.050 424.050 ;
        RECT 466.950 422.400 583.050 423.600 ;
        RECT 466.950 421.950 469.050 422.400 ;
        RECT 577.950 421.950 580.050 422.400 ;
        RECT 580.950 421.950 583.050 422.400 ;
        RECT 637.950 423.600 640.050 424.050 ;
        RECT 691.950 423.600 694.050 424.050 ;
        RECT 637.950 422.400 694.050 423.600 ;
        RECT 637.950 421.950 640.050 422.400 ;
        RECT 691.950 421.950 694.050 422.400 ;
        RECT 10.950 420.600 13.050 421.050 ;
        RECT 37.950 420.600 40.050 421.050 ;
        RECT 10.950 419.400 40.050 420.600 ;
        RECT 10.950 418.950 13.050 419.400 ;
        RECT 37.950 418.950 40.050 419.400 ;
        RECT 115.950 420.600 118.050 421.050 ;
        RECT 121.950 420.600 124.050 421.050 ;
        RECT 133.950 420.600 136.050 421.050 ;
        RECT 115.950 419.400 136.050 420.600 ;
        RECT 115.950 418.950 118.050 419.400 ;
        RECT 121.950 418.950 124.050 419.400 ;
        RECT 133.950 418.950 136.050 419.400 ;
        RECT 289.950 420.600 292.050 421.050 ;
        RECT 298.950 420.600 301.050 421.050 ;
        RECT 289.950 419.400 301.050 420.600 ;
        RECT 289.950 418.950 292.050 419.400 ;
        RECT 298.950 418.950 301.050 419.400 ;
        RECT 325.950 420.600 328.050 421.050 ;
        RECT 346.950 420.600 349.050 421.050 ;
        RECT 325.950 419.400 349.050 420.600 ;
        RECT 325.950 418.950 328.050 419.400 ;
        RECT 346.950 418.950 349.050 419.400 ;
        RECT 364.950 420.600 367.050 421.050 ;
        RECT 412.950 420.600 415.050 421.050 ;
        RECT 364.950 419.400 415.050 420.600 ;
        RECT 364.950 418.950 367.050 419.400 ;
        RECT 412.950 418.950 415.050 419.400 ;
        RECT 424.950 420.600 427.050 421.050 ;
        RECT 436.950 420.600 439.050 421.050 ;
        RECT 424.950 419.400 439.050 420.600 ;
        RECT 424.950 418.950 427.050 419.400 ;
        RECT 436.950 418.950 439.050 419.400 ;
        RECT 475.950 420.600 478.050 421.050 ;
        RECT 487.950 420.600 490.050 421.050 ;
        RECT 475.950 419.400 490.050 420.600 ;
        RECT 475.950 418.950 478.050 419.400 ;
        RECT 487.950 418.950 490.050 419.400 ;
        RECT 520.950 420.600 523.050 421.050 ;
        RECT 526.950 420.600 529.050 421.050 ;
        RECT 520.950 419.400 529.050 420.600 ;
        RECT 520.950 418.950 523.050 419.400 ;
        RECT 526.950 418.950 529.050 419.400 ;
        RECT 547.950 420.600 550.050 421.050 ;
        RECT 559.950 420.600 562.050 421.050 ;
        RECT 547.950 419.400 562.050 420.600 ;
        RECT 547.950 418.950 550.050 419.400 ;
        RECT 559.950 418.950 562.050 419.400 ;
        RECT 589.950 420.600 592.050 421.050 ;
        RECT 595.950 420.600 598.050 421.050 ;
        RECT 589.950 419.400 598.050 420.600 ;
        RECT 589.950 418.950 592.050 419.400 ;
        RECT 595.950 418.950 598.050 419.400 ;
        RECT 598.950 420.600 601.050 421.050 ;
        RECT 643.950 420.600 646.050 421.050 ;
        RECT 598.950 419.400 646.050 420.600 ;
        RECT 598.950 418.950 601.050 419.400 ;
        RECT 643.950 418.950 646.050 419.400 ;
        RECT 16.950 417.600 19.050 418.050 ;
        RECT 55.950 417.600 58.050 418.050 ;
        RECT 11.400 416.400 19.050 417.600 ;
        RECT 11.400 411.600 12.600 416.400 ;
        RECT 16.950 415.950 19.050 416.400 ;
        RECT 47.400 416.400 58.050 417.600 ;
        RECT 13.950 414.600 16.050 415.050 ;
        RECT 47.400 414.600 48.600 416.400 ;
        RECT 55.950 415.950 58.050 416.400 ;
        RECT 91.950 417.600 94.050 418.050 ;
        RECT 106.950 417.600 109.050 418.050 ;
        RECT 118.950 417.600 121.050 418.050 ;
        RECT 133.950 417.600 136.050 418.050 ;
        RECT 91.950 416.400 136.050 417.600 ;
        RECT 91.950 415.950 94.050 416.400 ;
        RECT 106.950 415.950 109.050 416.400 ;
        RECT 118.950 415.950 121.050 416.400 ;
        RECT 133.950 415.950 136.050 416.400 ;
        RECT 139.950 417.600 142.050 418.050 ;
        RECT 160.950 417.600 163.050 418.050 ;
        RECT 139.950 416.400 163.050 417.600 ;
        RECT 139.950 415.950 142.050 416.400 ;
        RECT 160.950 415.950 163.050 416.400 ;
        RECT 196.950 417.600 199.050 418.050 ;
        RECT 301.950 417.600 304.050 418.050 ;
        RECT 196.950 416.400 304.050 417.600 ;
        RECT 196.950 415.950 199.050 416.400 ;
        RECT 301.950 415.950 304.050 416.400 ;
        RECT 328.950 415.950 331.050 418.050 ;
        RECT 331.950 417.600 334.050 418.050 ;
        RECT 355.950 417.600 358.050 418.050 ;
        RECT 367.950 417.600 370.050 418.050 ;
        RECT 331.950 416.400 370.050 417.600 ;
        RECT 331.950 415.950 334.050 416.400 ;
        RECT 355.950 415.950 358.050 416.400 ;
        RECT 367.950 415.950 370.050 416.400 ;
        RECT 394.950 417.600 397.050 418.050 ;
        RECT 400.950 417.600 403.050 418.050 ;
        RECT 394.950 416.400 403.050 417.600 ;
        RECT 394.950 415.950 397.050 416.400 ;
        RECT 400.950 415.950 403.050 416.400 ;
        RECT 412.950 417.600 415.050 418.050 ;
        RECT 448.950 417.600 451.050 418.050 ;
        RECT 454.950 417.600 457.050 418.050 ;
        RECT 412.950 416.400 457.050 417.600 ;
        RECT 412.950 415.950 415.050 416.400 ;
        RECT 448.950 415.950 451.050 416.400 ;
        RECT 454.950 415.950 457.050 416.400 ;
        RECT 460.950 417.600 463.050 418.050 ;
        RECT 466.950 417.600 469.050 418.050 ;
        RECT 460.950 416.400 469.050 417.600 ;
        RECT 460.950 415.950 463.050 416.400 ;
        RECT 466.950 415.950 469.050 416.400 ;
        RECT 472.950 417.600 475.050 418.050 ;
        RECT 481.950 417.600 484.050 418.050 ;
        RECT 496.950 417.600 499.050 418.050 ;
        RECT 472.950 416.400 484.050 417.600 ;
        RECT 472.950 415.950 475.050 416.400 ;
        RECT 481.950 415.950 484.050 416.400 ;
        RECT 485.400 416.400 499.050 417.600 ;
        RECT 13.950 413.400 48.600 414.600 ;
        RECT 49.950 414.600 52.050 415.050 ;
        RECT 61.950 414.600 64.050 415.050 ;
        RECT 49.950 413.400 64.050 414.600 ;
        RECT 13.950 412.950 16.050 413.400 ;
        RECT 49.950 412.950 52.050 413.400 ;
        RECT 61.950 412.950 64.050 413.400 ;
        RECT 67.950 414.600 70.050 415.050 ;
        RECT 79.950 414.600 82.050 415.050 ;
        RECT 67.950 413.400 82.050 414.600 ;
        RECT 67.950 412.950 70.050 413.400 ;
        RECT 79.950 412.950 82.050 413.400 ;
        RECT 88.950 414.600 91.050 415.050 ;
        RECT 97.950 414.600 100.050 415.050 ;
        RECT 88.950 413.400 100.050 414.600 ;
        RECT 88.950 412.950 91.050 413.400 ;
        RECT 97.950 412.950 100.050 413.400 ;
        RECT 124.950 414.600 127.050 415.050 ;
        RECT 139.950 414.600 142.050 415.050 ;
        RECT 124.950 413.400 142.050 414.600 ;
        RECT 124.950 412.950 127.050 413.400 ;
        RECT 139.950 412.950 142.050 413.400 ;
        RECT 190.950 414.600 193.050 415.050 ;
        RECT 199.950 414.600 202.050 415.050 ;
        RECT 205.950 414.600 208.050 415.050 ;
        RECT 190.950 413.400 208.050 414.600 ;
        RECT 190.950 412.950 193.050 413.400 ;
        RECT 199.950 412.950 202.050 413.400 ;
        RECT 205.950 412.950 208.050 413.400 ;
        RECT 211.950 414.600 214.050 415.050 ;
        RECT 220.950 414.600 223.050 415.050 ;
        RECT 226.950 414.600 229.050 415.050 ;
        RECT 271.950 414.600 274.050 415.050 ;
        RECT 292.950 414.600 295.050 415.050 ;
        RECT 211.950 413.400 229.050 414.600 ;
        RECT 211.950 412.950 214.050 413.400 ;
        RECT 220.950 412.950 223.050 413.400 ;
        RECT 226.950 412.950 229.050 413.400 ;
        RECT 245.400 413.400 295.050 414.600 ;
        RECT 329.400 414.600 330.600 415.950 ;
        RECT 352.950 414.600 355.050 415.050 ;
        RECT 361.950 414.600 364.050 415.050 ;
        RECT 397.950 414.600 400.050 415.050 ;
        RECT 424.950 414.600 427.050 415.050 ;
        RECT 485.400 414.600 486.600 416.400 ;
        RECT 496.950 415.950 499.050 416.400 ;
        RECT 505.950 417.600 508.050 418.050 ;
        RECT 511.950 417.600 514.050 418.050 ;
        RECT 505.950 416.400 514.050 417.600 ;
        RECT 505.950 415.950 508.050 416.400 ;
        RECT 511.950 415.950 514.050 416.400 ;
        RECT 514.950 417.600 517.050 418.050 ;
        RECT 553.950 417.600 556.050 418.050 ;
        RECT 514.950 416.400 556.050 417.600 ;
        RECT 514.950 415.950 517.050 416.400 ;
        RECT 553.950 415.950 556.050 416.400 ;
        RECT 571.950 417.600 574.050 418.050 ;
        RECT 598.950 417.600 601.050 418.050 ;
        RECT 571.950 416.400 601.050 417.600 ;
        RECT 571.950 415.950 574.050 416.400 ;
        RECT 598.950 415.950 601.050 416.400 ;
        RECT 601.950 417.600 604.050 418.050 ;
        RECT 622.950 417.600 625.050 418.050 ;
        RECT 625.950 417.600 628.050 418.050 ;
        RECT 601.950 416.400 628.050 417.600 ;
        RECT 601.950 415.950 604.050 416.400 ;
        RECT 622.950 415.950 625.050 416.400 ;
        RECT 625.950 415.950 628.050 416.400 ;
        RECT 631.950 417.600 634.050 418.050 ;
        RECT 637.950 417.600 640.050 418.050 ;
        RECT 631.950 416.400 640.050 417.600 ;
        RECT 631.950 415.950 634.050 416.400 ;
        RECT 637.950 415.950 640.050 416.400 ;
        RECT 688.950 415.950 691.050 418.050 ;
        RECT 329.400 413.400 333.600 414.600 ;
        RECT 245.400 412.050 246.600 413.400 ;
        RECT 271.950 412.950 274.050 413.400 ;
        RECT 292.950 412.950 295.050 413.400 ;
        RECT 332.400 412.050 333.600 413.400 ;
        RECT 352.950 413.400 400.050 414.600 ;
        RECT 352.950 412.950 355.050 413.400 ;
        RECT 361.950 412.950 364.050 413.400 ;
        RECT 397.950 412.950 400.050 413.400 ;
        RECT 422.400 413.400 427.050 414.600 ;
        RECT 13.950 411.600 16.050 412.050 ;
        RECT 11.400 410.400 16.050 411.600 ;
        RECT 13.950 409.950 16.050 410.400 ;
        RECT 16.950 411.600 19.050 412.050 ;
        RECT 22.950 411.600 25.050 412.050 ;
        RECT 16.950 410.400 25.050 411.600 ;
        RECT 16.950 409.950 19.050 410.400 ;
        RECT 22.950 409.950 25.050 410.400 ;
        RECT 31.950 411.600 34.050 412.050 ;
        RECT 73.950 411.600 76.050 412.050 ;
        RECT 31.950 410.400 76.050 411.600 ;
        RECT 31.950 409.950 34.050 410.400 ;
        RECT 73.950 409.950 76.050 410.400 ;
        RECT 82.950 411.600 85.050 412.050 ;
        RECT 85.950 411.600 88.050 412.050 ;
        RECT 100.950 411.600 103.050 412.050 ;
        RECT 82.950 410.400 103.050 411.600 ;
        RECT 82.950 409.950 85.050 410.400 ;
        RECT 85.950 409.950 88.050 410.400 ;
        RECT 100.950 409.950 103.050 410.400 ;
        RECT 109.950 411.600 112.050 412.050 ;
        RECT 115.950 411.600 118.050 412.050 ;
        RECT 109.950 410.400 118.050 411.600 ;
        RECT 109.950 409.950 112.050 410.400 ;
        RECT 115.950 409.950 118.050 410.400 ;
        RECT 148.950 411.600 151.050 412.050 ;
        RECT 196.950 411.600 199.050 412.050 ;
        RECT 148.950 410.400 199.050 411.600 ;
        RECT 148.950 409.950 151.050 410.400 ;
        RECT 196.950 409.950 199.050 410.400 ;
        RECT 208.950 411.600 211.050 412.050 ;
        RECT 223.950 411.600 226.050 412.050 ;
        RECT 208.950 410.400 226.050 411.600 ;
        RECT 208.950 409.950 211.050 410.400 ;
        RECT 223.950 409.950 226.050 410.400 ;
        RECT 232.950 411.600 235.050 412.050 ;
        RECT 244.950 411.600 247.050 412.050 ;
        RECT 265.950 411.600 268.050 412.050 ;
        RECT 232.950 410.400 247.050 411.600 ;
        RECT 232.950 409.950 235.050 410.400 ;
        RECT 244.950 409.950 247.050 410.400 ;
        RECT 248.400 410.400 268.050 411.600 ;
        RECT 28.950 408.600 31.050 409.050 ;
        RECT 58.950 408.600 61.050 409.050 ;
        RECT 28.950 407.400 61.050 408.600 ;
        RECT 28.950 406.950 31.050 407.400 ;
        RECT 58.950 406.950 61.050 407.400 ;
        RECT 70.950 408.600 73.050 409.050 ;
        RECT 112.950 408.600 115.050 409.050 ;
        RECT 70.950 407.400 115.050 408.600 ;
        RECT 70.950 406.950 73.050 407.400 ;
        RECT 112.950 406.950 115.050 407.400 ;
        RECT 133.950 408.600 136.050 409.050 ;
        RECT 142.950 408.600 145.050 409.050 ;
        RECT 133.950 407.400 145.050 408.600 ;
        RECT 133.950 406.950 136.050 407.400 ;
        RECT 142.950 406.950 145.050 407.400 ;
        RECT 199.950 408.600 202.050 409.050 ;
        RECT 248.400 408.600 249.600 410.400 ;
        RECT 265.950 409.950 268.050 410.400 ;
        RECT 292.950 411.600 295.050 412.050 ;
        RECT 298.950 411.600 301.050 412.050 ;
        RECT 292.950 410.400 301.050 411.600 ;
        RECT 292.950 409.950 295.050 410.400 ;
        RECT 298.950 409.950 301.050 410.400 ;
        RECT 322.950 411.600 325.050 412.050 ;
        RECT 328.950 411.600 331.050 412.050 ;
        RECT 322.950 410.400 331.050 411.600 ;
        RECT 322.950 409.950 325.050 410.400 ;
        RECT 328.950 409.950 331.050 410.400 ;
        RECT 331.950 409.950 334.050 412.050 ;
        RECT 367.950 411.600 370.050 412.050 ;
        RECT 403.950 411.600 406.050 412.050 ;
        RECT 367.950 410.400 406.050 411.600 ;
        RECT 367.950 409.950 370.050 410.400 ;
        RECT 403.950 409.950 406.050 410.400 ;
        RECT 199.950 407.400 249.600 408.600 ;
        RECT 250.950 408.600 253.050 409.050 ;
        RECT 274.950 408.600 277.050 409.050 ;
        RECT 250.950 407.400 277.050 408.600 ;
        RECT 199.950 406.950 202.050 407.400 ;
        RECT 250.950 406.950 253.050 407.400 ;
        RECT 274.950 406.950 277.050 407.400 ;
        RECT 343.950 408.600 346.050 409.050 ;
        RECT 397.950 408.600 400.050 409.050 ;
        RECT 343.950 407.400 400.050 408.600 ;
        RECT 343.950 406.950 346.050 407.400 ;
        RECT 397.950 406.950 400.050 407.400 ;
        RECT 422.400 406.050 423.600 413.400 ;
        RECT 424.950 412.950 427.050 413.400 ;
        RECT 455.400 413.400 486.600 414.600 ;
        RECT 455.400 412.050 456.600 413.400 ;
        RECT 499.950 412.950 502.050 415.050 ;
        RECT 556.950 414.600 559.050 415.050 ;
        RECT 562.950 414.600 565.050 415.050 ;
        RECT 556.950 413.400 565.050 414.600 ;
        RECT 556.950 412.950 559.050 413.400 ;
        RECT 562.950 412.950 565.050 413.400 ;
        RECT 595.950 414.600 598.050 415.050 ;
        RECT 613.950 414.600 616.050 415.050 ;
        RECT 628.950 414.600 631.050 415.050 ;
        RECT 595.950 413.400 631.050 414.600 ;
        RECT 595.950 412.950 598.050 413.400 ;
        RECT 613.950 412.950 616.050 413.400 ;
        RECT 628.950 412.950 631.050 413.400 ;
        RECT 634.950 414.600 637.050 415.050 ;
        RECT 661.950 414.600 664.050 415.050 ;
        RECT 634.950 413.400 664.050 414.600 ;
        RECT 634.950 412.950 637.050 413.400 ;
        RECT 661.950 412.950 664.050 413.400 ;
        RECT 424.950 411.600 427.050 412.050 ;
        RECT 436.950 411.600 439.050 412.050 ;
        RECT 424.950 410.400 439.050 411.600 ;
        RECT 424.950 409.950 427.050 410.400 ;
        RECT 436.950 409.950 439.050 410.400 ;
        RECT 454.950 409.950 457.050 412.050 ;
        RECT 463.950 411.600 466.050 412.050 ;
        RECT 469.950 411.600 472.050 412.050 ;
        RECT 463.950 410.400 472.050 411.600 ;
        RECT 463.950 409.950 466.050 410.400 ;
        RECT 469.950 409.950 472.050 410.400 ;
        RECT 484.950 411.600 487.050 412.050 ;
        RECT 496.950 411.600 499.050 412.050 ;
        RECT 484.950 410.400 499.050 411.600 ;
        RECT 500.400 411.600 501.600 412.950 ;
        RECT 689.400 412.050 690.600 415.950 ;
        RECT 745.950 414.600 748.050 415.050 ;
        RECT 751.950 414.600 754.050 415.050 ;
        RECT 745.950 413.400 754.050 414.600 ;
        RECT 745.950 412.950 748.050 413.400 ;
        RECT 751.950 412.950 754.050 413.400 ;
        RECT 757.950 414.600 760.050 415.050 ;
        RECT 772.950 414.600 775.050 415.050 ;
        RECT 796.950 414.600 799.050 415.050 ;
        RECT 757.950 413.400 775.050 414.600 ;
        RECT 757.950 412.950 760.050 413.400 ;
        RECT 772.950 412.950 775.050 413.400 ;
        RECT 776.400 413.400 799.050 414.600 ;
        RECT 776.400 412.050 777.600 413.400 ;
        RECT 796.950 412.950 799.050 413.400 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 514.950 411.600 517.050 412.050 ;
        RECT 500.400 410.400 517.050 411.600 ;
        RECT 484.950 409.950 487.050 410.400 ;
        RECT 496.950 409.950 499.050 410.400 ;
        RECT 514.950 409.950 517.050 410.400 ;
        RECT 526.950 411.600 529.050 412.050 ;
        RECT 538.950 411.600 541.050 412.050 ;
        RECT 526.950 410.400 541.050 411.600 ;
        RECT 526.950 409.950 529.050 410.400 ;
        RECT 538.950 409.950 541.050 410.400 ;
        RECT 565.950 411.600 568.050 412.050 ;
        RECT 637.950 411.600 640.050 412.050 ;
        RECT 565.950 410.400 640.050 411.600 ;
        RECT 565.950 409.950 568.050 410.400 ;
        RECT 637.950 409.950 640.050 410.400 ;
        RECT 688.950 409.950 691.050 412.050 ;
        RECT 703.950 411.600 706.050 412.050 ;
        RECT 715.950 411.600 718.050 412.050 ;
        RECT 703.950 410.400 718.050 411.600 ;
        RECT 703.950 409.950 706.050 410.400 ;
        RECT 715.950 409.950 718.050 410.400 ;
        RECT 775.950 409.950 778.050 412.050 ;
        RECT 796.950 411.600 799.050 412.050 ;
        RECT 802.950 411.600 805.050 412.050 ;
        RECT 796.950 410.400 805.050 411.600 ;
        RECT 796.950 409.950 799.050 410.400 ;
        RECT 802.950 409.950 805.050 410.400 ;
        RECT 820.950 411.600 823.050 412.050 ;
        RECT 829.950 411.600 832.050 412.050 ;
        RECT 820.950 410.400 832.050 411.600 ;
        RECT 845.400 411.600 846.600 412.950 ;
        RECT 850.950 411.600 853.050 412.050 ;
        RECT 845.400 410.400 853.050 411.600 ;
        RECT 820.950 409.950 823.050 410.400 ;
        RECT 829.950 409.950 832.050 410.400 ;
        RECT 850.950 409.950 853.050 410.400 ;
        RECT 430.950 408.600 433.050 409.050 ;
        RECT 436.950 408.600 439.050 409.050 ;
        RECT 448.950 408.600 451.050 409.050 ;
        RECT 430.950 407.400 451.050 408.600 ;
        RECT 430.950 406.950 433.050 407.400 ;
        RECT 436.950 406.950 439.050 407.400 ;
        RECT 448.950 406.950 451.050 407.400 ;
        RECT 487.950 408.600 490.050 409.050 ;
        RECT 502.950 408.600 505.050 409.050 ;
        RECT 511.950 408.600 514.050 409.050 ;
        RECT 523.950 408.600 526.050 409.050 ;
        RECT 535.950 408.600 538.050 409.050 ;
        RECT 487.950 407.400 501.600 408.600 ;
        RECT 487.950 406.950 490.050 407.400 ;
        RECT 64.950 405.600 67.050 406.050 ;
        RECT 94.950 405.600 97.050 406.050 ;
        RECT 109.950 405.600 112.050 406.050 ;
        RECT 139.950 405.600 142.050 406.050 ;
        RECT 64.950 404.400 142.050 405.600 ;
        RECT 64.950 403.950 67.050 404.400 ;
        RECT 94.950 403.950 97.050 404.400 ;
        RECT 109.950 403.950 112.050 404.400 ;
        RECT 139.950 403.950 142.050 404.400 ;
        RECT 193.950 405.600 196.050 406.050 ;
        RECT 247.950 405.600 250.050 406.050 ;
        RECT 193.950 404.400 250.050 405.600 ;
        RECT 193.950 403.950 196.050 404.400 ;
        RECT 247.950 403.950 250.050 404.400 ;
        RECT 262.950 405.600 265.050 406.050 ;
        RECT 268.950 405.600 271.050 406.050 ;
        RECT 262.950 404.400 271.050 405.600 ;
        RECT 262.950 403.950 265.050 404.400 ;
        RECT 268.950 403.950 271.050 404.400 ;
        RECT 337.950 405.600 340.050 406.050 ;
        RECT 346.950 405.600 349.050 406.050 ;
        RECT 370.950 405.600 373.050 406.050 ;
        RECT 337.950 404.400 373.050 405.600 ;
        RECT 337.950 403.950 340.050 404.400 ;
        RECT 346.950 403.950 349.050 404.400 ;
        RECT 370.950 403.950 373.050 404.400 ;
        RECT 373.950 405.600 376.050 406.050 ;
        RECT 409.950 405.600 412.050 406.050 ;
        RECT 373.950 404.400 412.050 405.600 ;
        RECT 373.950 403.950 376.050 404.400 ;
        RECT 409.950 403.950 412.050 404.400 ;
        RECT 421.950 403.950 424.050 406.050 ;
        RECT 500.400 405.600 501.600 407.400 ;
        RECT 502.950 407.400 538.050 408.600 ;
        RECT 502.950 406.950 505.050 407.400 ;
        RECT 511.950 406.950 514.050 407.400 ;
        RECT 523.950 406.950 526.050 407.400 ;
        RECT 535.950 406.950 538.050 407.400 ;
        RECT 550.950 408.600 553.050 409.050 ;
        RECT 610.950 408.600 613.050 409.050 ;
        RECT 550.950 407.400 613.050 408.600 ;
        RECT 550.950 406.950 553.050 407.400 ;
        RECT 610.950 406.950 613.050 407.400 ;
        RECT 616.950 408.600 619.050 409.050 ;
        RECT 634.950 408.600 637.050 409.050 ;
        RECT 616.950 407.400 637.050 408.600 ;
        RECT 616.950 406.950 619.050 407.400 ;
        RECT 634.950 406.950 637.050 407.400 ;
        RECT 658.950 408.600 661.050 409.050 ;
        RECT 679.950 408.600 682.050 409.050 ;
        RECT 736.950 408.600 739.050 409.050 ;
        RECT 658.950 407.400 739.050 408.600 ;
        RECT 658.950 406.950 661.050 407.400 ;
        RECT 679.950 406.950 682.050 407.400 ;
        RECT 736.950 406.950 739.050 407.400 ;
        RECT 517.950 405.600 520.050 406.050 ;
        RECT 500.400 404.400 520.050 405.600 ;
        RECT 517.950 403.950 520.050 404.400 ;
        RECT 538.950 405.600 541.050 406.050 ;
        RECT 568.950 405.600 571.050 406.050 ;
        RECT 538.950 404.400 571.050 405.600 ;
        RECT 538.950 403.950 541.050 404.400 ;
        RECT 568.950 403.950 571.050 404.400 ;
        RECT 586.950 405.600 589.050 406.050 ;
        RECT 607.950 405.600 610.050 406.050 ;
        RECT 586.950 404.400 610.050 405.600 ;
        RECT 586.950 403.950 589.050 404.400 ;
        RECT 607.950 403.950 610.050 404.400 ;
        RECT 613.950 405.600 616.050 406.050 ;
        RECT 619.950 405.600 622.050 406.050 ;
        RECT 613.950 404.400 622.050 405.600 ;
        RECT 613.950 403.950 616.050 404.400 ;
        RECT 619.950 403.950 622.050 404.400 ;
        RECT 781.950 405.600 784.050 406.050 ;
        RECT 802.950 405.600 805.050 406.050 ;
        RECT 781.950 404.400 805.050 405.600 ;
        RECT 781.950 403.950 784.050 404.400 ;
        RECT 802.950 403.950 805.050 404.400 ;
        RECT 829.950 405.600 832.050 406.050 ;
        RECT 847.950 405.600 850.050 406.050 ;
        RECT 829.950 404.400 850.050 405.600 ;
        RECT 829.950 403.950 832.050 404.400 ;
        RECT 847.950 403.950 850.050 404.400 ;
        RECT 79.950 402.600 82.050 403.050 ;
        RECT 100.950 402.600 103.050 403.050 ;
        RECT 79.950 401.400 103.050 402.600 ;
        RECT 79.950 400.950 82.050 401.400 ;
        RECT 100.950 400.950 103.050 401.400 ;
        RECT 106.950 402.600 109.050 403.050 ;
        RECT 130.950 402.600 133.050 403.050 ;
        RECT 106.950 401.400 133.050 402.600 ;
        RECT 106.950 400.950 109.050 401.400 ;
        RECT 130.950 400.950 133.050 401.400 ;
        RECT 178.950 402.600 181.050 403.050 ;
        RECT 439.950 402.600 442.050 403.050 ;
        RECT 178.950 401.400 442.050 402.600 ;
        RECT 178.950 400.950 181.050 401.400 ;
        RECT 439.950 400.950 442.050 401.400 ;
        RECT 457.950 402.600 460.050 403.050 ;
        RECT 493.950 402.600 496.050 403.050 ;
        RECT 457.950 401.400 496.050 402.600 ;
        RECT 457.950 400.950 460.050 401.400 ;
        RECT 493.950 400.950 496.050 401.400 ;
        RECT 496.950 402.600 499.050 403.050 ;
        RECT 508.950 402.600 511.050 403.050 ;
        RECT 496.950 401.400 511.050 402.600 ;
        RECT 496.950 400.950 499.050 401.400 ;
        RECT 508.950 400.950 511.050 401.400 ;
        RECT 520.950 402.600 523.050 403.050 ;
        RECT 532.950 402.600 535.050 403.050 ;
        RECT 544.950 402.600 547.050 403.050 ;
        RECT 520.950 401.400 547.050 402.600 ;
        RECT 520.950 400.950 523.050 401.400 ;
        RECT 532.950 400.950 535.050 401.400 ;
        RECT 544.950 400.950 547.050 401.400 ;
        RECT 553.950 402.600 556.050 403.050 ;
        RECT 598.950 402.600 601.050 403.050 ;
        RECT 553.950 401.400 601.050 402.600 ;
        RECT 553.950 400.950 556.050 401.400 ;
        RECT 598.950 400.950 601.050 401.400 ;
        RECT 682.950 402.600 685.050 403.050 ;
        RECT 721.950 402.600 724.050 403.050 ;
        RECT 757.950 402.600 760.050 403.050 ;
        RECT 778.950 402.600 781.050 403.050 ;
        RECT 814.950 402.600 817.050 403.050 ;
        RECT 841.950 402.600 844.050 403.050 ;
        RECT 682.950 401.400 844.050 402.600 ;
        RECT 682.950 400.950 685.050 401.400 ;
        RECT 721.950 400.950 724.050 401.400 ;
        RECT 757.950 400.950 760.050 401.400 ;
        RECT 778.950 400.950 781.050 401.400 ;
        RECT 814.950 400.950 817.050 401.400 ;
        RECT 841.950 400.950 844.050 401.400 ;
        RECT 25.950 399.600 28.050 400.050 ;
        RECT 40.950 399.600 43.050 400.050 ;
        RECT 52.950 399.600 55.050 400.050 ;
        RECT 94.950 399.600 97.050 400.050 ;
        RECT 25.950 398.400 97.050 399.600 ;
        RECT 25.950 397.950 28.050 398.400 ;
        RECT 40.950 397.950 43.050 398.400 ;
        RECT 52.950 397.950 55.050 398.400 ;
        RECT 94.950 397.950 97.050 398.400 ;
        RECT 184.950 399.600 187.050 400.050 ;
        RECT 202.950 399.600 205.050 400.050 ;
        RECT 238.950 399.600 241.050 400.050 ;
        RECT 265.950 399.600 268.050 400.050 ;
        RECT 286.950 399.600 289.050 400.050 ;
        RECT 184.950 398.400 252.600 399.600 ;
        RECT 184.950 397.950 187.050 398.400 ;
        RECT 202.950 397.950 205.050 398.400 ;
        RECT 238.950 397.950 241.050 398.400 ;
        RECT 235.950 396.600 238.050 397.050 ;
        RECT 247.950 396.600 250.050 397.050 ;
        RECT 235.950 395.400 250.050 396.600 ;
        RECT 251.400 396.600 252.600 398.400 ;
        RECT 265.950 398.400 289.050 399.600 ;
        RECT 265.950 397.950 268.050 398.400 ;
        RECT 286.950 397.950 289.050 398.400 ;
        RECT 313.950 399.600 316.050 400.050 ;
        RECT 475.950 399.600 478.050 400.050 ;
        RECT 313.950 398.400 478.050 399.600 ;
        RECT 313.950 397.950 316.050 398.400 ;
        RECT 475.950 397.950 478.050 398.400 ;
        RECT 499.950 399.600 502.050 400.050 ;
        RECT 505.950 399.600 508.050 400.050 ;
        RECT 499.950 398.400 508.050 399.600 ;
        RECT 499.950 397.950 502.050 398.400 ;
        RECT 505.950 397.950 508.050 398.400 ;
        RECT 520.950 399.600 523.050 400.050 ;
        RECT 529.950 399.600 532.050 400.050 ;
        RECT 520.950 398.400 532.050 399.600 ;
        RECT 520.950 397.950 523.050 398.400 ;
        RECT 529.950 397.950 532.050 398.400 ;
        RECT 535.950 399.600 538.050 400.050 ;
        RECT 595.950 399.600 598.050 400.050 ;
        RECT 676.950 399.600 679.050 400.050 ;
        RECT 535.950 398.400 582.600 399.600 ;
        RECT 535.950 397.950 538.050 398.400 ;
        RECT 574.950 396.600 577.050 397.050 ;
        RECT 251.400 395.400 577.050 396.600 ;
        RECT 581.400 396.600 582.600 398.400 ;
        RECT 595.950 398.400 679.050 399.600 ;
        RECT 595.950 397.950 598.050 398.400 ;
        RECT 676.950 397.950 679.050 398.400 ;
        RECT 592.950 396.600 595.050 397.050 ;
        RECT 581.400 395.400 595.050 396.600 ;
        RECT 235.950 394.950 238.050 395.400 ;
        RECT 247.950 394.950 250.050 395.400 ;
        RECT 574.950 394.950 577.050 395.400 ;
        RECT 592.950 394.950 595.050 395.400 ;
        RECT 235.950 393.600 238.050 394.050 ;
        RECT 286.950 393.600 289.050 394.050 ;
        RECT 376.950 393.600 379.050 394.050 ;
        RECT 574.950 393.600 577.050 394.050 ;
        RECT 685.950 393.600 688.050 394.050 ;
        RECT 235.950 392.400 688.050 393.600 ;
        RECT 235.950 391.950 238.050 392.400 ;
        RECT 286.950 391.950 289.050 392.400 ;
        RECT 376.950 391.950 379.050 392.400 ;
        RECT 574.950 391.950 577.050 392.400 ;
        RECT 685.950 391.950 688.050 392.400 ;
        RECT 22.950 390.600 25.050 391.050 ;
        RECT 55.950 390.600 58.050 391.050 ;
        RECT 22.950 389.400 58.050 390.600 ;
        RECT 22.950 388.950 25.050 389.400 ;
        RECT 55.950 388.950 58.050 389.400 ;
        RECT 118.950 390.600 121.050 391.050 ;
        RECT 148.950 390.600 151.050 391.050 ;
        RECT 118.950 389.400 151.050 390.600 ;
        RECT 118.950 388.950 121.050 389.400 ;
        RECT 148.950 388.950 151.050 389.400 ;
        RECT 175.950 390.600 178.050 391.050 ;
        RECT 247.950 390.600 250.050 391.050 ;
        RECT 253.950 390.600 256.050 391.050 ;
        RECT 175.950 389.400 246.600 390.600 ;
        RECT 175.950 388.950 178.050 389.400 ;
        RECT 34.950 387.600 37.050 388.050 ;
        RECT 70.950 387.600 73.050 388.050 ;
        RECT 79.950 387.600 82.050 388.050 ;
        RECT 34.950 386.400 82.050 387.600 ;
        RECT 34.950 385.950 37.050 386.400 ;
        RECT 70.950 385.950 73.050 386.400 ;
        RECT 79.950 385.950 82.050 386.400 ;
        RECT 97.950 387.600 100.050 388.050 ;
        RECT 112.950 387.600 115.050 388.050 ;
        RECT 130.950 387.600 133.050 388.050 ;
        RECT 97.950 386.400 133.050 387.600 ;
        RECT 97.950 385.950 100.050 386.400 ;
        RECT 112.950 385.950 115.050 386.400 ;
        RECT 130.950 385.950 133.050 386.400 ;
        RECT 163.950 387.600 166.050 388.050 ;
        RECT 175.950 387.600 178.050 388.050 ;
        RECT 163.950 386.400 178.050 387.600 ;
        RECT 245.400 387.600 246.600 389.400 ;
        RECT 247.950 389.400 256.050 390.600 ;
        RECT 247.950 388.950 250.050 389.400 ;
        RECT 253.950 388.950 256.050 389.400 ;
        RECT 277.950 390.600 280.050 391.050 ;
        RECT 289.950 390.600 292.050 391.050 ;
        RECT 277.950 389.400 292.050 390.600 ;
        RECT 277.950 388.950 280.050 389.400 ;
        RECT 289.950 388.950 292.050 389.400 ;
        RECT 328.950 390.600 331.050 391.050 ;
        RECT 346.950 390.600 349.050 391.050 ;
        RECT 361.950 390.600 364.050 391.050 ;
        RECT 328.950 389.400 364.050 390.600 ;
        RECT 328.950 388.950 331.050 389.400 ;
        RECT 346.950 388.950 349.050 389.400 ;
        RECT 361.950 388.950 364.050 389.400 ;
        RECT 385.950 390.600 388.050 391.050 ;
        RECT 391.950 390.600 394.050 391.050 ;
        RECT 385.950 389.400 394.050 390.600 ;
        RECT 385.950 388.950 388.050 389.400 ;
        RECT 391.950 388.950 394.050 389.400 ;
        RECT 394.950 390.600 397.050 391.050 ;
        RECT 445.950 390.600 448.050 391.050 ;
        RECT 394.950 389.400 448.050 390.600 ;
        RECT 394.950 388.950 397.050 389.400 ;
        RECT 445.950 388.950 448.050 389.400 ;
        RECT 448.950 390.600 451.050 391.050 ;
        RECT 478.950 390.600 481.050 391.050 ;
        RECT 448.950 389.400 481.050 390.600 ;
        RECT 448.950 388.950 451.050 389.400 ;
        RECT 478.950 388.950 481.050 389.400 ;
        RECT 484.950 390.600 487.050 391.050 ;
        RECT 694.950 390.600 697.050 391.050 ;
        RECT 484.950 389.400 697.050 390.600 ;
        RECT 484.950 388.950 487.050 389.400 ;
        RECT 694.950 388.950 697.050 389.400 ;
        RECT 295.950 387.600 298.050 388.050 ;
        RECT 245.400 386.400 298.050 387.600 ;
        RECT 163.950 385.950 166.050 386.400 ;
        RECT 175.950 385.950 178.050 386.400 ;
        RECT 295.950 385.950 298.050 386.400 ;
        RECT 307.950 387.600 310.050 388.050 ;
        RECT 340.950 387.600 343.050 388.050 ;
        RECT 307.950 386.400 343.050 387.600 ;
        RECT 307.950 385.950 310.050 386.400 ;
        RECT 340.950 385.950 343.050 386.400 ;
        RECT 352.950 387.600 355.050 388.050 ;
        RECT 382.950 387.600 385.050 388.050 ;
        RECT 352.950 386.400 385.050 387.600 ;
        RECT 352.950 385.950 355.050 386.400 ;
        RECT 382.950 385.950 385.050 386.400 ;
        RECT 406.950 387.600 409.050 388.050 ;
        RECT 415.950 387.600 418.050 388.050 ;
        RECT 556.950 387.600 559.050 388.050 ;
        RECT 406.950 386.400 411.600 387.600 ;
        RECT 406.950 385.950 409.050 386.400 ;
        RECT 58.950 384.600 61.050 385.050 ;
        RECT 100.950 384.600 103.050 385.050 ;
        RECT 47.400 383.400 61.050 384.600 ;
        RECT 25.950 381.600 28.050 382.050 ;
        RECT 43.950 381.600 46.050 382.050 ;
        RECT 47.400 381.600 48.600 383.400 ;
        RECT 58.950 382.950 61.050 383.400 ;
        RECT 98.400 383.400 103.050 384.600 ;
        RECT 25.950 380.400 48.600 381.600 ;
        RECT 49.950 381.600 52.050 382.050 ;
        RECT 55.950 381.600 58.050 382.050 ;
        RECT 64.950 381.600 67.050 382.050 ;
        RECT 49.950 380.400 67.050 381.600 ;
        RECT 25.950 379.950 28.050 380.400 ;
        RECT 43.950 379.950 46.050 380.400 ;
        RECT 49.950 379.950 52.050 380.400 ;
        RECT 55.950 379.950 58.050 380.400 ;
        RECT 64.950 379.950 67.050 380.400 ;
        RECT 82.950 381.600 85.050 382.050 ;
        RECT 98.400 381.600 99.600 383.400 ;
        RECT 100.950 382.950 103.050 383.400 ;
        RECT 121.950 384.600 124.050 385.050 ;
        RECT 145.950 384.600 148.050 385.050 ;
        RECT 163.950 384.600 166.050 385.050 ;
        RECT 121.950 383.400 148.050 384.600 ;
        RECT 121.950 382.950 124.050 383.400 ;
        RECT 145.950 382.950 148.050 383.400 ;
        RECT 149.400 383.400 166.050 384.600 ;
        RECT 82.950 380.400 99.600 381.600 ;
        RECT 109.950 381.600 112.050 382.050 ;
        RECT 115.950 381.600 118.050 382.050 ;
        RECT 109.950 380.400 118.050 381.600 ;
        RECT 82.950 379.950 85.050 380.400 ;
        RECT 109.950 379.950 112.050 380.400 ;
        RECT 115.950 379.950 118.050 380.400 ;
        RECT 130.950 381.600 133.050 382.050 ;
        RECT 136.950 381.600 139.050 382.050 ;
        RECT 130.950 380.400 139.050 381.600 ;
        RECT 130.950 379.950 133.050 380.400 ;
        RECT 136.950 379.950 139.050 380.400 ;
        RECT 139.950 381.600 142.050 382.050 ;
        RECT 149.400 381.600 150.600 383.400 ;
        RECT 163.950 382.950 166.050 383.400 ;
        RECT 211.950 384.600 214.050 385.050 ;
        RECT 253.950 384.600 256.050 385.050 ;
        RECT 211.950 383.400 256.050 384.600 ;
        RECT 211.950 382.950 214.050 383.400 ;
        RECT 253.950 382.950 256.050 383.400 ;
        RECT 271.950 384.600 274.050 385.050 ;
        RECT 280.950 384.600 283.050 385.050 ;
        RECT 271.950 383.400 283.050 384.600 ;
        RECT 271.950 382.950 274.050 383.400 ;
        RECT 280.950 382.950 283.050 383.400 ;
        RECT 301.950 382.950 304.050 385.050 ;
        RECT 319.950 384.600 322.050 385.050 ;
        RECT 334.950 384.600 337.050 385.050 ;
        RECT 319.950 383.400 337.050 384.600 ;
        RECT 319.950 382.950 322.050 383.400 ;
        RECT 334.950 382.950 337.050 383.400 ;
        RECT 355.950 384.600 358.050 385.050 ;
        RECT 364.950 384.600 367.050 385.050 ;
        RECT 355.950 383.400 367.050 384.600 ;
        RECT 355.950 382.950 358.050 383.400 ;
        RECT 364.950 382.950 367.050 383.400 ;
        RECT 391.950 384.600 394.050 385.050 ;
        RECT 400.950 384.600 403.050 385.050 ;
        RECT 406.950 384.600 409.050 385.050 ;
        RECT 391.950 383.400 403.050 384.600 ;
        RECT 391.950 382.950 394.050 383.400 ;
        RECT 400.950 382.950 403.050 383.400 ;
        RECT 404.400 383.400 409.050 384.600 ;
        RECT 139.950 380.400 150.600 381.600 ;
        RECT 166.950 381.600 169.050 382.050 ;
        RECT 178.950 381.600 181.050 382.050 ;
        RECT 166.950 380.400 181.050 381.600 ;
        RECT 139.950 379.950 142.050 380.400 ;
        RECT 166.950 379.950 169.050 380.400 ;
        RECT 178.950 379.950 181.050 380.400 ;
        RECT 184.950 381.600 187.050 382.050 ;
        RECT 211.950 381.600 214.050 382.050 ;
        RECT 184.950 380.400 214.050 381.600 ;
        RECT 184.950 379.950 187.050 380.400 ;
        RECT 211.950 379.950 214.050 380.400 ;
        RECT 229.950 381.600 232.050 382.050 ;
        RECT 241.950 381.600 244.050 382.050 ;
        RECT 229.950 380.400 244.050 381.600 ;
        RECT 229.950 379.950 232.050 380.400 ;
        RECT 241.950 379.950 244.050 380.400 ;
        RECT 262.950 381.600 265.050 382.050 ;
        RECT 268.950 381.600 271.050 382.050 ;
        RECT 262.950 380.400 271.050 381.600 ;
        RECT 262.950 379.950 265.050 380.400 ;
        RECT 268.950 379.950 271.050 380.400 ;
        RECT 16.950 378.600 19.050 379.050 ;
        RECT 25.950 378.600 28.050 379.050 ;
        RECT 16.950 377.400 28.050 378.600 ;
        RECT 16.950 376.950 19.050 377.400 ;
        RECT 25.950 376.950 28.050 377.400 ;
        RECT 40.950 378.600 43.050 379.050 ;
        RECT 52.950 378.600 55.050 379.050 ;
        RECT 61.950 378.600 64.050 379.050 ;
        RECT 40.950 377.400 64.050 378.600 ;
        RECT 40.950 376.950 43.050 377.400 ;
        RECT 52.950 376.950 55.050 377.400 ;
        RECT 61.950 376.950 64.050 377.400 ;
        RECT 145.950 378.600 148.050 379.050 ;
        RECT 154.950 378.600 157.050 379.050 ;
        RECT 145.950 377.400 157.050 378.600 ;
        RECT 145.950 376.950 148.050 377.400 ;
        RECT 154.950 376.950 157.050 377.400 ;
        RECT 190.950 378.600 193.050 379.050 ;
        RECT 202.950 378.600 205.050 379.050 ;
        RECT 190.950 377.400 205.050 378.600 ;
        RECT 190.950 376.950 193.050 377.400 ;
        RECT 202.950 376.950 205.050 377.400 ;
        RECT 226.950 378.600 229.050 379.050 ;
        RECT 232.950 378.600 235.050 379.050 ;
        RECT 226.950 377.400 235.050 378.600 ;
        RECT 226.950 376.950 229.050 377.400 ;
        RECT 232.950 376.950 235.050 377.400 ;
        RECT 244.950 378.600 247.050 379.050 ;
        RECT 298.950 378.600 301.050 379.050 ;
        RECT 244.950 377.400 301.050 378.600 ;
        RECT 302.400 378.600 303.600 382.950 ;
        RECT 304.950 381.600 307.050 382.050 ;
        RECT 313.950 381.600 316.050 382.050 ;
        RECT 304.950 380.400 316.050 381.600 ;
        RECT 304.950 379.950 307.050 380.400 ;
        RECT 313.950 379.950 316.050 380.400 ;
        RECT 316.950 381.600 319.050 382.050 ;
        RECT 322.950 381.600 325.050 382.050 ;
        RECT 349.950 381.600 352.050 382.050 ;
        RECT 316.950 380.400 321.600 381.600 ;
        RECT 316.950 379.950 319.050 380.400 ;
        RECT 316.950 378.600 319.050 379.050 ;
        RECT 302.400 377.400 319.050 378.600 ;
        RECT 320.400 378.600 321.600 380.400 ;
        RECT 322.950 380.400 352.050 381.600 ;
        RECT 322.950 379.950 325.050 380.400 ;
        RECT 349.950 379.950 352.050 380.400 ;
        RECT 373.950 381.600 376.050 382.050 ;
        RECT 388.950 381.600 391.050 382.050 ;
        RECT 404.400 381.600 405.600 383.400 ;
        RECT 406.950 382.950 409.050 383.400 ;
        RECT 410.400 381.600 411.600 386.400 ;
        RECT 415.950 386.400 559.050 387.600 ;
        RECT 415.950 385.950 418.050 386.400 ;
        RECT 556.950 385.950 559.050 386.400 ;
        RECT 562.950 387.600 565.050 388.050 ;
        RECT 571.950 387.600 574.050 388.050 ;
        RECT 562.950 386.400 574.050 387.600 ;
        RECT 562.950 385.950 565.050 386.400 ;
        RECT 571.950 385.950 574.050 386.400 ;
        RECT 577.950 387.600 580.050 388.050 ;
        RECT 586.950 387.600 589.050 388.050 ;
        RECT 577.950 386.400 589.050 387.600 ;
        RECT 577.950 385.950 580.050 386.400 ;
        RECT 586.950 385.950 589.050 386.400 ;
        RECT 424.950 384.600 427.050 385.050 ;
        RECT 463.950 384.600 466.050 385.050 ;
        RECT 472.950 384.600 475.050 385.050 ;
        RECT 424.950 383.400 432.600 384.600 ;
        RECT 424.950 382.950 427.050 383.400 ;
        RECT 431.400 382.050 432.600 383.400 ;
        RECT 463.950 383.400 475.050 384.600 ;
        RECT 463.950 382.950 466.050 383.400 ;
        RECT 472.950 382.950 475.050 383.400 ;
        RECT 478.950 384.600 481.050 385.050 ;
        RECT 490.950 384.600 493.050 385.050 ;
        RECT 478.950 383.400 493.050 384.600 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 490.950 382.950 493.050 383.400 ;
        RECT 505.950 384.600 508.050 385.050 ;
        RECT 520.950 384.600 523.050 385.050 ;
        RECT 505.950 383.400 523.050 384.600 ;
        RECT 505.950 382.950 508.050 383.400 ;
        RECT 520.950 382.950 523.050 383.400 ;
        RECT 547.950 384.600 550.050 385.050 ;
        RECT 547.950 383.400 561.600 384.600 ;
        RECT 547.950 382.950 550.050 383.400 ;
        RECT 373.950 380.400 391.050 381.600 ;
        RECT 373.950 379.950 376.050 380.400 ;
        RECT 388.950 379.950 391.050 380.400 ;
        RECT 392.400 380.400 405.600 381.600 ;
        RECT 407.400 380.400 411.600 381.600 ;
        RECT 421.950 381.600 424.050 382.050 ;
        RECT 427.950 381.600 430.050 382.050 ;
        RECT 421.950 380.400 430.050 381.600 ;
        RECT 325.950 378.600 328.050 379.050 ;
        RECT 343.950 378.600 346.050 379.050 ;
        RECT 320.400 377.400 324.600 378.600 ;
        RECT 244.950 376.950 247.050 377.400 ;
        RECT 298.950 376.950 301.050 377.400 ;
        RECT 316.950 376.950 319.050 377.400 ;
        RECT 323.400 376.050 324.600 377.400 ;
        RECT 325.950 377.400 346.050 378.600 ;
        RECT 325.950 376.950 328.050 377.400 ;
        RECT 343.950 376.950 346.050 377.400 ;
        RECT 352.950 378.600 355.050 379.050 ;
        RECT 358.950 378.600 361.050 379.050 ;
        RECT 352.950 377.400 361.050 378.600 ;
        RECT 352.950 376.950 355.050 377.400 ;
        RECT 358.950 376.950 361.050 377.400 ;
        RECT 364.950 378.600 367.050 379.050 ;
        RECT 370.950 378.600 373.050 379.050 ;
        RECT 364.950 377.400 373.050 378.600 ;
        RECT 364.950 376.950 367.050 377.400 ;
        RECT 370.950 376.950 373.050 377.400 ;
        RECT 373.950 378.600 376.050 379.050 ;
        RECT 392.400 378.600 393.600 380.400 ;
        RECT 407.400 379.050 408.600 380.400 ;
        RECT 421.950 379.950 424.050 380.400 ;
        RECT 427.950 379.950 430.050 380.400 ;
        RECT 430.950 379.950 433.050 382.050 ;
        RECT 439.950 381.600 442.050 382.050 ;
        RECT 445.950 381.600 448.050 382.050 ;
        RECT 439.950 380.400 448.050 381.600 ;
        RECT 439.950 379.950 442.050 380.400 ;
        RECT 445.950 379.950 448.050 380.400 ;
        RECT 454.950 381.600 457.050 382.050 ;
        RECT 454.950 380.400 489.600 381.600 ;
        RECT 454.950 379.950 457.050 380.400 ;
        RECT 488.400 379.050 489.600 380.400 ;
        RECT 560.400 379.050 561.600 383.400 ;
        RECT 583.950 382.950 586.050 385.050 ;
        RECT 568.950 381.600 571.050 382.050 ;
        RECT 577.950 381.600 580.050 382.050 ;
        RECT 568.950 380.400 580.050 381.600 ;
        RECT 584.400 381.600 585.600 382.950 ;
        RECT 586.950 381.600 589.050 382.050 ;
        RECT 584.400 380.400 589.050 381.600 ;
        RECT 568.950 379.950 571.050 380.400 ;
        RECT 577.950 379.950 580.050 380.400 ;
        RECT 586.950 379.950 589.050 380.400 ;
        RECT 610.950 381.600 613.050 382.050 ;
        RECT 637.950 381.600 640.050 382.050 ;
        RECT 784.950 381.600 787.050 382.050 ;
        RECT 610.950 380.400 787.050 381.600 ;
        RECT 610.950 379.950 613.050 380.400 ;
        RECT 637.950 379.950 640.050 380.400 ;
        RECT 784.950 379.950 787.050 380.400 ;
        RECT 838.950 381.600 841.050 382.050 ;
        RECT 856.950 381.600 859.050 382.050 ;
        RECT 838.950 380.400 859.050 381.600 ;
        RECT 838.950 379.950 841.050 380.400 ;
        RECT 856.950 379.950 859.050 380.400 ;
        RECT 373.950 377.400 393.600 378.600 ;
        RECT 373.950 376.950 376.050 377.400 ;
        RECT 406.950 376.950 409.050 379.050 ;
        RECT 472.950 378.600 475.050 379.050 ;
        RECT 481.950 378.600 484.050 379.050 ;
        RECT 472.950 377.400 484.050 378.600 ;
        RECT 472.950 376.950 475.050 377.400 ;
        RECT 481.950 376.950 484.050 377.400 ;
        RECT 487.950 376.950 490.050 379.050 ;
        RECT 490.950 378.600 493.050 379.050 ;
        RECT 502.950 378.600 505.050 379.050 ;
        RECT 490.950 377.400 505.050 378.600 ;
        RECT 490.950 376.950 493.050 377.400 ;
        RECT 502.950 376.950 505.050 377.400 ;
        RECT 508.950 376.950 511.050 379.050 ;
        RECT 514.950 378.600 517.050 379.050 ;
        RECT 541.950 378.600 544.050 379.050 ;
        RECT 514.950 377.400 555.600 378.600 ;
        RECT 514.950 376.950 517.050 377.400 ;
        RECT 541.950 376.950 544.050 377.400 ;
        RECT 181.950 375.600 184.050 376.050 ;
        RECT 199.950 375.600 202.050 376.050 ;
        RECT 220.950 375.600 223.050 376.050 ;
        RECT 181.950 374.400 223.050 375.600 ;
        RECT 181.950 373.950 184.050 374.400 ;
        RECT 199.950 373.950 202.050 374.400 ;
        RECT 220.950 373.950 223.050 374.400 ;
        RECT 229.950 375.600 232.050 376.050 ;
        RECT 235.950 375.600 238.050 376.050 ;
        RECT 229.950 374.400 238.050 375.600 ;
        RECT 229.950 373.950 232.050 374.400 ;
        RECT 235.950 373.950 238.050 374.400 ;
        RECT 256.950 375.600 259.050 376.050 ;
        RECT 268.950 375.600 271.050 376.050 ;
        RECT 256.950 374.400 271.050 375.600 ;
        RECT 256.950 373.950 259.050 374.400 ;
        RECT 268.950 373.950 271.050 374.400 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 364.950 375.600 367.050 376.050 ;
        RECT 367.950 375.600 370.050 376.050 ;
        RECT 412.950 375.600 415.050 376.050 ;
        RECT 364.950 374.400 415.050 375.600 ;
        RECT 364.950 373.950 367.050 374.400 ;
        RECT 367.950 373.950 370.050 374.400 ;
        RECT 412.950 373.950 415.050 374.400 ;
        RECT 475.950 375.600 478.050 376.050 ;
        RECT 481.950 375.600 484.050 376.050 ;
        RECT 502.950 375.600 505.050 376.050 ;
        RECT 475.950 374.400 484.050 375.600 ;
        RECT 475.950 373.950 478.050 374.400 ;
        RECT 481.950 373.950 484.050 374.400 ;
        RECT 485.400 374.400 505.050 375.600 ;
        RECT 509.400 375.600 510.600 376.950 ;
        RECT 526.950 375.600 529.050 376.050 ;
        RECT 550.950 375.600 553.050 376.050 ;
        RECT 509.400 374.400 553.050 375.600 ;
        RECT 554.400 375.600 555.600 377.400 ;
        RECT 559.950 376.950 562.050 379.050 ;
        RECT 562.950 378.600 565.050 379.050 ;
        RECT 568.950 378.600 571.050 379.050 ;
        RECT 562.950 377.400 571.050 378.600 ;
        RECT 562.950 376.950 565.050 377.400 ;
        RECT 568.950 376.950 571.050 377.400 ;
        RECT 577.950 378.600 580.050 379.050 ;
        RECT 604.950 378.600 607.050 379.050 ;
        RECT 577.950 377.400 607.050 378.600 ;
        RECT 577.950 376.950 580.050 377.400 ;
        RECT 604.950 376.950 607.050 377.400 ;
        RECT 571.950 375.600 574.050 376.050 ;
        RECT 554.400 374.400 574.050 375.600 ;
        RECT 232.950 372.600 235.050 373.050 ;
        RECT 259.950 372.600 262.050 373.050 ;
        RECT 268.950 372.600 271.050 373.050 ;
        RECT 274.950 372.600 277.050 373.050 ;
        RECT 283.950 372.600 286.050 373.050 ;
        RECT 337.950 372.600 340.050 373.050 ;
        RECT 232.950 371.400 264.600 372.600 ;
        RECT 268.950 371.400 277.050 372.600 ;
        RECT 232.950 370.950 235.050 371.400 ;
        RECT 259.950 370.950 262.050 371.400 ;
        RECT 268.950 370.950 271.050 371.400 ;
        RECT 274.950 370.950 277.050 371.400 ;
        RECT 278.400 371.400 340.050 372.600 ;
        RECT 223.950 369.600 226.050 370.050 ;
        RECT 253.950 369.600 256.050 370.050 ;
        RECT 223.950 368.400 256.050 369.600 ;
        RECT 223.950 367.950 226.050 368.400 ;
        RECT 253.950 367.950 256.050 368.400 ;
        RECT 259.950 369.600 262.050 370.050 ;
        RECT 278.400 369.600 279.600 371.400 ;
        RECT 283.950 370.950 286.050 371.400 ;
        RECT 337.950 370.950 340.050 371.400 ;
        RECT 349.950 372.600 352.050 373.050 ;
        RECT 373.950 372.600 376.050 373.050 ;
        RECT 349.950 371.400 376.050 372.600 ;
        RECT 349.950 370.950 352.050 371.400 ;
        RECT 373.950 370.950 376.050 371.400 ;
        RECT 388.950 372.600 391.050 373.050 ;
        RECT 403.950 372.600 406.050 373.050 ;
        RECT 388.950 371.400 406.050 372.600 ;
        RECT 388.950 370.950 391.050 371.400 ;
        RECT 403.950 370.950 406.050 371.400 ;
        RECT 478.950 372.600 481.050 373.050 ;
        RECT 485.400 372.600 486.600 374.400 ;
        RECT 502.950 373.950 505.050 374.400 ;
        RECT 526.950 373.950 529.050 374.400 ;
        RECT 550.950 373.950 553.050 374.400 ;
        RECT 571.950 373.950 574.050 374.400 ;
        RECT 589.950 375.600 592.050 376.050 ;
        RECT 667.950 375.600 670.050 376.050 ;
        RECT 589.950 374.400 670.050 375.600 ;
        RECT 589.950 373.950 592.050 374.400 ;
        RECT 667.950 373.950 670.050 374.400 ;
        RECT 478.950 371.400 486.600 372.600 ;
        RECT 499.950 372.600 502.050 373.050 ;
        RECT 520.950 372.600 523.050 373.050 ;
        RECT 499.950 371.400 523.050 372.600 ;
        RECT 478.950 370.950 481.050 371.400 ;
        RECT 499.950 370.950 502.050 371.400 ;
        RECT 520.950 370.950 523.050 371.400 ;
        RECT 535.950 372.600 538.050 373.050 ;
        RECT 547.950 372.600 550.050 373.050 ;
        RECT 535.950 371.400 550.050 372.600 ;
        RECT 535.950 370.950 538.050 371.400 ;
        RECT 547.950 370.950 550.050 371.400 ;
        RECT 565.950 372.600 568.050 373.050 ;
        RECT 601.950 372.600 604.050 373.050 ;
        RECT 565.950 371.400 604.050 372.600 ;
        RECT 565.950 370.950 568.050 371.400 ;
        RECT 601.950 370.950 604.050 371.400 ;
        RECT 667.950 372.600 670.050 373.050 ;
        RECT 778.950 372.600 781.050 373.050 ;
        RECT 667.950 371.400 781.050 372.600 ;
        RECT 667.950 370.950 670.050 371.400 ;
        RECT 778.950 370.950 781.050 371.400 ;
        RECT 259.950 368.400 279.600 369.600 ;
        RECT 280.950 369.600 283.050 370.050 ;
        RECT 331.950 369.600 334.050 370.050 ;
        RECT 280.950 368.400 334.050 369.600 ;
        RECT 259.950 367.950 262.050 368.400 ;
        RECT 280.950 367.950 283.050 368.400 ;
        RECT 331.950 367.950 334.050 368.400 ;
        RECT 334.950 369.600 337.050 370.050 ;
        RECT 460.950 369.600 463.050 370.050 ;
        RECT 334.950 368.400 463.050 369.600 ;
        RECT 334.950 367.950 337.050 368.400 ;
        RECT 460.950 367.950 463.050 368.400 ;
        RECT 493.950 369.600 496.050 370.050 ;
        RECT 514.950 369.600 517.050 370.050 ;
        RECT 493.950 368.400 517.050 369.600 ;
        RECT 493.950 367.950 496.050 368.400 ;
        RECT 514.950 367.950 517.050 368.400 ;
        RECT 676.950 369.600 679.050 370.050 ;
        RECT 724.950 369.600 727.050 370.050 ;
        RECT 676.950 368.400 727.050 369.600 ;
        RECT 676.950 367.950 679.050 368.400 ;
        RECT 724.950 367.950 727.050 368.400 ;
        RECT 22.950 366.600 25.050 367.050 ;
        RECT 37.950 366.600 40.050 367.050 ;
        RECT 22.950 365.400 40.050 366.600 ;
        RECT 22.950 364.950 25.050 365.400 ;
        RECT 37.950 364.950 40.050 365.400 ;
        RECT 112.950 366.600 115.050 367.050 ;
        RECT 133.950 366.600 136.050 367.050 ;
        RECT 112.950 365.400 136.050 366.600 ;
        RECT 112.950 364.950 115.050 365.400 ;
        RECT 133.950 364.950 136.050 365.400 ;
        RECT 178.950 366.600 181.050 367.050 ;
        RECT 280.950 366.600 283.050 367.050 ;
        RECT 415.950 366.600 418.050 367.050 ;
        RECT 508.950 366.600 511.050 367.050 ;
        RECT 178.950 365.400 283.050 366.600 ;
        RECT 178.950 364.950 181.050 365.400 ;
        RECT 280.950 364.950 283.050 365.400 ;
        RECT 311.400 365.400 418.050 366.600 ;
        RECT 148.950 363.600 151.050 364.050 ;
        RECT 311.400 363.600 312.600 365.400 ;
        RECT 415.950 364.950 418.050 365.400 ;
        RECT 476.400 365.400 511.050 366.600 ;
        RECT 148.950 362.400 312.600 363.600 ;
        RECT 313.950 363.600 316.050 364.050 ;
        RECT 382.950 363.600 385.050 364.050 ;
        RECT 313.950 362.400 385.050 363.600 ;
        RECT 148.950 361.950 151.050 362.400 ;
        RECT 313.950 361.950 316.050 362.400 ;
        RECT 382.950 361.950 385.050 362.400 ;
        RECT 451.950 363.600 454.050 364.050 ;
        RECT 476.400 363.600 477.600 365.400 ;
        RECT 508.950 364.950 511.050 365.400 ;
        RECT 646.950 366.600 649.050 367.050 ;
        RECT 661.950 366.600 664.050 367.050 ;
        RECT 670.950 366.600 673.050 367.050 ;
        RECT 646.950 365.400 673.050 366.600 ;
        RECT 646.950 364.950 649.050 365.400 ;
        RECT 661.950 364.950 664.050 365.400 ;
        RECT 670.950 364.950 673.050 365.400 ;
        RECT 745.950 366.600 748.050 367.050 ;
        RECT 769.950 366.600 772.050 367.050 ;
        RECT 745.950 365.400 772.050 366.600 ;
        RECT 745.950 364.950 748.050 365.400 ;
        RECT 769.950 364.950 772.050 365.400 ;
        RECT 451.950 362.400 477.600 363.600 ;
        RECT 478.950 363.600 481.050 364.050 ;
        RECT 571.950 363.600 574.050 364.050 ;
        RECT 811.950 363.600 814.050 364.050 ;
        RECT 478.950 362.400 561.600 363.600 ;
        RECT 451.950 361.950 454.050 362.400 ;
        RECT 478.950 361.950 481.050 362.400 ;
        RECT 163.950 360.600 166.050 361.050 ;
        RECT 424.950 360.600 427.050 361.050 ;
        RECT 163.950 359.400 427.050 360.600 ;
        RECT 163.950 358.950 166.050 359.400 ;
        RECT 424.950 358.950 427.050 359.400 ;
        RECT 487.950 360.600 490.050 361.050 ;
        RECT 550.950 360.600 553.050 361.050 ;
        RECT 487.950 359.400 553.050 360.600 ;
        RECT 560.400 360.600 561.600 362.400 ;
        RECT 571.950 362.400 814.050 363.600 ;
        RECT 571.950 361.950 574.050 362.400 ;
        RECT 811.950 361.950 814.050 362.400 ;
        RECT 613.950 360.600 616.050 361.050 ;
        RECT 661.950 360.600 664.050 361.050 ;
        RECT 703.950 360.600 706.050 361.050 ;
        RECT 718.950 360.600 721.050 361.050 ;
        RECT 560.400 359.400 721.050 360.600 ;
        RECT 487.950 358.950 490.050 359.400 ;
        RECT 550.950 358.950 553.050 359.400 ;
        RECT 613.950 358.950 616.050 359.400 ;
        RECT 661.950 358.950 664.050 359.400 ;
        RECT 703.950 358.950 706.050 359.400 ;
        RECT 718.950 358.950 721.050 359.400 ;
        RECT 217.950 357.600 220.050 358.050 ;
        RECT 295.950 357.600 298.050 358.050 ;
        RECT 217.950 356.400 298.050 357.600 ;
        RECT 217.950 355.950 220.050 356.400 ;
        RECT 295.950 355.950 298.050 356.400 ;
        RECT 325.950 357.600 328.050 358.050 ;
        RECT 355.950 357.600 358.050 358.050 ;
        RECT 325.950 356.400 358.050 357.600 ;
        RECT 325.950 355.950 328.050 356.400 ;
        RECT 355.950 355.950 358.050 356.400 ;
        RECT 463.950 357.600 466.050 358.050 ;
        RECT 544.950 357.600 547.050 358.050 ;
        RECT 463.950 356.400 547.050 357.600 ;
        RECT 463.950 355.950 466.050 356.400 ;
        RECT 544.950 355.950 547.050 356.400 ;
        RECT 547.950 357.600 550.050 358.050 ;
        RECT 553.950 357.600 556.050 358.050 ;
        RECT 547.950 356.400 556.050 357.600 ;
        RECT 547.950 355.950 550.050 356.400 ;
        RECT 553.950 355.950 556.050 356.400 ;
        RECT 691.950 357.600 694.050 358.050 ;
        RECT 811.950 357.600 814.050 358.050 ;
        RECT 823.950 357.600 826.050 358.050 ;
        RECT 691.950 356.400 826.050 357.600 ;
        RECT 691.950 355.950 694.050 356.400 ;
        RECT 811.950 355.950 814.050 356.400 ;
        RECT 823.950 355.950 826.050 356.400 ;
        RECT 244.950 354.600 247.050 355.050 ;
        RECT 262.950 354.600 265.050 355.050 ;
        RECT 319.950 354.600 322.050 355.050 ;
        RECT 244.950 353.400 252.600 354.600 ;
        RECT 244.950 352.950 247.050 353.400 ;
        RECT 208.950 351.600 211.050 352.050 ;
        RECT 247.950 351.600 250.050 352.050 ;
        RECT 208.950 350.400 250.050 351.600 ;
        RECT 251.400 351.600 252.600 353.400 ;
        RECT 262.950 353.400 322.050 354.600 ;
        RECT 262.950 352.950 265.050 353.400 ;
        RECT 319.950 352.950 322.050 353.400 ;
        RECT 376.950 354.600 379.050 355.050 ;
        RECT 478.950 354.600 481.050 355.050 ;
        RECT 376.950 353.400 481.050 354.600 ;
        RECT 376.950 352.950 379.050 353.400 ;
        RECT 478.950 352.950 481.050 353.400 ;
        RECT 484.950 354.600 487.050 355.050 ;
        RECT 499.950 354.600 502.050 355.050 ;
        RECT 484.950 353.400 502.050 354.600 ;
        RECT 484.950 352.950 487.050 353.400 ;
        RECT 499.950 352.950 502.050 353.400 ;
        RECT 505.950 354.600 508.050 355.050 ;
        RECT 517.950 354.600 520.050 355.050 ;
        RECT 505.950 353.400 520.050 354.600 ;
        RECT 505.950 352.950 508.050 353.400 ;
        RECT 517.950 352.950 520.050 353.400 ;
        RECT 562.950 354.600 565.050 355.050 ;
        RECT 598.950 354.600 601.050 355.050 ;
        RECT 562.950 353.400 601.050 354.600 ;
        RECT 562.950 352.950 565.050 353.400 ;
        RECT 598.950 352.950 601.050 353.400 ;
        RECT 700.950 354.600 703.050 355.050 ;
        RECT 727.950 354.600 730.050 355.050 ;
        RECT 790.950 354.600 793.050 355.050 ;
        RECT 700.950 353.400 793.050 354.600 ;
        RECT 700.950 352.950 703.050 353.400 ;
        RECT 727.950 352.950 730.050 353.400 ;
        RECT 790.950 352.950 793.050 353.400 ;
        RECT 256.950 351.600 259.050 352.050 ;
        RECT 274.950 351.600 277.050 352.050 ;
        RECT 251.400 350.400 277.050 351.600 ;
        RECT 208.950 349.950 211.050 350.400 ;
        RECT 247.950 349.950 250.050 350.400 ;
        RECT 256.950 349.950 259.050 350.400 ;
        RECT 274.950 349.950 277.050 350.400 ;
        RECT 316.950 351.600 319.050 352.050 ;
        RECT 475.950 351.600 478.050 352.050 ;
        RECT 316.950 350.400 478.050 351.600 ;
        RECT 316.950 349.950 319.050 350.400 ;
        RECT 475.950 349.950 478.050 350.400 ;
        RECT 478.950 351.600 481.050 352.050 ;
        RECT 577.950 351.600 580.050 352.050 ;
        RECT 478.950 350.400 580.050 351.600 ;
        RECT 478.950 349.950 481.050 350.400 ;
        RECT 577.950 349.950 580.050 350.400 ;
        RECT 592.950 351.600 595.050 352.050 ;
        RECT 637.950 351.600 640.050 352.050 ;
        RECT 592.950 350.400 640.050 351.600 ;
        RECT 592.950 349.950 595.050 350.400 ;
        RECT 637.950 349.950 640.050 350.400 ;
        RECT 727.950 351.600 730.050 352.050 ;
        RECT 760.950 351.600 763.050 352.050 ;
        RECT 727.950 350.400 763.050 351.600 ;
        RECT 727.950 349.950 730.050 350.400 ;
        RECT 760.950 349.950 763.050 350.400 ;
        RECT 796.950 351.600 799.050 352.050 ;
        RECT 844.950 351.600 847.050 352.050 ;
        RECT 796.950 350.400 847.050 351.600 ;
        RECT 796.950 349.950 799.050 350.400 ;
        RECT 844.950 349.950 847.050 350.400 ;
        RECT 43.950 348.600 46.050 349.050 ;
        RECT 52.950 348.600 55.050 349.050 ;
        RECT 43.950 347.400 55.050 348.600 ;
        RECT 43.950 346.950 46.050 347.400 ;
        RECT 52.950 346.950 55.050 347.400 ;
        RECT 238.950 348.600 241.050 349.050 ;
        RECT 307.950 348.600 310.050 349.050 ;
        RECT 238.950 347.400 310.050 348.600 ;
        RECT 238.950 346.950 241.050 347.400 ;
        RECT 307.950 346.950 310.050 347.400 ;
        RECT 322.950 348.600 325.050 349.050 ;
        RECT 328.950 348.600 331.050 349.050 ;
        RECT 322.950 347.400 331.050 348.600 ;
        RECT 322.950 346.950 325.050 347.400 ;
        RECT 328.950 346.950 331.050 347.400 ;
        RECT 445.950 348.600 448.050 349.050 ;
        RECT 457.950 348.600 460.050 349.050 ;
        RECT 520.950 348.600 523.050 349.050 ;
        RECT 445.950 347.400 456.600 348.600 ;
        RECT 445.950 346.950 448.050 347.400 ;
        RECT 10.950 345.600 13.050 346.050 ;
        RECT 34.950 345.600 37.050 346.050 ;
        RECT 46.950 345.600 49.050 346.050 ;
        RECT 10.950 344.400 33.600 345.600 ;
        RECT 10.950 343.950 13.050 344.400 ;
        RECT 32.400 343.050 33.600 344.400 ;
        RECT 34.950 344.400 49.050 345.600 ;
        RECT 34.950 343.950 37.050 344.400 ;
        RECT 46.950 343.950 49.050 344.400 ;
        RECT 100.950 345.600 103.050 346.050 ;
        RECT 133.950 345.600 136.050 346.050 ;
        RECT 151.950 345.600 154.050 346.050 ;
        RECT 100.950 344.400 154.050 345.600 ;
        RECT 100.950 343.950 103.050 344.400 ;
        RECT 133.950 343.950 136.050 344.400 ;
        RECT 151.950 343.950 154.050 344.400 ;
        RECT 166.950 345.600 169.050 346.050 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 166.950 344.400 190.050 345.600 ;
        RECT 166.950 343.950 169.050 344.400 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 211.950 345.600 214.050 346.050 ;
        RECT 199.950 344.400 214.050 345.600 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 211.950 343.950 214.050 344.400 ;
        RECT 214.950 345.600 217.050 346.050 ;
        RECT 220.950 345.600 223.050 346.050 ;
        RECT 214.950 344.400 223.050 345.600 ;
        RECT 214.950 343.950 217.050 344.400 ;
        RECT 220.950 343.950 223.050 344.400 ;
        RECT 256.950 345.600 259.050 346.050 ;
        RECT 280.950 345.600 283.050 346.050 ;
        RECT 286.950 345.600 289.050 346.050 ;
        RECT 301.950 345.600 304.050 346.050 ;
        RECT 256.950 344.400 279.600 345.600 ;
        RECT 256.950 343.950 259.050 344.400 ;
        RECT 278.400 343.050 279.600 344.400 ;
        RECT 280.950 344.400 304.050 345.600 ;
        RECT 280.950 343.950 283.050 344.400 ;
        RECT 286.950 343.950 289.050 344.400 ;
        RECT 301.950 343.950 304.050 344.400 ;
        RECT 319.950 345.600 322.050 346.050 ;
        RECT 397.950 345.600 400.050 346.050 ;
        RECT 319.950 344.400 400.050 345.600 ;
        RECT 319.950 343.950 322.050 344.400 ;
        RECT 397.950 343.950 400.050 344.400 ;
        RECT 418.950 345.600 421.050 346.050 ;
        RECT 451.950 345.600 454.050 346.050 ;
        RECT 418.950 344.400 454.050 345.600 ;
        RECT 455.400 345.600 456.600 347.400 ;
        RECT 457.950 347.400 523.050 348.600 ;
        RECT 457.950 346.950 460.050 347.400 ;
        RECT 520.950 346.950 523.050 347.400 ;
        RECT 655.950 348.600 658.050 349.050 ;
        RECT 664.950 348.600 667.050 349.050 ;
        RECT 682.950 348.600 685.050 349.050 ;
        RECT 655.950 347.400 685.050 348.600 ;
        RECT 655.950 346.950 658.050 347.400 ;
        RECT 664.950 346.950 667.050 347.400 ;
        RECT 682.950 346.950 685.050 347.400 ;
        RECT 694.950 348.600 697.050 349.050 ;
        RECT 733.950 348.600 736.050 349.050 ;
        RECT 694.950 347.400 736.050 348.600 ;
        RECT 694.950 346.950 697.050 347.400 ;
        RECT 733.950 346.950 736.050 347.400 ;
        RECT 805.950 348.600 808.050 349.050 ;
        RECT 832.950 348.600 835.050 349.050 ;
        RECT 805.950 347.400 835.050 348.600 ;
        RECT 805.950 346.950 808.050 347.400 ;
        RECT 832.950 346.950 835.050 347.400 ;
        RECT 490.950 345.600 493.050 346.050 ;
        RECT 455.400 344.400 493.050 345.600 ;
        RECT 418.950 343.950 421.050 344.400 ;
        RECT 451.950 343.950 454.050 344.400 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 496.950 345.600 499.050 346.050 ;
        RECT 505.950 345.600 508.050 346.050 ;
        RECT 496.950 344.400 508.050 345.600 ;
        RECT 496.950 343.950 499.050 344.400 ;
        RECT 505.950 343.950 508.050 344.400 ;
        RECT 508.950 345.600 511.050 346.050 ;
        RECT 535.950 345.600 538.050 346.050 ;
        RECT 568.950 345.600 571.050 346.050 ;
        RECT 508.950 344.400 538.050 345.600 ;
        RECT 508.950 343.950 511.050 344.400 ;
        RECT 535.950 343.950 538.050 344.400 ;
        RECT 557.400 344.400 571.050 345.600 ;
        RECT 31.950 340.950 34.050 343.050 ;
        RECT 49.950 342.600 52.050 343.050 ;
        RECT 35.400 341.400 52.050 342.600 ;
        RECT 22.950 339.600 25.050 340.050 ;
        RECT 35.400 339.600 36.600 341.400 ;
        RECT 49.950 340.950 52.050 341.400 ;
        RECT 61.950 342.600 64.050 343.050 ;
        RECT 67.950 342.600 70.050 343.050 ;
        RECT 61.950 341.400 70.050 342.600 ;
        RECT 61.950 340.950 64.050 341.400 ;
        RECT 67.950 340.950 70.050 341.400 ;
        RECT 94.950 340.950 97.050 343.050 ;
        RECT 121.950 342.600 124.050 343.050 ;
        RECT 127.950 342.600 130.050 343.050 ;
        RECT 121.950 341.400 130.050 342.600 ;
        RECT 121.950 340.950 124.050 341.400 ;
        RECT 127.950 340.950 130.050 341.400 ;
        RECT 190.950 342.600 193.050 343.050 ;
        RECT 217.950 342.600 220.050 343.050 ;
        RECT 190.950 341.400 220.050 342.600 ;
        RECT 190.950 340.950 193.050 341.400 ;
        RECT 217.950 340.950 220.050 341.400 ;
        RECT 226.950 342.600 229.050 343.050 ;
        RECT 232.950 342.600 235.050 343.050 ;
        RECT 256.950 342.600 259.050 343.050 ;
        RECT 226.950 341.400 259.050 342.600 ;
        RECT 226.950 340.950 229.050 341.400 ;
        RECT 232.950 340.950 235.050 341.400 ;
        RECT 256.950 340.950 259.050 341.400 ;
        RECT 259.950 340.950 262.050 343.050 ;
        RECT 277.950 340.950 280.050 343.050 ;
        RECT 280.950 342.600 283.050 343.050 ;
        RECT 310.950 342.600 313.050 343.050 ;
        RECT 280.950 341.400 313.050 342.600 ;
        RECT 280.950 340.950 283.050 341.400 ;
        RECT 310.950 340.950 313.050 341.400 ;
        RECT 415.950 342.600 418.050 343.050 ;
        RECT 424.950 342.600 427.050 343.050 ;
        RECT 454.950 342.600 457.050 343.050 ;
        RECT 557.400 342.600 558.600 344.400 ;
        RECT 568.950 343.950 571.050 344.400 ;
        RECT 574.950 345.600 577.050 346.050 ;
        RECT 601.950 345.600 604.050 346.050 ;
        RECT 574.950 344.400 604.050 345.600 ;
        RECT 574.950 343.950 577.050 344.400 ;
        RECT 601.950 343.950 604.050 344.400 ;
        RECT 670.950 345.600 673.050 346.050 ;
        RECT 709.950 345.600 712.050 346.050 ;
        RECT 670.950 344.400 712.050 345.600 ;
        RECT 670.950 343.950 673.050 344.400 ;
        RECT 709.950 343.950 712.050 344.400 ;
        RECT 733.950 345.600 736.050 346.050 ;
        RECT 739.950 345.600 742.050 346.050 ;
        RECT 733.950 344.400 742.050 345.600 ;
        RECT 733.950 343.950 736.050 344.400 ;
        RECT 739.950 343.950 742.050 344.400 ;
        RECT 784.950 345.600 787.050 346.050 ;
        RECT 790.950 345.600 793.050 346.050 ;
        RECT 784.950 344.400 793.050 345.600 ;
        RECT 784.950 343.950 787.050 344.400 ;
        RECT 790.950 343.950 793.050 344.400 ;
        RECT 817.950 345.600 820.050 346.050 ;
        RECT 826.950 345.600 829.050 346.050 ;
        RECT 856.950 345.600 859.050 346.050 ;
        RECT 817.950 344.400 859.050 345.600 ;
        RECT 817.950 343.950 820.050 344.400 ;
        RECT 826.950 343.950 829.050 344.400 ;
        RECT 856.950 343.950 859.050 344.400 ;
        RECT 415.950 341.400 420.600 342.600 ;
        RECT 415.950 340.950 418.050 341.400 ;
        RECT 22.950 338.400 36.600 339.600 ;
        RECT 37.950 339.600 40.050 340.050 ;
        RECT 43.950 339.600 46.050 340.050 ;
        RECT 46.950 339.600 49.050 340.050 ;
        RECT 37.950 338.400 49.050 339.600 ;
        RECT 22.950 337.950 25.050 338.400 ;
        RECT 37.950 337.950 40.050 338.400 ;
        RECT 43.950 337.950 46.050 338.400 ;
        RECT 46.950 337.950 49.050 338.400 ;
        RECT 64.950 339.600 67.050 340.050 ;
        RECT 95.400 339.600 96.600 340.950 ;
        RECT 64.950 338.400 96.600 339.600 ;
        RECT 142.950 339.600 145.050 340.050 ;
        RECT 172.950 339.600 175.050 340.050 ;
        RECT 142.950 338.400 175.050 339.600 ;
        RECT 64.950 337.950 67.050 338.400 ;
        RECT 142.950 337.950 145.050 338.400 ;
        RECT 172.950 337.950 175.050 338.400 ;
        RECT 223.950 339.600 226.050 340.050 ;
        RECT 253.950 339.600 256.050 340.050 ;
        RECT 223.950 338.400 256.050 339.600 ;
        RECT 223.950 337.950 226.050 338.400 ;
        RECT 253.950 337.950 256.050 338.400 ;
        RECT 260.400 337.050 261.600 340.950 ;
        RECT 268.950 339.600 271.050 340.050 ;
        RECT 283.950 339.600 286.050 340.050 ;
        RECT 268.950 338.400 286.050 339.600 ;
        RECT 268.950 337.950 271.050 338.400 ;
        RECT 283.950 337.950 286.050 338.400 ;
        RECT 286.950 339.600 289.050 340.050 ;
        RECT 304.950 339.600 307.050 340.050 ;
        RECT 316.950 339.600 319.050 340.050 ;
        RECT 286.950 338.400 319.050 339.600 ;
        RECT 286.950 337.950 289.050 338.400 ;
        RECT 304.950 337.950 307.050 338.400 ;
        RECT 316.950 337.950 319.050 338.400 ;
        RECT 394.950 339.600 397.050 340.050 ;
        RECT 415.950 339.600 418.050 340.050 ;
        RECT 394.950 338.400 418.050 339.600 ;
        RECT 419.400 339.600 420.600 341.400 ;
        RECT 424.950 341.400 457.050 342.600 ;
        RECT 424.950 340.950 427.050 341.400 ;
        RECT 454.950 340.950 457.050 341.400 ;
        RECT 551.400 341.400 558.600 342.600 ;
        RECT 559.950 342.600 562.050 343.050 ;
        RECT 583.950 342.600 586.050 343.050 ;
        RECT 559.950 341.400 586.050 342.600 ;
        RECT 551.400 340.050 552.600 341.400 ;
        RECT 559.950 340.950 562.050 341.400 ;
        RECT 583.950 340.950 586.050 341.400 ;
        RECT 688.950 340.950 691.050 343.050 ;
        RECT 721.950 342.600 724.050 343.050 ;
        RECT 736.950 342.600 739.050 343.050 ;
        RECT 757.950 342.600 760.050 343.050 ;
        RECT 721.950 341.400 760.050 342.600 ;
        RECT 721.950 340.950 724.050 341.400 ;
        RECT 736.950 340.950 739.050 341.400 ;
        RECT 757.950 340.950 760.050 341.400 ;
        RECT 763.950 342.600 766.050 343.050 ;
        RECT 769.950 342.600 772.050 343.050 ;
        RECT 763.950 341.400 772.050 342.600 ;
        RECT 763.950 340.950 766.050 341.400 ;
        RECT 769.950 340.950 772.050 341.400 ;
        RECT 832.950 342.600 835.050 343.050 ;
        RECT 835.950 342.600 838.050 343.050 ;
        RECT 853.950 342.600 856.050 343.050 ;
        RECT 859.950 342.600 862.050 343.050 ;
        RECT 832.950 341.400 849.600 342.600 ;
        RECT 832.950 340.950 835.050 341.400 ;
        RECT 835.950 340.950 838.050 341.400 ;
        RECT 433.950 339.600 436.050 340.050 ;
        RECT 419.400 338.400 436.050 339.600 ;
        RECT 394.950 337.950 397.050 338.400 ;
        RECT 415.950 337.950 418.050 338.400 ;
        RECT 433.950 337.950 436.050 338.400 ;
        RECT 454.950 339.600 457.050 340.050 ;
        RECT 478.950 339.600 481.050 340.050 ;
        RECT 454.950 338.400 481.050 339.600 ;
        RECT 454.950 337.950 457.050 338.400 ;
        RECT 478.950 337.950 481.050 338.400 ;
        RECT 481.950 339.600 484.050 340.050 ;
        RECT 490.950 339.600 493.050 340.050 ;
        RECT 481.950 338.400 493.050 339.600 ;
        RECT 481.950 337.950 484.050 338.400 ;
        RECT 490.950 337.950 493.050 338.400 ;
        RECT 523.950 339.600 526.050 340.050 ;
        RECT 529.950 339.600 532.050 340.050 ;
        RECT 523.950 338.400 532.050 339.600 ;
        RECT 523.950 337.950 526.050 338.400 ;
        RECT 529.950 337.950 532.050 338.400 ;
        RECT 535.950 339.600 538.050 340.050 ;
        RECT 544.950 339.600 547.050 340.050 ;
        RECT 535.950 338.400 547.050 339.600 ;
        RECT 535.950 337.950 538.050 338.400 ;
        RECT 544.950 337.950 547.050 338.400 ;
        RECT 550.950 337.950 553.050 340.050 ;
        RECT 553.950 339.600 556.050 340.050 ;
        RECT 625.950 339.600 628.050 340.050 ;
        RECT 658.950 339.600 661.050 340.050 ;
        RECT 553.950 338.400 624.600 339.600 ;
        RECT 553.950 337.950 556.050 338.400 ;
        RECT 623.400 337.050 624.600 338.400 ;
        RECT 625.950 338.400 661.050 339.600 ;
        RECT 625.950 337.950 628.050 338.400 ;
        RECT 658.950 337.950 661.050 338.400 ;
        RECT 689.400 337.050 690.600 340.950 ;
        RECT 848.400 340.050 849.600 341.400 ;
        RECT 853.950 341.400 862.050 342.600 ;
        RECT 853.950 340.950 856.050 341.400 ;
        RECT 859.950 340.950 862.050 341.400 ;
        RECT 691.950 339.600 694.050 340.050 ;
        RECT 706.950 339.600 709.050 340.050 ;
        RECT 691.950 338.400 709.050 339.600 ;
        RECT 691.950 337.950 694.050 338.400 ;
        RECT 706.950 337.950 709.050 338.400 ;
        RECT 730.950 339.600 733.050 340.050 ;
        RECT 745.950 339.600 748.050 340.050 ;
        RECT 730.950 338.400 748.050 339.600 ;
        RECT 730.950 337.950 733.050 338.400 ;
        RECT 745.950 337.950 748.050 338.400 ;
        RECT 766.950 339.600 769.050 340.050 ;
        RECT 781.950 339.600 784.050 340.050 ;
        RECT 766.950 338.400 784.050 339.600 ;
        RECT 766.950 337.950 769.050 338.400 ;
        RECT 781.950 337.950 784.050 338.400 ;
        RECT 808.950 339.600 811.050 340.050 ;
        RECT 817.950 339.600 820.050 340.050 ;
        RECT 808.950 338.400 820.050 339.600 ;
        RECT 808.950 337.950 811.050 338.400 ;
        RECT 817.950 337.950 820.050 338.400 ;
        RECT 847.950 337.950 850.050 340.050 ;
        RECT 55.950 336.600 58.050 337.050 ;
        RECT 70.950 336.600 73.050 337.050 ;
        RECT 55.950 335.400 73.050 336.600 ;
        RECT 55.950 334.950 58.050 335.400 ;
        RECT 70.950 334.950 73.050 335.400 ;
        RECT 73.950 336.600 76.050 337.050 ;
        RECT 79.950 336.600 82.050 337.050 ;
        RECT 97.950 336.600 100.050 337.050 ;
        RECT 73.950 335.400 100.050 336.600 ;
        RECT 73.950 334.950 76.050 335.400 ;
        RECT 79.950 334.950 82.050 335.400 ;
        RECT 97.950 334.950 100.050 335.400 ;
        RECT 154.950 336.600 157.050 337.050 ;
        RECT 160.950 336.600 163.050 337.050 ;
        RECT 154.950 335.400 163.050 336.600 ;
        RECT 154.950 334.950 157.050 335.400 ;
        RECT 160.950 334.950 163.050 335.400 ;
        RECT 193.950 336.600 196.050 337.050 ;
        RECT 214.950 336.600 217.050 337.050 ;
        RECT 235.950 336.600 238.050 337.050 ;
        RECT 193.950 335.400 238.050 336.600 ;
        RECT 193.950 334.950 196.050 335.400 ;
        RECT 214.950 334.950 217.050 335.400 ;
        RECT 235.950 334.950 238.050 335.400 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 336.600 265.050 337.050 ;
        RECT 325.950 336.600 328.050 337.050 ;
        RECT 349.950 336.600 352.050 337.050 ;
        RECT 262.950 335.400 328.050 336.600 ;
        RECT 262.950 334.950 265.050 335.400 ;
        RECT 325.950 334.950 328.050 335.400 ;
        RECT 341.400 335.400 352.050 336.600 ;
        RECT 67.950 333.600 70.050 334.050 ;
        RECT 76.950 333.600 79.050 334.050 ;
        RECT 67.950 332.400 79.050 333.600 ;
        RECT 67.950 331.950 70.050 332.400 ;
        RECT 76.950 331.950 79.050 332.400 ;
        RECT 85.950 333.600 88.050 334.050 ;
        RECT 94.950 333.600 97.050 334.050 ;
        RECT 85.950 332.400 97.050 333.600 ;
        RECT 85.950 331.950 88.050 332.400 ;
        RECT 94.950 331.950 97.050 332.400 ;
        RECT 157.950 333.600 160.050 334.050 ;
        RECT 163.950 333.600 166.050 334.050 ;
        RECT 157.950 332.400 166.050 333.600 ;
        RECT 157.950 331.950 160.050 332.400 ;
        RECT 163.950 331.950 166.050 332.400 ;
        RECT 175.950 333.600 178.050 334.050 ;
        RECT 193.950 333.600 196.050 334.050 ;
        RECT 175.950 332.400 196.050 333.600 ;
        RECT 175.950 331.950 178.050 332.400 ;
        RECT 193.950 331.950 196.050 332.400 ;
        RECT 211.950 333.600 214.050 334.050 ;
        RECT 226.950 333.600 229.050 334.050 ;
        RECT 211.950 332.400 229.050 333.600 ;
        RECT 211.950 331.950 214.050 332.400 ;
        RECT 226.950 331.950 229.050 332.400 ;
        RECT 241.950 333.600 244.050 334.050 ;
        RECT 262.950 333.600 265.050 334.050 ;
        RECT 271.950 333.600 274.050 334.050 ;
        RECT 241.950 332.400 265.050 333.600 ;
        RECT 241.950 331.950 244.050 332.400 ;
        RECT 262.950 331.950 265.050 332.400 ;
        RECT 269.400 332.400 274.050 333.600 ;
        RECT 49.950 330.600 52.050 331.050 ;
        RECT 88.950 330.600 91.050 331.050 ;
        RECT 49.950 329.400 91.050 330.600 ;
        RECT 49.950 328.950 52.050 329.400 ;
        RECT 88.950 328.950 91.050 329.400 ;
        RECT 91.950 330.600 94.050 331.050 ;
        RECT 115.950 330.600 118.050 331.050 ;
        RECT 91.950 329.400 118.050 330.600 ;
        RECT 91.950 328.950 94.050 329.400 ;
        RECT 115.950 328.950 118.050 329.400 ;
        RECT 256.950 330.600 259.050 331.050 ;
        RECT 269.400 330.600 270.600 332.400 ;
        RECT 271.950 331.950 274.050 332.400 ;
        RECT 313.950 333.600 316.050 334.050 ;
        RECT 341.400 333.600 342.600 335.400 ;
        RECT 349.950 334.950 352.050 335.400 ;
        RECT 406.950 336.600 409.050 337.050 ;
        RECT 436.950 336.600 439.050 337.050 ;
        RECT 466.950 336.600 469.050 337.050 ;
        RECT 406.950 335.400 469.050 336.600 ;
        RECT 406.950 334.950 409.050 335.400 ;
        RECT 436.950 334.950 439.050 335.400 ;
        RECT 466.950 334.950 469.050 335.400 ;
        RECT 472.950 336.600 475.050 337.050 ;
        RECT 478.950 336.600 481.050 337.050 ;
        RECT 472.950 335.400 481.050 336.600 ;
        RECT 472.950 334.950 475.050 335.400 ;
        RECT 478.950 334.950 481.050 335.400 ;
        RECT 523.950 336.600 526.050 337.050 ;
        RECT 547.950 336.600 550.050 337.050 ;
        RECT 523.950 335.400 550.050 336.600 ;
        RECT 523.950 334.950 526.050 335.400 ;
        RECT 547.950 334.950 550.050 335.400 ;
        RECT 565.950 336.600 568.050 337.050 ;
        RECT 574.950 336.600 577.050 337.050 ;
        RECT 565.950 335.400 577.050 336.600 ;
        RECT 565.950 334.950 568.050 335.400 ;
        RECT 574.950 334.950 577.050 335.400 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 688.950 334.950 691.050 337.050 ;
        RECT 724.950 336.600 727.050 337.050 ;
        RECT 739.950 336.600 742.050 337.050 ;
        RECT 724.950 335.400 742.050 336.600 ;
        RECT 724.950 334.950 727.050 335.400 ;
        RECT 739.950 334.950 742.050 335.400 ;
        RECT 769.950 336.600 772.050 337.050 ;
        RECT 808.950 336.600 811.050 337.050 ;
        RECT 769.950 335.400 811.050 336.600 ;
        RECT 769.950 334.950 772.050 335.400 ;
        RECT 808.950 334.950 811.050 335.400 ;
        RECT 826.950 336.600 829.050 337.050 ;
        RECT 844.950 336.600 847.050 337.050 ;
        RECT 856.950 336.600 859.050 337.050 ;
        RECT 826.950 335.400 859.050 336.600 ;
        RECT 826.950 334.950 829.050 335.400 ;
        RECT 844.950 334.950 847.050 335.400 ;
        RECT 856.950 334.950 859.050 335.400 ;
        RECT 313.950 332.400 342.600 333.600 ;
        RECT 349.950 333.600 352.050 334.050 ;
        RECT 388.950 333.600 391.050 334.050 ;
        RECT 349.950 332.400 391.050 333.600 ;
        RECT 313.950 331.950 316.050 332.400 ;
        RECT 349.950 331.950 352.050 332.400 ;
        RECT 388.950 331.950 391.050 332.400 ;
        RECT 406.950 333.600 409.050 334.050 ;
        RECT 427.950 333.600 430.050 334.050 ;
        RECT 406.950 332.400 430.050 333.600 ;
        RECT 406.950 331.950 409.050 332.400 ;
        RECT 427.950 331.950 430.050 332.400 ;
        RECT 439.950 333.600 442.050 334.050 ;
        RECT 496.950 333.600 499.050 334.050 ;
        RECT 508.950 333.600 511.050 334.050 ;
        RECT 439.950 332.400 511.050 333.600 ;
        RECT 439.950 331.950 442.050 332.400 ;
        RECT 496.950 331.950 499.050 332.400 ;
        RECT 508.950 331.950 511.050 332.400 ;
        RECT 547.950 333.600 550.050 334.050 ;
        RECT 655.950 333.600 658.050 334.050 ;
        RECT 547.950 332.400 658.050 333.600 ;
        RECT 547.950 331.950 550.050 332.400 ;
        RECT 655.950 331.950 658.050 332.400 ;
        RECT 256.950 329.400 270.600 330.600 ;
        RECT 271.950 330.600 274.050 331.050 ;
        RECT 298.950 330.600 301.050 331.050 ;
        RECT 271.950 329.400 301.050 330.600 ;
        RECT 256.950 328.950 259.050 329.400 ;
        RECT 271.950 328.950 274.050 329.400 ;
        RECT 298.950 328.950 301.050 329.400 ;
        RECT 415.950 330.600 418.050 331.050 ;
        RECT 526.950 330.600 529.050 331.050 ;
        RECT 568.950 330.600 571.050 331.050 ;
        RECT 415.950 329.400 571.050 330.600 ;
        RECT 415.950 328.950 418.050 329.400 ;
        RECT 526.950 328.950 529.050 329.400 ;
        RECT 568.950 328.950 571.050 329.400 ;
        RECT 679.950 330.600 682.050 331.050 ;
        RECT 685.950 330.600 688.050 331.050 ;
        RECT 754.950 330.600 757.050 331.050 ;
        RECT 679.950 329.400 757.050 330.600 ;
        RECT 679.950 328.950 682.050 329.400 ;
        RECT 685.950 328.950 688.050 329.400 ;
        RECT 754.950 328.950 757.050 329.400 ;
        RECT 781.950 330.600 784.050 331.050 ;
        RECT 802.950 330.600 805.050 331.050 ;
        RECT 781.950 329.400 805.050 330.600 ;
        RECT 781.950 328.950 784.050 329.400 ;
        RECT 802.950 328.950 805.050 329.400 ;
        RECT 850.950 330.600 853.050 331.050 ;
        RECT 859.950 330.600 862.050 331.050 ;
        RECT 850.950 329.400 862.050 330.600 ;
        RECT 850.950 328.950 853.050 329.400 ;
        RECT 859.950 328.950 862.050 329.400 ;
        RECT 61.950 327.600 64.050 328.050 ;
        RECT 70.950 327.600 73.050 328.050 ;
        RECT 61.950 326.400 73.050 327.600 ;
        RECT 61.950 325.950 64.050 326.400 ;
        RECT 70.950 325.950 73.050 326.400 ;
        RECT 274.950 327.600 277.050 328.050 ;
        RECT 283.950 327.600 286.050 328.050 ;
        RECT 274.950 326.400 286.050 327.600 ;
        RECT 274.950 325.950 277.050 326.400 ;
        RECT 283.950 325.950 286.050 326.400 ;
        RECT 340.950 327.600 343.050 328.050 ;
        RECT 376.950 327.600 379.050 328.050 ;
        RECT 340.950 326.400 379.050 327.600 ;
        RECT 340.950 325.950 343.050 326.400 ;
        RECT 376.950 325.950 379.050 326.400 ;
        RECT 382.950 327.600 385.050 328.050 ;
        RECT 469.950 327.600 472.050 328.050 ;
        RECT 382.950 326.400 472.050 327.600 ;
        RECT 382.950 325.950 385.050 326.400 ;
        RECT 469.950 325.950 472.050 326.400 ;
        RECT 502.950 327.600 505.050 328.050 ;
        RECT 508.950 327.600 511.050 328.050 ;
        RECT 502.950 326.400 511.050 327.600 ;
        RECT 502.950 325.950 505.050 326.400 ;
        RECT 508.950 325.950 511.050 326.400 ;
        RECT 511.950 327.600 514.050 328.050 ;
        RECT 538.950 327.600 541.050 328.050 ;
        RECT 511.950 326.400 541.050 327.600 ;
        RECT 511.950 325.950 514.050 326.400 ;
        RECT 538.950 325.950 541.050 326.400 ;
        RECT 565.950 327.600 568.050 328.050 ;
        RECT 571.950 327.600 574.050 328.050 ;
        RECT 565.950 326.400 574.050 327.600 ;
        RECT 565.950 325.950 568.050 326.400 ;
        RECT 571.950 325.950 574.050 326.400 ;
        RECT 706.950 327.600 709.050 328.050 ;
        RECT 733.950 327.600 736.050 328.050 ;
        RECT 706.950 326.400 736.050 327.600 ;
        RECT 706.950 325.950 709.050 326.400 ;
        RECT 733.950 325.950 736.050 326.400 ;
        RECT 754.950 327.600 757.050 328.050 ;
        RECT 859.950 327.600 862.050 328.050 ;
        RECT 754.950 326.400 862.050 327.600 ;
        RECT 754.950 325.950 757.050 326.400 ;
        RECT 859.950 325.950 862.050 326.400 ;
        RECT 16.950 324.600 19.050 325.050 ;
        RECT 280.950 324.600 283.050 325.050 ;
        RECT 16.950 323.400 283.050 324.600 ;
        RECT 16.950 322.950 19.050 323.400 ;
        RECT 280.950 322.950 283.050 323.400 ;
        RECT 322.950 324.600 325.050 325.050 ;
        RECT 334.950 324.600 337.050 325.050 ;
        RECT 364.950 324.600 367.050 325.050 ;
        RECT 514.950 324.600 517.050 325.050 ;
        RECT 592.950 324.600 595.050 325.050 ;
        RECT 322.950 323.400 595.050 324.600 ;
        RECT 322.950 322.950 325.050 323.400 ;
        RECT 334.950 322.950 337.050 323.400 ;
        RECT 364.950 322.950 367.050 323.400 ;
        RECT 514.950 322.950 517.050 323.400 ;
        RECT 592.950 322.950 595.050 323.400 ;
        RECT 604.950 324.600 607.050 325.050 ;
        RECT 694.950 324.600 697.050 325.050 ;
        RECT 604.950 323.400 697.050 324.600 ;
        RECT 604.950 322.950 607.050 323.400 ;
        RECT 694.950 322.950 697.050 323.400 ;
        RECT 748.950 324.600 751.050 325.050 ;
        RECT 829.950 324.600 832.050 325.050 ;
        RECT 748.950 323.400 832.050 324.600 ;
        RECT 748.950 322.950 751.050 323.400 ;
        RECT 829.950 322.950 832.050 323.400 ;
        RECT 85.950 321.600 88.050 322.050 ;
        RECT 136.950 321.600 139.050 322.050 ;
        RECT 85.950 320.400 139.050 321.600 ;
        RECT 85.950 319.950 88.050 320.400 ;
        RECT 136.950 319.950 139.050 320.400 ;
        RECT 220.950 321.600 223.050 322.050 ;
        RECT 238.950 321.600 241.050 322.050 ;
        RECT 454.950 321.600 457.050 322.050 ;
        RECT 676.950 321.600 679.050 322.050 ;
        RECT 220.950 320.400 241.050 321.600 ;
        RECT 220.950 319.950 223.050 320.400 ;
        RECT 238.950 319.950 241.050 320.400 ;
        RECT 365.400 320.400 457.050 321.600 ;
        RECT 10.950 318.600 13.050 319.050 ;
        RECT 118.950 318.600 121.050 319.050 ;
        RECT 10.950 317.400 121.050 318.600 ;
        RECT 10.950 316.950 13.050 317.400 ;
        RECT 118.950 316.950 121.050 317.400 ;
        RECT 136.950 318.600 139.050 319.050 ;
        RECT 202.950 318.600 205.050 319.050 ;
        RECT 136.950 317.400 205.050 318.600 ;
        RECT 136.950 316.950 139.050 317.400 ;
        RECT 202.950 316.950 205.050 317.400 ;
        RECT 235.950 318.600 238.050 319.050 ;
        RECT 265.950 318.600 268.050 319.050 ;
        RECT 235.950 317.400 268.050 318.600 ;
        RECT 235.950 316.950 238.050 317.400 ;
        RECT 265.950 316.950 268.050 317.400 ;
        RECT 277.950 318.600 280.050 319.050 ;
        RECT 289.950 318.600 292.050 319.050 ;
        RECT 277.950 317.400 292.050 318.600 ;
        RECT 277.950 316.950 280.050 317.400 ;
        RECT 289.950 316.950 292.050 317.400 ;
        RECT 295.950 318.600 298.050 319.050 ;
        RECT 365.400 318.600 366.600 320.400 ;
        RECT 454.950 319.950 457.050 320.400 ;
        RECT 518.400 320.400 679.050 321.600 ;
        RECT 295.950 317.400 366.600 318.600 ;
        RECT 391.950 318.600 394.050 319.050 ;
        RECT 433.950 318.600 436.050 319.050 ;
        RECT 391.950 317.400 436.050 318.600 ;
        RECT 295.950 316.950 298.050 317.400 ;
        RECT 391.950 316.950 394.050 317.400 ;
        RECT 433.950 316.950 436.050 317.400 ;
        RECT 496.950 318.600 499.050 319.050 ;
        RECT 518.400 318.600 519.600 320.400 ;
        RECT 676.950 319.950 679.050 320.400 ;
        RECT 742.950 321.600 745.050 322.050 ;
        RECT 757.950 321.600 760.050 322.050 ;
        RECT 742.950 320.400 760.050 321.600 ;
        RECT 742.950 319.950 745.050 320.400 ;
        RECT 757.950 319.950 760.050 320.400 ;
        RECT 829.950 321.600 832.050 322.050 ;
        RECT 862.950 321.600 865.050 322.050 ;
        RECT 871.950 321.600 874.050 322.050 ;
        RECT 829.950 320.400 874.050 321.600 ;
        RECT 829.950 319.950 832.050 320.400 ;
        RECT 862.950 319.950 865.050 320.400 ;
        RECT 871.950 319.950 874.050 320.400 ;
        RECT 496.950 317.400 519.600 318.600 ;
        RECT 520.950 318.600 523.050 319.050 ;
        RECT 607.950 318.600 610.050 319.050 ;
        RECT 520.950 317.400 610.050 318.600 ;
        RECT 496.950 316.950 499.050 317.400 ;
        RECT 520.950 316.950 523.050 317.400 ;
        RECT 607.950 316.950 610.050 317.400 ;
        RECT 751.950 318.600 754.050 319.050 ;
        RECT 760.950 318.600 763.050 319.050 ;
        RECT 751.950 317.400 763.050 318.600 ;
        RECT 751.950 316.950 754.050 317.400 ;
        RECT 760.950 316.950 763.050 317.400 ;
        RECT 763.950 318.600 766.050 319.050 ;
        RECT 766.950 318.600 769.050 319.050 ;
        RECT 772.950 318.600 775.050 319.050 ;
        RECT 763.950 317.400 775.050 318.600 ;
        RECT 763.950 316.950 766.050 317.400 ;
        RECT 766.950 316.950 769.050 317.400 ;
        RECT 772.950 316.950 775.050 317.400 ;
        RECT 784.950 318.600 787.050 319.050 ;
        RECT 814.950 318.600 817.050 319.050 ;
        RECT 784.950 317.400 817.050 318.600 ;
        RECT 784.950 316.950 787.050 317.400 ;
        RECT 814.950 316.950 817.050 317.400 ;
        RECT 854.400 317.400 864.600 318.600 ;
        RECT 28.950 315.600 31.050 316.050 ;
        RECT 40.950 315.600 43.050 316.050 ;
        RECT 28.950 314.400 43.050 315.600 ;
        RECT 28.950 313.950 31.050 314.400 ;
        RECT 40.950 313.950 43.050 314.400 ;
        RECT 43.950 315.600 46.050 316.050 ;
        RECT 55.950 315.600 58.050 316.050 ;
        RECT 43.950 314.400 58.050 315.600 ;
        RECT 43.950 313.950 46.050 314.400 ;
        RECT 55.950 313.950 58.050 314.400 ;
        RECT 118.950 315.600 121.050 316.050 ;
        RECT 133.950 315.600 136.050 316.050 ;
        RECT 118.950 314.400 136.050 315.600 ;
        RECT 118.950 313.950 121.050 314.400 ;
        RECT 133.950 313.950 136.050 314.400 ;
        RECT 190.950 315.600 193.050 316.050 ;
        RECT 208.950 315.600 211.050 316.050 ;
        RECT 190.950 314.400 211.050 315.600 ;
        RECT 190.950 313.950 193.050 314.400 ;
        RECT 208.950 313.950 211.050 314.400 ;
        RECT 226.950 315.600 229.050 316.050 ;
        RECT 253.950 315.600 256.050 316.050 ;
        RECT 265.950 315.600 268.050 316.050 ;
        RECT 283.950 315.600 286.050 316.050 ;
        RECT 226.950 314.400 286.050 315.600 ;
        RECT 226.950 313.950 229.050 314.400 ;
        RECT 253.950 313.950 256.050 314.400 ;
        RECT 265.950 313.950 268.050 314.400 ;
        RECT 283.950 313.950 286.050 314.400 ;
        RECT 361.950 315.600 364.050 316.050 ;
        RECT 412.950 315.600 415.050 316.050 ;
        RECT 361.950 314.400 415.050 315.600 ;
        RECT 361.950 313.950 364.050 314.400 ;
        RECT 412.950 313.950 415.050 314.400 ;
        RECT 427.950 315.600 430.050 316.050 ;
        RECT 436.950 315.600 439.050 316.050 ;
        RECT 427.950 314.400 439.050 315.600 ;
        RECT 427.950 313.950 430.050 314.400 ;
        RECT 436.950 313.950 439.050 314.400 ;
        RECT 475.950 315.600 478.050 316.050 ;
        RECT 490.950 315.600 493.050 316.050 ;
        RECT 502.950 315.600 505.050 316.050 ;
        RECT 529.950 315.600 532.050 316.050 ;
        RECT 475.950 314.400 501.600 315.600 ;
        RECT 475.950 313.950 478.050 314.400 ;
        RECT 490.950 313.950 493.050 314.400 ;
        RECT 61.950 312.600 64.050 313.050 ;
        RECT 91.950 312.600 94.050 313.050 ;
        RECT 61.950 311.400 94.050 312.600 ;
        RECT 61.950 310.950 64.050 311.400 ;
        RECT 91.950 310.950 94.050 311.400 ;
        RECT 100.950 312.600 103.050 313.050 ;
        RECT 112.950 312.600 115.050 313.050 ;
        RECT 100.950 311.400 115.050 312.600 ;
        RECT 100.950 310.950 103.050 311.400 ;
        RECT 112.950 310.950 115.050 311.400 ;
        RECT 124.950 312.600 127.050 313.050 ;
        RECT 166.950 312.600 169.050 313.050 ;
        RECT 124.950 311.400 169.050 312.600 ;
        RECT 124.950 310.950 127.050 311.400 ;
        RECT 166.950 310.950 169.050 311.400 ;
        RECT 169.950 312.600 172.050 313.050 ;
        RECT 181.950 312.600 184.050 313.050 ;
        RECT 169.950 311.400 184.050 312.600 ;
        RECT 169.950 310.950 172.050 311.400 ;
        RECT 181.950 310.950 184.050 311.400 ;
        RECT 187.950 312.600 190.050 313.050 ;
        RECT 208.950 312.600 211.050 313.050 ;
        RECT 220.950 312.600 223.050 313.050 ;
        RECT 247.950 312.600 250.050 313.050 ;
        RECT 187.950 311.400 223.050 312.600 ;
        RECT 187.950 310.950 190.050 311.400 ;
        RECT 208.950 310.950 211.050 311.400 ;
        RECT 220.950 310.950 223.050 311.400 ;
        RECT 224.400 311.400 250.050 312.600 ;
        RECT 224.400 310.050 225.600 311.400 ;
        RECT 247.950 310.950 250.050 311.400 ;
        RECT 250.950 312.600 253.050 313.050 ;
        RECT 289.950 312.600 292.050 313.050 ;
        RECT 250.950 311.400 292.050 312.600 ;
        RECT 250.950 310.950 253.050 311.400 ;
        RECT 289.950 310.950 292.050 311.400 ;
        RECT 298.950 312.600 301.050 313.050 ;
        RECT 313.950 312.600 316.050 313.050 ;
        RECT 298.950 311.400 316.050 312.600 ;
        RECT 298.950 310.950 301.050 311.400 ;
        RECT 313.950 310.950 316.050 311.400 ;
        RECT 328.950 312.600 331.050 313.050 ;
        RECT 500.400 312.600 501.600 314.400 ;
        RECT 502.950 314.400 532.050 315.600 ;
        RECT 502.950 313.950 505.050 314.400 ;
        RECT 529.950 313.950 532.050 314.400 ;
        RECT 535.950 315.600 538.050 316.050 ;
        RECT 550.950 315.600 553.050 316.050 ;
        RECT 535.950 314.400 553.050 315.600 ;
        RECT 535.950 313.950 538.050 314.400 ;
        RECT 550.950 313.950 553.050 314.400 ;
        RECT 610.950 315.600 613.050 316.050 ;
        RECT 637.950 315.600 640.050 316.050 ;
        RECT 610.950 314.400 640.050 315.600 ;
        RECT 610.950 313.950 613.050 314.400 ;
        RECT 637.950 313.950 640.050 314.400 ;
        RECT 667.950 315.600 670.050 316.050 ;
        RECT 676.950 315.600 679.050 316.050 ;
        RECT 667.950 314.400 679.050 315.600 ;
        RECT 667.950 313.950 670.050 314.400 ;
        RECT 676.950 313.950 679.050 314.400 ;
        RECT 703.950 315.600 706.050 316.050 ;
        RECT 715.950 315.600 718.050 316.050 ;
        RECT 703.950 314.400 718.050 315.600 ;
        RECT 703.950 313.950 706.050 314.400 ;
        RECT 715.950 313.950 718.050 314.400 ;
        RECT 721.950 315.600 724.050 316.050 ;
        RECT 772.950 315.600 775.050 316.050 ;
        RECT 721.950 314.400 775.050 315.600 ;
        RECT 721.950 313.950 724.050 314.400 ;
        RECT 772.950 313.950 775.050 314.400 ;
        RECT 775.950 313.950 778.050 316.050 ;
        RECT 778.950 315.600 781.050 316.050 ;
        RECT 790.950 315.600 793.050 316.050 ;
        RECT 778.950 314.400 793.050 315.600 ;
        RECT 778.950 313.950 781.050 314.400 ;
        RECT 790.950 313.950 793.050 314.400 ;
        RECT 805.950 315.600 808.050 316.050 ;
        RECT 814.950 315.600 817.050 316.050 ;
        RECT 850.950 315.600 853.050 316.050 ;
        RECT 805.950 314.400 817.050 315.600 ;
        RECT 805.950 313.950 808.050 314.400 ;
        RECT 814.950 313.950 817.050 314.400 ;
        RECT 845.400 314.400 853.050 315.600 ;
        RECT 517.950 312.600 520.050 313.050 ;
        RECT 544.950 312.600 547.050 313.050 ;
        RECT 568.950 312.600 571.050 313.050 ;
        RECT 574.950 312.600 577.050 313.050 ;
        RECT 328.950 311.400 432.600 312.600 ;
        RECT 500.400 311.400 528.600 312.600 ;
        RECT 328.950 310.950 331.050 311.400 ;
        RECT 431.400 310.050 432.600 311.400 ;
        RECT 517.950 310.950 520.050 311.400 ;
        RECT 527.400 310.050 528.600 311.400 ;
        RECT 544.950 311.400 577.050 312.600 ;
        RECT 544.950 310.950 547.050 311.400 ;
        RECT 568.950 310.950 571.050 311.400 ;
        RECT 574.950 310.950 577.050 311.400 ;
        RECT 595.950 312.600 598.050 313.050 ;
        RECT 601.950 312.600 604.050 313.050 ;
        RECT 595.950 311.400 604.050 312.600 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 601.950 310.950 604.050 311.400 ;
        RECT 613.950 312.600 616.050 313.050 ;
        RECT 619.950 312.600 622.050 313.050 ;
        RECT 631.950 312.600 634.050 313.050 ;
        RECT 613.950 311.400 634.050 312.600 ;
        RECT 613.950 310.950 616.050 311.400 ;
        RECT 619.950 310.950 622.050 311.400 ;
        RECT 631.950 310.950 634.050 311.400 ;
        RECT 655.950 312.600 658.050 313.050 ;
        RECT 670.950 312.600 673.050 313.050 ;
        RECT 682.950 312.600 685.050 313.050 ;
        RECT 655.950 311.400 673.050 312.600 ;
        RECT 655.950 310.950 658.050 311.400 ;
        RECT 670.950 310.950 673.050 311.400 ;
        RECT 674.400 311.400 685.050 312.600 ;
        RECT 674.400 310.050 675.600 311.400 ;
        RECT 682.950 310.950 685.050 311.400 ;
        RECT 730.950 312.600 733.050 313.050 ;
        RECT 736.950 312.600 739.050 313.050 ;
        RECT 751.950 312.600 754.050 313.050 ;
        RECT 776.400 312.600 777.600 313.950 ;
        RECT 730.950 311.400 739.050 312.600 ;
        RECT 730.950 310.950 733.050 311.400 ;
        RECT 736.950 310.950 739.050 311.400 ;
        RECT 740.400 311.400 754.050 312.600 ;
        RECT 740.400 310.050 741.600 311.400 ;
        RECT 751.950 310.950 754.050 311.400 ;
        RECT 773.400 311.400 777.600 312.600 ;
        RECT 787.950 312.600 790.050 313.050 ;
        RECT 802.950 312.600 805.050 313.050 ;
        RECT 787.950 311.400 805.050 312.600 ;
        RECT 773.400 310.050 774.600 311.400 ;
        RECT 787.950 310.950 790.050 311.400 ;
        RECT 802.950 310.950 805.050 311.400 ;
        RECT 845.400 310.050 846.600 314.400 ;
        RECT 850.950 313.950 853.050 314.400 ;
        RECT 37.950 307.950 40.050 310.050 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 58.950 309.600 61.050 310.050 ;
        RECT 70.950 309.600 73.050 310.050 ;
        RECT 58.950 308.400 73.050 309.600 ;
        RECT 58.950 307.950 61.050 308.400 ;
        RECT 70.950 307.950 73.050 308.400 ;
        RECT 121.950 309.600 124.050 310.050 ;
        RECT 136.950 309.600 139.050 310.050 ;
        RECT 121.950 308.400 139.050 309.600 ;
        RECT 121.950 307.950 124.050 308.400 ;
        RECT 136.950 307.950 139.050 308.400 ;
        RECT 148.950 309.600 151.050 310.050 ;
        RECT 160.950 309.600 163.050 310.050 ;
        RECT 178.950 309.600 181.050 310.050 ;
        RECT 148.950 308.400 181.050 309.600 ;
        RECT 148.950 307.950 151.050 308.400 ;
        RECT 160.950 307.950 163.050 308.400 ;
        RECT 178.950 307.950 181.050 308.400 ;
        RECT 184.950 309.600 187.050 310.050 ;
        RECT 190.950 309.600 193.050 310.050 ;
        RECT 205.950 309.600 208.050 310.050 ;
        RECT 184.950 308.400 208.050 309.600 ;
        RECT 184.950 307.950 187.050 308.400 ;
        RECT 190.950 307.950 193.050 308.400 ;
        RECT 205.950 307.950 208.050 308.400 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 229.950 309.600 232.050 310.050 ;
        RECT 244.950 309.600 247.050 310.050 ;
        RECT 229.950 308.400 247.050 309.600 ;
        RECT 229.950 307.950 232.050 308.400 ;
        RECT 244.950 307.950 247.050 308.400 ;
        RECT 250.950 309.600 253.050 310.050 ;
        RECT 280.950 309.600 283.050 310.050 ;
        RECT 250.950 308.400 283.050 309.600 ;
        RECT 250.950 307.950 253.050 308.400 ;
        RECT 280.950 307.950 283.050 308.400 ;
        RECT 286.950 309.600 289.050 310.050 ;
        RECT 307.950 309.600 310.050 310.050 ;
        RECT 286.950 308.400 310.050 309.600 ;
        RECT 286.950 307.950 289.050 308.400 ;
        RECT 307.950 307.950 310.050 308.400 ;
        RECT 310.950 309.600 313.050 310.050 ;
        RECT 316.950 309.600 319.050 310.050 ;
        RECT 310.950 308.400 319.050 309.600 ;
        RECT 310.950 307.950 313.050 308.400 ;
        RECT 316.950 307.950 319.050 308.400 ;
        RECT 370.950 309.600 373.050 310.050 ;
        RECT 391.950 309.600 394.050 310.050 ;
        RECT 370.950 308.400 394.050 309.600 ;
        RECT 370.950 307.950 373.050 308.400 ;
        RECT 391.950 307.950 394.050 308.400 ;
        RECT 430.950 307.950 433.050 310.050 ;
        RECT 436.950 309.600 439.050 310.050 ;
        RECT 454.950 309.600 457.050 310.050 ;
        RECT 436.950 308.400 457.050 309.600 ;
        RECT 436.950 307.950 439.050 308.400 ;
        RECT 454.950 307.950 457.050 308.400 ;
        RECT 484.950 309.600 487.050 310.050 ;
        RECT 490.950 309.600 493.050 310.050 ;
        RECT 484.950 308.400 493.050 309.600 ;
        RECT 484.950 307.950 487.050 308.400 ;
        RECT 490.950 307.950 493.050 308.400 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 574.950 309.600 577.050 310.050 ;
        RECT 598.950 309.600 601.050 310.050 ;
        RECT 601.950 309.600 604.050 310.050 ;
        RECT 574.950 308.400 604.050 309.600 ;
        RECT 574.950 307.950 577.050 308.400 ;
        RECT 598.950 307.950 601.050 308.400 ;
        RECT 601.950 307.950 604.050 308.400 ;
        RECT 628.950 309.600 631.050 310.050 ;
        RECT 637.950 309.600 640.050 310.050 ;
        RECT 628.950 308.400 640.050 309.600 ;
        RECT 628.950 307.950 631.050 308.400 ;
        RECT 637.950 307.950 640.050 308.400 ;
        RECT 658.950 309.600 661.050 310.050 ;
        RECT 664.950 309.600 667.050 310.050 ;
        RECT 658.950 308.400 667.050 309.600 ;
        RECT 658.950 307.950 661.050 308.400 ;
        RECT 664.950 307.950 667.050 308.400 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 679.950 309.600 682.050 310.050 ;
        RECT 694.950 309.600 697.050 310.050 ;
        RECT 679.950 308.400 697.050 309.600 ;
        RECT 679.950 307.950 682.050 308.400 ;
        RECT 694.950 307.950 697.050 308.400 ;
        RECT 712.950 309.600 715.050 310.050 ;
        RECT 733.950 309.600 736.050 310.050 ;
        RECT 712.950 308.400 736.050 309.600 ;
        RECT 712.950 307.950 715.050 308.400 ;
        RECT 733.950 307.950 736.050 308.400 ;
        RECT 739.950 307.950 742.050 310.050 ;
        RECT 772.950 307.950 775.050 310.050 ;
        RECT 775.950 309.600 778.050 310.050 ;
        RECT 796.950 309.600 799.050 310.050 ;
        RECT 775.950 308.400 799.050 309.600 ;
        RECT 775.950 307.950 778.050 308.400 ;
        RECT 796.950 307.950 799.050 308.400 ;
        RECT 826.950 309.600 829.050 310.050 ;
        RECT 826.950 308.400 831.600 309.600 ;
        RECT 826.950 307.950 829.050 308.400 ;
        RECT 28.950 306.600 31.050 307.050 ;
        RECT 34.950 306.600 37.050 307.050 ;
        RECT 28.950 305.400 37.050 306.600 ;
        RECT 28.950 304.950 31.050 305.400 ;
        RECT 34.950 304.950 37.050 305.400 ;
        RECT 38.400 303.600 39.600 307.950 ;
        RECT 44.400 306.600 45.600 307.950 ;
        RECT 76.950 306.600 79.050 307.050 ;
        RECT 44.400 305.400 79.050 306.600 ;
        RECT 76.950 304.950 79.050 305.400 ;
        RECT 115.950 306.600 118.050 307.050 ;
        RECT 127.950 306.600 130.050 307.050 ;
        RECT 115.950 305.400 130.050 306.600 ;
        RECT 115.950 304.950 118.050 305.400 ;
        RECT 127.950 304.950 130.050 305.400 ;
        RECT 133.950 306.600 136.050 307.050 ;
        RECT 157.950 306.600 160.050 307.050 ;
        RECT 133.950 305.400 160.050 306.600 ;
        RECT 133.950 304.950 136.050 305.400 ;
        RECT 157.950 304.950 160.050 305.400 ;
        RECT 163.950 304.950 166.050 307.050 ;
        RECT 247.950 306.600 250.050 307.050 ;
        RECT 253.950 306.600 256.050 307.050 ;
        RECT 247.950 305.400 256.050 306.600 ;
        RECT 247.950 304.950 250.050 305.400 ;
        RECT 253.950 304.950 256.050 305.400 ;
        RECT 262.950 306.600 265.050 307.050 ;
        RECT 310.950 306.600 313.050 307.050 ;
        RECT 262.950 305.400 313.050 306.600 ;
        RECT 262.950 304.950 265.050 305.400 ;
        RECT 310.950 304.950 313.050 305.400 ;
        RECT 343.950 306.600 346.050 307.050 ;
        RECT 478.950 306.600 481.050 307.050 ;
        RECT 496.950 306.600 499.050 307.050 ;
        RECT 343.950 305.400 477.600 306.600 ;
        RECT 343.950 304.950 346.050 305.400 ;
        RECT 43.950 303.600 46.050 304.050 ;
        RECT 52.950 303.600 55.050 304.050 ;
        RECT 38.400 302.400 55.050 303.600 ;
        RECT 43.950 301.950 46.050 302.400 ;
        RECT 52.950 301.950 55.050 302.400 ;
        RECT 61.950 303.600 64.050 304.050 ;
        RECT 106.950 303.600 109.050 304.050 ;
        RECT 61.950 302.400 109.050 303.600 ;
        RECT 61.950 301.950 64.050 302.400 ;
        RECT 106.950 301.950 109.050 302.400 ;
        RECT 121.950 303.600 124.050 304.050 ;
        RECT 139.950 303.600 142.050 304.050 ;
        RECT 121.950 302.400 142.050 303.600 ;
        RECT 121.950 301.950 124.050 302.400 ;
        RECT 139.950 301.950 142.050 302.400 ;
        RECT 142.950 303.600 145.050 304.050 ;
        RECT 164.400 303.600 165.600 304.950 ;
        RECT 241.950 303.600 244.050 304.050 ;
        RECT 142.950 302.400 244.050 303.600 ;
        RECT 142.950 301.950 145.050 302.400 ;
        RECT 241.950 301.950 244.050 302.400 ;
        RECT 250.950 303.600 253.050 304.050 ;
        RECT 274.950 303.600 277.050 304.050 ;
        RECT 352.950 303.600 355.050 304.050 ;
        RECT 250.950 302.400 277.050 303.600 ;
        RECT 250.950 301.950 253.050 302.400 ;
        RECT 274.950 301.950 277.050 302.400 ;
        RECT 278.400 302.400 355.050 303.600 ;
        RECT 16.950 300.600 19.050 301.050 ;
        RECT 278.400 300.600 279.600 302.400 ;
        RECT 352.950 301.950 355.050 302.400 ;
        RECT 424.950 303.600 427.050 304.050 ;
        RECT 457.950 303.600 460.050 304.050 ;
        RECT 424.950 302.400 460.050 303.600 ;
        RECT 476.400 303.600 477.600 305.400 ;
        RECT 478.950 305.400 499.050 306.600 ;
        RECT 478.950 304.950 481.050 305.400 ;
        RECT 496.950 304.950 499.050 305.400 ;
        RECT 541.950 306.600 544.050 307.050 ;
        RECT 571.950 306.600 574.050 307.050 ;
        RECT 589.950 306.600 592.050 307.050 ;
        RECT 541.950 305.400 592.050 306.600 ;
        RECT 541.950 304.950 544.050 305.400 ;
        RECT 571.950 304.950 574.050 305.400 ;
        RECT 589.950 304.950 592.050 305.400 ;
        RECT 607.950 306.600 610.050 307.050 ;
        RECT 616.950 306.600 619.050 307.050 ;
        RECT 607.950 305.400 619.050 306.600 ;
        RECT 607.950 304.950 610.050 305.400 ;
        RECT 616.950 304.950 619.050 305.400 ;
        RECT 691.950 306.600 694.050 307.050 ;
        RECT 709.950 306.600 712.050 307.050 ;
        RECT 727.950 306.600 730.050 307.050 ;
        RECT 691.950 305.400 730.050 306.600 ;
        RECT 691.950 304.950 694.050 305.400 ;
        RECT 709.950 304.950 712.050 305.400 ;
        RECT 727.950 304.950 730.050 305.400 ;
        RECT 760.950 306.600 763.050 307.050 ;
        RECT 778.950 306.600 781.050 307.050 ;
        RECT 760.950 305.400 781.050 306.600 ;
        RECT 760.950 304.950 763.050 305.400 ;
        RECT 778.950 304.950 781.050 305.400 ;
        RECT 820.950 306.600 823.050 307.050 ;
        RECT 826.950 306.600 829.050 307.050 ;
        RECT 820.950 305.400 829.050 306.600 ;
        RECT 830.400 306.600 831.600 308.400 ;
        RECT 844.950 307.950 847.050 310.050 ;
        RECT 854.400 307.050 855.600 317.400 ;
        RECT 859.950 315.600 862.050 316.050 ;
        RECT 857.400 314.400 862.050 315.600 ;
        RECT 857.400 310.050 858.600 314.400 ;
        RECT 859.950 313.950 862.050 314.400 ;
        RECT 859.950 312.600 862.050 313.050 ;
        RECT 863.400 312.600 864.600 317.400 ;
        RECT 859.950 311.400 864.600 312.600 ;
        RECT 859.950 310.950 862.050 311.400 ;
        RECT 856.950 307.950 859.050 310.050 ;
        RECT 850.950 306.600 853.050 307.050 ;
        RECT 830.400 305.400 853.050 306.600 ;
        RECT 820.950 304.950 823.050 305.400 ;
        RECT 826.950 304.950 829.050 305.400 ;
        RECT 850.950 304.950 853.050 305.400 ;
        RECT 853.950 304.950 856.050 307.050 ;
        RECT 859.950 306.600 862.050 307.050 ;
        RECT 865.950 306.600 868.050 307.050 ;
        RECT 859.950 305.400 868.050 306.600 ;
        RECT 859.950 304.950 862.050 305.400 ;
        RECT 865.950 304.950 868.050 305.400 ;
        RECT 538.950 303.600 541.050 304.050 ;
        RECT 547.950 303.600 550.050 304.050 ;
        RECT 476.400 302.400 550.050 303.600 ;
        RECT 424.950 301.950 427.050 302.400 ;
        RECT 457.950 301.950 460.050 302.400 ;
        RECT 538.950 301.950 541.050 302.400 ;
        RECT 547.950 301.950 550.050 302.400 ;
        RECT 565.950 303.600 568.050 304.050 ;
        RECT 640.950 303.600 643.050 304.050 ;
        RECT 565.950 302.400 643.050 303.600 ;
        RECT 565.950 301.950 568.050 302.400 ;
        RECT 640.950 301.950 643.050 302.400 ;
        RECT 691.950 303.600 694.050 304.050 ;
        RECT 706.950 303.600 709.050 304.050 ;
        RECT 691.950 302.400 709.050 303.600 ;
        RECT 691.950 301.950 694.050 302.400 ;
        RECT 706.950 301.950 709.050 302.400 ;
        RECT 712.950 303.600 715.050 304.050 ;
        RECT 721.950 303.600 724.050 304.050 ;
        RECT 712.950 302.400 724.050 303.600 ;
        RECT 712.950 301.950 715.050 302.400 ;
        RECT 721.950 301.950 724.050 302.400 ;
        RECT 751.950 303.600 754.050 304.050 ;
        RECT 784.950 303.600 787.050 304.050 ;
        RECT 751.950 302.400 787.050 303.600 ;
        RECT 751.950 301.950 754.050 302.400 ;
        RECT 784.950 301.950 787.050 302.400 ;
        RECT 811.950 303.600 814.050 304.050 ;
        RECT 820.950 303.600 823.050 304.050 ;
        RECT 856.950 303.600 859.050 304.050 ;
        RECT 811.950 302.400 859.050 303.600 ;
        RECT 811.950 301.950 814.050 302.400 ;
        RECT 820.950 301.950 823.050 302.400 ;
        RECT 856.950 301.950 859.050 302.400 ;
        RECT 16.950 299.400 279.600 300.600 ;
        RECT 343.950 300.600 346.050 301.050 ;
        RECT 355.950 300.600 358.050 301.050 ;
        RECT 343.950 299.400 358.050 300.600 ;
        RECT 16.950 298.950 19.050 299.400 ;
        RECT 343.950 298.950 346.050 299.400 ;
        RECT 355.950 298.950 358.050 299.400 ;
        RECT 457.950 300.600 460.050 301.050 ;
        RECT 550.950 300.600 553.050 301.050 ;
        RECT 586.950 300.600 589.050 301.050 ;
        RECT 457.950 299.400 589.050 300.600 ;
        RECT 457.950 298.950 460.050 299.400 ;
        RECT 550.950 298.950 553.050 299.400 ;
        RECT 586.950 298.950 589.050 299.400 ;
        RECT 589.950 300.600 592.050 301.050 ;
        RECT 697.950 300.600 700.050 301.050 ;
        RECT 589.950 299.400 700.050 300.600 ;
        RECT 589.950 298.950 592.050 299.400 ;
        RECT 697.950 298.950 700.050 299.400 ;
        RECT 220.950 297.600 223.050 298.050 ;
        RECT 256.950 297.600 259.050 298.050 ;
        RECT 220.950 296.400 259.050 297.600 ;
        RECT 220.950 295.950 223.050 296.400 ;
        RECT 256.950 295.950 259.050 296.400 ;
        RECT 301.950 297.600 304.050 298.050 ;
        RECT 487.950 297.600 490.050 298.050 ;
        RECT 301.950 296.400 490.050 297.600 ;
        RECT 301.950 295.950 304.050 296.400 ;
        RECT 487.950 295.950 490.050 296.400 ;
        RECT 517.950 297.600 520.050 298.050 ;
        RECT 556.950 297.600 559.050 298.050 ;
        RECT 517.950 296.400 559.050 297.600 ;
        RECT 517.950 295.950 520.050 296.400 ;
        RECT 556.950 295.950 559.050 296.400 ;
        RECT 643.950 297.600 646.050 298.050 ;
        RECT 853.950 297.600 856.050 298.050 ;
        RECT 643.950 296.400 856.050 297.600 ;
        RECT 643.950 295.950 646.050 296.400 ;
        RECT 853.950 295.950 856.050 296.400 ;
        RECT 40.950 294.600 43.050 295.050 ;
        RECT 49.950 294.600 52.050 295.050 ;
        RECT 40.950 293.400 52.050 294.600 ;
        RECT 40.950 292.950 43.050 293.400 ;
        RECT 49.950 292.950 52.050 293.400 ;
        RECT 274.950 294.600 277.050 295.050 ;
        RECT 337.950 294.600 340.050 295.050 ;
        RECT 274.950 293.400 340.050 294.600 ;
        RECT 274.950 292.950 277.050 293.400 ;
        RECT 337.950 292.950 340.050 293.400 ;
        RECT 391.950 294.600 394.050 295.050 ;
        RECT 415.950 294.600 418.050 295.050 ;
        RECT 460.950 294.600 463.050 295.050 ;
        RECT 643.950 294.600 646.050 295.050 ;
        RECT 391.950 293.400 646.050 294.600 ;
        RECT 391.950 292.950 394.050 293.400 ;
        RECT 415.950 292.950 418.050 293.400 ;
        RECT 460.950 292.950 463.050 293.400 ;
        RECT 643.950 292.950 646.050 293.400 ;
        RECT 55.950 291.600 58.050 292.050 ;
        RECT 97.950 291.600 100.050 292.050 ;
        RECT 55.950 290.400 100.050 291.600 ;
        RECT 55.950 289.950 58.050 290.400 ;
        RECT 97.950 289.950 100.050 290.400 ;
        RECT 208.950 291.600 211.050 292.050 ;
        RECT 235.950 291.600 238.050 292.050 ;
        RECT 208.950 290.400 238.050 291.600 ;
        RECT 208.950 289.950 211.050 290.400 ;
        RECT 235.950 289.950 238.050 290.400 ;
        RECT 262.950 291.600 265.050 292.050 ;
        RECT 295.950 291.600 298.050 292.050 ;
        RECT 262.950 290.400 298.050 291.600 ;
        RECT 262.950 289.950 265.050 290.400 ;
        RECT 295.950 289.950 298.050 290.400 ;
        RECT 307.950 291.600 310.050 292.050 ;
        RECT 349.950 291.600 352.050 292.050 ;
        RECT 307.950 290.400 352.050 291.600 ;
        RECT 307.950 289.950 310.050 290.400 ;
        RECT 349.950 289.950 352.050 290.400 ;
        RECT 388.950 291.600 391.050 292.050 ;
        RECT 406.950 291.600 409.050 292.050 ;
        RECT 388.950 290.400 409.050 291.600 ;
        RECT 388.950 289.950 391.050 290.400 ;
        RECT 406.950 289.950 409.050 290.400 ;
        RECT 451.950 291.600 454.050 292.050 ;
        RECT 475.950 291.600 478.050 292.050 ;
        RECT 451.950 290.400 478.050 291.600 ;
        RECT 451.950 289.950 454.050 290.400 ;
        RECT 475.950 289.950 478.050 290.400 ;
        RECT 544.950 291.600 547.050 292.050 ;
        RECT 613.950 291.600 616.050 292.050 ;
        RECT 544.950 290.400 636.600 291.600 ;
        RECT 544.950 289.950 547.050 290.400 ;
        RECT 613.950 289.950 616.050 290.400 ;
        RECT 286.950 288.600 289.050 289.050 ;
        RECT 523.950 288.600 526.050 289.050 ;
        RECT 286.950 287.400 526.050 288.600 ;
        RECT 286.950 286.950 289.050 287.400 ;
        RECT 523.950 286.950 526.050 287.400 ;
        RECT 529.950 288.600 532.050 289.050 ;
        RECT 622.950 288.600 625.050 289.050 ;
        RECT 529.950 287.400 625.050 288.600 ;
        RECT 635.400 288.600 636.600 290.400 ;
        RECT 646.950 288.600 649.050 289.050 ;
        RECT 661.950 288.600 664.050 289.050 ;
        RECT 635.400 287.400 664.050 288.600 ;
        RECT 529.950 286.950 532.050 287.400 ;
        RECT 622.950 286.950 625.050 287.400 ;
        RECT 646.950 286.950 649.050 287.400 ;
        RECT 661.950 286.950 664.050 287.400 ;
        RECT 760.950 288.600 763.050 289.050 ;
        RECT 787.950 288.600 790.050 289.050 ;
        RECT 760.950 287.400 790.050 288.600 ;
        RECT 760.950 286.950 763.050 287.400 ;
        RECT 787.950 286.950 790.050 287.400 ;
        RECT 361.950 285.600 364.050 286.050 ;
        RECT 382.950 285.600 385.050 286.050 ;
        RECT 361.950 284.400 385.050 285.600 ;
        RECT 361.950 283.950 364.050 284.400 ;
        RECT 382.950 283.950 385.050 284.400 ;
        RECT 403.950 285.600 406.050 286.050 ;
        RECT 541.950 285.600 544.050 286.050 ;
        RECT 403.950 284.400 544.050 285.600 ;
        RECT 403.950 283.950 406.050 284.400 ;
        RECT 541.950 283.950 544.050 284.400 ;
        RECT 553.950 285.600 556.050 286.050 ;
        RECT 619.950 285.600 622.050 286.050 ;
        RECT 553.950 284.400 622.050 285.600 ;
        RECT 553.950 283.950 556.050 284.400 ;
        RECT 619.950 283.950 622.050 284.400 ;
        RECT 631.950 285.600 634.050 286.050 ;
        RECT 793.950 285.600 796.050 286.050 ;
        RECT 631.950 284.400 796.050 285.600 ;
        RECT 631.950 283.950 634.050 284.400 ;
        RECT 793.950 283.950 796.050 284.400 ;
        RECT 58.950 282.600 61.050 283.050 ;
        RECT 76.950 282.600 79.050 283.050 ;
        RECT 58.950 281.400 79.050 282.600 ;
        RECT 58.950 280.950 61.050 281.400 ;
        RECT 76.950 280.950 79.050 281.400 ;
        RECT 151.950 282.600 154.050 283.050 ;
        RECT 289.950 282.600 292.050 283.050 ;
        RECT 151.950 281.400 292.050 282.600 ;
        RECT 151.950 280.950 154.050 281.400 ;
        RECT 289.950 280.950 292.050 281.400 ;
        RECT 295.950 282.600 298.050 283.050 ;
        RECT 418.950 282.600 421.050 283.050 ;
        RECT 295.950 281.400 421.050 282.600 ;
        RECT 295.950 280.950 298.050 281.400 ;
        RECT 418.950 280.950 421.050 281.400 ;
        RECT 421.950 282.600 424.050 283.050 ;
        RECT 472.950 282.600 475.050 283.050 ;
        RECT 421.950 281.400 475.050 282.600 ;
        RECT 421.950 280.950 424.050 281.400 ;
        RECT 472.950 280.950 475.050 281.400 ;
        RECT 568.950 282.600 571.050 283.050 ;
        RECT 604.950 282.600 607.050 283.050 ;
        RECT 568.950 281.400 607.050 282.600 ;
        RECT 568.950 280.950 571.050 281.400 ;
        RECT 604.950 280.950 607.050 281.400 ;
        RECT 607.950 282.600 610.050 283.050 ;
        RECT 625.950 282.600 628.050 283.050 ;
        RECT 706.950 282.600 709.050 283.050 ;
        RECT 607.950 281.400 709.050 282.600 ;
        RECT 607.950 280.950 610.050 281.400 ;
        RECT 625.950 280.950 628.050 281.400 ;
        RECT 706.950 280.950 709.050 281.400 ;
        RECT 718.950 282.600 721.050 283.050 ;
        RECT 823.950 282.600 826.050 283.050 ;
        RECT 718.950 281.400 826.050 282.600 ;
        RECT 718.950 280.950 721.050 281.400 ;
        RECT 823.950 280.950 826.050 281.400 ;
        RECT 31.950 279.600 34.050 280.050 ;
        RECT 106.950 279.600 109.050 280.050 ;
        RECT 31.950 278.400 109.050 279.600 ;
        RECT 31.950 277.950 34.050 278.400 ;
        RECT 106.950 277.950 109.050 278.400 ;
        RECT 253.950 279.600 256.050 280.050 ;
        RECT 277.950 279.600 280.050 280.050 ;
        RECT 253.950 278.400 280.050 279.600 ;
        RECT 253.950 277.950 256.050 278.400 ;
        RECT 277.950 277.950 280.050 278.400 ;
        RECT 421.950 279.600 424.050 280.050 ;
        RECT 448.950 279.600 451.050 280.050 ;
        RECT 421.950 278.400 451.050 279.600 ;
        RECT 421.950 277.950 424.050 278.400 ;
        RECT 448.950 277.950 451.050 278.400 ;
        RECT 523.950 279.600 526.050 280.050 ;
        RECT 631.950 279.600 634.050 280.050 ;
        RECT 523.950 278.400 634.050 279.600 ;
        RECT 523.950 277.950 526.050 278.400 ;
        RECT 631.950 277.950 634.050 278.400 ;
        RECT 706.950 279.600 709.050 280.050 ;
        RECT 733.950 279.600 736.050 280.050 ;
        RECT 787.950 279.600 790.050 280.050 ;
        RECT 799.950 279.600 802.050 280.050 ;
        RECT 706.950 278.400 802.050 279.600 ;
        RECT 706.950 277.950 709.050 278.400 ;
        RECT 733.950 277.950 736.050 278.400 ;
        RECT 787.950 277.950 790.050 278.400 ;
        RECT 799.950 277.950 802.050 278.400 ;
        RECT 802.950 279.600 805.050 280.050 ;
        RECT 808.950 279.600 811.050 280.050 ;
        RECT 802.950 278.400 811.050 279.600 ;
        RECT 802.950 277.950 805.050 278.400 ;
        RECT 808.950 277.950 811.050 278.400 ;
        RECT 28.950 276.600 31.050 277.050 ;
        RECT 49.950 276.600 52.050 277.050 ;
        RECT 73.950 276.600 76.050 277.050 ;
        RECT 28.950 275.400 76.050 276.600 ;
        RECT 28.950 274.950 31.050 275.400 ;
        RECT 49.950 274.950 52.050 275.400 ;
        RECT 73.950 274.950 76.050 275.400 ;
        RECT 76.950 274.950 79.050 277.050 ;
        RECT 106.950 276.600 109.050 277.050 ;
        RECT 169.950 276.600 172.050 277.050 ;
        RECT 106.950 275.400 172.050 276.600 ;
        RECT 106.950 274.950 109.050 275.400 ;
        RECT 169.950 274.950 172.050 275.400 ;
        RECT 184.950 276.600 187.050 277.050 ;
        RECT 316.950 276.600 319.050 277.050 ;
        RECT 184.950 275.400 319.050 276.600 ;
        RECT 184.950 274.950 187.050 275.400 ;
        RECT 316.950 274.950 319.050 275.400 ;
        RECT 331.950 276.600 334.050 277.050 ;
        RECT 391.950 276.600 394.050 277.050 ;
        RECT 331.950 275.400 394.050 276.600 ;
        RECT 331.950 274.950 334.050 275.400 ;
        RECT 391.950 274.950 394.050 275.400 ;
        RECT 412.950 276.600 415.050 277.050 ;
        RECT 505.950 276.600 508.050 277.050 ;
        RECT 541.950 276.600 544.050 277.050 ;
        RECT 412.950 275.400 544.050 276.600 ;
        RECT 412.950 274.950 415.050 275.400 ;
        RECT 505.950 274.950 508.050 275.400 ;
        RECT 541.950 274.950 544.050 275.400 ;
        RECT 577.950 276.600 580.050 277.050 ;
        RECT 601.950 276.600 604.050 277.050 ;
        RECT 577.950 275.400 604.050 276.600 ;
        RECT 577.950 274.950 580.050 275.400 ;
        RECT 601.950 274.950 604.050 275.400 ;
        RECT 616.950 276.600 619.050 277.050 ;
        RECT 625.950 276.600 628.050 277.050 ;
        RECT 640.950 276.600 643.050 277.050 ;
        RECT 616.950 275.400 643.050 276.600 ;
        RECT 616.950 274.950 619.050 275.400 ;
        RECT 625.950 274.950 628.050 275.400 ;
        RECT 640.950 274.950 643.050 275.400 ;
        RECT 652.950 276.600 655.050 277.050 ;
        RECT 667.950 276.600 670.050 277.050 ;
        RECT 652.950 275.400 670.050 276.600 ;
        RECT 652.950 274.950 655.050 275.400 ;
        RECT 667.950 274.950 670.050 275.400 ;
        RECT 673.950 276.600 676.050 277.050 ;
        RECT 682.950 276.600 685.050 277.050 ;
        RECT 673.950 275.400 685.050 276.600 ;
        RECT 673.950 274.950 676.050 275.400 ;
        RECT 682.950 274.950 685.050 275.400 ;
        RECT 700.950 276.600 703.050 277.050 ;
        RECT 727.950 276.600 730.050 277.050 ;
        RECT 700.950 275.400 730.050 276.600 ;
        RECT 700.950 274.950 703.050 275.400 ;
        RECT 727.950 274.950 730.050 275.400 ;
        RECT 745.950 276.600 748.050 277.050 ;
        RECT 754.950 276.600 757.050 277.050 ;
        RECT 745.950 275.400 757.050 276.600 ;
        RECT 745.950 274.950 748.050 275.400 ;
        RECT 754.950 274.950 757.050 275.400 ;
        RECT 799.950 276.600 802.050 277.050 ;
        RECT 814.950 276.600 817.050 277.050 ;
        RECT 799.950 275.400 817.050 276.600 ;
        RECT 799.950 274.950 802.050 275.400 ;
        RECT 814.950 274.950 817.050 275.400 ;
        RECT 16.950 273.600 19.050 274.050 ;
        RECT 31.950 273.600 34.050 274.050 ;
        RECT 16.950 272.400 34.050 273.600 ;
        RECT 16.950 271.950 19.050 272.400 ;
        RECT 31.950 271.950 34.050 272.400 ;
        RECT 34.950 273.600 37.050 274.050 ;
        RECT 34.950 272.400 39.600 273.600 ;
        RECT 34.950 271.950 37.050 272.400 ;
        RECT 13.950 270.600 16.050 271.050 ;
        RECT 28.950 270.600 31.050 271.050 ;
        RECT 13.950 269.400 31.050 270.600 ;
        RECT 13.950 268.950 16.050 269.400 ;
        RECT 28.950 268.950 31.050 269.400 ;
        RECT 34.950 268.950 37.050 271.050 ;
        RECT 19.950 267.600 22.050 268.050 ;
        RECT 35.400 267.600 36.600 268.950 ;
        RECT 19.950 266.400 36.600 267.600 ;
        RECT 19.950 265.950 22.050 266.400 ;
        RECT 16.950 264.600 19.050 265.050 ;
        RECT 31.950 264.600 34.050 265.050 ;
        RECT 16.950 263.400 34.050 264.600 ;
        RECT 16.950 262.950 19.050 263.400 ;
        RECT 31.950 262.950 34.050 263.400 ;
        RECT 31.950 261.600 34.050 262.050 ;
        RECT 38.400 261.600 39.600 272.400 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 61.950 271.950 64.050 274.050 ;
        RECT 56.400 270.600 57.600 271.950 ;
        RECT 53.400 269.400 57.600 270.600 ;
        RECT 53.400 268.050 54.600 269.400 ;
        RECT 52.950 265.950 55.050 268.050 ;
        RECT 55.950 267.600 58.050 268.050 ;
        RECT 62.400 267.600 63.600 271.950 ;
        RECT 55.950 266.400 63.600 267.600 ;
        RECT 77.400 267.600 78.600 274.950 ;
        RECT 79.950 273.600 82.050 274.050 ;
        RECT 142.950 273.600 145.050 274.050 ;
        RECT 79.950 272.400 145.050 273.600 ;
        RECT 79.950 271.950 82.050 272.400 ;
        RECT 142.950 271.950 145.050 272.400 ;
        RECT 277.950 273.600 280.050 274.050 ;
        RECT 292.950 273.600 295.050 274.050 ;
        RECT 322.950 273.600 325.050 274.050 ;
        RECT 277.950 272.400 325.050 273.600 ;
        RECT 277.950 271.950 280.050 272.400 ;
        RECT 292.950 271.950 295.050 272.400 ;
        RECT 322.950 271.950 325.050 272.400 ;
        RECT 328.950 273.600 331.050 274.050 ;
        RECT 337.950 273.600 340.050 274.050 ;
        RECT 328.950 272.400 340.050 273.600 ;
        RECT 328.950 271.950 331.050 272.400 ;
        RECT 337.950 271.950 340.050 272.400 ;
        RECT 415.950 273.600 418.050 274.050 ;
        RECT 424.950 273.600 427.050 274.050 ;
        RECT 463.950 273.600 466.050 274.050 ;
        RECT 415.950 272.400 427.050 273.600 ;
        RECT 415.950 271.950 418.050 272.400 ;
        RECT 424.950 271.950 427.050 272.400 ;
        RECT 458.400 272.400 466.050 273.600 ;
        RECT 82.950 270.600 85.050 271.050 ;
        RECT 88.950 270.600 91.050 271.050 ;
        RECT 124.950 270.600 127.050 271.050 ;
        RECT 82.950 269.400 127.050 270.600 ;
        RECT 82.950 268.950 85.050 269.400 ;
        RECT 88.950 268.950 91.050 269.400 ;
        RECT 124.950 268.950 127.050 269.400 ;
        RECT 139.950 270.600 142.050 271.050 ;
        RECT 154.950 270.600 157.050 271.050 ;
        RECT 139.950 269.400 157.050 270.600 ;
        RECT 139.950 268.950 142.050 269.400 ;
        RECT 154.950 268.950 157.050 269.400 ;
        RECT 163.950 270.600 166.050 271.050 ;
        RECT 175.950 270.600 178.050 271.050 ;
        RECT 184.950 270.600 187.050 271.050 ;
        RECT 163.950 269.400 187.050 270.600 ;
        RECT 163.950 268.950 166.050 269.400 ;
        RECT 175.950 268.950 178.050 269.400 ;
        RECT 184.950 268.950 187.050 269.400 ;
        RECT 190.950 270.600 193.050 271.050 ;
        RECT 199.950 270.600 202.050 271.050 ;
        RECT 190.950 269.400 202.050 270.600 ;
        RECT 190.950 268.950 193.050 269.400 ;
        RECT 199.950 268.950 202.050 269.400 ;
        RECT 244.950 270.600 247.050 271.050 ;
        RECT 262.950 270.600 265.050 271.050 ;
        RECT 244.950 269.400 265.050 270.600 ;
        RECT 244.950 268.950 247.050 269.400 ;
        RECT 262.950 268.950 265.050 269.400 ;
        RECT 334.950 270.600 337.050 271.050 ;
        RECT 340.950 270.600 343.050 271.050 ;
        RECT 334.950 269.400 343.050 270.600 ;
        RECT 334.950 268.950 337.050 269.400 ;
        RECT 340.950 268.950 343.050 269.400 ;
        RECT 418.950 270.600 421.050 271.050 ;
        RECT 427.950 270.600 430.050 271.050 ;
        RECT 418.950 269.400 430.050 270.600 ;
        RECT 418.950 268.950 421.050 269.400 ;
        RECT 427.950 268.950 430.050 269.400 ;
        RECT 445.950 270.600 448.050 271.050 ;
        RECT 458.400 270.600 459.600 272.400 ;
        RECT 463.950 271.950 466.050 272.400 ;
        RECT 466.950 273.600 469.050 274.050 ;
        RECT 496.950 273.600 499.050 274.050 ;
        RECT 466.950 272.400 499.050 273.600 ;
        RECT 466.950 271.950 469.050 272.400 ;
        RECT 496.950 271.950 499.050 272.400 ;
        RECT 505.950 273.600 508.050 274.050 ;
        RECT 511.950 273.600 514.050 274.050 ;
        RECT 505.950 272.400 514.050 273.600 ;
        RECT 505.950 271.950 508.050 272.400 ;
        RECT 511.950 271.950 514.050 272.400 ;
        RECT 535.950 273.600 538.050 274.050 ;
        RECT 592.950 273.600 595.050 274.050 ;
        RECT 535.950 272.400 595.050 273.600 ;
        RECT 535.950 271.950 538.050 272.400 ;
        RECT 592.950 271.950 595.050 272.400 ;
        RECT 619.950 273.600 622.050 274.050 ;
        RECT 709.950 273.600 712.050 274.050 ;
        RECT 619.950 272.400 712.050 273.600 ;
        RECT 619.950 271.950 622.050 272.400 ;
        RECT 709.950 271.950 712.050 272.400 ;
        RECT 739.950 273.600 742.050 274.050 ;
        RECT 748.950 273.600 751.050 274.050 ;
        RECT 739.950 272.400 751.050 273.600 ;
        RECT 739.950 271.950 742.050 272.400 ;
        RECT 748.950 271.950 751.050 272.400 ;
        RECT 445.950 269.400 459.600 270.600 ;
        RECT 508.950 270.600 511.050 271.050 ;
        RECT 523.950 270.600 526.050 271.050 ;
        RECT 508.950 269.400 526.050 270.600 ;
        RECT 445.950 268.950 448.050 269.400 ;
        RECT 508.950 268.950 511.050 269.400 ;
        RECT 523.950 268.950 526.050 269.400 ;
        RECT 592.950 268.950 595.050 271.050 ;
        RECT 598.950 270.600 601.050 271.050 ;
        RECT 616.950 270.600 619.050 271.050 ;
        RECT 598.950 269.400 619.050 270.600 ;
        RECT 598.950 268.950 601.050 269.400 ;
        RECT 616.950 268.950 619.050 269.400 ;
        RECT 634.950 270.600 637.050 271.050 ;
        RECT 667.950 270.600 670.050 271.050 ;
        RECT 688.950 270.600 691.050 271.050 ;
        RECT 634.950 269.400 691.050 270.600 ;
        RECT 634.950 268.950 637.050 269.400 ;
        RECT 667.950 268.950 670.050 269.400 ;
        RECT 688.950 268.950 691.050 269.400 ;
        RECT 718.950 270.600 721.050 271.050 ;
        RECT 736.950 270.600 739.050 271.050 ;
        RECT 745.950 270.600 748.050 271.050 ;
        RECT 769.950 270.600 772.050 271.050 ;
        RECT 718.950 269.400 723.600 270.600 ;
        RECT 718.950 268.950 721.050 269.400 ;
        RECT 82.950 267.600 85.050 268.050 ;
        RECT 77.400 266.400 85.050 267.600 ;
        RECT 55.950 265.950 58.050 266.400 ;
        RECT 82.950 265.950 85.050 266.400 ;
        RECT 103.950 267.600 106.050 268.050 ;
        RECT 121.950 267.600 124.050 268.050 ;
        RECT 145.950 267.600 148.050 268.050 ;
        RECT 103.950 266.400 120.600 267.600 ;
        RECT 103.950 265.950 106.050 266.400 ;
        RECT 61.950 264.600 64.050 265.050 ;
        RECT 106.950 264.600 109.050 265.050 ;
        RECT 115.950 264.600 118.050 265.050 ;
        RECT 61.950 263.400 102.600 264.600 ;
        RECT 61.950 262.950 64.050 263.400 ;
        RECT 31.950 260.400 39.600 261.600 ;
        RECT 61.950 261.600 64.050 262.050 ;
        RECT 70.950 261.600 73.050 262.050 ;
        RECT 61.950 260.400 73.050 261.600 ;
        RECT 31.950 259.950 34.050 260.400 ;
        RECT 61.950 259.950 64.050 260.400 ;
        RECT 70.950 259.950 73.050 260.400 ;
        RECT 76.950 261.600 79.050 262.050 ;
        RECT 101.400 261.600 102.600 263.400 ;
        RECT 106.950 263.400 118.050 264.600 ;
        RECT 119.400 264.600 120.600 266.400 ;
        RECT 121.950 266.400 148.050 267.600 ;
        RECT 121.950 265.950 124.050 266.400 ;
        RECT 145.950 265.950 148.050 266.400 ;
        RECT 166.950 267.600 169.050 268.050 ;
        RECT 187.950 267.600 190.050 268.050 ;
        RECT 208.950 267.600 211.050 268.050 ;
        RECT 166.950 266.400 211.050 267.600 ;
        RECT 166.950 265.950 169.050 266.400 ;
        RECT 187.950 265.950 190.050 266.400 ;
        RECT 208.950 265.950 211.050 266.400 ;
        RECT 223.950 267.600 226.050 268.050 ;
        RECT 229.950 267.600 232.050 268.050 ;
        RECT 232.950 267.600 235.050 268.050 ;
        RECT 223.950 266.400 235.050 267.600 ;
        RECT 223.950 265.950 226.050 266.400 ;
        RECT 229.950 265.950 232.050 266.400 ;
        RECT 232.950 265.950 235.050 266.400 ;
        RECT 241.950 267.600 244.050 268.050 ;
        RECT 259.950 267.600 262.050 268.050 ;
        RECT 241.950 266.400 262.050 267.600 ;
        RECT 241.950 265.950 244.050 266.400 ;
        RECT 259.950 265.950 262.050 266.400 ;
        RECT 325.950 267.600 328.050 268.050 ;
        RECT 394.950 267.600 397.050 268.050 ;
        RECT 433.950 267.600 436.050 268.050 ;
        RECT 325.950 266.400 436.050 267.600 ;
        RECT 325.950 265.950 328.050 266.400 ;
        RECT 394.950 265.950 397.050 266.400 ;
        RECT 433.950 265.950 436.050 266.400 ;
        RECT 493.950 267.600 496.050 268.050 ;
        RECT 502.950 267.600 505.050 268.050 ;
        RECT 493.950 266.400 505.050 267.600 ;
        RECT 493.950 265.950 496.050 266.400 ;
        RECT 502.950 265.950 505.050 266.400 ;
        RECT 541.950 267.600 544.050 268.050 ;
        RECT 556.950 267.600 559.050 268.050 ;
        RECT 565.950 267.600 568.050 268.050 ;
        RECT 541.950 266.400 568.050 267.600 ;
        RECT 541.950 265.950 544.050 266.400 ;
        RECT 556.950 265.950 559.050 266.400 ;
        RECT 565.950 265.950 568.050 266.400 ;
        RECT 574.950 267.600 577.050 268.050 ;
        RECT 589.950 267.600 592.050 268.050 ;
        RECT 574.950 266.400 592.050 267.600 ;
        RECT 593.400 267.600 594.600 268.950 ;
        RECT 722.400 268.050 723.600 269.400 ;
        RECT 736.950 269.400 748.050 270.600 ;
        RECT 736.950 268.950 739.050 269.400 ;
        RECT 745.950 268.950 748.050 269.400 ;
        RECT 752.400 269.400 772.050 270.600 ;
        RECT 752.400 268.050 753.600 269.400 ;
        RECT 769.950 268.950 772.050 269.400 ;
        RECT 775.950 270.600 778.050 271.050 ;
        RECT 793.950 270.600 796.050 271.050 ;
        RECT 823.950 270.600 826.050 271.050 ;
        RECT 829.950 270.600 832.050 271.050 ;
        RECT 775.950 269.400 792.600 270.600 ;
        RECT 775.950 268.950 778.050 269.400 ;
        RECT 791.400 268.050 792.600 269.400 ;
        RECT 793.950 269.400 807.600 270.600 ;
        RECT 793.950 268.950 796.050 269.400 ;
        RECT 806.400 268.050 807.600 269.400 ;
        RECT 823.950 269.400 832.050 270.600 ;
        RECT 823.950 268.950 826.050 269.400 ;
        RECT 829.950 268.950 832.050 269.400 ;
        RECT 598.950 267.600 601.050 268.050 ;
        RECT 593.400 266.400 601.050 267.600 ;
        RECT 574.950 265.950 577.050 266.400 ;
        RECT 589.950 265.950 592.050 266.400 ;
        RECT 598.950 265.950 601.050 266.400 ;
        RECT 622.950 267.600 625.050 268.050 ;
        RECT 637.950 267.600 640.050 268.050 ;
        RECT 622.950 266.400 640.050 267.600 ;
        RECT 622.950 265.950 625.050 266.400 ;
        RECT 637.950 265.950 640.050 266.400 ;
        RECT 664.950 267.600 667.050 268.050 ;
        RECT 670.950 267.600 673.050 268.050 ;
        RECT 664.950 266.400 673.050 267.600 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 670.950 265.950 673.050 266.400 ;
        RECT 682.950 267.600 685.050 268.050 ;
        RECT 694.950 267.600 697.050 268.050 ;
        RECT 682.950 266.400 697.050 267.600 ;
        RECT 682.950 265.950 685.050 266.400 ;
        RECT 694.950 265.950 697.050 266.400 ;
        RECT 721.950 265.950 724.050 268.050 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 757.950 267.600 760.050 268.050 ;
        RECT 769.950 267.600 772.050 268.050 ;
        RECT 757.950 266.400 772.050 267.600 ;
        RECT 757.950 265.950 760.050 266.400 ;
        RECT 769.950 265.950 772.050 266.400 ;
        RECT 790.950 265.950 793.050 268.050 ;
        RECT 805.950 265.950 808.050 268.050 ;
        RECT 811.950 267.600 814.050 268.050 ;
        RECT 829.950 267.600 832.050 268.050 ;
        RECT 811.950 266.400 832.050 267.600 ;
        RECT 811.950 265.950 814.050 266.400 ;
        RECT 829.950 265.950 832.050 266.400 ;
        RECT 148.950 264.600 151.050 265.050 ;
        RECT 119.400 263.400 151.050 264.600 ;
        RECT 106.950 262.950 109.050 263.400 ;
        RECT 115.950 262.950 118.050 263.400 ;
        RECT 148.950 262.950 151.050 263.400 ;
        RECT 154.950 264.600 157.050 265.050 ;
        RECT 169.950 264.600 172.050 265.050 ;
        RECT 178.950 264.600 181.050 265.050 ;
        RECT 154.950 263.400 181.050 264.600 ;
        RECT 154.950 262.950 157.050 263.400 ;
        RECT 169.950 262.950 172.050 263.400 ;
        RECT 178.950 262.950 181.050 263.400 ;
        RECT 214.950 264.600 217.050 265.050 ;
        RECT 226.950 264.600 229.050 265.050 ;
        RECT 265.950 264.600 268.050 265.050 ;
        RECT 274.950 264.600 277.050 265.050 ;
        RECT 214.950 263.400 277.050 264.600 ;
        RECT 214.950 262.950 217.050 263.400 ;
        RECT 226.950 262.950 229.050 263.400 ;
        RECT 265.950 262.950 268.050 263.400 ;
        RECT 274.950 262.950 277.050 263.400 ;
        RECT 367.950 264.600 370.050 265.050 ;
        RECT 382.950 264.600 385.050 265.050 ;
        RECT 367.950 263.400 385.050 264.600 ;
        RECT 367.950 262.950 370.050 263.400 ;
        RECT 382.950 262.950 385.050 263.400 ;
        RECT 403.950 264.600 406.050 265.050 ;
        RECT 412.950 264.600 415.050 265.050 ;
        RECT 403.950 263.400 415.050 264.600 ;
        RECT 403.950 262.950 406.050 263.400 ;
        RECT 412.950 262.950 415.050 263.400 ;
        RECT 421.950 264.600 424.050 265.050 ;
        RECT 448.950 264.600 451.050 265.050 ;
        RECT 421.950 263.400 451.050 264.600 ;
        RECT 421.950 262.950 424.050 263.400 ;
        RECT 448.950 262.950 451.050 263.400 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 466.950 264.600 469.050 265.050 ;
        RECT 454.950 263.400 469.050 264.600 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 466.950 262.950 469.050 263.400 ;
        RECT 508.950 264.600 511.050 265.050 ;
        RECT 544.950 264.600 547.050 265.050 ;
        RECT 508.950 263.400 547.050 264.600 ;
        RECT 508.950 262.950 511.050 263.400 ;
        RECT 544.950 262.950 547.050 263.400 ;
        RECT 547.950 264.600 550.050 265.050 ;
        RECT 571.950 264.600 574.050 265.050 ;
        RECT 649.950 264.600 652.050 265.050 ;
        RECT 547.950 263.400 652.050 264.600 ;
        RECT 547.950 262.950 550.050 263.400 ;
        RECT 571.950 262.950 574.050 263.400 ;
        RECT 649.950 262.950 652.050 263.400 ;
        RECT 703.950 264.600 706.050 265.050 ;
        RECT 712.950 264.600 715.050 265.050 ;
        RECT 703.950 263.400 715.050 264.600 ;
        RECT 703.950 262.950 706.050 263.400 ;
        RECT 712.950 262.950 715.050 263.400 ;
        RECT 748.950 264.600 751.050 265.050 ;
        RECT 757.950 264.600 760.050 265.050 ;
        RECT 763.950 264.600 766.050 265.050 ;
        RECT 748.950 263.400 766.050 264.600 ;
        RECT 748.950 262.950 751.050 263.400 ;
        RECT 757.950 262.950 760.050 263.400 ;
        RECT 763.950 262.950 766.050 263.400 ;
        RECT 796.950 264.600 799.050 265.050 ;
        RECT 802.950 264.600 805.050 265.050 ;
        RECT 811.950 264.600 814.050 265.050 ;
        RECT 838.950 264.600 841.050 265.050 ;
        RECT 796.950 263.400 841.050 264.600 ;
        RECT 796.950 262.950 799.050 263.400 ;
        RECT 802.950 262.950 805.050 263.400 ;
        RECT 811.950 262.950 814.050 263.400 ;
        RECT 838.950 262.950 841.050 263.400 ;
        RECT 127.950 261.600 130.050 262.050 ;
        RECT 76.950 260.400 99.600 261.600 ;
        RECT 101.400 260.400 130.050 261.600 ;
        RECT 76.950 259.950 79.050 260.400 ;
        RECT 37.950 258.600 40.050 259.050 ;
        RECT 52.950 258.600 55.050 259.050 ;
        RECT 37.950 257.400 55.050 258.600 ;
        RECT 37.950 256.950 40.050 257.400 ;
        RECT 52.950 256.950 55.050 257.400 ;
        RECT 76.950 258.600 79.050 259.050 ;
        RECT 82.950 258.600 85.050 259.050 ;
        RECT 76.950 257.400 85.050 258.600 ;
        RECT 98.400 258.600 99.600 260.400 ;
        RECT 127.950 259.950 130.050 260.400 ;
        RECT 142.950 261.600 145.050 262.050 ;
        RECT 157.950 261.600 160.050 262.050 ;
        RECT 142.950 260.400 160.050 261.600 ;
        RECT 142.950 259.950 145.050 260.400 ;
        RECT 157.950 259.950 160.050 260.400 ;
        RECT 202.950 261.600 205.050 262.050 ;
        RECT 211.950 261.600 214.050 262.050 ;
        RECT 202.950 260.400 214.050 261.600 ;
        RECT 202.950 259.950 205.050 260.400 ;
        RECT 211.950 259.950 214.050 260.400 ;
        RECT 223.950 261.600 226.050 262.050 ;
        RECT 271.950 261.600 274.050 262.050 ;
        RECT 223.950 260.400 274.050 261.600 ;
        RECT 223.950 259.950 226.050 260.400 ;
        RECT 271.950 259.950 274.050 260.400 ;
        RECT 289.950 261.600 292.050 262.050 ;
        RECT 385.950 261.600 388.050 262.050 ;
        RECT 289.950 260.400 388.050 261.600 ;
        RECT 289.950 259.950 292.050 260.400 ;
        RECT 385.950 259.950 388.050 260.400 ;
        RECT 406.950 261.600 409.050 262.050 ;
        RECT 436.950 261.600 439.050 262.050 ;
        RECT 406.950 260.400 439.050 261.600 ;
        RECT 406.950 259.950 409.050 260.400 ;
        RECT 436.950 259.950 439.050 260.400 ;
        RECT 460.950 261.600 463.050 262.050 ;
        RECT 493.950 261.600 496.050 262.050 ;
        RECT 460.950 260.400 496.050 261.600 ;
        RECT 460.950 259.950 463.050 260.400 ;
        RECT 493.950 259.950 496.050 260.400 ;
        RECT 520.950 261.600 523.050 262.050 ;
        RECT 547.950 261.600 550.050 262.050 ;
        RECT 520.950 260.400 550.050 261.600 ;
        RECT 520.950 259.950 523.050 260.400 ;
        RECT 547.950 259.950 550.050 260.400 ;
        RECT 565.950 261.600 568.050 262.050 ;
        RECT 592.950 261.600 595.050 262.050 ;
        RECT 565.950 260.400 595.050 261.600 ;
        RECT 565.950 259.950 568.050 260.400 ;
        RECT 592.950 259.950 595.050 260.400 ;
        RECT 649.950 261.600 652.050 262.050 ;
        RECT 679.950 261.600 682.050 262.050 ;
        RECT 715.950 261.600 718.050 262.050 ;
        RECT 736.950 261.600 739.050 262.050 ;
        RECT 784.950 261.600 787.050 262.050 ;
        RECT 814.950 261.600 817.050 262.050 ;
        RECT 835.950 261.600 838.050 262.050 ;
        RECT 649.950 260.400 838.050 261.600 ;
        RECT 649.950 259.950 652.050 260.400 ;
        RECT 679.950 259.950 682.050 260.400 ;
        RECT 715.950 259.950 718.050 260.400 ;
        RECT 736.950 259.950 739.050 260.400 ;
        RECT 784.950 259.950 787.050 260.400 ;
        RECT 814.950 259.950 817.050 260.400 ;
        RECT 835.950 259.950 838.050 260.400 ;
        RECT 196.950 258.600 199.050 259.050 ;
        RECT 98.400 257.400 199.050 258.600 ;
        RECT 76.950 256.950 79.050 257.400 ;
        RECT 82.950 256.950 85.050 257.400 ;
        RECT 196.950 256.950 199.050 257.400 ;
        RECT 205.950 258.600 208.050 259.050 ;
        RECT 280.950 258.600 283.050 259.050 ;
        RECT 205.950 257.400 283.050 258.600 ;
        RECT 205.950 256.950 208.050 257.400 ;
        RECT 280.950 256.950 283.050 257.400 ;
        RECT 388.950 258.600 391.050 259.050 ;
        RECT 421.950 258.600 424.050 259.050 ;
        RECT 388.950 257.400 424.050 258.600 ;
        RECT 388.950 256.950 391.050 257.400 ;
        RECT 421.950 256.950 424.050 257.400 ;
        RECT 436.950 258.600 439.050 259.050 ;
        RECT 475.950 258.600 478.050 259.050 ;
        RECT 436.950 257.400 478.050 258.600 ;
        RECT 436.950 256.950 439.050 257.400 ;
        RECT 475.950 256.950 478.050 257.400 ;
        RECT 487.950 258.600 490.050 259.050 ;
        RECT 544.950 258.600 547.050 259.050 ;
        RECT 553.950 258.600 556.050 259.050 ;
        RECT 682.950 258.600 685.050 259.050 ;
        RECT 487.950 257.400 556.050 258.600 ;
        RECT 487.950 256.950 490.050 257.400 ;
        RECT 544.950 256.950 547.050 257.400 ;
        RECT 553.950 256.950 556.050 257.400 ;
        RECT 650.400 257.400 685.050 258.600 ;
        RECT 650.400 256.050 651.600 257.400 ;
        RECT 682.950 256.950 685.050 257.400 ;
        RECT 775.950 258.600 778.050 259.050 ;
        RECT 784.950 258.600 787.050 259.050 ;
        RECT 805.950 258.600 808.050 259.050 ;
        RECT 775.950 257.400 808.050 258.600 ;
        RECT 775.950 256.950 778.050 257.400 ;
        RECT 784.950 256.950 787.050 257.400 ;
        RECT 805.950 256.950 808.050 257.400 ;
        RECT 808.950 258.600 811.050 259.050 ;
        RECT 817.950 258.600 820.050 259.050 ;
        RECT 808.950 257.400 820.050 258.600 ;
        RECT 808.950 256.950 811.050 257.400 ;
        RECT 817.950 256.950 820.050 257.400 ;
        RECT 19.950 255.600 22.050 256.050 ;
        RECT 109.950 255.600 112.050 256.050 ;
        RECT 19.950 254.400 112.050 255.600 ;
        RECT 19.950 253.950 22.050 254.400 ;
        RECT 109.950 253.950 112.050 254.400 ;
        RECT 277.950 255.600 280.050 256.050 ;
        RECT 334.950 255.600 337.050 256.050 ;
        RECT 277.950 254.400 337.050 255.600 ;
        RECT 277.950 253.950 280.050 254.400 ;
        RECT 334.950 253.950 337.050 254.400 ;
        RECT 358.950 255.600 361.050 256.050 ;
        RECT 370.950 255.600 373.050 256.050 ;
        RECT 358.950 254.400 373.050 255.600 ;
        RECT 358.950 253.950 361.050 254.400 ;
        RECT 370.950 253.950 373.050 254.400 ;
        RECT 511.950 255.600 514.050 256.050 ;
        RECT 520.950 255.600 523.050 256.050 ;
        RECT 583.950 255.600 586.050 256.050 ;
        RECT 511.950 254.400 586.050 255.600 ;
        RECT 511.950 253.950 514.050 254.400 ;
        RECT 520.950 253.950 523.050 254.400 ;
        RECT 583.950 253.950 586.050 254.400 ;
        RECT 595.950 255.600 598.050 256.050 ;
        RECT 613.950 255.600 616.050 256.050 ;
        RECT 595.950 254.400 616.050 255.600 ;
        RECT 595.950 253.950 598.050 254.400 ;
        RECT 613.950 253.950 616.050 254.400 ;
        RECT 649.950 253.950 652.050 256.050 ;
        RECT 667.950 255.600 670.050 256.050 ;
        RECT 682.950 255.600 685.050 256.050 ;
        RECT 667.950 254.400 685.050 255.600 ;
        RECT 667.950 253.950 670.050 254.400 ;
        RECT 682.950 253.950 685.050 254.400 ;
        RECT 691.950 255.600 694.050 256.050 ;
        RECT 721.950 255.600 724.050 256.050 ;
        RECT 814.950 255.600 817.050 256.050 ;
        RECT 691.950 254.400 724.050 255.600 ;
        RECT 691.950 253.950 694.050 254.400 ;
        RECT 721.950 253.950 724.050 254.400 ;
        RECT 788.400 254.400 817.050 255.600 ;
        RECT 28.950 252.600 31.050 253.050 ;
        RECT 43.950 252.600 46.050 253.050 ;
        RECT 28.950 251.400 46.050 252.600 ;
        RECT 28.950 250.950 31.050 251.400 ;
        RECT 43.950 250.950 46.050 251.400 ;
        RECT 169.950 252.600 172.050 253.050 ;
        RECT 196.950 252.600 199.050 253.050 ;
        RECT 169.950 251.400 199.050 252.600 ;
        RECT 169.950 250.950 172.050 251.400 ;
        RECT 196.950 250.950 199.050 251.400 ;
        RECT 214.950 252.600 217.050 253.050 ;
        RECT 238.950 252.600 241.050 253.050 ;
        RECT 214.950 251.400 241.050 252.600 ;
        RECT 214.950 250.950 217.050 251.400 ;
        RECT 238.950 250.950 241.050 251.400 ;
        RECT 268.950 252.600 271.050 253.050 ;
        RECT 286.950 252.600 289.050 253.050 ;
        RECT 298.950 252.600 301.050 253.050 ;
        RECT 268.950 251.400 289.050 252.600 ;
        RECT 268.950 250.950 271.050 251.400 ;
        RECT 286.950 250.950 289.050 251.400 ;
        RECT 290.400 251.400 301.050 252.600 ;
        RECT 139.950 249.600 142.050 250.050 ;
        RECT 163.950 249.600 166.050 250.050 ;
        RECT 290.400 249.600 291.600 251.400 ;
        RECT 298.950 250.950 301.050 251.400 ;
        RECT 376.950 252.600 379.050 253.050 ;
        RECT 478.950 252.600 481.050 253.050 ;
        RECT 496.950 252.600 499.050 253.050 ;
        RECT 376.950 251.400 481.050 252.600 ;
        RECT 376.950 250.950 379.050 251.400 ;
        RECT 478.950 250.950 481.050 251.400 ;
        RECT 491.400 251.400 499.050 252.600 ;
        RECT 139.950 248.400 291.600 249.600 ;
        RECT 433.950 249.600 436.050 250.050 ;
        RECT 481.950 249.600 484.050 250.050 ;
        RECT 433.950 248.400 484.050 249.600 ;
        RECT 139.950 247.950 142.050 248.400 ;
        RECT 163.950 247.950 166.050 248.400 ;
        RECT 433.950 247.950 436.050 248.400 ;
        RECT 481.950 247.950 484.050 248.400 ;
        RECT 484.950 249.600 487.050 250.050 ;
        RECT 484.950 248.400 489.600 249.600 ;
        RECT 484.950 247.950 487.050 248.400 ;
        RECT 10.950 246.600 13.050 247.050 ;
        RECT 85.950 246.600 88.050 247.050 ;
        RECT 91.950 246.600 94.050 247.050 ;
        RECT 10.950 245.400 94.050 246.600 ;
        RECT 10.950 244.950 13.050 245.400 ;
        RECT 85.950 244.950 88.050 245.400 ;
        RECT 91.950 244.950 94.050 245.400 ;
        RECT 193.950 246.600 196.050 247.050 ;
        RECT 337.950 246.600 340.050 247.050 ;
        RECT 193.950 245.400 340.050 246.600 ;
        RECT 193.950 244.950 196.050 245.400 ;
        RECT 337.950 244.950 340.050 245.400 ;
        RECT 373.950 246.600 376.050 247.050 ;
        RECT 427.950 246.600 430.050 247.050 ;
        RECT 373.950 245.400 430.050 246.600 ;
        RECT 373.950 244.950 376.050 245.400 ;
        RECT 427.950 244.950 430.050 245.400 ;
        RECT 448.950 246.600 451.050 247.050 ;
        RECT 484.950 246.600 487.050 247.050 ;
        RECT 448.950 245.400 487.050 246.600 ;
        RECT 448.950 244.950 451.050 245.400 ;
        RECT 484.950 244.950 487.050 245.400 ;
        RECT 46.950 243.600 49.050 244.050 ;
        RECT 55.950 243.600 58.050 244.050 ;
        RECT 46.950 242.400 58.050 243.600 ;
        RECT 46.950 241.950 49.050 242.400 ;
        RECT 55.950 241.950 58.050 242.400 ;
        RECT 82.950 243.600 85.050 244.050 ;
        RECT 103.950 243.600 106.050 244.050 ;
        RECT 82.950 242.400 106.050 243.600 ;
        RECT 82.950 241.950 85.050 242.400 ;
        RECT 103.950 241.950 106.050 242.400 ;
        RECT 109.950 243.600 112.050 244.050 ;
        RECT 112.950 243.600 115.050 244.050 ;
        RECT 133.950 243.600 136.050 244.050 ;
        RECT 109.950 242.400 136.050 243.600 ;
        RECT 109.950 241.950 112.050 242.400 ;
        RECT 112.950 241.950 115.050 242.400 ;
        RECT 133.950 241.950 136.050 242.400 ;
        RECT 145.950 243.600 148.050 244.050 ;
        RECT 193.950 243.600 196.050 244.050 ;
        RECT 145.950 242.400 196.050 243.600 ;
        RECT 145.950 241.950 148.050 242.400 ;
        RECT 193.950 241.950 196.050 242.400 ;
        RECT 199.950 243.600 202.050 244.050 ;
        RECT 217.950 243.600 220.050 244.050 ;
        RECT 199.950 242.400 220.050 243.600 ;
        RECT 199.950 241.950 202.050 242.400 ;
        RECT 217.950 241.950 220.050 242.400 ;
        RECT 235.950 243.600 238.050 244.050 ;
        RECT 244.950 243.600 247.050 244.050 ;
        RECT 235.950 242.400 247.050 243.600 ;
        RECT 235.950 241.950 238.050 242.400 ;
        RECT 244.950 241.950 247.050 242.400 ;
        RECT 259.950 243.600 262.050 244.050 ;
        RECT 274.950 243.600 277.050 244.050 ;
        RECT 259.950 242.400 277.050 243.600 ;
        RECT 259.950 241.950 262.050 242.400 ;
        RECT 274.950 241.950 277.050 242.400 ;
        RECT 304.950 243.600 307.050 244.050 ;
        RECT 349.950 243.600 352.050 244.050 ;
        RECT 304.950 242.400 352.050 243.600 ;
        RECT 304.950 241.950 307.050 242.400 ;
        RECT 349.950 241.950 352.050 242.400 ;
        RECT 379.950 243.600 382.050 244.050 ;
        RECT 406.950 243.600 409.050 244.050 ;
        RECT 379.950 242.400 409.050 243.600 ;
        RECT 379.950 241.950 382.050 242.400 ;
        RECT 406.950 241.950 409.050 242.400 ;
        RECT 418.950 243.600 421.050 244.050 ;
        RECT 454.950 243.600 457.050 244.050 ;
        RECT 457.950 243.600 460.050 244.050 ;
        RECT 418.950 242.400 460.050 243.600 ;
        RECT 418.950 241.950 421.050 242.400 ;
        RECT 454.950 241.950 457.050 242.400 ;
        RECT 457.950 241.950 460.050 242.400 ;
        RECT 40.950 240.600 43.050 241.050 ;
        RECT 130.950 240.600 133.050 241.050 ;
        RECT 154.950 240.600 157.050 241.050 ;
        RECT 40.950 239.400 57.600 240.600 ;
        RECT 40.950 238.950 43.050 239.400 ;
        RECT 56.400 238.050 57.600 239.400 ;
        RECT 130.950 239.400 157.050 240.600 ;
        RECT 130.950 238.950 133.050 239.400 ;
        RECT 154.950 238.950 157.050 239.400 ;
        RECT 172.950 240.600 175.050 241.050 ;
        RECT 205.950 240.600 208.050 241.050 ;
        RECT 172.950 239.400 208.050 240.600 ;
        RECT 172.950 238.950 175.050 239.400 ;
        RECT 205.950 238.950 208.050 239.400 ;
        RECT 238.950 240.600 241.050 241.050 ;
        RECT 244.950 240.600 247.050 241.050 ;
        RECT 238.950 239.400 247.050 240.600 ;
        RECT 238.950 238.950 241.050 239.400 ;
        RECT 244.950 238.950 247.050 239.400 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 343.950 240.600 346.050 241.050 ;
        RECT 361.950 240.600 364.050 241.050 ;
        RECT 343.950 239.400 364.050 240.600 ;
        RECT 343.950 238.950 346.050 239.400 ;
        RECT 361.950 238.950 364.050 239.400 ;
        RECT 388.950 240.600 391.050 241.050 ;
        RECT 466.950 240.600 469.050 241.050 ;
        RECT 388.950 239.400 408.600 240.600 ;
        RECT 388.950 238.950 391.050 239.400 ;
        RECT 4.950 237.600 7.050 238.050 ;
        RECT 16.950 237.600 19.050 238.050 ;
        RECT 4.950 236.400 19.050 237.600 ;
        RECT 4.950 235.950 7.050 236.400 ;
        RECT 16.950 235.950 19.050 236.400 ;
        RECT 37.950 235.950 40.050 238.050 ;
        RECT 40.950 237.600 43.050 238.050 ;
        RECT 52.950 237.600 55.050 238.050 ;
        RECT 40.950 236.400 55.050 237.600 ;
        RECT 40.950 235.950 43.050 236.400 ;
        RECT 52.950 235.950 55.050 236.400 ;
        RECT 55.950 235.950 58.050 238.050 ;
        RECT 73.950 237.600 76.050 238.050 ;
        RECT 79.950 237.600 82.050 238.050 ;
        RECT 73.950 236.400 82.050 237.600 ;
        RECT 73.950 235.950 76.050 236.400 ;
        RECT 79.950 235.950 82.050 236.400 ;
        RECT 115.950 237.600 118.050 238.050 ;
        RECT 127.950 237.600 130.050 238.050 ;
        RECT 115.950 236.400 130.050 237.600 ;
        RECT 115.950 235.950 118.050 236.400 ;
        RECT 127.950 235.950 130.050 236.400 ;
        RECT 136.950 237.600 139.050 238.050 ;
        RECT 145.950 237.600 148.050 238.050 ;
        RECT 136.950 236.400 148.050 237.600 ;
        RECT 136.950 235.950 139.050 236.400 ;
        RECT 145.950 235.950 148.050 236.400 ;
        RECT 154.950 237.600 157.050 238.050 ;
        RECT 175.950 237.600 178.050 238.050 ;
        RECT 154.950 236.400 178.050 237.600 ;
        RECT 154.950 235.950 157.050 236.400 ;
        RECT 175.950 235.950 178.050 236.400 ;
        RECT 232.950 237.600 235.050 238.050 ;
        RECT 247.950 237.600 250.050 238.050 ;
        RECT 232.950 236.400 250.050 237.600 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 247.950 235.950 250.050 236.400 ;
        RECT 304.950 237.600 307.050 238.050 ;
        RECT 320.400 237.600 321.600 238.950 ;
        RECT 304.950 236.400 321.600 237.600 ;
        RECT 337.950 237.600 340.050 238.050 ;
        RECT 346.950 237.600 349.050 238.050 ;
        RECT 337.950 236.400 349.050 237.600 ;
        RECT 304.950 235.950 307.050 236.400 ;
        RECT 337.950 235.950 340.050 236.400 ;
        RECT 346.950 235.950 349.050 236.400 ;
        RECT 352.950 237.600 355.050 238.050 ;
        RECT 367.950 237.600 370.050 238.050 ;
        RECT 352.950 236.400 370.050 237.600 ;
        RECT 352.950 235.950 355.050 236.400 ;
        RECT 367.950 235.950 370.050 236.400 ;
        RECT 13.950 232.950 16.050 235.050 ;
        RECT 19.950 234.600 22.050 235.050 ;
        RECT 31.950 234.600 34.050 235.050 ;
        RECT 19.950 233.400 34.050 234.600 ;
        RECT 38.400 234.600 39.600 235.950 ;
        RECT 407.400 235.050 408.600 239.400 ;
        RECT 464.400 239.400 469.050 240.600 ;
        RECT 409.950 237.600 412.050 238.050 ;
        RECT 445.950 237.600 448.050 238.050 ;
        RECT 409.950 236.400 448.050 237.600 ;
        RECT 409.950 235.950 412.050 236.400 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 58.950 234.600 61.050 235.050 ;
        RECT 38.400 233.400 61.050 234.600 ;
        RECT 19.950 232.950 22.050 233.400 ;
        RECT 31.950 232.950 34.050 233.400 ;
        RECT 58.950 232.950 61.050 233.400 ;
        RECT 88.950 234.600 91.050 235.050 ;
        RECT 94.950 234.600 97.050 235.050 ;
        RECT 88.950 233.400 97.050 234.600 ;
        RECT 88.950 232.950 91.050 233.400 ;
        RECT 94.950 232.950 97.050 233.400 ;
        RECT 178.950 234.600 181.050 235.050 ;
        RECT 187.950 234.600 190.050 235.050 ;
        RECT 196.950 234.600 199.050 235.050 ;
        RECT 178.950 233.400 199.050 234.600 ;
        RECT 178.950 232.950 181.050 233.400 ;
        RECT 187.950 232.950 190.050 233.400 ;
        RECT 196.950 232.950 199.050 233.400 ;
        RECT 220.950 234.600 223.050 235.050 ;
        RECT 265.950 234.600 268.050 235.050 ;
        RECT 220.950 233.400 268.050 234.600 ;
        RECT 220.950 232.950 223.050 233.400 ;
        RECT 265.950 232.950 268.050 233.400 ;
        RECT 406.950 232.950 409.050 235.050 ;
        RECT 464.400 234.600 465.600 239.400 ;
        RECT 466.950 238.950 469.050 239.400 ;
        RECT 464.400 233.400 468.600 234.600 ;
        RECT 14.400 231.600 15.600 232.950 ;
        RECT 467.400 232.050 468.600 233.400 ;
        RECT 16.950 231.600 19.050 232.050 ;
        RECT 14.400 230.400 19.050 231.600 ;
        RECT 16.950 229.950 19.050 230.400 ;
        RECT 28.950 231.600 31.050 232.050 ;
        RECT 34.950 231.600 37.050 232.050 ;
        RECT 28.950 230.400 37.050 231.600 ;
        RECT 28.950 229.950 31.050 230.400 ;
        RECT 34.950 229.950 37.050 230.400 ;
        RECT 52.950 231.600 55.050 232.050 ;
        RECT 112.950 231.600 115.050 232.050 ;
        RECT 52.950 230.400 115.050 231.600 ;
        RECT 52.950 229.950 55.050 230.400 ;
        RECT 112.950 229.950 115.050 230.400 ;
        RECT 364.950 231.600 367.050 232.050 ;
        RECT 412.950 231.600 415.050 232.050 ;
        RECT 418.950 231.600 421.050 232.050 ;
        RECT 364.950 230.400 421.050 231.600 ;
        RECT 364.950 229.950 367.050 230.400 ;
        RECT 412.950 229.950 415.050 230.400 ;
        RECT 418.950 229.950 421.050 230.400 ;
        RECT 436.950 231.600 439.050 232.050 ;
        RECT 445.950 231.600 448.050 232.050 ;
        RECT 436.950 230.400 448.050 231.600 ;
        RECT 436.950 229.950 439.050 230.400 ;
        RECT 445.950 229.950 448.050 230.400 ;
        RECT 466.950 229.950 469.050 232.050 ;
        RECT 10.950 228.600 13.050 229.050 ;
        RECT 55.950 228.600 58.050 229.050 ;
        RECT 10.950 227.400 58.050 228.600 ;
        RECT 10.950 226.950 13.050 227.400 ;
        RECT 55.950 226.950 58.050 227.400 ;
        RECT 142.950 228.600 145.050 229.050 ;
        RECT 187.950 228.600 190.050 229.050 ;
        RECT 142.950 227.400 190.050 228.600 ;
        RECT 142.950 226.950 145.050 227.400 ;
        RECT 187.950 226.950 190.050 227.400 ;
        RECT 397.950 228.600 400.050 229.050 ;
        RECT 427.950 228.600 430.050 229.050 ;
        RECT 397.950 227.400 430.050 228.600 ;
        RECT 397.950 226.950 400.050 227.400 ;
        RECT 427.950 226.950 430.050 227.400 ;
        RECT 451.950 228.600 454.050 229.050 ;
        RECT 469.950 228.600 472.050 229.050 ;
        RECT 451.950 227.400 472.050 228.600 ;
        RECT 451.950 226.950 454.050 227.400 ;
        RECT 469.950 226.950 472.050 227.400 ;
        RECT 488.400 223.050 489.600 248.400 ;
        RECT 491.400 223.050 492.600 251.400 ;
        RECT 496.950 250.950 499.050 251.400 ;
        RECT 532.950 252.600 535.050 253.050 ;
        RECT 550.950 252.600 553.050 253.050 ;
        RECT 532.950 251.400 553.050 252.600 ;
        RECT 532.950 250.950 535.050 251.400 ;
        RECT 550.950 250.950 553.050 251.400 ;
        RECT 610.950 252.600 613.050 253.050 ;
        RECT 634.950 252.600 637.050 253.050 ;
        RECT 610.950 251.400 637.050 252.600 ;
        RECT 610.950 250.950 613.050 251.400 ;
        RECT 634.950 250.950 637.050 251.400 ;
        RECT 715.950 252.600 718.050 253.050 ;
        RECT 751.950 252.600 754.050 253.050 ;
        RECT 715.950 251.400 754.050 252.600 ;
        RECT 715.950 250.950 718.050 251.400 ;
        RECT 751.950 250.950 754.050 251.400 ;
        RECT 778.950 252.600 781.050 253.050 ;
        RECT 788.400 252.600 789.600 254.400 ;
        RECT 814.950 253.950 817.050 254.400 ;
        RECT 778.950 251.400 789.600 252.600 ;
        RECT 790.950 252.600 793.050 253.050 ;
        RECT 799.950 252.600 802.050 253.050 ;
        RECT 790.950 251.400 802.050 252.600 ;
        RECT 778.950 250.950 781.050 251.400 ;
        RECT 790.950 250.950 793.050 251.400 ;
        RECT 799.950 250.950 802.050 251.400 ;
        RECT 559.950 249.600 562.050 250.050 ;
        RECT 586.950 249.600 589.050 250.050 ;
        RECT 559.950 248.400 589.050 249.600 ;
        RECT 559.950 247.950 562.050 248.400 ;
        RECT 586.950 247.950 589.050 248.400 ;
        RECT 598.950 249.600 601.050 250.050 ;
        RECT 643.950 249.600 646.050 250.050 ;
        RECT 598.950 248.400 646.050 249.600 ;
        RECT 598.950 247.950 601.050 248.400 ;
        RECT 643.950 247.950 646.050 248.400 ;
        RECT 652.950 249.600 655.050 250.050 ;
        RECT 724.950 249.600 727.050 250.050 ;
        RECT 652.950 248.400 727.050 249.600 ;
        RECT 652.950 247.950 655.050 248.400 ;
        RECT 724.950 247.950 727.050 248.400 ;
        RECT 760.950 249.600 763.050 250.050 ;
        RECT 778.950 249.600 781.050 250.050 ;
        RECT 787.950 249.600 790.050 250.050 ;
        RECT 760.950 248.400 790.050 249.600 ;
        RECT 760.950 247.950 763.050 248.400 ;
        RECT 778.950 247.950 781.050 248.400 ;
        RECT 787.950 247.950 790.050 248.400 ;
        RECT 793.950 249.600 796.050 250.050 ;
        RECT 820.950 249.600 823.050 250.050 ;
        RECT 793.950 248.400 823.050 249.600 ;
        RECT 793.950 247.950 796.050 248.400 ;
        RECT 820.950 247.950 823.050 248.400 ;
        RECT 562.950 246.600 565.050 247.050 ;
        RECT 610.950 246.600 613.050 247.050 ;
        RECT 718.950 246.600 721.050 247.050 ;
        RECT 562.950 245.400 613.050 246.600 ;
        RECT 562.950 244.950 565.050 245.400 ;
        RECT 610.950 244.950 613.050 245.400 ;
        RECT 614.400 245.400 721.050 246.600 ;
        RECT 532.950 243.600 535.050 244.050 ;
        RECT 538.950 243.600 541.050 244.050 ;
        RECT 532.950 242.400 541.050 243.600 ;
        RECT 532.950 241.950 535.050 242.400 ;
        RECT 538.950 241.950 541.050 242.400 ;
        RECT 550.950 243.600 553.050 244.050 ;
        RECT 562.950 243.600 565.050 244.050 ;
        RECT 550.950 242.400 565.050 243.600 ;
        RECT 550.950 241.950 553.050 242.400 ;
        RECT 562.950 241.950 565.050 242.400 ;
        RECT 595.950 243.600 598.050 244.050 ;
        RECT 614.400 243.600 615.600 245.400 ;
        RECT 718.950 244.950 721.050 245.400 ;
        RECT 766.950 246.600 769.050 247.050 ;
        RECT 805.950 246.600 808.050 247.050 ;
        RECT 766.950 245.400 808.050 246.600 ;
        RECT 766.950 244.950 769.050 245.400 ;
        RECT 805.950 244.950 808.050 245.400 ;
        RECT 835.950 246.600 838.050 247.050 ;
        RECT 862.950 246.600 865.050 247.050 ;
        RECT 835.950 245.400 865.050 246.600 ;
        RECT 835.950 244.950 838.050 245.400 ;
        RECT 862.950 244.950 865.050 245.400 ;
        RECT 595.950 242.400 615.600 243.600 ;
        RECT 667.950 243.600 670.050 244.050 ;
        RECT 670.950 243.600 673.050 244.050 ;
        RECT 667.950 242.400 673.050 243.600 ;
        RECT 595.950 241.950 598.050 242.400 ;
        RECT 667.950 241.950 670.050 242.400 ;
        RECT 670.950 241.950 673.050 242.400 ;
        RECT 679.950 243.600 682.050 244.050 ;
        RECT 691.950 243.600 694.050 244.050 ;
        RECT 679.950 242.400 694.050 243.600 ;
        RECT 679.950 241.950 682.050 242.400 ;
        RECT 691.950 241.950 694.050 242.400 ;
        RECT 718.950 243.600 721.050 244.050 ;
        RECT 727.950 243.600 730.050 244.050 ;
        RECT 718.950 242.400 730.050 243.600 ;
        RECT 718.950 241.950 721.050 242.400 ;
        RECT 727.950 241.950 730.050 242.400 ;
        RECT 730.950 243.600 733.050 244.050 ;
        RECT 739.950 243.600 742.050 244.050 ;
        RECT 730.950 242.400 742.050 243.600 ;
        RECT 730.950 241.950 733.050 242.400 ;
        RECT 739.950 241.950 742.050 242.400 ;
        RECT 751.950 243.600 754.050 244.050 ;
        RECT 844.950 243.600 847.050 244.050 ;
        RECT 856.950 243.600 859.050 244.050 ;
        RECT 751.950 242.400 804.600 243.600 ;
        RECT 751.950 241.950 754.050 242.400 ;
        RECT 529.950 240.600 532.050 241.050 ;
        RECT 538.950 240.600 541.050 241.050 ;
        RECT 556.950 240.600 559.050 241.050 ;
        RECT 529.950 239.400 541.050 240.600 ;
        RECT 529.950 238.950 532.050 239.400 ;
        RECT 538.950 238.950 541.050 239.400 ;
        RECT 551.400 239.400 559.050 240.600 ;
        RECT 547.950 237.600 550.050 238.050 ;
        RECT 551.400 237.600 552.600 239.400 ;
        RECT 556.950 238.950 559.050 239.400 ;
        RECT 598.950 240.600 601.050 241.050 ;
        RECT 601.950 240.600 604.050 241.050 ;
        RECT 619.950 240.600 622.050 241.050 ;
        RECT 637.950 240.600 640.050 241.050 ;
        RECT 598.950 239.400 618.600 240.600 ;
        RECT 598.950 238.950 601.050 239.400 ;
        RECT 601.950 238.950 604.050 239.400 ;
        RECT 547.950 236.400 552.600 237.600 ;
        RECT 553.950 237.600 556.050 238.050 ;
        RECT 559.950 237.600 562.050 238.050 ;
        RECT 553.950 236.400 562.050 237.600 ;
        RECT 547.950 235.950 550.050 236.400 ;
        RECT 553.950 235.950 556.050 236.400 ;
        RECT 559.950 235.950 562.050 236.400 ;
        RECT 565.950 237.600 568.050 238.050 ;
        RECT 583.950 237.600 586.050 238.050 ;
        RECT 565.950 236.400 586.050 237.600 ;
        RECT 565.950 235.950 568.050 236.400 ;
        RECT 583.950 235.950 586.050 236.400 ;
        RECT 514.950 234.600 517.050 235.050 ;
        RECT 520.950 234.600 523.050 235.050 ;
        RECT 514.950 233.400 523.050 234.600 ;
        RECT 514.950 232.950 517.050 233.400 ;
        RECT 520.950 232.950 523.050 233.400 ;
        RECT 541.950 234.600 544.050 235.050 ;
        RECT 550.950 234.600 553.050 235.050 ;
        RECT 541.950 233.400 553.050 234.600 ;
        RECT 617.400 234.600 618.600 239.400 ;
        RECT 619.950 239.400 640.050 240.600 ;
        RECT 619.950 238.950 622.050 239.400 ;
        RECT 637.950 238.950 640.050 239.400 ;
        RECT 649.950 240.600 652.050 241.050 ;
        RECT 673.950 240.600 676.050 241.050 ;
        RECT 685.950 240.600 688.050 241.050 ;
        RECT 649.950 239.400 688.050 240.600 ;
        RECT 649.950 238.950 652.050 239.400 ;
        RECT 673.950 238.950 676.050 239.400 ;
        RECT 685.950 238.950 688.050 239.400 ;
        RECT 697.950 240.600 700.050 241.050 ;
        RECT 712.950 240.600 715.050 241.050 ;
        RECT 697.950 239.400 715.050 240.600 ;
        RECT 697.950 238.950 700.050 239.400 ;
        RECT 712.950 238.950 715.050 239.400 ;
        RECT 715.950 238.950 718.050 241.050 ;
        RECT 733.950 240.600 736.050 241.050 ;
        RECT 728.400 239.400 736.050 240.600 ;
        RECT 640.950 237.600 643.050 238.050 ;
        RECT 664.950 237.600 667.050 238.050 ;
        RECT 682.950 237.600 685.050 238.050 ;
        RECT 694.950 237.600 697.050 238.050 ;
        RECT 716.400 237.600 717.600 238.950 ;
        RECT 640.950 236.400 717.600 237.600 ;
        RECT 640.950 235.950 643.050 236.400 ;
        RECT 664.950 235.950 667.050 236.400 ;
        RECT 682.950 235.950 685.050 236.400 ;
        RECT 694.950 235.950 697.050 236.400 ;
        RECT 728.400 235.050 729.600 239.400 ;
        RECT 733.950 238.950 736.050 239.400 ;
        RECT 790.950 240.600 793.050 241.050 ;
        RECT 799.950 240.600 802.050 241.050 ;
        RECT 790.950 239.400 802.050 240.600 ;
        RECT 790.950 238.950 793.050 239.400 ;
        RECT 799.950 238.950 802.050 239.400 ;
        RECT 803.400 238.050 804.600 242.400 ;
        RECT 844.950 242.400 859.050 243.600 ;
        RECT 844.950 241.950 847.050 242.400 ;
        RECT 856.950 241.950 859.050 242.400 ;
        RECT 820.950 240.600 823.050 241.050 ;
        RECT 829.950 240.600 832.050 241.050 ;
        RECT 820.950 239.400 832.050 240.600 ;
        RECT 820.950 238.950 823.050 239.400 ;
        RECT 829.950 238.950 832.050 239.400 ;
        RECT 847.950 240.600 850.050 241.050 ;
        RECT 868.950 240.600 871.050 241.050 ;
        RECT 847.950 239.400 871.050 240.600 ;
        RECT 847.950 238.950 850.050 239.400 ;
        RECT 868.950 238.950 871.050 239.400 ;
        RECT 796.950 237.600 799.050 238.050 ;
        RECT 796.950 236.400 801.600 237.600 ;
        RECT 796.950 235.950 799.050 236.400 ;
        RECT 800.400 235.050 801.600 236.400 ;
        RECT 802.950 235.950 805.050 238.050 ;
        RECT 835.950 237.600 838.050 238.050 ;
        RECT 818.400 236.400 838.050 237.600 ;
        RECT 818.400 235.050 819.600 236.400 ;
        RECT 835.950 235.950 838.050 236.400 ;
        RECT 841.950 237.600 844.050 238.050 ;
        RECT 868.950 237.600 871.050 238.050 ;
        RECT 841.950 236.400 871.050 237.600 ;
        RECT 841.950 235.950 844.050 236.400 ;
        RECT 868.950 235.950 871.050 236.400 ;
        RECT 622.950 234.600 625.050 235.050 ;
        RECT 617.400 233.400 625.050 234.600 ;
        RECT 541.950 232.950 544.050 233.400 ;
        RECT 550.950 232.950 553.050 233.400 ;
        RECT 622.950 232.950 625.050 233.400 ;
        RECT 709.950 234.600 712.050 235.050 ;
        RECT 724.950 234.600 727.050 235.050 ;
        RECT 709.950 233.400 727.050 234.600 ;
        RECT 709.950 232.950 712.050 233.400 ;
        RECT 724.950 232.950 727.050 233.400 ;
        RECT 727.950 232.950 730.050 235.050 ;
        RECT 760.950 234.600 763.050 235.050 ;
        RECT 775.950 234.600 778.050 235.050 ;
        RECT 760.950 233.400 778.050 234.600 ;
        RECT 760.950 232.950 763.050 233.400 ;
        RECT 775.950 232.950 778.050 233.400 ;
        RECT 799.950 234.600 802.050 235.050 ;
        RECT 814.950 234.600 817.050 235.050 ;
        RECT 799.950 233.400 817.050 234.600 ;
        RECT 799.950 232.950 802.050 233.400 ;
        RECT 814.950 232.950 817.050 233.400 ;
        RECT 817.950 232.950 820.050 235.050 ;
        RECT 823.950 234.600 826.050 235.050 ;
        RECT 832.950 234.600 835.050 235.050 ;
        RECT 838.950 234.600 841.050 235.050 ;
        RECT 823.950 233.400 841.050 234.600 ;
        RECT 823.950 232.950 826.050 233.400 ;
        RECT 832.950 232.950 835.050 233.400 ;
        RECT 838.950 232.950 841.050 233.400 ;
        RECT 520.950 231.600 523.050 232.050 ;
        RECT 526.950 231.600 529.050 232.050 ;
        RECT 520.950 230.400 529.050 231.600 ;
        RECT 520.950 229.950 523.050 230.400 ;
        RECT 526.950 229.950 529.050 230.400 ;
        RECT 529.950 231.600 532.050 232.050 ;
        RECT 538.950 231.600 541.050 232.050 ;
        RECT 529.950 230.400 541.050 231.600 ;
        RECT 529.950 229.950 532.050 230.400 ;
        RECT 538.950 229.950 541.050 230.400 ;
        RECT 559.950 231.600 562.050 232.050 ;
        RECT 688.950 231.600 691.050 232.050 ;
        RECT 721.950 231.600 724.050 232.050 ;
        RECT 754.950 231.600 757.050 232.050 ;
        RECT 559.950 230.400 757.050 231.600 ;
        RECT 559.950 229.950 562.050 230.400 ;
        RECT 688.950 229.950 691.050 230.400 ;
        RECT 721.950 229.950 724.050 230.400 ;
        RECT 754.950 229.950 757.050 230.400 ;
        RECT 778.950 231.600 781.050 232.050 ;
        RECT 787.950 231.600 790.050 232.050 ;
        RECT 778.950 230.400 790.050 231.600 ;
        RECT 778.950 229.950 781.050 230.400 ;
        RECT 787.950 229.950 790.050 230.400 ;
        RECT 808.950 231.600 811.050 232.050 ;
        RECT 817.950 231.600 820.050 232.050 ;
        RECT 808.950 230.400 820.050 231.600 ;
        RECT 808.950 229.950 811.050 230.400 ;
        RECT 817.950 229.950 820.050 230.400 ;
        RECT 841.950 231.600 844.050 232.050 ;
        RECT 850.950 231.600 853.050 232.050 ;
        RECT 841.950 230.400 853.050 231.600 ;
        RECT 841.950 229.950 844.050 230.400 ;
        RECT 850.950 229.950 853.050 230.400 ;
        RECT 526.950 228.600 529.050 229.050 ;
        RECT 577.950 228.600 580.050 229.050 ;
        RECT 616.950 228.600 619.050 229.050 ;
        RECT 526.950 227.400 619.050 228.600 ;
        RECT 526.950 226.950 529.050 227.400 ;
        RECT 577.950 226.950 580.050 227.400 ;
        RECT 616.950 226.950 619.050 227.400 ;
        RECT 715.950 228.600 718.050 229.050 ;
        RECT 730.950 228.600 733.050 229.050 ;
        RECT 748.950 228.600 751.050 229.050 ;
        RECT 715.950 227.400 751.050 228.600 ;
        RECT 715.950 226.950 718.050 227.400 ;
        RECT 730.950 226.950 733.050 227.400 ;
        RECT 748.950 226.950 751.050 227.400 ;
        RECT 766.950 228.600 769.050 229.050 ;
        RECT 781.950 228.600 784.050 229.050 ;
        RECT 766.950 227.400 784.050 228.600 ;
        RECT 766.950 226.950 769.050 227.400 ;
        RECT 781.950 226.950 784.050 227.400 ;
        RECT 796.950 228.600 799.050 229.050 ;
        RECT 865.950 228.600 868.050 229.050 ;
        RECT 796.950 227.400 868.050 228.600 ;
        RECT 796.950 226.950 799.050 227.400 ;
        RECT 865.950 226.950 868.050 227.400 ;
        RECT 514.950 225.600 517.050 226.050 ;
        RECT 709.950 225.600 712.050 226.050 ;
        RECT 514.950 224.400 712.050 225.600 ;
        RECT 514.950 223.950 517.050 224.400 ;
        RECT 709.950 223.950 712.050 224.400 ;
        RECT 811.950 225.600 814.050 226.050 ;
        RECT 865.950 225.600 868.050 226.050 ;
        RECT 811.950 224.400 868.050 225.600 ;
        RECT 811.950 223.950 814.050 224.400 ;
        RECT 865.950 223.950 868.050 224.400 ;
        RECT 43.950 222.600 46.050 223.050 ;
        RECT 58.950 222.600 61.050 223.050 ;
        RECT 43.950 221.400 61.050 222.600 ;
        RECT 43.950 220.950 46.050 221.400 ;
        RECT 58.950 220.950 61.050 221.400 ;
        RECT 304.950 222.600 307.050 223.050 ;
        RECT 316.950 222.600 319.050 223.050 ;
        RECT 304.950 221.400 319.050 222.600 ;
        RECT 304.950 220.950 307.050 221.400 ;
        RECT 316.950 220.950 319.050 221.400 ;
        RECT 487.950 220.950 490.050 223.050 ;
        RECT 490.950 220.950 493.050 223.050 ;
        RECT 529.950 222.600 532.050 223.050 ;
        RECT 601.950 222.600 604.050 223.050 ;
        RECT 640.950 222.600 643.050 223.050 ;
        RECT 646.950 222.600 649.050 223.050 ;
        RECT 670.950 222.600 673.050 223.050 ;
        RECT 529.950 221.400 673.050 222.600 ;
        RECT 529.950 220.950 532.050 221.400 ;
        RECT 601.950 220.950 604.050 221.400 ;
        RECT 640.950 220.950 643.050 221.400 ;
        RECT 646.950 220.950 649.050 221.400 ;
        RECT 670.950 220.950 673.050 221.400 ;
        RECT 814.950 222.600 817.050 223.050 ;
        RECT 826.950 222.600 829.050 223.050 ;
        RECT 814.950 221.400 829.050 222.600 ;
        RECT 814.950 220.950 817.050 221.400 ;
        RECT 826.950 220.950 829.050 221.400 ;
        RECT 46.950 219.600 49.050 220.050 ;
        RECT 52.950 219.600 55.050 220.050 ;
        RECT 46.950 218.400 55.050 219.600 ;
        RECT 46.950 217.950 49.050 218.400 ;
        RECT 52.950 217.950 55.050 218.400 ;
        RECT 379.950 219.600 382.050 220.050 ;
        RECT 517.950 219.600 520.050 220.050 ;
        RECT 754.950 219.600 757.050 220.050 ;
        RECT 760.950 219.600 763.050 220.050 ;
        RECT 799.950 219.600 802.050 220.050 ;
        RECT 379.950 218.400 802.050 219.600 ;
        RECT 379.950 217.950 382.050 218.400 ;
        RECT 517.950 217.950 520.050 218.400 ;
        RECT 754.950 217.950 757.050 218.400 ;
        RECT 760.950 217.950 763.050 218.400 ;
        RECT 799.950 217.950 802.050 218.400 ;
        RECT 343.950 216.600 346.050 217.050 ;
        RECT 529.950 216.600 532.050 217.050 ;
        RECT 343.950 215.400 532.050 216.600 ;
        RECT 343.950 214.950 346.050 215.400 ;
        RECT 529.950 214.950 532.050 215.400 ;
        RECT 775.950 216.600 778.050 217.050 ;
        RECT 784.950 216.600 787.050 217.050 ;
        RECT 775.950 215.400 787.050 216.600 ;
        RECT 775.950 214.950 778.050 215.400 ;
        RECT 784.950 214.950 787.050 215.400 ;
        RECT 16.950 213.600 19.050 214.050 ;
        RECT 46.950 213.600 49.050 214.050 ;
        RECT 16.950 212.400 49.050 213.600 ;
        RECT 16.950 211.950 19.050 212.400 ;
        RECT 46.950 211.950 49.050 212.400 ;
        RECT 205.950 213.600 208.050 214.050 ;
        RECT 388.950 213.600 391.050 214.050 ;
        RECT 409.950 213.600 412.050 214.050 ;
        RECT 439.950 213.600 442.050 214.050 ;
        RECT 205.950 212.400 442.050 213.600 ;
        RECT 205.950 211.950 208.050 212.400 ;
        RECT 388.950 211.950 391.050 212.400 ;
        RECT 409.950 211.950 412.050 212.400 ;
        RECT 439.950 211.950 442.050 212.400 ;
        RECT 568.950 213.600 571.050 214.050 ;
        RECT 574.950 213.600 577.050 214.050 ;
        RECT 568.950 212.400 577.050 213.600 ;
        RECT 568.950 211.950 571.050 212.400 ;
        RECT 574.950 211.950 577.050 212.400 ;
        RECT 592.950 213.600 595.050 214.050 ;
        RECT 712.950 213.600 715.050 214.050 ;
        RECT 592.950 212.400 715.050 213.600 ;
        RECT 592.950 211.950 595.050 212.400 ;
        RECT 712.950 211.950 715.050 212.400 ;
        RECT 763.950 213.600 766.050 214.050 ;
        RECT 784.950 213.600 787.050 214.050 ;
        RECT 763.950 212.400 787.050 213.600 ;
        RECT 763.950 211.950 766.050 212.400 ;
        RECT 784.950 211.950 787.050 212.400 ;
        RECT 382.950 210.600 385.050 211.050 ;
        RECT 391.950 210.600 394.050 211.050 ;
        RECT 382.950 209.400 394.050 210.600 ;
        RECT 382.950 208.950 385.050 209.400 ;
        RECT 391.950 208.950 394.050 209.400 ;
        RECT 424.950 210.600 427.050 211.050 ;
        RECT 430.950 210.600 433.050 211.050 ;
        RECT 424.950 209.400 433.050 210.600 ;
        RECT 424.950 208.950 427.050 209.400 ;
        RECT 430.950 208.950 433.050 209.400 ;
        RECT 466.950 210.600 469.050 211.050 ;
        RECT 493.950 210.600 496.050 211.050 ;
        RECT 466.950 209.400 496.050 210.600 ;
        RECT 466.950 208.950 469.050 209.400 ;
        RECT 493.950 208.950 496.050 209.400 ;
        RECT 547.950 210.600 550.050 211.050 ;
        RECT 553.950 210.600 556.050 211.050 ;
        RECT 652.950 210.600 655.050 211.050 ;
        RECT 547.950 209.400 655.050 210.600 ;
        RECT 547.950 208.950 550.050 209.400 ;
        RECT 553.950 208.950 556.050 209.400 ;
        RECT 652.950 208.950 655.050 209.400 ;
        RECT 721.950 210.600 724.050 211.050 ;
        RECT 727.950 210.600 730.050 211.050 ;
        RECT 721.950 209.400 730.050 210.600 ;
        RECT 721.950 208.950 724.050 209.400 ;
        RECT 727.950 208.950 730.050 209.400 ;
        RECT 835.950 210.600 838.050 211.050 ;
        RECT 847.950 210.600 850.050 211.050 ;
        RECT 835.950 209.400 850.050 210.600 ;
        RECT 835.950 208.950 838.050 209.400 ;
        RECT 847.950 208.950 850.050 209.400 ;
        RECT 253.950 207.600 256.050 208.050 ;
        RECT 262.950 207.600 265.050 208.050 ;
        RECT 268.950 207.600 271.050 208.050 ;
        RECT 310.950 207.600 313.050 208.050 ;
        RECT 253.950 206.400 313.050 207.600 ;
        RECT 253.950 205.950 256.050 206.400 ;
        RECT 262.950 205.950 265.050 206.400 ;
        RECT 268.950 205.950 271.050 206.400 ;
        RECT 310.950 205.950 313.050 206.400 ;
        RECT 319.950 207.600 322.050 208.050 ;
        RECT 334.950 207.600 337.050 208.050 ;
        RECT 319.950 206.400 337.050 207.600 ;
        RECT 319.950 205.950 322.050 206.400 ;
        RECT 334.950 205.950 337.050 206.400 ;
        RECT 436.950 207.600 439.050 208.050 ;
        RECT 454.950 207.600 457.050 208.050 ;
        RECT 436.950 206.400 457.050 207.600 ;
        RECT 436.950 205.950 439.050 206.400 ;
        RECT 454.950 205.950 457.050 206.400 ;
        RECT 517.950 207.600 520.050 208.050 ;
        RECT 523.950 207.600 526.050 208.050 ;
        RECT 517.950 206.400 526.050 207.600 ;
        RECT 517.950 205.950 520.050 206.400 ;
        RECT 523.950 205.950 526.050 206.400 ;
        RECT 559.950 207.600 562.050 208.050 ;
        RECT 565.950 207.600 568.050 208.050 ;
        RECT 625.950 207.600 628.050 208.050 ;
        RECT 559.950 206.400 628.050 207.600 ;
        RECT 559.950 205.950 562.050 206.400 ;
        RECT 565.950 205.950 568.050 206.400 ;
        RECT 625.950 205.950 628.050 206.400 ;
        RECT 679.950 207.600 682.050 208.050 ;
        RECT 727.950 207.600 730.050 208.050 ;
        RECT 679.950 206.400 730.050 207.600 ;
        RECT 679.950 205.950 682.050 206.400 ;
        RECT 727.950 205.950 730.050 206.400 ;
        RECT 769.950 207.600 772.050 208.050 ;
        RECT 781.950 207.600 784.050 208.050 ;
        RECT 769.950 206.400 784.050 207.600 ;
        RECT 769.950 205.950 772.050 206.400 ;
        RECT 781.950 205.950 784.050 206.400 ;
        RECT 829.950 207.600 832.050 208.050 ;
        RECT 847.950 207.600 850.050 208.050 ;
        RECT 829.950 206.400 850.050 207.600 ;
        RECT 829.950 205.950 832.050 206.400 ;
        RECT 847.950 205.950 850.050 206.400 ;
        RECT 121.950 204.600 124.050 205.050 ;
        RECT 136.950 204.600 139.050 205.050 ;
        RECT 151.950 204.600 154.050 205.050 ;
        RECT 259.950 204.600 262.050 205.050 ;
        RECT 394.950 204.600 397.050 205.050 ;
        RECT 427.950 204.600 430.050 205.050 ;
        RECT 436.950 204.600 439.050 205.050 ;
        RECT 121.950 203.400 154.050 204.600 ;
        RECT 121.950 202.950 124.050 203.400 ;
        RECT 136.950 202.950 139.050 203.400 ;
        RECT 151.950 202.950 154.050 203.400 ;
        RECT 257.400 203.400 297.600 204.600 ;
        RECT 257.400 202.050 258.600 203.400 ;
        RECT 259.950 202.950 262.050 203.400 ;
        RECT 296.400 202.050 297.600 203.400 ;
        RECT 394.950 203.400 439.050 204.600 ;
        RECT 394.950 202.950 397.050 203.400 ;
        RECT 427.950 202.950 430.050 203.400 ;
        RECT 436.950 202.950 439.050 203.400 ;
        RECT 448.950 204.600 451.050 205.050 ;
        RECT 457.950 204.600 460.050 205.050 ;
        RECT 448.950 203.400 460.050 204.600 ;
        RECT 448.950 202.950 451.050 203.400 ;
        RECT 457.950 202.950 460.050 203.400 ;
        RECT 478.950 204.600 481.050 205.050 ;
        RECT 586.950 204.600 589.050 205.050 ;
        RECT 478.950 203.400 589.050 204.600 ;
        RECT 478.950 202.950 481.050 203.400 ;
        RECT 586.950 202.950 589.050 203.400 ;
        RECT 610.950 204.600 613.050 205.050 ;
        RECT 619.950 204.600 622.050 205.050 ;
        RECT 610.950 203.400 622.050 204.600 ;
        RECT 610.950 202.950 613.050 203.400 ;
        RECT 619.950 202.950 622.050 203.400 ;
        RECT 769.950 204.600 772.050 205.050 ;
        RECT 787.950 204.600 790.050 205.050 ;
        RECT 832.950 204.600 835.050 205.050 ;
        RECT 769.950 203.400 835.050 204.600 ;
        RECT 769.950 202.950 772.050 203.400 ;
        RECT 787.950 202.950 790.050 203.400 ;
        RECT 832.950 202.950 835.050 203.400 ;
        RECT 853.950 204.600 856.050 205.050 ;
        RECT 862.950 204.600 865.050 205.050 ;
        RECT 853.950 203.400 865.050 204.600 ;
        RECT 853.950 202.950 856.050 203.400 ;
        RECT 862.950 202.950 865.050 203.400 ;
        RECT 28.950 201.600 31.050 202.050 ;
        RECT 70.950 201.600 73.050 202.050 ;
        RECT 79.950 201.600 82.050 202.050 ;
        RECT 28.950 200.400 73.050 201.600 ;
        RECT 28.950 199.950 31.050 200.400 ;
        RECT 70.950 199.950 73.050 200.400 ;
        RECT 77.400 200.400 82.050 201.600 ;
        RECT 13.950 198.600 16.050 199.050 ;
        RECT 28.950 198.600 31.050 199.050 ;
        RECT 13.950 197.400 31.050 198.600 ;
        RECT 13.950 196.950 16.050 197.400 ;
        RECT 28.950 196.950 31.050 197.400 ;
        RECT 34.950 198.600 37.050 199.050 ;
        RECT 40.950 198.600 43.050 199.050 ;
        RECT 34.950 197.400 43.050 198.600 ;
        RECT 34.950 196.950 37.050 197.400 ;
        RECT 40.950 196.950 43.050 197.400 ;
        RECT 58.950 198.600 61.050 199.050 ;
        RECT 73.950 198.600 76.050 199.050 ;
        RECT 58.950 197.400 76.050 198.600 ;
        RECT 58.950 196.950 61.050 197.400 ;
        RECT 73.950 196.950 76.050 197.400 ;
        RECT 77.400 196.050 78.600 200.400 ;
        RECT 79.950 199.950 82.050 200.400 ;
        RECT 130.950 201.600 133.050 202.050 ;
        RECT 142.950 201.600 145.050 202.050 ;
        RECT 178.950 201.600 181.050 202.050 ;
        RECT 130.950 200.400 181.050 201.600 ;
        RECT 130.950 199.950 133.050 200.400 ;
        RECT 142.950 199.950 145.050 200.400 ;
        RECT 178.950 199.950 181.050 200.400 ;
        RECT 217.950 201.600 220.050 202.050 ;
        RECT 250.950 201.600 253.050 202.050 ;
        RECT 217.950 200.400 253.050 201.600 ;
        RECT 217.950 199.950 220.050 200.400 ;
        RECT 250.950 199.950 253.050 200.400 ;
        RECT 256.950 199.950 259.050 202.050 ;
        RECT 280.950 201.600 283.050 202.050 ;
        RECT 289.950 201.600 292.050 202.050 ;
        RECT 280.950 200.400 292.050 201.600 ;
        RECT 280.950 199.950 283.050 200.400 ;
        RECT 289.950 199.950 292.050 200.400 ;
        RECT 295.950 199.950 298.050 202.050 ;
        RECT 301.950 201.600 304.050 202.050 ;
        RECT 328.950 201.600 331.050 202.050 ;
        RECT 301.950 200.400 331.050 201.600 ;
        RECT 301.950 199.950 304.050 200.400 ;
        RECT 328.950 199.950 331.050 200.400 ;
        RECT 334.950 201.600 337.050 202.050 ;
        RECT 343.950 201.600 346.050 202.050 ;
        RECT 334.950 200.400 346.050 201.600 ;
        RECT 334.950 199.950 337.050 200.400 ;
        RECT 343.950 199.950 346.050 200.400 ;
        RECT 355.950 201.600 358.050 202.050 ;
        RECT 673.950 201.600 676.050 202.050 ;
        RECT 697.950 201.600 700.050 202.050 ;
        RECT 700.950 201.600 703.050 202.050 ;
        RECT 355.950 200.400 703.050 201.600 ;
        RECT 355.950 199.950 358.050 200.400 ;
        RECT 673.950 199.950 676.050 200.400 ;
        RECT 697.950 199.950 700.050 200.400 ;
        RECT 700.950 199.950 703.050 200.400 ;
        RECT 706.950 201.600 709.050 202.050 ;
        RECT 763.950 201.600 766.050 202.050 ;
        RECT 790.950 201.600 793.050 202.050 ;
        RECT 796.950 201.600 799.050 202.050 ;
        RECT 706.950 200.400 799.050 201.600 ;
        RECT 706.950 199.950 709.050 200.400 ;
        RECT 763.950 199.950 766.050 200.400 ;
        RECT 790.950 199.950 793.050 200.400 ;
        RECT 796.950 199.950 799.050 200.400 ;
        RECT 808.950 201.600 811.050 202.050 ;
        RECT 823.950 201.600 826.050 202.050 ;
        RECT 808.950 200.400 826.050 201.600 ;
        RECT 808.950 199.950 811.050 200.400 ;
        RECT 823.950 199.950 826.050 200.400 ;
        RECT 838.950 201.600 841.050 202.050 ;
        RECT 844.950 201.600 847.050 202.050 ;
        RECT 838.950 200.400 847.050 201.600 ;
        RECT 838.950 199.950 841.050 200.400 ;
        RECT 844.950 199.950 847.050 200.400 ;
        RECT 79.950 198.600 82.050 199.050 ;
        RECT 85.950 198.600 88.050 199.050 ;
        RECT 100.950 198.600 103.050 199.050 ;
        RECT 79.950 197.400 103.050 198.600 ;
        RECT 79.950 196.950 82.050 197.400 ;
        RECT 85.950 196.950 88.050 197.400 ;
        RECT 100.950 196.950 103.050 197.400 ;
        RECT 157.950 198.600 160.050 199.050 ;
        RECT 169.950 198.600 172.050 199.050 ;
        RECT 157.950 197.400 172.050 198.600 ;
        RECT 157.950 196.950 160.050 197.400 ;
        RECT 169.950 196.950 172.050 197.400 ;
        RECT 175.950 198.600 178.050 199.050 ;
        RECT 181.950 198.600 184.050 199.050 ;
        RECT 175.950 197.400 184.050 198.600 ;
        RECT 175.950 196.950 178.050 197.400 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 232.950 198.600 235.050 199.050 ;
        RECT 253.950 198.600 256.050 199.050 ;
        RECT 292.950 198.600 295.050 199.050 ;
        RECT 232.950 197.400 295.050 198.600 ;
        RECT 232.950 196.950 235.050 197.400 ;
        RECT 253.950 196.950 256.050 197.400 ;
        RECT 292.950 196.950 295.050 197.400 ;
        RECT 307.950 198.600 310.050 199.050 ;
        RECT 337.950 198.600 340.050 199.050 ;
        RECT 307.950 197.400 340.050 198.600 ;
        RECT 307.950 196.950 310.050 197.400 ;
        RECT 337.950 196.950 340.050 197.400 ;
        RECT 358.950 198.600 361.050 199.050 ;
        RECT 400.950 198.600 403.050 199.050 ;
        RECT 358.950 197.400 403.050 198.600 ;
        RECT 358.950 196.950 361.050 197.400 ;
        RECT 400.950 196.950 403.050 197.400 ;
        RECT 409.950 198.600 412.050 199.050 ;
        RECT 430.950 198.600 433.050 199.050 ;
        RECT 451.950 198.600 454.050 199.050 ;
        RECT 472.950 198.600 475.050 199.050 ;
        RECT 409.950 197.400 475.050 198.600 ;
        RECT 409.950 196.950 412.050 197.400 ;
        RECT 430.950 196.950 433.050 197.400 ;
        RECT 451.950 196.950 454.050 197.400 ;
        RECT 472.950 196.950 475.050 197.400 ;
        RECT 553.950 198.600 556.050 199.050 ;
        RECT 553.950 197.400 564.600 198.600 ;
        RECT 553.950 196.950 556.050 197.400 ;
        RECT 563.400 196.050 564.600 197.400 ;
        RECT 607.950 196.950 610.050 199.050 ;
        RECT 613.950 198.600 616.050 199.050 ;
        RECT 622.950 198.600 625.050 199.050 ;
        RECT 613.950 197.400 625.050 198.600 ;
        RECT 613.950 196.950 616.050 197.400 ;
        RECT 622.950 196.950 625.050 197.400 ;
        RECT 628.950 196.950 631.050 199.050 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 682.950 198.600 685.050 199.050 ;
        RECT 688.950 198.600 691.050 199.050 ;
        RECT 682.950 197.400 691.050 198.600 ;
        RECT 682.950 196.950 685.050 197.400 ;
        RECT 688.950 196.950 691.050 197.400 ;
        RECT 694.950 198.600 697.050 199.050 ;
        RECT 709.950 198.600 712.050 199.050 ;
        RECT 694.950 197.400 712.050 198.600 ;
        RECT 694.950 196.950 697.050 197.400 ;
        RECT 709.950 196.950 712.050 197.400 ;
        RECT 733.950 198.600 736.050 199.050 ;
        RECT 766.950 198.600 769.050 199.050 ;
        RECT 733.950 197.400 769.050 198.600 ;
        RECT 733.950 196.950 736.050 197.400 ;
        RECT 766.950 196.950 769.050 197.400 ;
        RECT 787.950 198.600 790.050 199.050 ;
        RECT 802.950 198.600 805.050 199.050 ;
        RECT 823.950 198.600 826.050 199.050 ;
        RECT 787.950 197.400 805.050 198.600 ;
        RECT 787.950 196.950 790.050 197.400 ;
        RECT 802.950 196.950 805.050 197.400 ;
        RECT 806.400 197.400 826.050 198.600 ;
        RECT 37.950 195.600 40.050 196.050 ;
        RECT 64.950 195.600 67.050 196.050 ;
        RECT 37.950 194.400 67.050 195.600 ;
        RECT 37.950 193.950 40.050 194.400 ;
        RECT 64.950 193.950 67.050 194.400 ;
        RECT 76.950 193.950 79.050 196.050 ;
        RECT 82.950 195.600 85.050 196.050 ;
        RECT 94.950 195.600 97.050 196.050 ;
        RECT 118.950 195.600 121.050 196.050 ;
        RECT 82.950 194.400 121.050 195.600 ;
        RECT 82.950 193.950 85.050 194.400 ;
        RECT 94.950 193.950 97.050 194.400 ;
        RECT 118.950 193.950 121.050 194.400 ;
        RECT 172.950 195.600 175.050 196.050 ;
        RECT 193.950 195.600 196.050 196.050 ;
        RECT 172.950 194.400 196.050 195.600 ;
        RECT 172.950 193.950 175.050 194.400 ;
        RECT 193.950 193.950 196.050 194.400 ;
        RECT 331.950 195.600 334.050 196.050 ;
        RECT 352.950 195.600 355.050 196.050 ;
        RECT 331.950 194.400 355.050 195.600 ;
        RECT 331.950 193.950 334.050 194.400 ;
        RECT 352.950 193.950 355.050 194.400 ;
        RECT 382.950 195.600 385.050 196.050 ;
        RECT 391.950 195.600 394.050 196.050 ;
        RECT 382.950 194.400 394.050 195.600 ;
        RECT 382.950 193.950 385.050 194.400 ;
        RECT 391.950 193.950 394.050 194.400 ;
        RECT 415.950 195.600 418.050 196.050 ;
        RECT 421.950 195.600 424.050 196.050 ;
        RECT 415.950 194.400 424.050 195.600 ;
        RECT 415.950 193.950 418.050 194.400 ;
        RECT 421.950 193.950 424.050 194.400 ;
        RECT 424.950 195.600 427.050 196.050 ;
        RECT 433.950 195.600 436.050 196.050 ;
        RECT 424.950 194.400 436.050 195.600 ;
        RECT 424.950 193.950 427.050 194.400 ;
        RECT 433.950 193.950 436.050 194.400 ;
        RECT 445.950 195.600 448.050 196.050 ;
        RECT 454.950 195.600 457.050 196.050 ;
        RECT 445.950 194.400 457.050 195.600 ;
        RECT 445.950 193.950 448.050 194.400 ;
        RECT 454.950 193.950 457.050 194.400 ;
        RECT 469.950 195.600 472.050 196.050 ;
        RECT 511.950 195.600 514.050 196.050 ;
        RECT 469.950 194.400 514.050 195.600 ;
        RECT 469.950 193.950 472.050 194.400 ;
        RECT 511.950 193.950 514.050 194.400 ;
        RECT 517.950 195.600 520.050 196.050 ;
        RECT 529.950 195.600 532.050 196.050 ;
        RECT 517.950 194.400 532.050 195.600 ;
        RECT 517.950 193.950 520.050 194.400 ;
        RECT 529.950 193.950 532.050 194.400 ;
        RECT 562.950 193.950 565.050 196.050 ;
        RECT 608.400 195.600 609.600 196.950 ;
        RECT 629.400 195.600 630.600 196.950 ;
        RECT 643.950 195.600 646.050 196.050 ;
        RECT 608.400 194.400 646.050 195.600 ;
        RECT 647.400 195.600 648.600 196.950 ;
        RECT 667.950 195.600 670.050 196.050 ;
        RECT 647.400 194.400 670.050 195.600 ;
        RECT 643.950 193.950 646.050 194.400 ;
        RECT 667.950 193.950 670.050 194.400 ;
        RECT 676.950 195.600 679.050 196.050 ;
        RECT 685.950 195.600 688.050 196.050 ;
        RECT 676.950 194.400 688.050 195.600 ;
        RECT 676.950 193.950 679.050 194.400 ;
        RECT 685.950 193.950 688.050 194.400 ;
        RECT 751.950 195.600 754.050 196.050 ;
        RECT 806.400 195.600 807.600 197.400 ;
        RECT 823.950 196.950 826.050 197.400 ;
        RECT 751.950 194.400 807.600 195.600 ;
        RECT 751.950 193.950 754.050 194.400 ;
        RECT 55.950 192.600 58.050 193.050 ;
        RECT 82.950 192.600 85.050 193.050 ;
        RECT 55.950 191.400 85.050 192.600 ;
        RECT 55.950 190.950 58.050 191.400 ;
        RECT 82.950 190.950 85.050 191.400 ;
        RECT 187.950 192.600 190.050 193.050 ;
        RECT 196.950 192.600 199.050 193.050 ;
        RECT 187.950 191.400 199.050 192.600 ;
        RECT 187.950 190.950 190.050 191.400 ;
        RECT 196.950 190.950 199.050 191.400 ;
        RECT 298.950 192.600 301.050 193.050 ;
        RECT 313.950 192.600 316.050 193.050 ;
        RECT 346.950 192.600 349.050 193.050 ;
        RECT 298.950 191.400 349.050 192.600 ;
        RECT 298.950 190.950 301.050 191.400 ;
        RECT 313.950 190.950 316.050 191.400 ;
        RECT 346.950 190.950 349.050 191.400 ;
        RECT 349.950 192.600 352.050 193.050 ;
        RECT 367.950 192.600 370.050 193.050 ;
        RECT 379.950 192.600 382.050 193.050 ;
        RECT 349.950 191.400 382.050 192.600 ;
        RECT 349.950 190.950 352.050 191.400 ;
        RECT 367.950 190.950 370.050 191.400 ;
        RECT 379.950 190.950 382.050 191.400 ;
        RECT 415.950 192.600 418.050 193.050 ;
        RECT 427.950 192.600 430.050 193.050 ;
        RECT 415.950 191.400 430.050 192.600 ;
        RECT 415.950 190.950 418.050 191.400 ;
        RECT 427.950 190.950 430.050 191.400 ;
        RECT 454.950 192.600 457.050 193.050 ;
        RECT 490.950 192.600 493.050 193.050 ;
        RECT 454.950 191.400 493.050 192.600 ;
        RECT 454.950 190.950 457.050 191.400 ;
        RECT 490.950 190.950 493.050 191.400 ;
        RECT 496.950 192.600 499.050 193.050 ;
        RECT 517.950 192.600 520.050 193.050 ;
        RECT 496.950 191.400 520.050 192.600 ;
        RECT 496.950 190.950 499.050 191.400 ;
        RECT 517.950 190.950 520.050 191.400 ;
        RECT 550.950 192.600 553.050 193.050 ;
        RECT 559.950 192.600 562.050 193.050 ;
        RECT 550.950 191.400 562.050 192.600 ;
        RECT 550.950 190.950 553.050 191.400 ;
        RECT 559.950 190.950 562.050 191.400 ;
        RECT 601.950 192.600 604.050 193.050 ;
        RECT 625.950 192.600 628.050 193.050 ;
        RECT 601.950 191.400 628.050 192.600 ;
        RECT 601.950 190.950 604.050 191.400 ;
        RECT 625.950 190.950 628.050 191.400 ;
        RECT 640.950 192.600 643.050 193.050 ;
        RECT 649.950 192.600 652.050 193.050 ;
        RECT 640.950 191.400 652.050 192.600 ;
        RECT 640.950 190.950 643.050 191.400 ;
        RECT 649.950 190.950 652.050 191.400 ;
        RECT 685.950 192.600 688.050 193.050 ;
        RECT 703.950 192.600 706.050 193.050 ;
        RECT 685.950 191.400 706.050 192.600 ;
        RECT 685.950 190.950 688.050 191.400 ;
        RECT 703.950 190.950 706.050 191.400 ;
        RECT 718.950 192.600 721.050 193.050 ;
        RECT 733.950 192.600 736.050 193.050 ;
        RECT 751.950 192.600 754.050 193.050 ;
        RECT 718.950 191.400 754.050 192.600 ;
        RECT 718.950 190.950 721.050 191.400 ;
        RECT 733.950 190.950 736.050 191.400 ;
        RECT 751.950 190.950 754.050 191.400 ;
        RECT 781.950 192.600 784.050 193.050 ;
        RECT 844.950 192.600 847.050 193.050 ;
        RECT 781.950 191.400 847.050 192.600 ;
        RECT 781.950 190.950 784.050 191.400 ;
        RECT 844.950 190.950 847.050 191.400 ;
        RECT 25.950 189.600 28.050 190.050 ;
        RECT 34.950 189.600 37.050 190.050 ;
        RECT 25.950 188.400 37.050 189.600 ;
        RECT 25.950 187.950 28.050 188.400 ;
        RECT 34.950 187.950 37.050 188.400 ;
        RECT 46.950 189.600 49.050 190.050 ;
        RECT 55.950 189.600 58.050 190.050 ;
        RECT 46.950 188.400 58.050 189.600 ;
        RECT 46.950 187.950 49.050 188.400 ;
        RECT 55.950 187.950 58.050 188.400 ;
        RECT 67.950 189.600 70.050 190.050 ;
        RECT 76.950 189.600 79.050 190.050 ;
        RECT 67.950 188.400 79.050 189.600 ;
        RECT 67.950 187.950 70.050 188.400 ;
        RECT 76.950 187.950 79.050 188.400 ;
        RECT 79.950 189.600 82.050 190.050 ;
        RECT 97.950 189.600 100.050 190.050 ;
        RECT 79.950 188.400 100.050 189.600 ;
        RECT 79.950 187.950 82.050 188.400 ;
        RECT 97.950 187.950 100.050 188.400 ;
        RECT 313.950 189.600 316.050 190.050 ;
        RECT 340.950 189.600 343.050 190.050 ;
        RECT 313.950 188.400 343.050 189.600 ;
        RECT 313.950 187.950 316.050 188.400 ;
        RECT 340.950 187.950 343.050 188.400 ;
        RECT 352.950 189.600 355.050 190.050 ;
        RECT 535.950 189.600 538.050 190.050 ;
        RECT 352.950 188.400 538.050 189.600 ;
        RECT 352.950 187.950 355.050 188.400 ;
        RECT 535.950 187.950 538.050 188.400 ;
        RECT 556.950 189.600 559.050 190.050 ;
        RECT 568.950 189.600 571.050 190.050 ;
        RECT 556.950 188.400 571.050 189.600 ;
        RECT 556.950 187.950 559.050 188.400 ;
        RECT 568.950 187.950 571.050 188.400 ;
        RECT 664.950 189.600 667.050 190.050 ;
        RECT 670.950 189.600 673.050 190.050 ;
        RECT 718.950 189.600 721.050 190.050 ;
        RECT 664.950 188.400 721.050 189.600 ;
        RECT 664.950 187.950 667.050 188.400 ;
        RECT 670.950 187.950 673.050 188.400 ;
        RECT 718.950 187.950 721.050 188.400 ;
        RECT 793.950 189.600 796.050 190.050 ;
        RECT 811.950 189.600 814.050 190.050 ;
        RECT 793.950 188.400 814.050 189.600 ;
        RECT 793.950 187.950 796.050 188.400 ;
        RECT 811.950 187.950 814.050 188.400 ;
        RECT 16.950 186.600 19.050 187.050 ;
        RECT 40.950 186.600 43.050 187.050 ;
        RECT 70.950 186.600 73.050 187.050 ;
        RECT 16.950 185.400 73.050 186.600 ;
        RECT 16.950 184.950 19.050 185.400 ;
        RECT 40.950 184.950 43.050 185.400 ;
        RECT 70.950 184.950 73.050 185.400 ;
        RECT 268.950 186.600 271.050 187.050 ;
        RECT 355.950 186.600 358.050 187.050 ;
        RECT 268.950 185.400 358.050 186.600 ;
        RECT 268.950 184.950 271.050 185.400 ;
        RECT 355.950 184.950 358.050 185.400 ;
        RECT 478.950 186.600 481.050 187.050 ;
        RECT 505.950 186.600 508.050 187.050 ;
        RECT 478.950 185.400 508.050 186.600 ;
        RECT 478.950 184.950 481.050 185.400 ;
        RECT 505.950 184.950 508.050 185.400 ;
        RECT 631.950 186.600 634.050 187.050 ;
        RECT 748.950 186.600 751.050 187.050 ;
        RECT 631.950 185.400 751.050 186.600 ;
        RECT 631.950 184.950 634.050 185.400 ;
        RECT 748.950 184.950 751.050 185.400 ;
        RECT 19.950 183.600 22.050 184.050 ;
        RECT 31.950 183.600 34.050 184.050 ;
        RECT 79.950 183.600 82.050 184.050 ;
        RECT 19.950 182.400 82.050 183.600 ;
        RECT 19.950 181.950 22.050 182.400 ;
        RECT 31.950 181.950 34.050 182.400 ;
        RECT 79.950 181.950 82.050 182.400 ;
        RECT 376.950 183.600 379.050 184.050 ;
        RECT 409.950 183.600 412.050 184.050 ;
        RECT 376.950 182.400 412.050 183.600 ;
        RECT 376.950 181.950 379.050 182.400 ;
        RECT 409.950 181.950 412.050 182.400 ;
        RECT 418.950 183.600 421.050 184.050 ;
        RECT 475.950 183.600 478.050 184.050 ;
        RECT 418.950 182.400 478.050 183.600 ;
        RECT 418.950 181.950 421.050 182.400 ;
        RECT 475.950 181.950 478.050 182.400 ;
        RECT 571.950 183.600 574.050 184.050 ;
        RECT 583.950 183.600 586.050 184.050 ;
        RECT 664.950 183.600 667.050 184.050 ;
        RECT 571.950 182.400 667.050 183.600 ;
        RECT 571.950 181.950 574.050 182.400 ;
        RECT 583.950 181.950 586.050 182.400 ;
        RECT 664.950 181.950 667.050 182.400 ;
        RECT 346.950 180.600 349.050 181.050 ;
        RECT 403.950 180.600 406.050 181.050 ;
        RECT 346.950 179.400 406.050 180.600 ;
        RECT 346.950 178.950 349.050 179.400 ;
        RECT 403.950 178.950 406.050 179.400 ;
        RECT 412.950 180.600 415.050 181.050 ;
        RECT 514.950 180.600 517.050 181.050 ;
        RECT 412.950 179.400 517.050 180.600 ;
        RECT 412.950 178.950 415.050 179.400 ;
        RECT 514.950 178.950 517.050 179.400 ;
        RECT 520.950 180.600 523.050 181.050 ;
        RECT 544.950 180.600 547.050 181.050 ;
        RECT 556.950 180.600 559.050 181.050 ;
        RECT 520.950 179.400 559.050 180.600 ;
        RECT 520.950 178.950 523.050 179.400 ;
        RECT 544.950 178.950 547.050 179.400 ;
        RECT 556.950 178.950 559.050 179.400 ;
        RECT 565.950 180.600 568.050 181.050 ;
        RECT 631.950 180.600 634.050 181.050 ;
        RECT 565.950 179.400 634.050 180.600 ;
        RECT 565.950 178.950 568.050 179.400 ;
        RECT 631.950 178.950 634.050 179.400 ;
        RECT 661.950 180.600 664.050 181.050 ;
        RECT 730.950 180.600 733.050 181.050 ;
        RECT 661.950 179.400 733.050 180.600 ;
        RECT 661.950 178.950 664.050 179.400 ;
        RECT 730.950 178.950 733.050 179.400 ;
        RECT 838.950 180.600 841.050 181.050 ;
        RECT 844.950 180.600 847.050 181.050 ;
        RECT 838.950 179.400 847.050 180.600 ;
        RECT 838.950 178.950 841.050 179.400 ;
        RECT 844.950 178.950 847.050 179.400 ;
        RECT 13.950 177.600 16.050 178.050 ;
        RECT 64.950 177.600 67.050 178.050 ;
        RECT 13.950 176.400 67.050 177.600 ;
        RECT 13.950 175.950 16.050 176.400 ;
        RECT 64.950 175.950 67.050 176.400 ;
        RECT 232.950 177.600 235.050 178.050 ;
        RECT 241.950 177.600 244.050 178.050 ;
        RECT 301.950 177.600 304.050 178.050 ;
        RECT 232.950 176.400 304.050 177.600 ;
        RECT 232.950 175.950 235.050 176.400 ;
        RECT 241.950 175.950 244.050 176.400 ;
        RECT 301.950 175.950 304.050 176.400 ;
        RECT 310.950 177.600 313.050 178.050 ;
        RECT 373.950 177.600 376.050 178.050 ;
        RECT 310.950 176.400 376.050 177.600 ;
        RECT 310.950 175.950 313.050 176.400 ;
        RECT 373.950 175.950 376.050 176.400 ;
        RECT 523.950 177.600 526.050 178.050 ;
        RECT 538.950 177.600 541.050 178.050 ;
        RECT 550.950 177.600 553.050 178.050 ;
        RECT 523.950 176.400 553.050 177.600 ;
        RECT 523.950 175.950 526.050 176.400 ;
        RECT 538.950 175.950 541.050 176.400 ;
        RECT 550.950 175.950 553.050 176.400 ;
        RECT 637.950 177.600 640.050 178.050 ;
        RECT 655.950 177.600 658.050 178.050 ;
        RECT 637.950 176.400 658.050 177.600 ;
        RECT 637.950 175.950 640.050 176.400 ;
        RECT 655.950 175.950 658.050 176.400 ;
        RECT 697.950 177.600 700.050 178.050 ;
        RECT 703.950 177.600 706.050 178.050 ;
        RECT 697.950 176.400 706.050 177.600 ;
        RECT 697.950 175.950 700.050 176.400 ;
        RECT 703.950 175.950 706.050 176.400 ;
        RECT 769.950 177.600 772.050 178.050 ;
        RECT 820.950 177.600 823.050 178.050 ;
        RECT 769.950 176.400 823.050 177.600 ;
        RECT 769.950 175.950 772.050 176.400 ;
        RECT 820.950 175.950 823.050 176.400 ;
        RECT 838.950 177.600 841.050 178.050 ;
        RECT 850.950 177.600 853.050 178.050 ;
        RECT 838.950 176.400 853.050 177.600 ;
        RECT 838.950 175.950 841.050 176.400 ;
        RECT 850.950 175.950 853.050 176.400 ;
        RECT 31.950 174.600 34.050 175.050 ;
        RECT 43.950 174.600 46.050 175.050 ;
        RECT 31.950 173.400 46.050 174.600 ;
        RECT 31.950 172.950 34.050 173.400 ;
        RECT 43.950 172.950 46.050 173.400 ;
        RECT 97.950 174.600 100.050 175.050 ;
        RECT 115.950 174.600 118.050 175.050 ;
        RECT 139.950 174.600 142.050 175.050 ;
        RECT 97.950 173.400 142.050 174.600 ;
        RECT 97.950 172.950 100.050 173.400 ;
        RECT 115.950 172.950 118.050 173.400 ;
        RECT 139.950 172.950 142.050 173.400 ;
        RECT 169.950 174.600 172.050 175.050 ;
        RECT 214.950 174.600 217.050 175.050 ;
        RECT 169.950 173.400 217.050 174.600 ;
        RECT 169.950 172.950 172.050 173.400 ;
        RECT 214.950 172.950 217.050 173.400 ;
        RECT 226.950 174.600 229.050 175.050 ;
        RECT 244.950 174.600 247.050 175.050 ;
        RECT 226.950 173.400 247.050 174.600 ;
        RECT 226.950 172.950 229.050 173.400 ;
        RECT 244.950 172.950 247.050 173.400 ;
        RECT 472.950 174.600 475.050 175.050 ;
        RECT 505.950 174.600 508.050 175.050 ;
        RECT 472.950 173.400 508.050 174.600 ;
        RECT 472.950 172.950 475.050 173.400 ;
        RECT 505.950 172.950 508.050 173.400 ;
        RECT 532.950 174.600 535.050 175.050 ;
        RECT 652.950 174.600 655.050 175.050 ;
        RECT 532.950 173.400 655.050 174.600 ;
        RECT 532.950 172.950 535.050 173.400 ;
        RECT 652.950 172.950 655.050 173.400 ;
        RECT 658.950 174.600 661.050 175.050 ;
        RECT 673.950 174.600 676.050 175.050 ;
        RECT 679.950 174.600 682.050 175.050 ;
        RECT 706.950 174.600 709.050 175.050 ;
        RECT 658.950 173.400 709.050 174.600 ;
        RECT 658.950 172.950 661.050 173.400 ;
        RECT 673.950 172.950 676.050 173.400 ;
        RECT 679.950 172.950 682.050 173.400 ;
        RECT 706.950 172.950 709.050 173.400 ;
        RECT 799.950 174.600 802.050 175.050 ;
        RECT 805.950 174.600 808.050 175.050 ;
        RECT 799.950 173.400 808.050 174.600 ;
        RECT 799.950 172.950 802.050 173.400 ;
        RECT 805.950 172.950 808.050 173.400 ;
        RECT 850.950 174.600 853.050 175.050 ;
        RECT 862.950 174.600 865.050 175.050 ;
        RECT 850.950 173.400 865.050 174.600 ;
        RECT 850.950 172.950 853.050 173.400 ;
        RECT 862.950 172.950 865.050 173.400 ;
        RECT 4.950 171.600 7.050 172.050 ;
        RECT 25.950 171.600 28.050 172.050 ;
        RECT 4.950 170.400 28.050 171.600 ;
        RECT 4.950 169.950 7.050 170.400 ;
        RECT 25.950 169.950 28.050 170.400 ;
        RECT 64.950 171.600 67.050 172.050 ;
        RECT 91.950 171.600 94.050 172.050 ;
        RECT 64.950 170.400 94.050 171.600 ;
        RECT 64.950 169.950 67.050 170.400 ;
        RECT 91.950 169.950 94.050 170.400 ;
        RECT 100.950 171.600 103.050 172.050 ;
        RECT 133.950 171.600 136.050 172.050 ;
        RECT 100.950 170.400 136.050 171.600 ;
        RECT 100.950 169.950 103.050 170.400 ;
        RECT 133.950 169.950 136.050 170.400 ;
        RECT 139.950 171.600 142.050 172.050 ;
        RECT 148.950 171.600 151.050 172.050 ;
        RECT 139.950 170.400 151.050 171.600 ;
        RECT 139.950 169.950 142.050 170.400 ;
        RECT 148.950 169.950 151.050 170.400 ;
        RECT 178.950 171.600 181.050 172.050 ;
        RECT 190.950 171.600 193.050 172.050 ;
        RECT 199.950 171.600 202.050 172.050 ;
        RECT 178.950 170.400 202.050 171.600 ;
        RECT 178.950 169.950 181.050 170.400 ;
        RECT 190.950 169.950 193.050 170.400 ;
        RECT 199.950 169.950 202.050 170.400 ;
        RECT 205.950 171.600 208.050 172.050 ;
        RECT 229.950 171.600 232.050 172.050 ;
        RECT 205.950 170.400 232.050 171.600 ;
        RECT 205.950 169.950 208.050 170.400 ;
        RECT 229.950 169.950 232.050 170.400 ;
        RECT 274.950 171.600 277.050 172.050 ;
        RECT 331.950 171.600 334.050 172.050 ;
        RECT 337.950 171.600 340.050 172.050 ;
        RECT 274.950 170.400 340.050 171.600 ;
        RECT 274.950 169.950 277.050 170.400 ;
        RECT 331.950 169.950 334.050 170.400 ;
        RECT 337.950 169.950 340.050 170.400 ;
        RECT 364.950 171.600 367.050 172.050 ;
        RECT 382.950 171.600 385.050 172.050 ;
        RECT 364.950 170.400 385.050 171.600 ;
        RECT 364.950 169.950 367.050 170.400 ;
        RECT 382.950 169.950 385.050 170.400 ;
        RECT 442.950 171.600 445.050 172.050 ;
        RECT 457.950 171.600 460.050 172.050 ;
        RECT 487.950 171.600 490.050 172.050 ;
        RECT 442.950 170.400 460.050 171.600 ;
        RECT 442.950 169.950 445.050 170.400 ;
        RECT 457.950 169.950 460.050 170.400 ;
        RECT 485.400 170.400 490.050 171.600 ;
        RECT 52.950 168.600 55.050 169.050 ;
        RECT 26.400 167.400 55.050 168.600 ;
        RECT 10.950 165.600 13.050 166.050 ;
        RECT 22.950 165.600 25.050 166.050 ;
        RECT 26.400 165.600 27.600 167.400 ;
        RECT 52.950 166.950 55.050 167.400 ;
        RECT 58.950 168.600 61.050 169.050 ;
        RECT 91.950 168.600 94.050 169.050 ;
        RECT 58.950 167.400 94.050 168.600 ;
        RECT 58.950 166.950 61.050 167.400 ;
        RECT 91.950 166.950 94.050 167.400 ;
        RECT 124.950 168.600 127.050 169.050 ;
        RECT 157.950 168.600 160.050 169.050 ;
        RECT 124.950 167.400 160.050 168.600 ;
        RECT 124.950 166.950 127.050 167.400 ;
        RECT 157.950 166.950 160.050 167.400 ;
        RECT 181.950 168.600 184.050 169.050 ;
        RECT 304.950 168.600 307.050 169.050 ;
        RECT 181.950 167.400 307.050 168.600 ;
        RECT 181.950 166.950 184.050 167.400 ;
        RECT 304.950 166.950 307.050 167.400 ;
        RECT 325.950 168.600 328.050 169.050 ;
        RECT 346.950 168.600 349.050 169.050 ;
        RECT 325.950 167.400 349.050 168.600 ;
        RECT 325.950 166.950 328.050 167.400 ;
        RECT 346.950 166.950 349.050 167.400 ;
        RECT 355.950 168.600 358.050 169.050 ;
        RECT 367.950 168.600 370.050 169.050 ;
        RECT 355.950 167.400 370.050 168.600 ;
        RECT 355.950 166.950 358.050 167.400 ;
        RECT 367.950 166.950 370.050 167.400 ;
        RECT 388.950 168.600 391.050 169.050 ;
        RECT 412.950 168.600 415.050 169.050 ;
        RECT 388.950 167.400 415.050 168.600 ;
        RECT 388.950 166.950 391.050 167.400 ;
        RECT 412.950 166.950 415.050 167.400 ;
        RECT 433.950 168.600 436.050 169.050 ;
        RECT 439.950 168.600 442.050 169.050 ;
        RECT 433.950 167.400 442.050 168.600 ;
        RECT 433.950 166.950 436.050 167.400 ;
        RECT 439.950 166.950 442.050 167.400 ;
        RECT 460.950 168.600 463.050 169.050 ;
        RECT 466.950 168.600 469.050 169.050 ;
        RECT 460.950 167.400 469.050 168.600 ;
        RECT 460.950 166.950 463.050 167.400 ;
        RECT 466.950 166.950 469.050 167.400 ;
        RECT 485.400 166.050 486.600 170.400 ;
        RECT 487.950 169.950 490.050 170.400 ;
        RECT 508.950 171.600 511.050 172.050 ;
        RECT 514.950 171.600 517.050 172.050 ;
        RECT 508.950 170.400 517.050 171.600 ;
        RECT 508.950 169.950 511.050 170.400 ;
        RECT 514.950 169.950 517.050 170.400 ;
        RECT 529.950 171.600 532.050 172.050 ;
        RECT 577.950 171.600 580.050 172.050 ;
        RECT 529.950 170.400 580.050 171.600 ;
        RECT 529.950 169.950 532.050 170.400 ;
        RECT 577.950 169.950 580.050 170.400 ;
        RECT 601.950 171.600 604.050 172.050 ;
        RECT 613.950 171.600 616.050 172.050 ;
        RECT 601.950 170.400 616.050 171.600 ;
        RECT 601.950 169.950 604.050 170.400 ;
        RECT 613.950 169.950 616.050 170.400 ;
        RECT 652.950 171.600 655.050 172.050 ;
        RECT 667.950 171.600 670.050 172.050 ;
        RECT 652.950 170.400 670.050 171.600 ;
        RECT 652.950 169.950 655.050 170.400 ;
        RECT 667.950 169.950 670.050 170.400 ;
        RECT 691.950 171.600 694.050 172.050 ;
        RECT 706.950 171.600 709.050 172.050 ;
        RECT 709.950 171.600 712.050 172.050 ;
        RECT 736.950 171.600 739.050 172.050 ;
        RECT 745.950 171.600 748.050 172.050 ;
        RECT 691.950 170.400 699.600 171.600 ;
        RECT 691.950 169.950 694.050 170.400 ;
        RECT 496.950 168.600 499.050 169.050 ;
        RECT 538.950 168.600 541.050 169.050 ;
        RECT 496.950 167.400 541.050 168.600 ;
        RECT 496.950 166.950 499.050 167.400 ;
        RECT 538.950 166.950 541.050 167.400 ;
        RECT 553.950 168.600 556.050 169.050 ;
        RECT 559.950 168.600 562.050 169.050 ;
        RECT 553.950 167.400 562.050 168.600 ;
        RECT 553.950 166.950 556.050 167.400 ;
        RECT 559.950 166.950 562.050 167.400 ;
        RECT 583.950 168.600 586.050 169.050 ;
        RECT 595.950 168.600 598.050 169.050 ;
        RECT 583.950 167.400 598.050 168.600 ;
        RECT 583.950 166.950 586.050 167.400 ;
        RECT 595.950 166.950 598.050 167.400 ;
        RECT 616.950 168.600 619.050 169.050 ;
        RECT 622.950 168.600 625.050 169.050 ;
        RECT 616.950 167.400 625.050 168.600 ;
        RECT 616.950 166.950 619.050 167.400 ;
        RECT 622.950 166.950 625.050 167.400 ;
        RECT 625.950 168.600 628.050 169.050 ;
        RECT 646.950 168.600 649.050 169.050 ;
        RECT 673.950 168.600 676.050 169.050 ;
        RECT 625.950 167.400 649.050 168.600 ;
        RECT 625.950 166.950 628.050 167.400 ;
        RECT 646.950 166.950 649.050 167.400 ;
        RECT 650.400 167.400 676.050 168.600 ;
        RECT 650.400 166.050 651.600 167.400 ;
        RECT 673.950 166.950 676.050 167.400 ;
        RECT 698.400 166.050 699.600 170.400 ;
        RECT 706.950 170.400 748.050 171.600 ;
        RECT 706.950 169.950 709.050 170.400 ;
        RECT 709.950 169.950 712.050 170.400 ;
        RECT 736.950 169.950 739.050 170.400 ;
        RECT 745.950 169.950 748.050 170.400 ;
        RECT 748.950 171.600 751.050 172.050 ;
        RECT 784.950 171.600 787.050 172.050 ;
        RECT 748.950 170.400 787.050 171.600 ;
        RECT 748.950 169.950 751.050 170.400 ;
        RECT 784.950 169.950 787.050 170.400 ;
        RECT 793.950 171.600 796.050 172.050 ;
        RECT 796.950 171.600 799.050 172.050 ;
        RECT 811.950 171.600 814.050 172.050 ;
        RECT 820.950 171.600 823.050 172.050 ;
        RECT 793.950 170.400 823.050 171.600 ;
        RECT 793.950 169.950 796.050 170.400 ;
        RECT 796.950 169.950 799.050 170.400 ;
        RECT 811.950 169.950 814.050 170.400 ;
        RECT 820.950 169.950 823.050 170.400 ;
        RECT 823.950 171.600 826.050 172.050 ;
        RECT 829.950 171.600 832.050 172.050 ;
        RECT 823.950 170.400 832.050 171.600 ;
        RECT 823.950 169.950 826.050 170.400 ;
        RECT 829.950 169.950 832.050 170.400 ;
        RECT 856.950 171.600 859.050 172.050 ;
        RECT 856.950 170.400 867.600 171.600 ;
        RECT 856.950 169.950 859.050 170.400 ;
        RECT 715.950 168.600 718.050 169.050 ;
        RECT 721.950 168.600 724.050 169.050 ;
        RECT 715.950 167.400 724.050 168.600 ;
        RECT 715.950 166.950 718.050 167.400 ;
        RECT 721.950 166.950 724.050 167.400 ;
        RECT 790.950 168.600 793.050 169.050 ;
        RECT 805.950 168.600 808.050 169.050 ;
        RECT 826.950 168.600 829.050 169.050 ;
        RECT 790.950 167.400 808.050 168.600 ;
        RECT 790.950 166.950 793.050 167.400 ;
        RECT 805.950 166.950 808.050 167.400 ;
        RECT 809.400 167.400 829.050 168.600 ;
        RECT 809.400 166.050 810.600 167.400 ;
        RECT 826.950 166.950 829.050 167.400 ;
        RECT 841.950 168.600 844.050 169.050 ;
        RECT 841.950 167.400 861.600 168.600 ;
        RECT 841.950 166.950 844.050 167.400 ;
        RECT 10.950 164.400 27.600 165.600 ;
        RECT 28.950 165.600 31.050 166.050 ;
        RECT 40.950 165.600 43.050 166.050 ;
        RECT 55.950 165.600 58.050 166.050 ;
        RECT 73.950 165.600 76.050 166.050 ;
        RECT 28.950 164.400 43.050 165.600 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 22.950 163.950 25.050 164.400 ;
        RECT 28.950 163.950 31.050 164.400 ;
        RECT 40.950 163.950 43.050 164.400 ;
        RECT 44.400 164.400 76.050 165.600 ;
        RECT 10.950 162.600 13.050 163.050 ;
        RECT 44.400 162.600 45.600 164.400 ;
        RECT 55.950 163.950 58.050 164.400 ;
        RECT 73.950 163.950 76.050 164.400 ;
        RECT 115.950 165.600 118.050 166.050 ;
        RECT 130.950 165.600 133.050 166.050 ;
        RECT 115.950 164.400 133.050 165.600 ;
        RECT 115.950 163.950 118.050 164.400 ;
        RECT 130.950 163.950 133.050 164.400 ;
        RECT 154.950 163.950 157.050 166.050 ;
        RECT 166.950 165.600 169.050 166.050 ;
        RECT 193.950 165.600 196.050 166.050 ;
        RECT 205.950 165.600 208.050 166.050 ;
        RECT 166.950 164.400 208.050 165.600 ;
        RECT 166.950 163.950 169.050 164.400 ;
        RECT 193.950 163.950 196.050 164.400 ;
        RECT 205.950 163.950 208.050 164.400 ;
        RECT 229.950 165.600 232.050 166.050 ;
        RECT 286.950 165.600 289.050 166.050 ;
        RECT 229.950 164.400 289.050 165.600 ;
        RECT 229.950 163.950 232.050 164.400 ;
        RECT 286.950 163.950 289.050 164.400 ;
        RECT 301.950 163.950 304.050 166.050 ;
        RECT 307.950 165.600 310.050 166.050 ;
        RECT 316.950 165.600 319.050 166.050 ;
        RECT 307.950 164.400 319.050 165.600 ;
        RECT 307.950 163.950 310.050 164.400 ;
        RECT 316.950 163.950 319.050 164.400 ;
        RECT 340.950 165.600 343.050 166.050 ;
        RECT 349.950 165.600 352.050 166.050 ;
        RECT 340.950 164.400 352.050 165.600 ;
        RECT 340.950 163.950 343.050 164.400 ;
        RECT 349.950 163.950 352.050 164.400 ;
        RECT 352.950 165.600 355.050 166.050 ;
        RECT 358.950 165.600 361.050 166.050 ;
        RECT 352.950 164.400 361.050 165.600 ;
        RECT 352.950 163.950 355.050 164.400 ;
        RECT 358.950 163.950 361.050 164.400 ;
        RECT 370.950 165.600 373.050 166.050 ;
        RECT 379.950 165.600 382.050 166.050 ;
        RECT 370.950 164.400 382.050 165.600 ;
        RECT 370.950 163.950 373.050 164.400 ;
        RECT 379.950 163.950 382.050 164.400 ;
        RECT 394.950 165.600 397.050 166.050 ;
        RECT 400.950 165.600 403.050 166.050 ;
        RECT 394.950 164.400 403.050 165.600 ;
        RECT 394.950 163.950 397.050 164.400 ;
        RECT 400.950 163.950 403.050 164.400 ;
        RECT 409.950 165.600 412.050 166.050 ;
        RECT 415.950 165.600 418.050 166.050 ;
        RECT 409.950 164.400 418.050 165.600 ;
        RECT 409.950 163.950 412.050 164.400 ;
        RECT 415.950 163.950 418.050 164.400 ;
        RECT 484.950 163.950 487.050 166.050 ;
        RECT 535.950 163.950 538.050 166.050 ;
        RECT 541.950 165.600 544.050 166.050 ;
        RECT 547.950 165.600 550.050 166.050 ;
        RECT 541.950 164.400 550.050 165.600 ;
        RECT 541.950 163.950 544.050 164.400 ;
        RECT 547.950 163.950 550.050 164.400 ;
        RECT 586.950 165.600 589.050 166.050 ;
        RECT 595.950 165.600 598.050 166.050 ;
        RECT 586.950 164.400 598.050 165.600 ;
        RECT 586.950 163.950 589.050 164.400 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 649.950 163.950 652.050 166.050 ;
        RECT 667.950 165.600 670.050 166.050 ;
        RECT 676.950 165.600 679.050 166.050 ;
        RECT 667.950 164.400 679.050 165.600 ;
        RECT 667.950 163.950 670.050 164.400 ;
        RECT 676.950 163.950 679.050 164.400 ;
        RECT 697.950 163.950 700.050 166.050 ;
        RECT 700.950 165.600 703.050 166.050 ;
        RECT 706.950 165.600 709.050 166.050 ;
        RECT 700.950 164.400 709.050 165.600 ;
        RECT 700.950 163.950 703.050 164.400 ;
        RECT 706.950 163.950 709.050 164.400 ;
        RECT 808.950 163.950 811.050 166.050 ;
        RECT 850.950 165.600 853.050 166.050 ;
        RECT 853.950 165.600 856.050 166.050 ;
        RECT 856.950 165.600 859.050 166.050 ;
        RECT 850.950 164.400 859.050 165.600 ;
        RECT 860.400 165.600 861.600 167.400 ;
        RECT 866.400 166.050 867.600 170.400 ;
        RECT 862.950 165.600 865.050 166.050 ;
        RECT 860.400 164.400 865.050 165.600 ;
        RECT 850.950 163.950 853.050 164.400 ;
        RECT 853.950 163.950 856.050 164.400 ;
        RECT 856.950 163.950 859.050 164.400 ;
        RECT 862.950 163.950 865.050 164.400 ;
        RECT 865.950 163.950 868.050 166.050 ;
        RECT 10.950 161.400 45.600 162.600 ;
        RECT 46.950 162.600 49.050 163.050 ;
        RECT 67.950 162.600 70.050 163.050 ;
        RECT 46.950 161.400 70.050 162.600 ;
        RECT 10.950 160.950 13.050 161.400 ;
        RECT 46.950 160.950 49.050 161.400 ;
        RECT 67.950 160.950 70.050 161.400 ;
        RECT 79.950 162.600 82.050 163.050 ;
        RECT 88.950 162.600 91.050 163.050 ;
        RECT 79.950 161.400 91.050 162.600 ;
        RECT 79.950 160.950 82.050 161.400 ;
        RECT 88.950 160.950 91.050 161.400 ;
        RECT 94.950 162.600 97.050 163.050 ;
        RECT 100.950 162.600 103.050 163.050 ;
        RECT 94.950 161.400 103.050 162.600 ;
        RECT 94.950 160.950 97.050 161.400 ;
        RECT 100.950 160.950 103.050 161.400 ;
        RECT 103.950 162.600 106.050 163.050 ;
        RECT 133.950 162.600 136.050 163.050 ;
        RECT 103.950 161.400 136.050 162.600 ;
        RECT 155.400 162.600 156.600 163.950 ;
        RECT 187.950 162.600 190.050 163.050 ;
        RECT 211.950 162.600 214.050 163.050 ;
        RECT 155.400 161.400 214.050 162.600 ;
        RECT 103.950 160.950 106.050 161.400 ;
        RECT 133.950 160.950 136.050 161.400 ;
        RECT 187.950 160.950 190.050 161.400 ;
        RECT 211.950 160.950 214.050 161.400 ;
        RECT 217.950 162.600 220.050 163.050 ;
        RECT 262.950 162.600 265.050 163.050 ;
        RECT 217.950 161.400 265.050 162.600 ;
        RECT 217.950 160.950 220.050 161.400 ;
        RECT 262.950 160.950 265.050 161.400 ;
        RECT 280.950 162.600 283.050 163.050 ;
        RECT 289.950 162.600 292.050 163.050 ;
        RECT 280.950 161.400 292.050 162.600 ;
        RECT 280.950 160.950 283.050 161.400 ;
        RECT 289.950 160.950 292.050 161.400 ;
        RECT 292.950 162.600 295.050 163.050 ;
        RECT 302.400 162.600 303.600 163.950 ;
        RECT 322.950 162.600 325.050 163.050 ;
        RECT 292.950 161.400 325.050 162.600 ;
        RECT 292.950 160.950 295.050 161.400 ;
        RECT 322.950 160.950 325.050 161.400 ;
        RECT 328.950 162.600 331.050 163.050 ;
        RECT 391.950 162.600 394.050 163.050 ;
        RECT 445.950 162.600 448.050 163.050 ;
        RECT 328.950 161.400 448.050 162.600 ;
        RECT 328.950 160.950 331.050 161.400 ;
        RECT 391.950 160.950 394.050 161.400 ;
        RECT 445.950 160.950 448.050 161.400 ;
        RECT 463.950 162.600 466.050 163.050 ;
        RECT 472.950 162.600 475.050 163.050 ;
        RECT 463.950 161.400 475.050 162.600 ;
        RECT 536.400 162.600 537.600 163.950 ;
        RECT 538.950 162.600 541.050 163.050 ;
        RECT 553.950 162.600 556.050 163.050 ;
        RECT 536.400 161.400 556.050 162.600 ;
        RECT 463.950 160.950 466.050 161.400 ;
        RECT 472.950 160.950 475.050 161.400 ;
        RECT 538.950 160.950 541.050 161.400 ;
        RECT 553.950 160.950 556.050 161.400 ;
        RECT 568.950 162.600 571.050 163.050 ;
        RECT 574.950 162.600 577.050 163.050 ;
        RECT 568.950 161.400 577.050 162.600 ;
        RECT 568.950 160.950 571.050 161.400 ;
        RECT 574.950 160.950 577.050 161.400 ;
        RECT 580.950 162.600 583.050 163.050 ;
        RECT 661.950 162.600 664.050 163.050 ;
        RECT 580.950 161.400 664.050 162.600 ;
        RECT 580.950 160.950 583.050 161.400 ;
        RECT 661.950 160.950 664.050 161.400 ;
        RECT 703.950 162.600 706.050 163.050 ;
        RECT 712.950 162.600 715.050 163.050 ;
        RECT 703.950 161.400 715.050 162.600 ;
        RECT 703.950 160.950 706.050 161.400 ;
        RECT 712.950 160.950 715.050 161.400 ;
        RECT 715.950 162.600 718.050 163.050 ;
        RECT 721.950 162.600 724.050 163.050 ;
        RECT 715.950 161.400 724.050 162.600 ;
        RECT 715.950 160.950 718.050 161.400 ;
        RECT 721.950 160.950 724.050 161.400 ;
        RECT 727.950 162.600 730.050 163.050 ;
        RECT 736.950 162.600 739.050 163.050 ;
        RECT 742.950 162.600 745.050 163.050 ;
        RECT 727.950 161.400 745.050 162.600 ;
        RECT 727.950 160.950 730.050 161.400 ;
        RECT 736.950 160.950 739.050 161.400 ;
        RECT 742.950 160.950 745.050 161.400 ;
        RECT 835.950 162.600 838.050 163.050 ;
        RECT 847.950 162.600 850.050 163.050 ;
        RECT 835.950 161.400 850.050 162.600 ;
        RECT 835.950 160.950 838.050 161.400 ;
        RECT 847.950 160.950 850.050 161.400 ;
        RECT 187.950 159.600 190.050 160.050 ;
        RECT 223.950 159.600 226.050 160.050 ;
        RECT 187.950 158.400 226.050 159.600 ;
        RECT 187.950 157.950 190.050 158.400 ;
        RECT 223.950 157.950 226.050 158.400 ;
        RECT 277.950 159.600 280.050 160.050 ;
        RECT 283.950 159.600 286.050 160.050 ;
        RECT 277.950 158.400 286.050 159.600 ;
        RECT 277.950 157.950 280.050 158.400 ;
        RECT 283.950 157.950 286.050 158.400 ;
        RECT 310.950 159.600 313.050 160.050 ;
        RECT 469.950 159.600 472.050 160.050 ;
        RECT 310.950 158.400 472.050 159.600 ;
        RECT 310.950 157.950 313.050 158.400 ;
        RECT 469.950 157.950 472.050 158.400 ;
        RECT 490.950 159.600 493.050 160.050 ;
        RECT 607.950 159.600 610.050 160.050 ;
        RECT 751.950 159.600 754.050 160.050 ;
        RECT 490.950 158.400 754.050 159.600 ;
        RECT 490.950 157.950 493.050 158.400 ;
        RECT 607.950 157.950 610.050 158.400 ;
        RECT 751.950 157.950 754.050 158.400 ;
        RECT 193.950 156.600 196.050 157.050 ;
        RECT 202.950 156.600 205.050 157.050 ;
        RECT 193.950 155.400 205.050 156.600 ;
        RECT 193.950 154.950 196.050 155.400 ;
        RECT 202.950 154.950 205.050 155.400 ;
        RECT 361.950 156.600 364.050 157.050 ;
        RECT 376.950 156.600 379.050 157.050 ;
        RECT 361.950 155.400 379.050 156.600 ;
        RECT 361.950 154.950 364.050 155.400 ;
        RECT 376.950 154.950 379.050 155.400 ;
        RECT 430.950 156.600 433.050 157.050 ;
        RECT 499.950 156.600 502.050 157.050 ;
        RECT 430.950 155.400 502.050 156.600 ;
        RECT 430.950 154.950 433.050 155.400 ;
        RECT 499.950 154.950 502.050 155.400 ;
        RECT 547.950 156.600 550.050 157.050 ;
        RECT 562.950 156.600 565.050 157.050 ;
        RECT 547.950 155.400 565.050 156.600 ;
        RECT 547.950 154.950 550.050 155.400 ;
        RECT 562.950 154.950 565.050 155.400 ;
        RECT 52.950 153.600 55.050 154.050 ;
        RECT 58.950 153.600 61.050 154.050 ;
        RECT 52.950 152.400 61.050 153.600 ;
        RECT 52.950 151.950 55.050 152.400 ;
        RECT 58.950 151.950 61.050 152.400 ;
        RECT 61.950 153.600 64.050 154.050 ;
        RECT 94.950 153.600 97.050 154.050 ;
        RECT 100.950 153.600 103.050 154.050 ;
        RECT 61.950 152.400 103.050 153.600 ;
        RECT 61.950 151.950 64.050 152.400 ;
        RECT 94.950 151.950 97.050 152.400 ;
        RECT 100.950 151.950 103.050 152.400 ;
        RECT 514.950 153.600 517.050 154.050 ;
        RECT 586.950 153.600 589.050 154.050 ;
        RECT 514.950 152.400 589.050 153.600 ;
        RECT 514.950 151.950 517.050 152.400 ;
        RECT 586.950 151.950 589.050 152.400 ;
        RECT 271.950 150.600 274.050 151.050 ;
        RECT 526.950 150.600 529.050 151.050 ;
        RECT 271.950 149.400 529.050 150.600 ;
        RECT 271.950 148.950 274.050 149.400 ;
        RECT 526.950 148.950 529.050 149.400 ;
        RECT 436.950 147.600 439.050 148.050 ;
        RECT 523.950 147.600 526.050 148.050 ;
        RECT 553.950 147.600 556.050 148.050 ;
        RECT 436.950 146.400 556.050 147.600 ;
        RECT 436.950 145.950 439.050 146.400 ;
        RECT 523.950 145.950 526.050 146.400 ;
        RECT 553.950 145.950 556.050 146.400 ;
        RECT 70.950 144.600 73.050 145.050 ;
        RECT 76.950 144.600 79.050 145.050 ;
        RECT 751.950 144.600 754.050 145.050 ;
        RECT 757.950 144.600 760.050 145.050 ;
        RECT 70.950 143.400 79.050 144.600 ;
        RECT 70.950 142.950 73.050 143.400 ;
        RECT 76.950 142.950 79.050 143.400 ;
        RECT 527.400 143.400 760.050 144.600 ;
        RECT 445.950 141.600 448.050 142.050 ;
        RECT 527.400 141.600 528.600 143.400 ;
        RECT 751.950 142.950 754.050 143.400 ;
        RECT 757.950 142.950 760.050 143.400 ;
        RECT 445.950 140.400 528.600 141.600 ;
        RECT 445.950 139.950 448.050 140.400 ;
        RECT 334.950 138.600 337.050 139.050 ;
        RECT 343.950 138.600 346.050 139.050 ;
        RECT 334.950 137.400 346.050 138.600 ;
        RECT 334.950 136.950 337.050 137.400 ;
        RECT 343.950 136.950 346.050 137.400 ;
        RECT 487.950 138.600 490.050 139.050 ;
        RECT 529.950 138.600 532.050 139.050 ;
        RECT 487.950 137.400 532.050 138.600 ;
        RECT 487.950 136.950 490.050 137.400 ;
        RECT 529.950 136.950 532.050 137.400 ;
        RECT 547.950 138.600 550.050 139.050 ;
        RECT 631.950 138.600 634.050 139.050 ;
        RECT 547.950 137.400 634.050 138.600 ;
        RECT 547.950 136.950 550.050 137.400 ;
        RECT 631.950 136.950 634.050 137.400 ;
        RECT 823.950 138.600 826.050 139.050 ;
        RECT 829.950 138.600 832.050 139.050 ;
        RECT 823.950 137.400 832.050 138.600 ;
        RECT 823.950 136.950 826.050 137.400 ;
        RECT 829.950 136.950 832.050 137.400 ;
        RECT 85.950 135.600 88.050 136.050 ;
        RECT 91.950 135.600 94.050 136.050 ;
        RECT 109.950 135.600 112.050 136.050 ;
        RECT 85.950 134.400 112.050 135.600 ;
        RECT 85.950 133.950 88.050 134.400 ;
        RECT 91.950 133.950 94.050 134.400 ;
        RECT 109.950 133.950 112.050 134.400 ;
        RECT 319.950 135.600 322.050 136.050 ;
        RECT 331.950 135.600 334.050 136.050 ;
        RECT 319.950 134.400 334.050 135.600 ;
        RECT 319.950 133.950 322.050 134.400 ;
        RECT 331.950 133.950 334.050 134.400 ;
        RECT 343.950 135.600 346.050 136.050 ;
        RECT 382.950 135.600 385.050 136.050 ;
        RECT 343.950 134.400 385.050 135.600 ;
        RECT 343.950 133.950 346.050 134.400 ;
        RECT 382.950 133.950 385.050 134.400 ;
        RECT 571.950 135.600 574.050 136.050 ;
        RECT 580.950 135.600 583.050 136.050 ;
        RECT 598.950 135.600 601.050 136.050 ;
        RECT 634.950 135.600 637.050 136.050 ;
        RECT 571.950 134.400 583.050 135.600 ;
        RECT 571.950 133.950 574.050 134.400 ;
        RECT 580.950 133.950 583.050 134.400 ;
        RECT 584.400 134.400 637.050 135.600 ;
        RECT 19.950 132.600 22.050 133.050 ;
        RECT 25.950 132.600 28.050 133.050 ;
        RECT 19.950 131.400 28.050 132.600 ;
        RECT 19.950 130.950 22.050 131.400 ;
        RECT 25.950 130.950 28.050 131.400 ;
        RECT 130.950 132.600 133.050 133.050 ;
        RECT 181.950 132.600 184.050 133.050 ;
        RECT 130.950 131.400 184.050 132.600 ;
        RECT 130.950 130.950 133.050 131.400 ;
        RECT 181.950 130.950 184.050 131.400 ;
        RECT 199.950 132.600 202.050 133.050 ;
        RECT 214.950 132.600 217.050 133.050 ;
        RECT 277.950 132.600 280.050 133.050 ;
        RECT 340.950 132.600 343.050 133.050 ;
        RECT 199.950 131.400 204.600 132.600 ;
        RECT 199.950 130.950 202.050 131.400 ;
        RECT 34.950 129.600 37.050 130.050 ;
        RECT 14.400 128.400 37.050 129.600 ;
        RECT 14.400 127.050 15.600 128.400 ;
        RECT 34.950 127.950 37.050 128.400 ;
        RECT 64.950 129.600 67.050 130.050 ;
        RECT 82.950 129.600 85.050 130.050 ;
        RECT 64.950 128.400 85.050 129.600 ;
        RECT 64.950 127.950 67.050 128.400 ;
        RECT 82.950 127.950 85.050 128.400 ;
        RECT 100.950 129.600 103.050 130.050 ;
        RECT 106.950 129.600 109.050 130.050 ;
        RECT 118.950 129.600 121.050 130.050 ;
        RECT 169.950 129.600 172.050 130.050 ;
        RECT 100.950 128.400 121.050 129.600 ;
        RECT 100.950 127.950 103.050 128.400 ;
        RECT 106.950 127.950 109.050 128.400 ;
        RECT 118.950 127.950 121.050 128.400 ;
        RECT 137.400 128.400 172.050 129.600 ;
        RECT 203.400 129.600 204.600 131.400 ;
        RECT 214.950 131.400 280.050 132.600 ;
        RECT 214.950 130.950 217.050 131.400 ;
        RECT 277.950 130.950 280.050 131.400 ;
        RECT 302.400 131.400 343.050 132.600 ;
        RECT 205.950 129.600 208.050 130.050 ;
        RECT 203.400 128.400 208.050 129.600 ;
        RECT 137.400 127.050 138.600 128.400 ;
        RECT 169.950 127.950 172.050 128.400 ;
        RECT 205.950 127.950 208.050 128.400 ;
        RECT 211.950 129.600 214.050 130.050 ;
        RECT 217.950 129.600 220.050 130.050 ;
        RECT 211.950 128.400 220.050 129.600 ;
        RECT 211.950 127.950 214.050 128.400 ;
        RECT 217.950 127.950 220.050 128.400 ;
        RECT 220.950 129.600 223.050 130.050 ;
        RECT 232.950 129.600 235.050 130.050 ;
        RECT 220.950 128.400 235.050 129.600 ;
        RECT 220.950 127.950 223.050 128.400 ;
        RECT 232.950 127.950 235.050 128.400 ;
        RECT 244.950 129.600 247.050 130.050 ;
        RECT 256.950 129.600 259.050 130.050 ;
        RECT 244.950 128.400 259.050 129.600 ;
        RECT 244.950 127.950 247.050 128.400 ;
        RECT 256.950 127.950 259.050 128.400 ;
        RECT 283.950 129.600 286.050 130.050 ;
        RECT 302.400 129.600 303.600 131.400 ;
        RECT 340.950 130.950 343.050 131.400 ;
        RECT 439.950 132.600 442.050 133.050 ;
        RECT 466.950 132.600 469.050 133.050 ;
        RECT 584.400 132.600 585.600 134.400 ;
        RECT 598.950 133.950 601.050 134.400 ;
        RECT 634.950 133.950 637.050 134.400 ;
        RECT 754.950 135.600 757.050 136.050 ;
        RECT 769.950 135.600 772.050 136.050 ;
        RECT 754.950 134.400 772.050 135.600 ;
        RECT 754.950 133.950 757.050 134.400 ;
        RECT 769.950 133.950 772.050 134.400 ;
        RECT 811.950 135.600 814.050 136.050 ;
        RECT 841.950 135.600 844.050 136.050 ;
        RECT 811.950 134.400 844.050 135.600 ;
        RECT 811.950 133.950 814.050 134.400 ;
        RECT 841.950 133.950 844.050 134.400 ;
        RECT 439.950 131.400 585.600 132.600 ;
        RECT 613.950 132.600 616.050 133.050 ;
        RECT 619.950 132.600 622.050 133.050 ;
        RECT 613.950 131.400 622.050 132.600 ;
        RECT 439.950 130.950 442.050 131.400 ;
        RECT 466.950 130.950 469.050 131.400 ;
        RECT 613.950 130.950 616.050 131.400 ;
        RECT 619.950 130.950 622.050 131.400 ;
        RECT 688.950 132.600 691.050 133.050 ;
        RECT 718.950 132.600 721.050 133.050 ;
        RECT 688.950 131.400 721.050 132.600 ;
        RECT 688.950 130.950 691.050 131.400 ;
        RECT 718.950 130.950 721.050 131.400 ;
        RECT 730.950 132.600 733.050 133.050 ;
        RECT 739.950 132.600 742.050 133.050 ;
        RECT 730.950 131.400 742.050 132.600 ;
        RECT 730.950 130.950 733.050 131.400 ;
        RECT 739.950 130.950 742.050 131.400 ;
        RECT 784.950 132.600 787.050 133.050 ;
        RECT 796.950 132.600 799.050 133.050 ;
        RECT 784.950 131.400 799.050 132.600 ;
        RECT 784.950 130.950 787.050 131.400 ;
        RECT 796.950 130.950 799.050 131.400 ;
        RECT 829.950 132.600 832.050 133.050 ;
        RECT 853.950 132.600 856.050 133.050 ;
        RECT 862.950 132.600 865.050 133.050 ;
        RECT 829.950 131.400 852.600 132.600 ;
        RECT 829.950 130.950 832.050 131.400 ;
        RECT 283.950 128.400 303.600 129.600 ;
        RECT 304.950 129.600 307.050 130.050 ;
        RECT 307.950 129.600 310.050 130.050 ;
        RECT 319.950 129.600 322.050 130.050 ;
        RECT 304.950 128.400 322.050 129.600 ;
        RECT 283.950 127.950 286.050 128.400 ;
        RECT 304.950 127.950 307.050 128.400 ;
        RECT 307.950 127.950 310.050 128.400 ;
        RECT 319.950 127.950 322.050 128.400 ;
        RECT 376.950 129.600 379.050 130.050 ;
        RECT 394.950 129.600 397.050 130.050 ;
        RECT 376.950 128.400 397.050 129.600 ;
        RECT 376.950 127.950 379.050 128.400 ;
        RECT 394.950 127.950 397.050 128.400 ;
        RECT 427.950 129.600 430.050 130.050 ;
        RECT 433.950 129.600 436.050 130.050 ;
        RECT 427.950 128.400 436.050 129.600 ;
        RECT 427.950 127.950 430.050 128.400 ;
        RECT 433.950 127.950 436.050 128.400 ;
        RECT 493.950 129.600 496.050 130.050 ;
        RECT 520.950 129.600 523.050 130.050 ;
        RECT 493.950 128.400 523.050 129.600 ;
        RECT 493.950 127.950 496.050 128.400 ;
        RECT 520.950 127.950 523.050 128.400 ;
        RECT 556.950 129.600 559.050 130.050 ;
        RECT 583.950 129.600 586.050 130.050 ;
        RECT 556.950 128.400 586.050 129.600 ;
        RECT 556.950 127.950 559.050 128.400 ;
        RECT 583.950 127.950 586.050 128.400 ;
        RECT 604.950 129.600 607.050 130.050 ;
        RECT 616.950 129.600 619.050 130.050 ;
        RECT 622.950 129.600 625.050 130.050 ;
        RECT 604.950 128.400 625.050 129.600 ;
        RECT 604.950 127.950 607.050 128.400 ;
        RECT 616.950 127.950 619.050 128.400 ;
        RECT 622.950 127.950 625.050 128.400 ;
        RECT 691.950 129.600 694.050 130.050 ;
        RECT 697.950 129.600 700.050 130.050 ;
        RECT 715.950 129.600 718.050 130.050 ;
        RECT 691.950 128.400 718.050 129.600 ;
        RECT 691.950 127.950 694.050 128.400 ;
        RECT 697.950 127.950 700.050 128.400 ;
        RECT 715.950 127.950 718.050 128.400 ;
        RECT 733.950 129.600 736.050 130.050 ;
        RECT 841.950 129.600 844.050 130.050 ;
        RECT 847.950 129.600 850.050 130.050 ;
        RECT 733.950 128.400 850.050 129.600 ;
        RECT 851.400 129.600 852.600 131.400 ;
        RECT 853.950 131.400 865.050 132.600 ;
        RECT 853.950 130.950 856.050 131.400 ;
        RECT 862.950 130.950 865.050 131.400 ;
        RECT 851.400 128.400 858.600 129.600 ;
        RECT 733.950 127.950 736.050 128.400 ;
        RECT 841.950 127.950 844.050 128.400 ;
        RECT 847.950 127.950 850.050 128.400 ;
        RECT 13.950 124.950 16.050 127.050 ;
        RECT 19.950 126.600 22.050 127.050 ;
        RECT 28.950 126.600 31.050 127.050 ;
        RECT 19.950 125.400 31.050 126.600 ;
        RECT 19.950 124.950 22.050 125.400 ;
        RECT 28.950 124.950 31.050 125.400 ;
        RECT 55.950 126.600 58.050 127.050 ;
        RECT 76.950 126.600 79.050 127.050 ;
        RECT 55.950 125.400 79.050 126.600 ;
        RECT 55.950 124.950 58.050 125.400 ;
        RECT 76.950 124.950 79.050 125.400 ;
        RECT 82.950 126.600 85.050 127.050 ;
        RECT 127.950 126.600 130.050 127.050 ;
        RECT 82.950 125.400 130.050 126.600 ;
        RECT 82.950 124.950 85.050 125.400 ;
        RECT 127.950 124.950 130.050 125.400 ;
        RECT 136.950 124.950 139.050 127.050 ;
        RECT 142.950 126.600 145.050 127.050 ;
        RECT 151.950 126.600 154.050 127.050 ;
        RECT 142.950 125.400 154.050 126.600 ;
        RECT 142.950 124.950 145.050 125.400 ;
        RECT 151.950 124.950 154.050 125.400 ;
        RECT 160.950 126.600 163.050 127.050 ;
        RECT 169.950 126.600 172.050 127.050 ;
        RECT 160.950 125.400 172.050 126.600 ;
        RECT 160.950 124.950 163.050 125.400 ;
        RECT 169.950 124.950 172.050 125.400 ;
        RECT 178.950 124.950 181.050 127.050 ;
        RECT 202.950 126.600 205.050 127.050 ;
        RECT 235.950 126.600 238.050 127.050 ;
        RECT 202.950 125.400 238.050 126.600 ;
        RECT 202.950 124.950 205.050 125.400 ;
        RECT 235.950 124.950 238.050 125.400 ;
        RECT 265.950 126.600 268.050 127.050 ;
        RECT 274.950 126.600 277.050 127.050 ;
        RECT 286.950 126.600 289.050 127.050 ;
        RECT 295.950 126.600 298.050 127.050 ;
        RECT 265.950 125.400 298.050 126.600 ;
        RECT 265.950 124.950 268.050 125.400 ;
        RECT 274.950 124.950 277.050 125.400 ;
        RECT 286.950 124.950 289.050 125.400 ;
        RECT 295.950 124.950 298.050 125.400 ;
        RECT 385.950 126.600 388.050 127.050 ;
        RECT 415.950 126.600 418.050 127.050 ;
        RECT 385.950 125.400 418.050 126.600 ;
        RECT 385.950 124.950 388.050 125.400 ;
        RECT 415.950 124.950 418.050 125.400 ;
        RECT 451.950 126.600 454.050 127.050 ;
        RECT 457.950 126.600 460.050 127.050 ;
        RECT 451.950 125.400 460.050 126.600 ;
        RECT 451.950 124.950 454.050 125.400 ;
        RECT 457.950 124.950 460.050 125.400 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 475.950 126.600 478.050 127.050 ;
        RECT 469.950 125.400 478.050 126.600 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 550.950 126.600 553.050 127.050 ;
        RECT 559.950 126.600 562.050 127.050 ;
        RECT 550.950 125.400 562.050 126.600 ;
        RECT 550.950 124.950 553.050 125.400 ;
        RECT 559.950 124.950 562.050 125.400 ;
        RECT 568.950 126.600 571.050 127.050 ;
        RECT 574.950 126.600 577.050 127.050 ;
        RECT 568.950 125.400 577.050 126.600 ;
        RECT 568.950 124.950 571.050 125.400 ;
        RECT 574.950 124.950 577.050 125.400 ;
        RECT 586.950 126.600 589.050 127.050 ;
        RECT 601.950 126.600 604.050 127.050 ;
        RECT 586.950 125.400 604.050 126.600 ;
        RECT 586.950 124.950 589.050 125.400 ;
        RECT 601.950 124.950 604.050 125.400 ;
        RECT 625.950 126.600 628.050 127.050 ;
        RECT 646.950 126.600 649.050 127.050 ;
        RECT 625.950 125.400 649.050 126.600 ;
        RECT 625.950 124.950 628.050 125.400 ;
        RECT 646.950 124.950 649.050 125.400 ;
        RECT 658.950 126.600 661.050 127.050 ;
        RECT 664.950 126.600 667.050 127.050 ;
        RECT 658.950 125.400 667.050 126.600 ;
        RECT 658.950 124.950 661.050 125.400 ;
        RECT 664.950 124.950 667.050 125.400 ;
        RECT 676.950 126.600 679.050 127.050 ;
        RECT 685.950 126.600 688.050 127.050 ;
        RECT 676.950 125.400 688.050 126.600 ;
        RECT 676.950 124.950 679.050 125.400 ;
        RECT 685.950 124.950 688.050 125.400 ;
        RECT 703.950 126.600 706.050 127.050 ;
        RECT 709.950 126.600 712.050 127.050 ;
        RECT 733.950 126.600 736.050 127.050 ;
        RECT 739.950 126.600 742.050 127.050 ;
        RECT 703.950 125.400 712.050 126.600 ;
        RECT 703.950 124.950 706.050 125.400 ;
        RECT 709.950 124.950 712.050 125.400 ;
        RECT 713.400 125.400 742.050 126.600 ;
        RECT 37.950 123.600 40.050 124.050 ;
        RECT 46.950 123.600 49.050 124.050 ;
        RECT 37.950 122.400 49.050 123.600 ;
        RECT 37.950 121.950 40.050 122.400 ;
        RECT 46.950 121.950 49.050 122.400 ;
        RECT 73.950 123.600 76.050 124.050 ;
        RECT 91.950 123.600 94.050 124.050 ;
        RECT 73.950 122.400 94.050 123.600 ;
        RECT 73.950 121.950 76.050 122.400 ;
        RECT 91.950 121.950 94.050 122.400 ;
        RECT 121.950 123.600 124.050 124.050 ;
        RECT 133.950 123.600 136.050 124.050 ;
        RECT 121.950 122.400 136.050 123.600 ;
        RECT 121.950 121.950 124.050 122.400 ;
        RECT 133.950 121.950 136.050 122.400 ;
        RECT 151.950 123.600 154.050 124.050 ;
        RECT 179.400 123.600 180.600 124.950 ;
        RECT 151.950 122.400 180.600 123.600 ;
        RECT 181.950 123.600 184.050 124.050 ;
        RECT 193.950 123.600 196.050 124.050 ;
        RECT 181.950 122.400 196.050 123.600 ;
        RECT 151.950 121.950 154.050 122.400 ;
        RECT 181.950 121.950 184.050 122.400 ;
        RECT 193.950 121.950 196.050 122.400 ;
        RECT 259.950 123.600 262.050 124.050 ;
        RECT 271.950 123.600 274.050 124.050 ;
        RECT 259.950 122.400 274.050 123.600 ;
        RECT 259.950 121.950 262.050 122.400 ;
        RECT 271.950 121.950 274.050 122.400 ;
        RECT 280.950 123.600 283.050 124.050 ;
        RECT 301.950 123.600 304.050 124.050 ;
        RECT 310.950 123.600 313.050 124.050 ;
        RECT 280.950 122.400 313.050 123.600 ;
        RECT 280.950 121.950 283.050 122.400 ;
        RECT 301.950 121.950 304.050 122.400 ;
        RECT 310.950 121.950 313.050 122.400 ;
        RECT 322.950 123.600 325.050 124.050 ;
        RECT 364.950 123.600 367.050 124.050 ;
        RECT 322.950 122.400 367.050 123.600 ;
        RECT 322.950 121.950 325.050 122.400 ;
        RECT 364.950 121.950 367.050 122.400 ;
        RECT 400.950 123.600 403.050 124.050 ;
        RECT 409.950 123.600 412.050 124.050 ;
        RECT 400.950 122.400 412.050 123.600 ;
        RECT 400.950 121.950 403.050 122.400 ;
        RECT 409.950 121.950 412.050 122.400 ;
        RECT 508.950 123.600 511.050 124.050 ;
        RECT 526.950 123.600 529.050 124.050 ;
        RECT 583.950 123.600 586.050 124.050 ;
        RECT 508.950 122.400 516.600 123.600 ;
        RECT 508.950 121.950 511.050 122.400 ;
        RECT 16.950 120.600 19.050 121.050 ;
        RECT 31.950 120.600 34.050 121.050 ;
        RECT 16.950 119.400 34.050 120.600 ;
        RECT 16.950 118.950 19.050 119.400 ;
        RECT 31.950 118.950 34.050 119.400 ;
        RECT 34.950 120.600 37.050 121.050 ;
        RECT 40.950 120.600 43.050 121.050 ;
        RECT 34.950 119.400 43.050 120.600 ;
        RECT 34.950 118.950 37.050 119.400 ;
        RECT 40.950 118.950 43.050 119.400 ;
        RECT 49.950 120.600 52.050 121.050 ;
        RECT 55.950 120.600 58.050 121.050 ;
        RECT 49.950 119.400 58.050 120.600 ;
        RECT 49.950 118.950 52.050 119.400 ;
        RECT 55.950 118.950 58.050 119.400 ;
        RECT 58.950 120.600 61.050 121.050 ;
        RECT 79.950 120.600 82.050 121.050 ;
        RECT 139.950 120.600 142.050 121.050 ;
        RECT 58.950 119.400 142.050 120.600 ;
        RECT 58.950 118.950 61.050 119.400 ;
        RECT 79.950 118.950 82.050 119.400 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 163.950 120.600 166.050 121.050 ;
        RECT 184.950 120.600 187.050 121.050 ;
        RECT 163.950 119.400 187.050 120.600 ;
        RECT 163.950 118.950 166.050 119.400 ;
        RECT 184.950 118.950 187.050 119.400 ;
        RECT 217.950 120.600 220.050 121.050 ;
        RECT 241.950 120.600 244.050 121.050 ;
        RECT 217.950 119.400 244.050 120.600 ;
        RECT 217.950 118.950 220.050 119.400 ;
        RECT 241.950 118.950 244.050 119.400 ;
        RECT 265.950 120.600 268.050 121.050 ;
        RECT 316.950 120.600 319.050 121.050 ;
        RECT 346.950 120.600 349.050 121.050 ;
        RECT 265.950 119.400 349.050 120.600 ;
        RECT 265.950 118.950 268.050 119.400 ;
        RECT 316.950 118.950 319.050 119.400 ;
        RECT 346.950 118.950 349.050 119.400 ;
        RECT 466.950 120.600 469.050 121.050 ;
        RECT 472.950 120.600 475.050 121.050 ;
        RECT 466.950 119.400 475.050 120.600 ;
        RECT 466.950 118.950 469.050 119.400 ;
        RECT 472.950 118.950 475.050 119.400 ;
        RECT 499.950 120.600 502.050 121.050 ;
        RECT 511.950 120.600 514.050 121.050 ;
        RECT 499.950 119.400 514.050 120.600 ;
        RECT 515.400 120.600 516.600 122.400 ;
        RECT 526.950 122.400 586.050 123.600 ;
        RECT 526.950 121.950 529.050 122.400 ;
        RECT 583.950 121.950 586.050 122.400 ;
        RECT 628.950 123.600 631.050 124.050 ;
        RECT 637.950 123.600 640.050 124.050 ;
        RECT 628.950 122.400 640.050 123.600 ;
        RECT 628.950 121.950 631.050 122.400 ;
        RECT 637.950 121.950 640.050 122.400 ;
        RECT 679.950 123.600 682.050 124.050 ;
        RECT 713.400 123.600 714.600 125.400 ;
        RECT 733.950 124.950 736.050 125.400 ;
        RECT 739.950 124.950 742.050 125.400 ;
        RECT 745.950 126.600 748.050 127.050 ;
        RECT 760.950 126.600 763.050 127.050 ;
        RECT 745.950 125.400 763.050 126.600 ;
        RECT 745.950 124.950 748.050 125.400 ;
        RECT 679.950 122.400 714.600 123.600 ;
        RECT 742.950 123.600 745.050 124.050 ;
        RECT 754.950 123.600 757.050 124.050 ;
        RECT 742.950 122.400 757.050 123.600 ;
        RECT 679.950 121.950 682.050 122.400 ;
        RECT 742.950 121.950 745.050 122.400 ;
        RECT 754.950 121.950 757.050 122.400 ;
        RECT 529.950 120.600 532.050 121.050 ;
        RECT 515.400 119.400 532.050 120.600 ;
        RECT 499.950 118.950 502.050 119.400 ;
        RECT 511.950 118.950 514.050 119.400 ;
        RECT 529.950 118.950 532.050 119.400 ;
        RECT 532.950 120.600 535.050 121.050 ;
        RECT 550.950 120.600 553.050 121.050 ;
        RECT 562.950 120.600 565.050 121.050 ;
        RECT 532.950 119.400 565.050 120.600 ;
        RECT 532.950 118.950 535.050 119.400 ;
        RECT 550.950 118.950 553.050 119.400 ;
        RECT 562.950 118.950 565.050 119.400 ;
        RECT 568.950 120.600 571.050 121.050 ;
        RECT 598.950 120.600 601.050 121.050 ;
        RECT 607.950 120.600 610.050 121.050 ;
        RECT 568.950 119.400 610.050 120.600 ;
        RECT 568.950 118.950 571.050 119.400 ;
        RECT 598.950 118.950 601.050 119.400 ;
        RECT 607.950 118.950 610.050 119.400 ;
        RECT 619.950 120.600 622.050 121.050 ;
        RECT 643.950 120.600 646.050 121.050 ;
        RECT 661.950 120.600 664.050 121.050 ;
        RECT 619.950 119.400 664.050 120.600 ;
        RECT 619.950 118.950 622.050 119.400 ;
        RECT 643.950 118.950 646.050 119.400 ;
        RECT 661.950 118.950 664.050 119.400 ;
        RECT 682.950 120.600 685.050 121.050 ;
        RECT 709.950 120.600 712.050 121.050 ;
        RECT 682.950 119.400 712.050 120.600 ;
        RECT 682.950 118.950 685.050 119.400 ;
        RECT 709.950 118.950 712.050 119.400 ;
        RECT 715.950 120.600 718.050 121.050 ;
        RECT 721.950 120.600 724.050 121.050 ;
        RECT 758.400 120.600 759.600 125.400 ;
        RECT 760.950 124.950 763.050 125.400 ;
        RECT 796.950 126.600 799.050 127.050 ;
        RECT 805.950 126.600 808.050 127.050 ;
        RECT 823.950 126.600 826.050 127.050 ;
        RECT 796.950 125.400 808.050 126.600 ;
        RECT 796.950 124.950 799.050 125.400 ;
        RECT 805.950 124.950 808.050 125.400 ;
        RECT 809.400 125.400 826.050 126.600 ;
        RECT 787.950 123.600 790.050 124.050 ;
        RECT 796.950 123.600 799.050 124.050 ;
        RECT 787.950 122.400 799.050 123.600 ;
        RECT 787.950 121.950 790.050 122.400 ;
        RECT 796.950 121.950 799.050 122.400 ;
        RECT 809.400 121.050 810.600 125.400 ;
        RECT 823.950 124.950 826.050 125.400 ;
        RECT 835.950 126.600 838.050 127.050 ;
        RECT 853.950 126.600 856.050 127.050 ;
        RECT 835.950 125.400 856.050 126.600 ;
        RECT 835.950 124.950 838.050 125.400 ;
        RECT 853.950 124.950 856.050 125.400 ;
        RECT 811.950 123.600 814.050 124.050 ;
        RECT 820.950 123.600 823.050 124.050 ;
        RECT 811.950 122.400 823.050 123.600 ;
        RECT 811.950 121.950 814.050 122.400 ;
        RECT 820.950 121.950 823.050 122.400 ;
        RECT 832.950 123.600 835.050 124.050 ;
        RECT 838.950 123.600 841.050 124.050 ;
        RECT 832.950 122.400 841.050 123.600 ;
        RECT 832.950 121.950 835.050 122.400 ;
        RECT 838.950 121.950 841.050 122.400 ;
        RECT 850.950 123.600 853.050 124.050 ;
        RECT 857.400 123.600 858.600 128.400 ;
        RECT 850.950 122.400 858.600 123.600 ;
        RECT 850.950 121.950 853.050 122.400 ;
        RECT 760.950 120.600 763.050 121.050 ;
        RECT 715.950 119.400 763.050 120.600 ;
        RECT 715.950 118.950 718.050 119.400 ;
        RECT 721.950 118.950 724.050 119.400 ;
        RECT 760.950 118.950 763.050 119.400 ;
        RECT 766.950 120.600 769.050 121.050 ;
        RECT 787.950 120.600 790.050 121.050 ;
        RECT 766.950 119.400 790.050 120.600 ;
        RECT 766.950 118.950 769.050 119.400 ;
        RECT 787.950 118.950 790.050 119.400 ;
        RECT 790.950 120.600 793.050 121.050 ;
        RECT 799.950 120.600 802.050 121.050 ;
        RECT 790.950 119.400 802.050 120.600 ;
        RECT 790.950 118.950 793.050 119.400 ;
        RECT 799.950 118.950 802.050 119.400 ;
        RECT 808.950 118.950 811.050 121.050 ;
        RECT 97.950 117.600 100.050 118.050 ;
        RECT 109.950 117.600 112.050 118.050 ;
        RECT 142.950 117.600 145.050 118.050 ;
        RECT 97.950 116.400 145.050 117.600 ;
        RECT 97.950 115.950 100.050 116.400 ;
        RECT 109.950 115.950 112.050 116.400 ;
        RECT 142.950 115.950 145.050 116.400 ;
        RECT 262.950 117.600 265.050 118.050 ;
        RECT 298.950 117.600 301.050 118.050 ;
        RECT 262.950 116.400 301.050 117.600 ;
        RECT 262.950 115.950 265.050 116.400 ;
        RECT 298.950 115.950 301.050 116.400 ;
        RECT 403.950 117.600 406.050 118.050 ;
        RECT 421.950 117.600 424.050 118.050 ;
        RECT 490.950 117.600 493.050 118.050 ;
        RECT 403.950 116.400 493.050 117.600 ;
        RECT 403.950 115.950 406.050 116.400 ;
        RECT 421.950 115.950 424.050 116.400 ;
        RECT 490.950 115.950 493.050 116.400 ;
        RECT 514.950 117.600 517.050 118.050 ;
        RECT 610.950 117.600 613.050 118.050 ;
        RECT 514.950 116.400 613.050 117.600 ;
        RECT 514.950 115.950 517.050 116.400 ;
        RECT 610.950 115.950 613.050 116.400 ;
        RECT 727.950 117.600 730.050 118.050 ;
        RECT 736.950 117.600 739.050 118.050 ;
        RECT 766.950 117.600 769.050 118.050 ;
        RECT 727.950 116.400 769.050 117.600 ;
        RECT 727.950 115.950 730.050 116.400 ;
        RECT 736.950 115.950 739.050 116.400 ;
        RECT 766.950 115.950 769.050 116.400 ;
        RECT 793.950 117.600 796.050 118.050 ;
        RECT 823.950 117.600 826.050 118.050 ;
        RECT 793.950 116.400 826.050 117.600 ;
        RECT 793.950 115.950 796.050 116.400 ;
        RECT 823.950 115.950 826.050 116.400 ;
        RECT 100.950 114.600 103.050 115.050 ;
        RECT 115.950 114.600 118.050 115.050 ;
        RECT 154.950 114.600 157.050 115.050 ;
        RECT 100.950 113.400 157.050 114.600 ;
        RECT 100.950 112.950 103.050 113.400 ;
        RECT 115.950 112.950 118.050 113.400 ;
        RECT 154.950 112.950 157.050 113.400 ;
        RECT 295.950 114.600 298.050 115.050 ;
        RECT 313.950 114.600 316.050 115.050 ;
        RECT 295.950 113.400 316.050 114.600 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 313.950 112.950 316.050 113.400 ;
        RECT 364.950 114.600 367.050 115.050 ;
        RECT 397.950 114.600 400.050 115.050 ;
        RECT 364.950 113.400 400.050 114.600 ;
        RECT 364.950 112.950 367.050 113.400 ;
        RECT 397.950 112.950 400.050 113.400 ;
        RECT 577.950 114.600 580.050 115.050 ;
        RECT 649.950 114.600 652.050 115.050 ;
        RECT 715.950 114.600 718.050 115.050 ;
        RECT 577.950 113.400 718.050 114.600 ;
        RECT 577.950 112.950 580.050 113.400 ;
        RECT 649.950 112.950 652.050 113.400 ;
        RECT 715.950 112.950 718.050 113.400 ;
        RECT 199.950 111.600 202.050 112.050 ;
        RECT 292.950 111.600 295.050 112.050 ;
        RECT 199.950 110.400 295.050 111.600 ;
        RECT 199.950 109.950 202.050 110.400 ;
        RECT 292.950 109.950 295.050 110.400 ;
        RECT 298.950 111.600 301.050 112.050 ;
        RECT 676.950 111.600 679.050 112.050 ;
        RECT 700.950 111.600 703.050 112.050 ;
        RECT 298.950 110.400 703.050 111.600 ;
        RECT 298.950 109.950 301.050 110.400 ;
        RECT 676.950 109.950 679.050 110.400 ;
        RECT 700.950 109.950 703.050 110.400 ;
        RECT 787.950 111.600 790.050 112.050 ;
        RECT 814.950 111.600 817.050 112.050 ;
        RECT 820.950 111.600 823.050 112.050 ;
        RECT 847.950 111.600 850.050 112.050 ;
        RECT 787.950 110.400 850.050 111.600 ;
        RECT 787.950 109.950 790.050 110.400 ;
        RECT 814.950 109.950 817.050 110.400 ;
        RECT 820.950 109.950 823.050 110.400 ;
        RECT 847.950 109.950 850.050 110.400 ;
        RECT 19.950 108.600 22.050 109.050 ;
        RECT 52.950 108.600 55.050 109.050 ;
        RECT 19.950 107.400 55.050 108.600 ;
        RECT 19.950 106.950 22.050 107.400 ;
        RECT 52.950 106.950 55.050 107.400 ;
        RECT 799.950 108.600 802.050 109.050 ;
        RECT 850.950 108.600 853.050 109.050 ;
        RECT 799.950 107.400 853.050 108.600 ;
        RECT 799.950 106.950 802.050 107.400 ;
        RECT 850.950 106.950 853.050 107.400 ;
        RECT 217.950 105.600 220.050 106.050 ;
        RECT 271.950 105.600 274.050 106.050 ;
        RECT 217.950 104.400 274.050 105.600 ;
        RECT 217.950 103.950 220.050 104.400 ;
        RECT 271.950 103.950 274.050 104.400 ;
        RECT 277.950 105.600 280.050 106.050 ;
        RECT 355.950 105.600 358.050 106.050 ;
        RECT 277.950 104.400 358.050 105.600 ;
        RECT 277.950 103.950 280.050 104.400 ;
        RECT 355.950 103.950 358.050 104.400 ;
        RECT 580.950 105.600 583.050 106.050 ;
        RECT 604.950 105.600 607.050 106.050 ;
        RECT 664.950 105.600 667.050 106.050 ;
        RECT 580.950 104.400 667.050 105.600 ;
        RECT 580.950 103.950 583.050 104.400 ;
        RECT 604.950 103.950 607.050 104.400 ;
        RECT 664.950 103.950 667.050 104.400 ;
        RECT 727.950 105.600 730.050 106.050 ;
        RECT 802.950 105.600 805.050 106.050 ;
        RECT 805.950 105.600 808.050 106.050 ;
        RECT 727.950 104.400 808.050 105.600 ;
        RECT 727.950 103.950 730.050 104.400 ;
        RECT 802.950 103.950 805.050 104.400 ;
        RECT 805.950 103.950 808.050 104.400 ;
        RECT 814.950 105.600 817.050 106.050 ;
        RECT 838.950 105.600 841.050 106.050 ;
        RECT 814.950 104.400 841.050 105.600 ;
        RECT 814.950 103.950 817.050 104.400 ;
        RECT 838.950 103.950 841.050 104.400 ;
        RECT 139.950 102.600 142.050 103.050 ;
        RECT 166.950 102.600 169.050 103.050 ;
        RECT 181.950 102.600 184.050 103.050 ;
        RECT 229.950 102.600 232.050 103.050 ;
        RECT 139.950 101.400 232.050 102.600 ;
        RECT 139.950 100.950 142.050 101.400 ;
        RECT 166.950 100.950 169.050 101.400 ;
        RECT 181.950 100.950 184.050 101.400 ;
        RECT 229.950 100.950 232.050 101.400 ;
        RECT 271.950 102.600 274.050 103.050 ;
        RECT 325.950 102.600 328.050 103.050 ;
        RECT 271.950 101.400 328.050 102.600 ;
        RECT 271.950 100.950 274.050 101.400 ;
        RECT 325.950 100.950 328.050 101.400 ;
        RECT 532.950 102.600 535.050 103.050 ;
        RECT 652.950 102.600 655.050 103.050 ;
        RECT 688.950 102.600 691.050 103.050 ;
        RECT 532.950 101.400 691.050 102.600 ;
        RECT 532.950 100.950 535.050 101.400 ;
        RECT 652.950 100.950 655.050 101.400 ;
        RECT 688.950 100.950 691.050 101.400 ;
        RECT 706.950 102.600 709.050 103.050 ;
        RECT 724.950 102.600 727.050 103.050 ;
        RECT 748.950 102.600 751.050 103.050 ;
        RECT 706.950 101.400 751.050 102.600 ;
        RECT 706.950 100.950 709.050 101.400 ;
        RECT 724.950 100.950 727.050 101.400 ;
        RECT 748.950 100.950 751.050 101.400 ;
        RECT 772.950 102.600 775.050 103.050 ;
        RECT 781.950 102.600 784.050 103.050 ;
        RECT 772.950 101.400 784.050 102.600 ;
        RECT 772.950 100.950 775.050 101.400 ;
        RECT 781.950 100.950 784.050 101.400 ;
        RECT 790.950 102.600 793.050 103.050 ;
        RECT 832.950 102.600 835.050 103.050 ;
        RECT 790.950 101.400 835.050 102.600 ;
        RECT 790.950 100.950 793.050 101.400 ;
        RECT 832.950 100.950 835.050 101.400 ;
        RECT 22.950 99.600 25.050 100.050 ;
        RECT 40.950 99.600 43.050 100.050 ;
        RECT 22.950 98.400 43.050 99.600 ;
        RECT 22.950 97.950 25.050 98.400 ;
        RECT 40.950 97.950 43.050 98.400 ;
        RECT 67.950 99.600 70.050 100.050 ;
        RECT 97.950 99.600 100.050 100.050 ;
        RECT 67.950 98.400 100.050 99.600 ;
        RECT 67.950 97.950 70.050 98.400 ;
        RECT 97.950 97.950 100.050 98.400 ;
        RECT 145.950 99.600 148.050 100.050 ;
        RECT 148.950 99.600 151.050 100.050 ;
        RECT 208.950 99.600 211.050 100.050 ;
        RECT 226.950 99.600 229.050 100.050 ;
        RECT 145.950 98.400 177.600 99.600 ;
        RECT 145.950 97.950 148.050 98.400 ;
        RECT 148.950 97.950 151.050 98.400 ;
        RECT 16.950 96.600 19.050 97.050 ;
        RECT 79.950 96.600 82.050 97.050 ;
        RECT 16.950 95.400 82.050 96.600 ;
        RECT 16.950 94.950 19.050 95.400 ;
        RECT 44.400 94.050 45.600 95.400 ;
        RECT 79.950 94.950 82.050 95.400 ;
        RECT 163.950 96.600 166.050 97.050 ;
        RECT 172.950 96.600 175.050 97.050 ;
        RECT 163.950 95.400 175.050 96.600 ;
        RECT 176.400 96.600 177.600 98.400 ;
        RECT 208.950 98.400 229.050 99.600 ;
        RECT 208.950 97.950 211.050 98.400 ;
        RECT 226.950 97.950 229.050 98.400 ;
        RECT 247.950 99.600 250.050 100.050 ;
        RECT 289.950 99.600 292.050 100.050 ;
        RECT 247.950 98.400 292.050 99.600 ;
        RECT 247.950 97.950 250.050 98.400 ;
        RECT 289.950 97.950 292.050 98.400 ;
        RECT 298.950 99.600 301.050 100.050 ;
        RECT 313.950 99.600 316.050 100.050 ;
        RECT 298.950 98.400 316.050 99.600 ;
        RECT 298.950 97.950 301.050 98.400 ;
        RECT 313.950 97.950 316.050 98.400 ;
        RECT 316.950 99.600 319.050 100.050 ;
        RECT 337.950 99.600 340.050 100.050 ;
        RECT 316.950 98.400 340.050 99.600 ;
        RECT 316.950 97.950 319.050 98.400 ;
        RECT 337.950 97.950 340.050 98.400 ;
        RECT 409.950 99.600 412.050 100.050 ;
        RECT 430.950 99.600 433.050 100.050 ;
        RECT 463.950 99.600 466.050 100.050 ;
        RECT 478.950 99.600 481.050 100.050 ;
        RECT 505.950 99.600 508.050 100.050 ;
        RECT 409.950 98.400 426.600 99.600 ;
        RECT 409.950 97.950 412.050 98.400 ;
        RECT 202.950 96.600 205.050 97.050 ;
        RECT 176.400 95.400 205.050 96.600 ;
        RECT 163.950 94.950 166.050 95.400 ;
        RECT 172.950 94.950 175.050 95.400 ;
        RECT 185.400 94.050 186.600 95.400 ;
        RECT 202.950 94.950 205.050 95.400 ;
        RECT 226.950 96.600 229.050 97.050 ;
        RECT 250.950 96.600 253.050 97.050 ;
        RECT 226.950 95.400 253.050 96.600 ;
        RECT 226.950 94.950 229.050 95.400 ;
        RECT 250.950 94.950 253.050 95.400 ;
        RECT 256.950 96.600 259.050 97.050 ;
        RECT 259.950 96.600 262.050 97.050 ;
        RECT 298.950 96.600 301.050 97.050 ;
        RECT 256.950 95.400 301.050 96.600 ;
        RECT 256.950 94.950 259.050 95.400 ;
        RECT 259.950 94.950 262.050 95.400 ;
        RECT 298.950 94.950 301.050 95.400 ;
        RECT 310.950 96.600 313.050 97.050 ;
        RECT 334.950 96.600 337.050 97.050 ;
        RECT 340.950 96.600 343.050 97.050 ;
        RECT 310.950 95.400 343.050 96.600 ;
        RECT 310.950 94.950 313.050 95.400 ;
        RECT 334.950 94.950 337.050 95.400 ;
        RECT 340.950 94.950 343.050 95.400 ;
        RECT 425.400 94.050 426.600 98.400 ;
        RECT 430.950 98.400 508.050 99.600 ;
        RECT 430.950 97.950 433.050 98.400 ;
        RECT 463.950 97.950 466.050 98.400 ;
        RECT 478.950 97.950 481.050 98.400 ;
        RECT 505.950 97.950 508.050 98.400 ;
        RECT 511.950 99.600 514.050 100.050 ;
        RECT 544.950 99.600 547.050 100.050 ;
        RECT 511.950 98.400 547.050 99.600 ;
        RECT 511.950 97.950 514.050 98.400 ;
        RECT 544.950 97.950 547.050 98.400 ;
        RECT 571.950 99.600 574.050 100.050 ;
        RECT 589.950 99.600 592.050 100.050 ;
        RECT 571.950 98.400 592.050 99.600 ;
        RECT 571.950 97.950 574.050 98.400 ;
        RECT 589.950 97.950 592.050 98.400 ;
        RECT 625.950 99.600 628.050 100.050 ;
        RECT 631.950 99.600 634.050 100.050 ;
        RECT 625.950 98.400 634.050 99.600 ;
        RECT 625.950 97.950 628.050 98.400 ;
        RECT 631.950 97.950 634.050 98.400 ;
        RECT 655.950 99.600 658.050 100.050 ;
        RECT 670.950 99.600 673.050 100.050 ;
        RECT 655.950 98.400 673.050 99.600 ;
        RECT 655.950 97.950 658.050 98.400 ;
        RECT 670.950 97.950 673.050 98.400 ;
        RECT 697.950 99.600 700.050 100.050 ;
        RECT 718.950 99.600 721.050 100.050 ;
        RECT 697.950 98.400 721.050 99.600 ;
        RECT 697.950 97.950 700.050 98.400 ;
        RECT 718.950 97.950 721.050 98.400 ;
        RECT 730.950 99.600 733.050 100.050 ;
        RECT 736.950 99.600 739.050 100.050 ;
        RECT 742.950 99.600 745.050 100.050 ;
        RECT 730.950 98.400 745.050 99.600 ;
        RECT 730.950 97.950 733.050 98.400 ;
        RECT 736.950 97.950 739.050 98.400 ;
        RECT 742.950 97.950 745.050 98.400 ;
        RECT 763.950 99.600 766.050 100.050 ;
        RECT 769.950 99.600 772.050 100.050 ;
        RECT 763.950 98.400 772.050 99.600 ;
        RECT 763.950 97.950 766.050 98.400 ;
        RECT 769.950 97.950 772.050 98.400 ;
        RECT 772.950 99.600 775.050 100.050 ;
        RECT 817.950 99.600 820.050 100.050 ;
        RECT 844.950 99.600 847.050 100.050 ;
        RECT 772.950 98.400 847.050 99.600 ;
        RECT 772.950 97.950 775.050 98.400 ;
        RECT 817.950 97.950 820.050 98.400 ;
        RECT 844.950 97.950 847.050 98.400 ;
        RECT 454.950 96.600 457.050 97.050 ;
        RECT 469.950 96.600 472.050 97.050 ;
        RECT 454.950 95.400 472.050 96.600 ;
        RECT 454.950 94.950 457.050 95.400 ;
        RECT 469.950 94.950 472.050 95.400 ;
        RECT 472.950 96.600 475.050 97.050 ;
        RECT 526.950 96.600 529.050 97.050 ;
        RECT 472.950 95.400 529.050 96.600 ;
        RECT 472.950 94.950 475.050 95.400 ;
        RECT 526.950 94.950 529.050 95.400 ;
        RECT 532.950 96.600 535.050 97.050 ;
        RECT 538.950 96.600 541.050 97.050 ;
        RECT 532.950 95.400 541.050 96.600 ;
        RECT 532.950 94.950 535.050 95.400 ;
        RECT 538.950 94.950 541.050 95.400 ;
        RECT 541.950 94.950 544.050 97.050 ;
        RECT 550.950 96.600 553.050 97.050 ;
        RECT 565.950 96.600 568.050 97.050 ;
        RECT 550.950 95.400 568.050 96.600 ;
        RECT 550.950 94.950 553.050 95.400 ;
        RECT 565.950 94.950 568.050 95.400 ;
        RECT 586.950 94.950 589.050 97.050 ;
        RECT 610.950 96.600 613.050 97.050 ;
        RECT 610.950 95.400 630.600 96.600 ;
        RECT 610.950 94.950 613.050 95.400 ;
        RECT 7.950 93.600 10.050 94.050 ;
        RECT 13.950 93.600 16.050 94.050 ;
        RECT 37.950 93.600 40.050 94.050 ;
        RECT 7.950 92.400 40.050 93.600 ;
        RECT 7.950 91.950 10.050 92.400 ;
        RECT 13.950 91.950 16.050 92.400 ;
        RECT 37.950 91.950 40.050 92.400 ;
        RECT 43.950 91.950 46.050 94.050 ;
        RECT 46.950 93.600 49.050 94.050 ;
        RECT 58.950 93.600 61.050 94.050 ;
        RECT 46.950 92.400 61.050 93.600 ;
        RECT 46.950 91.950 49.050 92.400 ;
        RECT 58.950 91.950 61.050 92.400 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 88.950 93.600 91.050 94.050 ;
        RECT 100.950 93.600 103.050 94.050 ;
        RECT 118.950 93.600 121.050 94.050 ;
        RECT 88.950 92.400 103.050 93.600 ;
        RECT 88.950 91.950 91.050 92.400 ;
        RECT 100.950 91.950 103.050 92.400 ;
        RECT 104.400 92.400 121.050 93.600 ;
        RECT 4.950 90.600 7.050 91.050 ;
        RECT 10.950 90.600 13.050 91.050 ;
        RECT 4.950 89.400 13.050 90.600 ;
        RECT 4.950 88.950 7.050 89.400 ;
        RECT 10.950 88.950 13.050 89.400 ;
        RECT 61.950 90.600 64.050 91.050 ;
        RECT 77.400 90.600 78.600 91.950 ;
        RECT 94.950 90.600 97.050 91.050 ;
        RECT 104.400 90.600 105.600 92.400 ;
        RECT 118.950 91.950 121.050 92.400 ;
        RECT 145.950 93.600 148.050 94.050 ;
        RECT 151.950 93.600 154.050 94.050 ;
        RECT 145.950 92.400 154.050 93.600 ;
        RECT 145.950 91.950 148.050 92.400 ;
        RECT 151.950 91.950 154.050 92.400 ;
        RECT 169.950 93.600 172.050 94.050 ;
        RECT 178.950 93.600 181.050 94.050 ;
        RECT 169.950 92.400 181.050 93.600 ;
        RECT 169.950 91.950 172.050 92.400 ;
        RECT 178.950 91.950 181.050 92.400 ;
        RECT 184.950 91.950 187.050 94.050 ;
        RECT 211.950 93.600 214.050 94.050 ;
        RECT 229.950 93.600 232.050 94.050 ;
        RECT 211.950 92.400 232.050 93.600 ;
        RECT 211.950 91.950 214.050 92.400 ;
        RECT 229.950 91.950 232.050 92.400 ;
        RECT 238.950 93.600 241.050 94.050 ;
        RECT 247.950 93.600 250.050 94.050 ;
        RECT 238.950 92.400 250.050 93.600 ;
        RECT 238.950 91.950 241.050 92.400 ;
        RECT 247.950 91.950 250.050 92.400 ;
        RECT 253.950 93.600 256.050 94.050 ;
        RECT 265.950 93.600 268.050 94.050 ;
        RECT 253.950 92.400 268.050 93.600 ;
        RECT 253.950 91.950 256.050 92.400 ;
        RECT 265.950 91.950 268.050 92.400 ;
        RECT 277.950 93.600 280.050 94.050 ;
        RECT 286.950 93.600 289.050 94.050 ;
        RECT 277.950 92.400 289.050 93.600 ;
        RECT 277.950 91.950 280.050 92.400 ;
        RECT 286.950 91.950 289.050 92.400 ;
        RECT 292.950 93.600 295.050 94.050 ;
        RECT 298.950 93.600 301.050 94.050 ;
        RECT 370.950 93.600 373.050 94.050 ;
        RECT 292.950 92.400 301.050 93.600 ;
        RECT 292.950 91.950 295.050 92.400 ;
        RECT 298.950 91.950 301.050 92.400 ;
        RECT 353.400 92.400 373.050 93.600 ;
        RECT 353.400 91.050 354.600 92.400 ;
        RECT 370.950 91.950 373.050 92.400 ;
        RECT 391.950 93.600 394.050 94.050 ;
        RECT 409.950 93.600 412.050 94.050 ;
        RECT 391.950 92.400 423.600 93.600 ;
        RECT 391.950 91.950 394.050 92.400 ;
        RECT 409.950 91.950 412.050 92.400 ;
        RECT 61.950 89.400 105.600 90.600 ;
        RECT 127.950 90.600 130.050 91.050 ;
        RECT 160.950 90.600 163.050 91.050 ;
        RECT 127.950 89.400 163.050 90.600 ;
        RECT 61.950 88.950 64.050 89.400 ;
        RECT 94.950 88.950 97.050 89.400 ;
        RECT 127.950 88.950 130.050 89.400 ;
        RECT 160.950 88.950 163.050 89.400 ;
        RECT 178.950 90.600 181.050 91.050 ;
        RECT 232.950 90.600 235.050 91.050 ;
        RECT 178.950 89.400 235.050 90.600 ;
        RECT 178.950 88.950 181.050 89.400 ;
        RECT 232.950 88.950 235.050 89.400 ;
        RECT 256.950 90.600 259.050 91.050 ;
        RECT 274.950 90.600 277.050 91.050 ;
        RECT 307.950 90.600 310.050 91.050 ;
        RECT 256.950 89.400 310.050 90.600 ;
        RECT 256.950 88.950 259.050 89.400 ;
        RECT 274.950 88.950 277.050 89.400 ;
        RECT 307.950 88.950 310.050 89.400 ;
        RECT 352.950 88.950 355.050 91.050 ;
        RECT 422.400 90.600 423.600 92.400 ;
        RECT 424.950 91.950 427.050 94.050 ;
        RECT 448.950 93.600 451.050 94.050 ;
        RECT 460.950 93.600 463.050 94.050 ;
        RECT 448.950 92.400 463.050 93.600 ;
        RECT 448.950 91.950 451.050 92.400 ;
        RECT 460.950 91.950 463.050 92.400 ;
        RECT 466.950 93.600 469.050 94.050 ;
        RECT 475.950 93.600 478.050 94.050 ;
        RECT 466.950 92.400 478.050 93.600 ;
        RECT 466.950 91.950 469.050 92.400 ;
        RECT 475.950 91.950 478.050 92.400 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 493.950 93.600 496.050 94.050 ;
        RECT 499.950 93.600 502.050 94.050 ;
        RECT 523.950 93.600 526.050 94.050 ;
        RECT 493.950 92.400 526.050 93.600 ;
        RECT 493.950 91.950 496.050 92.400 ;
        RECT 499.950 91.950 502.050 92.400 ;
        RECT 523.950 91.950 526.050 92.400 ;
        RECT 529.950 93.600 532.050 94.050 ;
        RECT 542.400 93.600 543.600 94.950 ;
        RECT 553.950 93.600 556.050 94.050 ;
        RECT 568.950 93.600 571.050 94.050 ;
        RECT 583.950 93.600 586.050 94.050 ;
        RECT 529.950 92.400 549.600 93.600 ;
        RECT 529.950 91.950 532.050 92.400 ;
        RECT 445.950 90.600 448.050 91.050 ;
        RECT 422.400 89.400 448.050 90.600 ;
        RECT 445.950 88.950 448.050 89.400 ;
        RECT 451.950 90.600 454.050 91.050 ;
        RECT 484.950 90.600 487.050 91.050 ;
        RECT 451.950 89.400 487.050 90.600 ;
        RECT 488.400 90.600 489.600 91.950 ;
        RECT 502.950 90.600 505.050 91.050 ;
        RECT 488.400 89.400 505.050 90.600 ;
        RECT 451.950 88.950 454.050 89.400 ;
        RECT 484.950 88.950 487.050 89.400 ;
        RECT 502.950 88.950 505.050 89.400 ;
        RECT 10.950 87.600 13.050 88.050 ;
        RECT 22.950 87.600 25.050 88.050 ;
        RECT 10.950 86.400 25.050 87.600 ;
        RECT 10.950 85.950 13.050 86.400 ;
        RECT 22.950 85.950 25.050 86.400 ;
        RECT 100.950 87.600 103.050 88.050 ;
        RECT 115.950 87.600 118.050 88.050 ;
        RECT 196.950 87.600 199.050 88.050 ;
        RECT 100.950 86.400 199.050 87.600 ;
        RECT 100.950 85.950 103.050 86.400 ;
        RECT 115.950 85.950 118.050 86.400 ;
        RECT 196.950 85.950 199.050 86.400 ;
        RECT 211.950 87.600 214.050 88.050 ;
        RECT 268.950 87.600 271.050 88.050 ;
        RECT 211.950 86.400 271.050 87.600 ;
        RECT 211.950 85.950 214.050 86.400 ;
        RECT 268.950 85.950 271.050 86.400 ;
        RECT 325.950 87.600 328.050 88.050 ;
        RECT 418.950 87.600 421.050 88.050 ;
        RECT 463.950 87.600 466.050 88.050 ;
        RECT 325.950 86.400 466.050 87.600 ;
        RECT 524.400 87.600 525.600 91.950 ;
        RECT 548.400 91.050 549.600 92.400 ;
        RECT 553.950 92.400 586.050 93.600 ;
        RECT 553.950 91.950 556.050 92.400 ;
        RECT 568.950 91.950 571.050 92.400 ;
        RECT 583.950 91.950 586.050 92.400 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 559.950 90.600 562.050 91.050 ;
        RECT 587.400 90.600 588.600 94.950 ;
        RECT 629.400 94.050 630.600 95.400 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 694.950 96.600 697.050 97.050 ;
        RECT 706.950 96.600 709.050 97.050 ;
        RECT 694.950 95.400 709.050 96.600 ;
        RECT 694.950 94.950 697.050 95.400 ;
        RECT 706.950 94.950 709.050 95.400 ;
        RECT 709.950 94.950 712.050 97.050 ;
        RECT 715.950 96.600 718.050 97.050 ;
        RECT 727.950 96.600 730.050 97.050 ;
        RECT 715.950 95.400 730.050 96.600 ;
        RECT 715.950 94.950 718.050 95.400 ;
        RECT 727.950 94.950 730.050 95.400 ;
        RECT 733.950 94.950 736.050 97.050 ;
        RECT 769.950 96.600 772.050 97.050 ;
        RECT 790.950 96.600 793.050 97.050 ;
        RECT 811.950 96.600 814.050 97.050 ;
        RECT 829.950 96.600 832.050 97.050 ;
        RECT 769.950 95.400 793.050 96.600 ;
        RECT 769.950 94.950 772.050 95.400 ;
        RECT 790.950 94.950 793.050 95.400 ;
        RECT 794.400 95.400 832.050 96.600 ;
        RECT 598.950 93.600 601.050 94.050 ;
        RECT 607.950 93.600 610.050 94.050 ;
        RECT 598.950 92.400 610.050 93.600 ;
        RECT 598.950 91.950 601.050 92.400 ;
        RECT 607.950 91.950 610.050 92.400 ;
        RECT 628.950 91.950 631.050 94.050 ;
        RECT 632.400 91.050 633.600 94.950 ;
        RECT 634.950 93.600 637.050 94.050 ;
        RECT 649.950 93.600 652.050 94.050 ;
        RECT 634.950 92.400 652.050 93.600 ;
        RECT 634.950 91.950 637.050 92.400 ;
        RECT 649.950 91.950 652.050 92.400 ;
        RECT 658.950 93.600 661.050 94.050 ;
        RECT 667.950 93.600 670.050 94.050 ;
        RECT 658.950 92.400 670.050 93.600 ;
        RECT 658.950 91.950 661.050 92.400 ;
        RECT 667.950 91.950 670.050 92.400 ;
        RECT 685.950 91.950 688.050 94.050 ;
        RECT 691.950 93.600 694.050 94.050 ;
        RECT 697.950 93.600 700.050 94.050 ;
        RECT 710.400 93.600 711.600 94.950 ;
        RECT 691.950 92.400 700.050 93.600 ;
        RECT 691.950 91.950 694.050 92.400 ;
        RECT 697.950 91.950 700.050 92.400 ;
        RECT 701.400 92.400 711.600 93.600 ;
        RECT 712.950 93.600 715.050 94.050 ;
        RECT 718.950 93.600 721.050 94.050 ;
        RECT 712.950 92.400 721.050 93.600 ;
        RECT 559.950 89.400 588.600 90.600 ;
        RECT 559.950 88.950 562.050 89.400 ;
        RECT 631.950 88.950 634.050 91.050 ;
        RECT 686.400 90.600 687.600 91.950 ;
        RECT 701.400 90.600 702.600 92.400 ;
        RECT 712.950 91.950 715.050 92.400 ;
        RECT 718.950 91.950 721.050 92.400 ;
        RECT 724.950 93.600 727.050 94.050 ;
        RECT 730.950 93.600 733.050 94.050 ;
        RECT 724.950 92.400 733.050 93.600 ;
        RECT 724.950 91.950 727.050 92.400 ;
        RECT 730.950 91.950 733.050 92.400 ;
        RECT 635.400 89.400 702.600 90.600 ;
        RECT 721.950 90.600 724.050 91.050 ;
        RECT 734.400 90.600 735.600 94.950 ;
        RECT 787.950 93.600 790.050 94.050 ;
        RECT 794.400 93.600 795.600 95.400 ;
        RECT 811.950 94.950 814.050 95.400 ;
        RECT 829.950 94.950 832.050 95.400 ;
        RECT 838.950 96.600 841.050 97.050 ;
        RECT 853.950 96.600 856.050 97.050 ;
        RECT 838.950 95.400 856.050 96.600 ;
        RECT 838.950 94.950 841.050 95.400 ;
        RECT 853.950 94.950 856.050 95.400 ;
        RECT 787.950 92.400 795.600 93.600 ;
        RECT 808.950 93.600 811.050 94.050 ;
        RECT 820.950 93.600 823.050 94.050 ;
        RECT 835.950 93.600 838.050 94.050 ;
        RECT 808.950 92.400 838.050 93.600 ;
        RECT 787.950 91.950 790.050 92.400 ;
        RECT 808.950 91.950 811.050 92.400 ;
        RECT 820.950 91.950 823.050 92.400 ;
        RECT 835.950 91.950 838.050 92.400 ;
        RECT 721.950 89.400 735.600 90.600 ;
        RECT 793.950 90.600 796.050 91.050 ;
        RECT 799.950 90.600 802.050 91.050 ;
        RECT 793.950 89.400 802.050 90.600 ;
        RECT 635.400 87.600 636.600 89.400 ;
        RECT 721.950 88.950 724.050 89.400 ;
        RECT 793.950 88.950 796.050 89.400 ;
        RECT 799.950 88.950 802.050 89.400 ;
        RECT 847.950 90.600 850.050 91.050 ;
        RECT 859.950 90.600 862.050 91.050 ;
        RECT 847.950 89.400 862.050 90.600 ;
        RECT 847.950 88.950 850.050 89.400 ;
        RECT 859.950 88.950 862.050 89.400 ;
        RECT 524.400 86.400 636.600 87.600 ;
        RECT 325.950 85.950 328.050 86.400 ;
        RECT 418.950 85.950 421.050 86.400 ;
        RECT 463.950 85.950 466.050 86.400 ;
        RECT 184.950 84.600 187.050 85.050 ;
        RECT 205.950 84.600 208.050 85.050 ;
        RECT 220.950 84.600 223.050 85.050 ;
        RECT 184.950 83.400 223.050 84.600 ;
        RECT 184.950 82.950 187.050 83.400 ;
        RECT 205.950 82.950 208.050 83.400 ;
        RECT 220.950 82.950 223.050 83.400 ;
        RECT 274.950 84.600 277.050 85.050 ;
        RECT 373.950 84.600 376.050 85.050 ;
        RECT 274.950 83.400 376.050 84.600 ;
        RECT 274.950 82.950 277.050 83.400 ;
        RECT 373.950 82.950 376.050 83.400 ;
        RECT 487.950 84.600 490.050 85.050 ;
        RECT 502.950 84.600 505.050 85.050 ;
        RECT 631.950 84.600 634.050 85.050 ;
        RECT 487.950 83.400 634.050 84.600 ;
        RECT 487.950 82.950 490.050 83.400 ;
        RECT 502.950 82.950 505.050 83.400 ;
        RECT 631.950 82.950 634.050 83.400 ;
        RECT 22.950 81.600 25.050 82.050 ;
        RECT 67.950 81.600 70.050 82.050 ;
        RECT 76.950 81.600 79.050 82.050 ;
        RECT 22.950 80.400 79.050 81.600 ;
        RECT 22.950 79.950 25.050 80.400 ;
        RECT 67.950 79.950 70.050 80.400 ;
        RECT 76.950 79.950 79.050 80.400 ;
        RECT 166.950 81.600 169.050 82.050 ;
        RECT 172.950 81.600 175.050 82.050 ;
        RECT 166.950 80.400 175.050 81.600 ;
        RECT 166.950 79.950 169.050 80.400 ;
        RECT 172.950 79.950 175.050 80.400 ;
        RECT 349.950 81.600 352.050 82.050 ;
        RECT 388.950 81.600 391.050 82.050 ;
        RECT 403.950 81.600 406.050 82.050 ;
        RECT 445.950 81.600 448.050 82.050 ;
        RECT 472.950 81.600 475.050 82.050 ;
        RECT 349.950 80.400 475.050 81.600 ;
        RECT 349.950 79.950 352.050 80.400 ;
        RECT 388.950 79.950 391.050 80.400 ;
        RECT 403.950 79.950 406.050 80.400 ;
        RECT 445.950 79.950 448.050 80.400 ;
        RECT 472.950 79.950 475.050 80.400 ;
        RECT 586.950 81.600 589.050 82.050 ;
        RECT 592.950 81.600 595.050 82.050 ;
        RECT 586.950 80.400 595.050 81.600 ;
        RECT 586.950 79.950 589.050 80.400 ;
        RECT 592.950 79.950 595.050 80.400 ;
        RECT 823.950 81.600 826.050 82.050 ;
        RECT 850.950 81.600 853.050 82.050 ;
        RECT 823.950 80.400 853.050 81.600 ;
        RECT 823.950 79.950 826.050 80.400 ;
        RECT 850.950 79.950 853.050 80.400 ;
        RECT 394.950 78.600 397.050 79.050 ;
        RECT 415.950 78.600 418.050 79.050 ;
        RECT 418.950 78.600 421.050 79.050 ;
        RECT 394.950 77.400 421.050 78.600 ;
        RECT 394.950 76.950 397.050 77.400 ;
        RECT 415.950 76.950 418.050 77.400 ;
        RECT 418.950 76.950 421.050 77.400 ;
        RECT 571.950 78.600 574.050 79.050 ;
        RECT 601.950 78.600 604.050 79.050 ;
        RECT 571.950 77.400 604.050 78.600 ;
        RECT 571.950 76.950 574.050 77.400 ;
        RECT 601.950 76.950 604.050 77.400 ;
        RECT 781.950 78.600 784.050 79.050 ;
        RECT 808.950 78.600 811.050 79.050 ;
        RECT 781.950 77.400 811.050 78.600 ;
        RECT 781.950 76.950 784.050 77.400 ;
        RECT 808.950 76.950 811.050 77.400 ;
        RECT 310.950 75.600 313.050 76.050 ;
        RECT 343.950 75.600 346.050 76.050 ;
        RECT 310.950 74.400 346.050 75.600 ;
        RECT 310.950 73.950 313.050 74.400 ;
        RECT 343.950 73.950 346.050 74.400 ;
        RECT 718.950 75.600 721.050 76.050 ;
        RECT 826.950 75.600 829.050 76.050 ;
        RECT 718.950 74.400 829.050 75.600 ;
        RECT 718.950 73.950 721.050 74.400 ;
        RECT 826.950 73.950 829.050 74.400 ;
        RECT 763.950 72.600 766.050 73.050 ;
        RECT 811.950 72.600 814.050 73.050 ;
        RECT 838.950 72.600 841.050 73.050 ;
        RECT 763.950 71.400 841.050 72.600 ;
        RECT 763.950 70.950 766.050 71.400 ;
        RECT 811.950 70.950 814.050 71.400 ;
        RECT 838.950 70.950 841.050 71.400 ;
        RECT 397.950 69.600 400.050 70.050 ;
        RECT 436.950 69.600 439.050 70.050 ;
        RECT 397.950 68.400 439.050 69.600 ;
        RECT 397.950 67.950 400.050 68.400 ;
        RECT 436.950 67.950 439.050 68.400 ;
        RECT 475.950 69.600 478.050 70.050 ;
        RECT 553.950 69.600 556.050 70.050 ;
        RECT 475.950 68.400 556.050 69.600 ;
        RECT 475.950 67.950 478.050 68.400 ;
        RECT 553.950 67.950 556.050 68.400 ;
        RECT 673.950 69.600 676.050 70.050 ;
        RECT 679.950 69.600 682.050 70.050 ;
        RECT 673.950 68.400 682.050 69.600 ;
        RECT 673.950 67.950 676.050 68.400 ;
        RECT 679.950 67.950 682.050 68.400 ;
        RECT 787.950 69.600 790.050 70.050 ;
        RECT 802.950 69.600 805.050 70.050 ;
        RECT 787.950 68.400 805.050 69.600 ;
        RECT 787.950 67.950 790.050 68.400 ;
        RECT 802.950 67.950 805.050 68.400 ;
        RECT 388.950 66.600 391.050 67.050 ;
        RECT 523.950 66.600 526.050 67.050 ;
        RECT 388.950 65.400 526.050 66.600 ;
        RECT 388.950 64.950 391.050 65.400 ;
        RECT 523.950 64.950 526.050 65.400 ;
        RECT 616.950 66.600 619.050 67.050 ;
        RECT 628.950 66.600 631.050 67.050 ;
        RECT 616.950 65.400 631.050 66.600 ;
        RECT 616.950 64.950 619.050 65.400 ;
        RECT 628.950 64.950 631.050 65.400 ;
        RECT 772.950 66.600 775.050 67.050 ;
        RECT 841.950 66.600 844.050 67.050 ;
        RECT 772.950 65.400 844.050 66.600 ;
        RECT 772.950 64.950 775.050 65.400 ;
        RECT 841.950 64.950 844.050 65.400 ;
        RECT 43.950 63.600 46.050 64.050 ;
        RECT 82.950 63.600 85.050 64.050 ;
        RECT 43.950 62.400 85.050 63.600 ;
        RECT 43.950 61.950 46.050 62.400 ;
        RECT 82.950 61.950 85.050 62.400 ;
        RECT 151.950 63.600 154.050 64.050 ;
        RECT 244.950 63.600 247.050 64.050 ;
        RECT 151.950 62.400 247.050 63.600 ;
        RECT 151.950 61.950 154.050 62.400 ;
        RECT 244.950 61.950 247.050 62.400 ;
        RECT 337.950 63.600 340.050 64.050 ;
        RECT 379.950 63.600 382.050 64.050 ;
        RECT 337.950 62.400 382.050 63.600 ;
        RECT 337.950 61.950 340.050 62.400 ;
        RECT 379.950 61.950 382.050 62.400 ;
        RECT 424.950 63.600 427.050 64.050 ;
        RECT 469.950 63.600 472.050 64.050 ;
        RECT 496.950 63.600 499.050 64.050 ;
        RECT 424.950 62.400 499.050 63.600 ;
        RECT 424.950 61.950 427.050 62.400 ;
        RECT 469.950 61.950 472.050 62.400 ;
        RECT 496.950 61.950 499.050 62.400 ;
        RECT 769.950 63.600 772.050 64.050 ;
        RECT 802.950 63.600 805.050 64.050 ;
        RECT 769.950 62.400 805.050 63.600 ;
        RECT 769.950 61.950 772.050 62.400 ;
        RECT 802.950 61.950 805.050 62.400 ;
        RECT 109.950 60.600 112.050 61.050 ;
        RECT 121.950 60.600 124.050 61.050 ;
        RECT 109.950 59.400 124.050 60.600 ;
        RECT 109.950 58.950 112.050 59.400 ;
        RECT 121.950 58.950 124.050 59.400 ;
        RECT 220.950 60.600 223.050 61.050 ;
        RECT 286.950 60.600 289.050 61.050 ;
        RECT 220.950 59.400 289.050 60.600 ;
        RECT 220.950 58.950 223.050 59.400 ;
        RECT 286.950 58.950 289.050 59.400 ;
        RECT 352.950 60.600 355.050 61.050 ;
        RECT 394.950 60.600 397.050 61.050 ;
        RECT 352.950 59.400 397.050 60.600 ;
        RECT 352.950 58.950 355.050 59.400 ;
        RECT 394.950 58.950 397.050 59.400 ;
        RECT 406.950 60.600 409.050 61.050 ;
        RECT 457.950 60.600 460.050 61.050 ;
        RECT 406.950 59.400 460.050 60.600 ;
        RECT 406.950 58.950 409.050 59.400 ;
        RECT 457.950 58.950 460.050 59.400 ;
        RECT 481.950 60.600 484.050 61.050 ;
        RECT 511.950 60.600 514.050 61.050 ;
        RECT 481.950 59.400 514.050 60.600 ;
        RECT 481.950 58.950 484.050 59.400 ;
        RECT 511.950 58.950 514.050 59.400 ;
        RECT 523.950 60.600 526.050 61.050 ;
        RECT 535.950 60.600 538.050 61.050 ;
        RECT 523.950 59.400 538.050 60.600 ;
        RECT 523.950 58.950 526.050 59.400 ;
        RECT 535.950 58.950 538.050 59.400 ;
        RECT 538.950 60.600 541.050 61.050 ;
        RECT 559.950 60.600 562.050 61.050 ;
        RECT 538.950 59.400 562.050 60.600 ;
        RECT 538.950 58.950 541.050 59.400 ;
        RECT 559.950 58.950 562.050 59.400 ;
        RECT 568.950 60.600 571.050 61.050 ;
        RECT 574.950 60.600 577.050 61.050 ;
        RECT 622.950 60.600 625.050 61.050 ;
        RECT 568.950 59.400 577.050 60.600 ;
        RECT 568.950 58.950 571.050 59.400 ;
        RECT 574.950 58.950 577.050 59.400 ;
        RECT 620.400 59.400 625.050 60.600 ;
        RECT 620.400 58.050 621.600 59.400 ;
        RECT 622.950 58.950 625.050 59.400 ;
        RECT 625.950 60.600 628.050 61.050 ;
        RECT 676.950 60.600 679.050 61.050 ;
        RECT 625.950 59.400 679.050 60.600 ;
        RECT 625.950 58.950 628.050 59.400 ;
        RECT 676.950 58.950 679.050 59.400 ;
        RECT 760.950 60.600 763.050 61.050 ;
        RECT 793.950 60.600 796.050 61.050 ;
        RECT 760.950 59.400 796.050 60.600 ;
        RECT 760.950 58.950 763.050 59.400 ;
        RECT 793.950 58.950 796.050 59.400 ;
        RECT 805.950 60.600 808.050 61.050 ;
        RECT 826.950 60.600 829.050 61.050 ;
        RECT 832.950 60.600 835.050 61.050 ;
        RECT 844.950 60.600 847.050 61.050 ;
        RECT 805.950 59.400 847.050 60.600 ;
        RECT 805.950 58.950 808.050 59.400 ;
        RECT 826.950 58.950 829.050 59.400 ;
        RECT 832.950 58.950 835.050 59.400 ;
        RECT 844.950 58.950 847.050 59.400 ;
        RECT 856.950 60.600 859.050 61.050 ;
        RECT 862.950 60.600 865.050 61.050 ;
        RECT 856.950 59.400 865.050 60.600 ;
        RECT 856.950 58.950 859.050 59.400 ;
        RECT 862.950 58.950 865.050 59.400 ;
        RECT 61.950 57.600 64.050 58.050 ;
        RECT 118.950 57.600 121.050 58.050 ;
        RECT 32.400 56.400 64.050 57.600 ;
        RECT 32.400 55.050 33.600 56.400 ;
        RECT 61.950 55.950 64.050 56.400 ;
        RECT 83.400 56.400 121.050 57.600 ;
        RECT 13.950 54.600 16.050 55.050 ;
        RECT 31.950 54.600 34.050 55.050 ;
        RECT 13.950 53.400 34.050 54.600 ;
        RECT 13.950 52.950 16.050 53.400 ;
        RECT 31.950 52.950 34.050 53.400 ;
        RECT 37.950 54.600 40.050 55.050 ;
        RECT 43.950 54.600 46.050 55.050 ;
        RECT 37.950 53.400 46.050 54.600 ;
        RECT 37.950 52.950 40.050 53.400 ;
        RECT 43.950 52.950 46.050 53.400 ;
        RECT 61.950 52.950 64.050 55.050 ;
        RECT 67.950 54.600 70.050 55.050 ;
        RECT 79.950 54.600 82.050 55.050 ;
        RECT 83.400 54.600 84.600 56.400 ;
        RECT 118.950 55.950 121.050 56.400 ;
        RECT 142.950 57.600 145.050 58.050 ;
        RECT 154.950 57.600 157.050 58.050 ;
        RECT 160.950 57.600 163.050 58.050 ;
        RECT 202.950 57.600 205.050 58.050 ;
        RECT 142.950 56.400 163.050 57.600 ;
        RECT 142.950 55.950 145.050 56.400 ;
        RECT 154.950 55.950 157.050 56.400 ;
        RECT 160.950 55.950 163.050 56.400 ;
        RECT 167.400 56.400 205.050 57.600 ;
        RECT 67.950 53.400 84.600 54.600 ;
        RECT 67.950 52.950 70.050 53.400 ;
        RECT 79.950 52.950 82.050 53.400 ;
        RECT 145.950 52.950 148.050 55.050 ;
        RECT 148.950 54.600 151.050 55.050 ;
        RECT 163.950 54.600 166.050 55.050 ;
        RECT 167.400 54.600 168.600 56.400 ;
        RECT 202.950 55.950 205.050 56.400 ;
        RECT 208.950 57.600 211.050 58.050 ;
        RECT 226.950 57.600 229.050 58.050 ;
        RECT 238.950 57.600 241.050 58.050 ;
        RECT 208.950 56.400 241.050 57.600 ;
        RECT 208.950 55.950 211.050 56.400 ;
        RECT 226.950 55.950 229.050 56.400 ;
        RECT 238.950 55.950 241.050 56.400 ;
        RECT 247.950 57.600 250.050 58.050 ;
        RECT 253.950 57.600 256.050 58.050 ;
        RECT 247.950 56.400 256.050 57.600 ;
        RECT 247.950 55.950 250.050 56.400 ;
        RECT 253.950 55.950 256.050 56.400 ;
        RECT 265.950 57.600 268.050 58.050 ;
        RECT 277.950 57.600 280.050 58.050 ;
        RECT 298.950 57.600 301.050 58.050 ;
        RECT 382.950 57.600 385.050 58.050 ;
        RECT 430.950 57.600 433.050 58.050 ;
        RECT 529.950 57.600 532.050 58.050 ;
        RECT 550.950 57.600 553.050 58.050 ;
        RECT 265.950 56.400 553.050 57.600 ;
        RECT 265.950 55.950 268.050 56.400 ;
        RECT 277.950 55.950 280.050 56.400 ;
        RECT 298.950 55.950 301.050 56.400 ;
        RECT 382.950 55.950 385.050 56.400 ;
        RECT 430.950 55.950 433.050 56.400 ;
        RECT 529.950 55.950 532.050 56.400 ;
        RECT 550.950 55.950 553.050 56.400 ;
        RECT 577.950 57.600 580.050 58.050 ;
        RECT 589.950 57.600 592.050 58.050 ;
        RECT 613.950 57.600 616.050 58.050 ;
        RECT 577.950 56.400 616.050 57.600 ;
        RECT 577.950 55.950 580.050 56.400 ;
        RECT 589.950 55.950 592.050 56.400 ;
        RECT 613.950 55.950 616.050 56.400 ;
        RECT 619.950 57.600 622.050 58.050 ;
        RECT 661.950 57.600 664.050 58.050 ;
        RECT 619.950 56.400 664.050 57.600 ;
        RECT 619.950 55.950 622.050 56.400 ;
        RECT 661.950 55.950 664.050 56.400 ;
        RECT 676.950 57.600 679.050 58.050 ;
        RECT 721.950 57.600 724.050 58.050 ;
        RECT 676.950 56.400 724.050 57.600 ;
        RECT 676.950 55.950 679.050 56.400 ;
        RECT 721.950 55.950 724.050 56.400 ;
        RECT 751.950 57.600 754.050 58.050 ;
        RECT 751.950 56.400 771.600 57.600 ;
        RECT 751.950 55.950 754.050 56.400 ;
        RECT 770.400 55.050 771.600 56.400 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 775.950 57.600 778.050 58.050 ;
        RECT 814.950 57.600 817.050 58.050 ;
        RECT 775.950 56.400 817.050 57.600 ;
        RECT 775.950 55.950 778.050 56.400 ;
        RECT 814.950 55.950 817.050 56.400 ;
        RECT 841.950 57.600 844.050 58.050 ;
        RECT 841.950 56.400 846.600 57.600 ;
        RECT 841.950 55.950 844.050 56.400 ;
        RECT 148.950 53.400 168.600 54.600 ;
        RECT 205.950 54.600 208.050 55.050 ;
        RECT 217.950 54.600 220.050 55.050 ;
        RECT 205.950 53.400 220.050 54.600 ;
        RECT 148.950 52.950 151.050 53.400 ;
        RECT 163.950 52.950 166.050 53.400 ;
        RECT 205.950 52.950 208.050 53.400 ;
        RECT 217.950 52.950 220.050 53.400 ;
        RECT 241.950 54.600 244.050 55.050 ;
        RECT 256.950 54.600 259.050 55.050 ;
        RECT 241.950 53.400 259.050 54.600 ;
        RECT 241.950 52.950 244.050 53.400 ;
        RECT 256.950 52.950 259.050 53.400 ;
        RECT 304.950 54.600 307.050 55.050 ;
        RECT 319.950 54.600 322.050 55.050 ;
        RECT 304.950 53.400 322.050 54.600 ;
        RECT 304.950 52.950 307.050 53.400 ;
        RECT 319.950 52.950 322.050 53.400 ;
        RECT 331.950 54.600 334.050 55.050 ;
        RECT 343.950 54.600 346.050 55.050 ;
        RECT 361.950 54.600 364.050 55.050 ;
        RECT 331.950 53.400 364.050 54.600 ;
        RECT 331.950 52.950 334.050 53.400 ;
        RECT 343.950 52.950 346.050 53.400 ;
        RECT 361.950 52.950 364.050 53.400 ;
        RECT 379.950 54.600 382.050 55.050 ;
        RECT 409.950 54.600 412.050 55.050 ;
        RECT 379.950 53.400 412.050 54.600 ;
        RECT 379.950 52.950 382.050 53.400 ;
        RECT 409.950 52.950 412.050 53.400 ;
        RECT 451.950 54.600 454.050 55.050 ;
        RECT 472.950 54.600 475.050 55.050 ;
        RECT 451.950 53.400 475.050 54.600 ;
        RECT 451.950 52.950 454.050 53.400 ;
        RECT 472.950 52.950 475.050 53.400 ;
        RECT 475.950 54.600 478.050 55.050 ;
        RECT 487.950 54.600 490.050 55.050 ;
        RECT 475.950 53.400 490.050 54.600 ;
        RECT 475.950 52.950 478.050 53.400 ;
        RECT 487.950 52.950 490.050 53.400 ;
        RECT 517.950 54.600 520.050 55.050 ;
        RECT 544.950 54.600 547.050 55.050 ;
        RECT 517.950 53.400 547.050 54.600 ;
        RECT 517.950 52.950 520.050 53.400 ;
        RECT 544.950 52.950 547.050 53.400 ;
        RECT 586.950 54.600 589.050 55.050 ;
        RECT 592.950 54.600 595.050 55.050 ;
        RECT 586.950 53.400 595.050 54.600 ;
        RECT 586.950 52.950 589.050 53.400 ;
        RECT 592.950 52.950 595.050 53.400 ;
        RECT 601.950 54.600 604.050 55.050 ;
        RECT 616.950 54.600 619.050 55.050 ;
        RECT 601.950 53.400 619.050 54.600 ;
        RECT 601.950 52.950 604.050 53.400 ;
        RECT 616.950 52.950 619.050 53.400 ;
        RECT 628.950 54.600 631.050 55.050 ;
        RECT 628.950 53.400 636.600 54.600 ;
        RECT 628.950 52.950 631.050 53.400 ;
        RECT 16.950 51.600 19.050 52.050 ;
        RECT 46.950 51.600 49.050 52.050 ;
        RECT 55.950 51.600 58.050 52.050 ;
        RECT 16.950 50.400 58.050 51.600 ;
        RECT 62.400 51.600 63.600 52.950 ;
        RECT 97.950 51.600 100.050 52.050 ;
        RECT 62.400 50.400 100.050 51.600 ;
        RECT 16.950 49.950 19.050 50.400 ;
        RECT 46.950 49.950 49.050 50.400 ;
        RECT 55.950 49.950 58.050 50.400 ;
        RECT 97.950 49.950 100.050 50.400 ;
        RECT 139.950 51.600 142.050 52.050 ;
        RECT 146.400 51.600 147.600 52.950 ;
        RECT 139.950 50.400 147.600 51.600 ;
        RECT 187.950 51.600 190.050 52.050 ;
        RECT 199.950 51.600 202.050 52.050 ;
        RECT 187.950 50.400 202.050 51.600 ;
        RECT 139.950 49.950 142.050 50.400 ;
        RECT 187.950 49.950 190.050 50.400 ;
        RECT 199.950 49.950 202.050 50.400 ;
        RECT 250.950 51.600 253.050 52.050 ;
        RECT 259.950 51.600 262.050 52.050 ;
        RECT 250.950 50.400 262.050 51.600 ;
        RECT 250.950 49.950 253.050 50.400 ;
        RECT 259.950 49.950 262.050 50.400 ;
        RECT 271.950 51.600 274.050 52.050 ;
        RECT 286.950 51.600 289.050 52.050 ;
        RECT 340.950 51.600 343.050 52.050 ;
        RECT 271.950 50.400 343.050 51.600 ;
        RECT 271.950 49.950 274.050 50.400 ;
        RECT 286.950 49.950 289.050 50.400 ;
        RECT 340.950 49.950 343.050 50.400 ;
        RECT 367.950 51.600 370.050 52.050 ;
        RECT 400.950 51.600 403.050 52.050 ;
        RECT 367.950 50.400 403.050 51.600 ;
        RECT 367.950 49.950 370.050 50.400 ;
        RECT 400.950 49.950 403.050 50.400 ;
        RECT 403.950 51.600 406.050 52.050 ;
        RECT 412.950 51.600 415.050 52.050 ;
        RECT 403.950 50.400 415.050 51.600 ;
        RECT 403.950 49.950 406.050 50.400 ;
        RECT 412.950 49.950 415.050 50.400 ;
        RECT 430.950 51.600 433.050 52.050 ;
        RECT 439.950 51.600 442.050 52.050 ;
        RECT 430.950 50.400 442.050 51.600 ;
        RECT 430.950 49.950 433.050 50.400 ;
        RECT 439.950 49.950 442.050 50.400 ;
        RECT 556.950 51.600 559.050 52.050 ;
        RECT 574.950 51.600 577.050 52.050 ;
        RECT 556.950 50.400 577.050 51.600 ;
        RECT 556.950 49.950 559.050 50.400 ;
        RECT 574.950 49.950 577.050 50.400 ;
        RECT 580.950 51.600 583.050 52.050 ;
        RECT 598.950 51.600 601.050 52.050 ;
        RECT 631.950 51.600 634.050 52.050 ;
        RECT 580.950 50.400 634.050 51.600 ;
        RECT 635.400 51.600 636.600 53.400 ;
        RECT 640.950 52.950 643.050 55.050 ;
        RECT 655.950 54.600 658.050 55.050 ;
        RECT 673.950 54.600 676.050 55.050 ;
        RECT 679.950 54.600 682.050 55.050 ;
        RECT 655.950 53.400 672.600 54.600 ;
        RECT 655.950 52.950 658.050 53.400 ;
        RECT 637.950 51.600 640.050 52.050 ;
        RECT 635.400 50.400 640.050 51.600 ;
        RECT 580.950 49.950 583.050 50.400 ;
        RECT 598.950 49.950 601.050 50.400 ;
        RECT 631.950 49.950 634.050 50.400 ;
        RECT 637.950 49.950 640.050 50.400 ;
        RECT 37.950 48.600 40.050 49.050 ;
        RECT 43.950 48.600 46.050 49.050 ;
        RECT 64.950 48.600 67.050 49.050 ;
        RECT 37.950 47.400 67.050 48.600 ;
        RECT 37.950 46.950 40.050 47.400 ;
        RECT 43.950 46.950 46.050 47.400 ;
        RECT 64.950 46.950 67.050 47.400 ;
        RECT 229.950 48.600 232.050 49.050 ;
        RECT 241.950 48.600 244.050 49.050 ;
        RECT 229.950 47.400 244.050 48.600 ;
        RECT 229.950 46.950 232.050 47.400 ;
        RECT 241.950 46.950 244.050 47.400 ;
        RECT 346.950 48.600 349.050 49.050 ;
        RECT 352.950 48.600 355.050 49.050 ;
        RECT 346.950 47.400 355.050 48.600 ;
        RECT 346.950 46.950 349.050 47.400 ;
        RECT 352.950 46.950 355.050 47.400 ;
        RECT 364.950 48.600 367.050 49.050 ;
        RECT 385.950 48.600 388.050 49.050 ;
        RECT 364.950 47.400 388.050 48.600 ;
        RECT 364.950 46.950 367.050 47.400 ;
        RECT 385.950 46.950 388.050 47.400 ;
        RECT 424.950 48.600 427.050 49.050 ;
        RECT 433.950 48.600 436.050 49.050 ;
        RECT 424.950 47.400 436.050 48.600 ;
        RECT 424.950 46.950 427.050 47.400 ;
        RECT 433.950 46.950 436.050 47.400 ;
        RECT 436.950 48.600 439.050 49.050 ;
        RECT 448.950 48.600 451.050 49.050 ;
        RECT 436.950 47.400 451.050 48.600 ;
        RECT 436.950 46.950 439.050 47.400 ;
        RECT 448.950 46.950 451.050 47.400 ;
        RECT 472.950 48.600 475.050 49.050 ;
        RECT 490.950 48.600 493.050 49.050 ;
        RECT 499.950 48.600 502.050 49.050 ;
        RECT 472.950 47.400 502.050 48.600 ;
        RECT 472.950 46.950 475.050 47.400 ;
        RECT 490.950 46.950 493.050 47.400 ;
        RECT 499.950 46.950 502.050 47.400 ;
        RECT 625.950 48.600 628.050 49.050 ;
        RECT 641.400 48.600 642.600 52.950 ;
        RECT 671.400 51.600 672.600 53.400 ;
        RECT 673.950 53.400 682.050 54.600 ;
        RECT 673.950 52.950 676.050 53.400 ;
        RECT 679.950 52.950 682.050 53.400 ;
        RECT 685.950 54.600 688.050 55.050 ;
        RECT 694.950 54.600 697.050 55.050 ;
        RECT 685.950 53.400 697.050 54.600 ;
        RECT 685.950 52.950 688.050 53.400 ;
        RECT 694.950 52.950 697.050 53.400 ;
        RECT 700.950 54.600 703.050 55.050 ;
        RECT 709.950 54.600 712.050 55.050 ;
        RECT 742.950 54.600 745.050 55.050 ;
        RECT 700.950 53.400 712.050 54.600 ;
        RECT 700.950 52.950 703.050 53.400 ;
        RECT 709.950 52.950 712.050 53.400 ;
        RECT 734.400 53.400 745.050 54.600 ;
        RECT 734.400 52.050 735.600 53.400 ;
        RECT 742.950 52.950 745.050 53.400 ;
        RECT 769.950 52.950 772.050 55.050 ;
        RECT 773.400 54.600 774.600 55.950 ;
        RECT 845.400 55.050 846.600 56.400 ;
        RECT 775.950 54.600 778.050 55.050 ;
        RECT 773.400 53.400 778.050 54.600 ;
        RECT 775.950 52.950 778.050 53.400 ;
        RECT 784.950 54.600 787.050 55.050 ;
        RECT 799.950 54.600 802.050 55.050 ;
        RECT 784.950 53.400 802.050 54.600 ;
        RECT 784.950 52.950 787.050 53.400 ;
        RECT 799.950 52.950 802.050 53.400 ;
        RECT 820.950 52.950 823.050 55.050 ;
        RECT 844.950 52.950 847.050 55.050 ;
        RECT 859.950 54.600 862.050 55.050 ;
        RECT 868.950 54.600 871.050 55.050 ;
        RECT 859.950 53.400 871.050 54.600 ;
        RECT 859.950 52.950 862.050 53.400 ;
        RECT 868.950 52.950 871.050 53.400 ;
        RECT 688.950 51.600 691.050 52.050 ;
        RECT 671.400 50.400 691.050 51.600 ;
        RECT 688.950 49.950 691.050 50.400 ;
        RECT 733.950 49.950 736.050 52.050 ;
        RECT 754.950 51.600 757.050 52.050 ;
        RECT 772.950 51.600 775.050 52.050 ;
        RECT 754.950 50.400 775.050 51.600 ;
        RECT 754.950 49.950 757.050 50.400 ;
        RECT 772.950 49.950 775.050 50.400 ;
        RECT 778.950 51.600 781.050 52.050 ;
        RECT 805.950 51.600 808.050 52.050 ;
        RECT 778.950 50.400 808.050 51.600 ;
        RECT 821.400 51.600 822.600 52.950 ;
        RECT 841.950 51.600 844.050 52.050 ;
        RECT 821.400 50.400 844.050 51.600 ;
        RECT 778.950 49.950 781.050 50.400 ;
        RECT 805.950 49.950 808.050 50.400 ;
        RECT 841.950 49.950 844.050 50.400 ;
        RECT 625.950 47.400 642.600 48.600 ;
        RECT 646.950 48.600 649.050 49.050 ;
        RECT 691.950 48.600 694.050 49.050 ;
        RECT 646.950 47.400 694.050 48.600 ;
        RECT 625.950 46.950 628.050 47.400 ;
        RECT 646.950 46.950 649.050 47.400 ;
        RECT 691.950 46.950 694.050 47.400 ;
        RECT 712.950 48.600 715.050 49.050 ;
        RECT 721.950 48.600 724.050 49.050 ;
        RECT 712.950 47.400 724.050 48.600 ;
        RECT 712.950 46.950 715.050 47.400 ;
        RECT 721.950 46.950 724.050 47.400 ;
        RECT 745.950 48.600 748.050 49.050 ;
        RECT 769.950 48.600 772.050 49.050 ;
        RECT 745.950 47.400 772.050 48.600 ;
        RECT 745.950 46.950 748.050 47.400 ;
        RECT 769.950 46.950 772.050 47.400 ;
        RECT 811.950 48.600 814.050 49.050 ;
        RECT 823.950 48.600 826.050 49.050 ;
        RECT 811.950 47.400 826.050 48.600 ;
        RECT 811.950 46.950 814.050 47.400 ;
        RECT 823.950 46.950 826.050 47.400 ;
        RECT 49.950 45.600 52.050 46.050 ;
        RECT 58.950 45.600 61.050 46.050 ;
        RECT 49.950 44.400 61.050 45.600 ;
        RECT 49.950 43.950 52.050 44.400 ;
        RECT 58.950 43.950 61.050 44.400 ;
        RECT 145.950 45.600 148.050 46.050 ;
        RECT 157.950 45.600 160.050 46.050 ;
        RECT 244.950 45.600 247.050 46.050 ;
        RECT 145.950 44.400 247.050 45.600 ;
        RECT 145.950 43.950 148.050 44.400 ;
        RECT 157.950 43.950 160.050 44.400 ;
        RECT 244.950 43.950 247.050 44.400 ;
        RECT 355.950 45.600 358.050 46.050 ;
        RECT 394.950 45.600 397.050 46.050 ;
        RECT 355.950 44.400 397.050 45.600 ;
        RECT 355.950 43.950 358.050 44.400 ;
        RECT 394.950 43.950 397.050 44.400 ;
        RECT 514.950 45.600 517.050 46.050 ;
        RECT 550.950 45.600 553.050 46.050 ;
        RECT 634.950 45.600 637.050 46.050 ;
        RECT 661.950 45.600 664.050 46.050 ;
        RECT 514.950 44.400 664.050 45.600 ;
        RECT 514.950 43.950 517.050 44.400 ;
        RECT 550.950 43.950 553.050 44.400 ;
        RECT 634.950 43.950 637.050 44.400 ;
        RECT 661.950 43.950 664.050 44.400 ;
        RECT 121.950 42.600 124.050 43.050 ;
        RECT 160.950 42.600 163.050 43.050 ;
        RECT 178.950 42.600 181.050 43.050 ;
        RECT 121.950 41.400 181.050 42.600 ;
        RECT 121.950 40.950 124.050 41.400 ;
        RECT 160.950 40.950 163.050 41.400 ;
        RECT 178.950 40.950 181.050 41.400 ;
        RECT 625.950 42.600 628.050 43.050 ;
        RECT 685.950 42.600 688.050 43.050 ;
        RECT 625.950 41.400 688.050 42.600 ;
        RECT 625.950 40.950 628.050 41.400 ;
        RECT 685.950 40.950 688.050 41.400 ;
        RECT 40.950 39.600 43.050 40.050 ;
        RECT 55.950 39.600 58.050 40.050 ;
        RECT 88.950 39.600 91.050 40.050 ;
        RECT 40.950 38.400 91.050 39.600 ;
        RECT 40.950 37.950 43.050 38.400 ;
        RECT 55.950 37.950 58.050 38.400 ;
        RECT 88.950 37.950 91.050 38.400 ;
        RECT 601.950 39.600 604.050 40.050 ;
        RECT 667.950 39.600 670.050 40.050 ;
        RECT 601.950 38.400 670.050 39.600 ;
        RECT 601.950 37.950 604.050 38.400 ;
        RECT 667.950 37.950 670.050 38.400 ;
        RECT 70.950 36.600 73.050 37.050 ;
        RECT 85.950 36.600 88.050 37.050 ;
        RECT 70.950 35.400 88.050 36.600 ;
        RECT 70.950 34.950 73.050 35.400 ;
        RECT 85.950 34.950 88.050 35.400 ;
        RECT 694.950 36.600 697.050 37.050 ;
        RECT 727.950 36.600 730.050 37.050 ;
        RECT 694.950 35.400 730.050 36.600 ;
        RECT 694.950 34.950 697.050 35.400 ;
        RECT 727.950 34.950 730.050 35.400 ;
        RECT 778.950 36.600 781.050 37.050 ;
        RECT 802.950 36.600 805.050 37.050 ;
        RECT 778.950 35.400 805.050 36.600 ;
        RECT 778.950 34.950 781.050 35.400 ;
        RECT 802.950 34.950 805.050 35.400 ;
        RECT 76.950 33.600 79.050 34.050 ;
        RECT 124.950 33.600 127.050 34.050 ;
        RECT 136.950 33.600 139.050 34.050 ;
        RECT 151.950 33.600 154.050 34.050 ;
        RECT 76.950 32.400 154.050 33.600 ;
        RECT 76.950 31.950 79.050 32.400 ;
        RECT 124.950 31.950 127.050 32.400 ;
        RECT 136.950 31.950 139.050 32.400 ;
        RECT 151.950 31.950 154.050 32.400 ;
        RECT 688.950 33.600 691.050 34.050 ;
        RECT 703.950 33.600 706.050 34.050 ;
        RECT 742.950 33.600 745.050 34.050 ;
        RECT 796.950 33.600 799.050 34.050 ;
        RECT 688.950 32.400 799.050 33.600 ;
        RECT 688.950 31.950 691.050 32.400 ;
        RECT 703.950 31.950 706.050 32.400 ;
        RECT 742.950 31.950 745.050 32.400 ;
        RECT 796.950 31.950 799.050 32.400 ;
        RECT 61.950 30.600 64.050 31.050 ;
        RECT 82.950 30.600 85.050 31.050 ;
        RECT 100.950 30.600 103.050 31.050 ;
        RECT 61.950 29.400 103.050 30.600 ;
        RECT 61.950 28.950 64.050 29.400 ;
        RECT 82.950 28.950 85.050 29.400 ;
        RECT 100.950 28.950 103.050 29.400 ;
        RECT 127.950 30.600 130.050 31.050 ;
        RECT 169.950 30.600 172.050 31.050 ;
        RECT 127.950 29.400 172.050 30.600 ;
        RECT 127.950 28.950 130.050 29.400 ;
        RECT 169.950 28.950 172.050 29.400 ;
        RECT 238.950 30.600 241.050 31.050 ;
        RECT 325.950 30.600 328.050 31.050 ;
        RECT 238.950 29.400 328.050 30.600 ;
        RECT 238.950 28.950 241.050 29.400 ;
        RECT 325.950 28.950 328.050 29.400 ;
        RECT 376.950 30.600 379.050 31.050 ;
        RECT 406.950 30.600 409.050 31.050 ;
        RECT 376.950 29.400 409.050 30.600 ;
        RECT 376.950 28.950 379.050 29.400 ;
        RECT 406.950 28.950 409.050 29.400 ;
        RECT 496.950 30.600 499.050 31.050 ;
        RECT 505.950 30.600 508.050 31.050 ;
        RECT 532.950 30.600 535.050 31.050 ;
        RECT 496.950 29.400 535.050 30.600 ;
        RECT 496.950 28.950 499.050 29.400 ;
        RECT 505.950 28.950 508.050 29.400 ;
        RECT 532.950 28.950 535.050 29.400 ;
        RECT 607.950 30.600 610.050 31.050 ;
        RECT 619.950 30.600 622.050 31.050 ;
        RECT 649.950 30.600 652.050 31.050 ;
        RECT 748.950 30.600 751.050 31.050 ;
        RECT 763.950 30.600 766.050 31.050 ;
        RECT 607.950 29.400 751.050 30.600 ;
        RECT 607.950 28.950 610.050 29.400 ;
        RECT 619.950 28.950 622.050 29.400 ;
        RECT 649.950 28.950 652.050 29.400 ;
        RECT 748.950 28.950 751.050 29.400 ;
        RECT 752.400 29.400 766.050 30.600 ;
        RECT 22.950 27.600 25.050 28.050 ;
        RECT 31.950 27.600 34.050 28.050 ;
        RECT 79.950 27.600 82.050 28.050 ;
        RECT 22.950 26.400 82.050 27.600 ;
        RECT 22.950 25.950 25.050 26.400 ;
        RECT 31.950 25.950 34.050 26.400 ;
        RECT 79.950 25.950 82.050 26.400 ;
        RECT 85.950 27.600 88.050 28.050 ;
        RECT 94.950 27.600 97.050 28.050 ;
        RECT 130.950 27.600 133.050 28.050 ;
        RECT 85.950 26.400 133.050 27.600 ;
        RECT 85.950 25.950 88.050 26.400 ;
        RECT 94.950 25.950 97.050 26.400 ;
        RECT 130.950 25.950 133.050 26.400 ;
        RECT 133.950 27.600 136.050 28.050 ;
        RECT 175.950 27.600 178.050 28.050 ;
        RECT 133.950 26.400 178.050 27.600 ;
        RECT 133.950 25.950 136.050 26.400 ;
        RECT 175.950 25.950 178.050 26.400 ;
        RECT 184.950 27.600 187.050 28.050 ;
        RECT 196.950 27.600 199.050 28.050 ;
        RECT 184.950 26.400 199.050 27.600 ;
        RECT 184.950 25.950 187.050 26.400 ;
        RECT 196.950 25.950 199.050 26.400 ;
        RECT 199.950 27.600 202.050 28.050 ;
        RECT 214.950 27.600 217.050 28.050 ;
        RECT 199.950 26.400 217.050 27.600 ;
        RECT 199.950 25.950 202.050 26.400 ;
        RECT 214.950 25.950 217.050 26.400 ;
        RECT 259.950 27.600 262.050 28.050 ;
        RECT 283.950 27.600 286.050 28.050 ;
        RECT 259.950 26.400 286.050 27.600 ;
        RECT 259.950 25.950 262.050 26.400 ;
        RECT 283.950 25.950 286.050 26.400 ;
        RECT 325.950 27.600 328.050 28.050 ;
        RECT 337.950 27.600 340.050 28.050 ;
        RECT 325.950 26.400 340.050 27.600 ;
        RECT 325.950 25.950 328.050 26.400 ;
        RECT 337.950 25.950 340.050 26.400 ;
        RECT 397.950 27.600 400.050 28.050 ;
        RECT 454.950 27.600 457.050 28.050 ;
        RECT 397.950 26.400 457.050 27.600 ;
        RECT 397.950 25.950 400.050 26.400 ;
        RECT 454.950 25.950 457.050 26.400 ;
        RECT 478.950 27.600 481.050 28.050 ;
        RECT 532.950 27.600 535.050 28.050 ;
        RECT 559.950 27.600 562.050 28.050 ;
        RECT 478.950 26.400 562.050 27.600 ;
        RECT 478.950 25.950 481.050 26.400 ;
        RECT 532.950 25.950 535.050 26.400 ;
        RECT 559.950 25.950 562.050 26.400 ;
        RECT 712.950 27.600 715.050 28.050 ;
        RECT 752.400 27.600 753.600 29.400 ;
        RECT 763.950 28.950 766.050 29.400 ;
        RECT 781.950 30.600 784.050 31.050 ;
        RECT 799.950 30.600 802.050 31.050 ;
        RECT 781.950 29.400 802.050 30.600 ;
        RECT 781.950 28.950 784.050 29.400 ;
        RECT 799.950 28.950 802.050 29.400 ;
        RECT 712.950 26.400 753.600 27.600 ;
        RECT 754.950 27.600 757.050 28.050 ;
        RECT 760.950 27.600 763.050 28.050 ;
        RECT 817.950 27.600 820.050 28.050 ;
        RECT 754.950 26.400 820.050 27.600 ;
        RECT 712.950 25.950 715.050 26.400 ;
        RECT 754.950 25.950 757.050 26.400 ;
        RECT 760.950 25.950 763.050 26.400 ;
        RECT 817.950 25.950 820.050 26.400 ;
        RECT 841.950 27.600 844.050 28.050 ;
        RECT 850.950 27.600 853.050 28.050 ;
        RECT 859.950 27.600 862.050 28.050 ;
        RECT 841.950 26.400 862.050 27.600 ;
        RECT 841.950 25.950 844.050 26.400 ;
        RECT 850.950 25.950 853.050 26.400 ;
        RECT 859.950 25.950 862.050 26.400 ;
        RECT 13.950 24.600 16.050 25.050 ;
        RECT 25.950 24.600 28.050 25.050 ;
        RECT 142.950 24.600 145.050 25.050 ;
        RECT 13.950 23.400 28.050 24.600 ;
        RECT 13.950 22.950 16.050 23.400 ;
        RECT 25.950 22.950 28.050 23.400 ;
        RECT 98.400 23.400 145.050 24.600 ;
        RECT 98.400 22.050 99.600 23.400 ;
        RECT 142.950 22.950 145.050 23.400 ;
        RECT 190.950 24.600 193.050 25.050 ;
        RECT 193.950 24.600 196.050 25.050 ;
        RECT 211.950 24.600 214.050 25.050 ;
        RECT 190.950 23.400 214.050 24.600 ;
        RECT 190.950 22.950 193.050 23.400 ;
        RECT 193.950 22.950 196.050 23.400 ;
        RECT 211.950 22.950 214.050 23.400 ;
        RECT 253.950 24.600 256.050 25.050 ;
        RECT 268.950 24.600 271.050 25.050 ;
        RECT 286.950 24.600 289.050 25.050 ;
        RECT 253.950 23.400 289.050 24.600 ;
        RECT 253.950 22.950 256.050 23.400 ;
        RECT 268.950 22.950 271.050 23.400 ;
        RECT 286.950 22.950 289.050 23.400 ;
        RECT 316.950 24.600 319.050 25.050 ;
        RECT 322.950 24.600 325.050 25.050 ;
        RECT 349.950 24.600 352.050 25.050 ;
        RECT 367.950 24.600 370.050 25.050 ;
        RECT 391.950 24.600 394.050 25.050 ;
        RECT 436.950 24.600 439.050 25.050 ;
        RECT 511.950 24.600 514.050 25.050 ;
        RECT 316.950 23.400 370.050 24.600 ;
        RECT 316.950 22.950 319.050 23.400 ;
        RECT 322.950 22.950 325.050 23.400 ;
        RECT 349.950 22.950 352.050 23.400 ;
        RECT 367.950 22.950 370.050 23.400 ;
        RECT 371.400 23.400 394.050 24.600 ;
        RECT 16.950 21.600 19.050 22.050 ;
        RECT 14.400 20.400 19.050 21.600 ;
        RECT 10.950 18.600 13.050 19.050 ;
        RECT 14.400 18.600 15.600 20.400 ;
        RECT 16.950 19.950 19.050 20.400 ;
        RECT 19.950 21.600 22.050 22.050 ;
        RECT 28.950 21.600 31.050 22.050 ;
        RECT 19.950 20.400 31.050 21.600 ;
        RECT 19.950 19.950 22.050 20.400 ;
        RECT 28.950 19.950 31.050 20.400 ;
        RECT 58.950 21.600 61.050 22.050 ;
        RECT 70.950 21.600 73.050 22.050 ;
        RECT 58.950 20.400 73.050 21.600 ;
        RECT 58.950 19.950 61.050 20.400 ;
        RECT 70.950 19.950 73.050 20.400 ;
        RECT 82.950 21.600 85.050 22.050 ;
        RECT 97.950 21.600 100.050 22.050 ;
        RECT 82.950 20.400 100.050 21.600 ;
        RECT 82.950 19.950 85.050 20.400 ;
        RECT 97.950 19.950 100.050 20.400 ;
        RECT 103.950 21.600 106.050 22.050 ;
        RECT 124.950 21.600 127.050 22.050 ;
        RECT 103.950 20.400 127.050 21.600 ;
        RECT 103.950 19.950 106.050 20.400 ;
        RECT 124.950 19.950 127.050 20.400 ;
        RECT 130.950 21.600 133.050 22.050 ;
        RECT 178.950 21.600 181.050 22.050 ;
        RECT 184.950 21.600 187.050 22.050 ;
        RECT 130.950 20.400 187.050 21.600 ;
        RECT 130.950 19.950 133.050 20.400 ;
        RECT 178.950 19.950 181.050 20.400 ;
        RECT 184.950 19.950 187.050 20.400 ;
        RECT 235.950 21.600 238.050 22.050 ;
        RECT 250.950 21.600 253.050 22.050 ;
        RECT 235.950 20.400 253.050 21.600 ;
        RECT 235.950 19.950 238.050 20.400 ;
        RECT 250.950 19.950 253.050 20.400 ;
        RECT 256.950 21.600 259.050 22.050 ;
        RECT 262.950 21.600 265.050 22.050 ;
        RECT 256.950 20.400 265.050 21.600 ;
        RECT 256.950 19.950 259.050 20.400 ;
        RECT 262.950 19.950 265.050 20.400 ;
        RECT 292.950 21.600 295.050 22.050 ;
        RECT 371.400 21.600 372.600 23.400 ;
        RECT 391.950 22.950 394.050 23.400 ;
        RECT 395.400 23.400 439.050 24.600 ;
        RECT 395.400 22.050 396.600 23.400 ;
        RECT 436.950 22.950 439.050 23.400 ;
        RECT 440.400 23.400 514.050 24.600 ;
        RECT 292.950 20.400 372.600 21.600 ;
        RECT 292.950 19.950 295.050 20.400 ;
        RECT 394.950 19.950 397.050 22.050 ;
        RECT 400.950 21.600 403.050 22.050 ;
        RECT 406.950 21.600 409.050 22.050 ;
        RECT 400.950 20.400 409.050 21.600 ;
        RECT 400.950 19.950 403.050 20.400 ;
        RECT 406.950 19.950 409.050 20.400 ;
        RECT 424.950 21.600 427.050 22.050 ;
        RECT 440.400 21.600 441.600 23.400 ;
        RECT 511.950 22.950 514.050 23.400 ;
        RECT 577.950 24.600 580.050 25.050 ;
        RECT 610.950 24.600 613.050 25.050 ;
        RECT 577.950 23.400 613.050 24.600 ;
        RECT 577.950 22.950 580.050 23.400 ;
        RECT 610.950 22.950 613.050 23.400 ;
        RECT 613.950 24.600 616.050 25.050 ;
        RECT 616.950 24.600 619.050 25.050 ;
        RECT 643.950 24.600 646.050 25.050 ;
        RECT 706.950 24.600 709.050 25.050 ;
        RECT 613.950 23.400 709.050 24.600 ;
        RECT 613.950 22.950 616.050 23.400 ;
        RECT 616.950 22.950 619.050 23.400 ;
        RECT 643.950 22.950 646.050 23.400 ;
        RECT 706.950 22.950 709.050 23.400 ;
        RECT 730.950 24.600 733.050 25.050 ;
        RECT 745.950 24.600 748.050 25.050 ;
        RECT 730.950 23.400 748.050 24.600 ;
        RECT 730.950 22.950 733.050 23.400 ;
        RECT 745.950 22.950 748.050 23.400 ;
        RECT 751.950 24.600 754.050 25.050 ;
        RECT 766.950 24.600 769.050 25.050 ;
        RECT 784.950 24.600 787.050 25.050 ;
        RECT 793.950 24.600 796.050 25.050 ;
        RECT 751.950 23.400 796.050 24.600 ;
        RECT 751.950 22.950 754.050 23.400 ;
        RECT 766.950 22.950 769.050 23.400 ;
        RECT 784.950 22.950 787.050 23.400 ;
        RECT 793.950 22.950 796.050 23.400 ;
        RECT 424.950 20.400 441.600 21.600 ;
        RECT 424.950 19.950 427.050 20.400 ;
        RECT 440.400 19.050 441.600 20.400 ;
        RECT 457.950 21.600 460.050 22.050 ;
        RECT 475.950 21.600 478.050 22.050 ;
        RECT 457.950 20.400 478.050 21.600 ;
        RECT 457.950 19.950 460.050 20.400 ;
        RECT 475.950 19.950 478.050 20.400 ;
        RECT 481.950 21.600 484.050 22.050 ;
        RECT 493.950 21.600 496.050 22.050 ;
        RECT 481.950 20.400 496.050 21.600 ;
        RECT 481.950 19.950 484.050 20.400 ;
        RECT 493.950 19.950 496.050 20.400 ;
        RECT 499.950 21.600 502.050 22.050 ;
        RECT 508.950 21.600 511.050 22.050 ;
        RECT 499.950 20.400 511.050 21.600 ;
        RECT 499.950 19.950 502.050 20.400 ;
        RECT 508.950 19.950 511.050 20.400 ;
        RECT 514.950 21.600 517.050 22.050 ;
        RECT 529.950 21.600 532.050 22.050 ;
        RECT 601.950 21.600 604.050 22.050 ;
        RECT 514.950 20.400 532.050 21.600 ;
        RECT 514.950 19.950 517.050 20.400 ;
        RECT 529.950 19.950 532.050 20.400 ;
        RECT 551.400 20.400 604.050 21.600 ;
        RECT 551.400 19.050 552.600 20.400 ;
        RECT 601.950 19.950 604.050 20.400 ;
        RECT 667.950 21.600 670.050 22.050 ;
        RECT 682.950 21.600 685.050 22.050 ;
        RECT 691.950 21.600 694.050 22.050 ;
        RECT 724.950 21.600 727.050 22.050 ;
        RECT 667.950 20.400 690.600 21.600 ;
        RECT 667.950 19.950 670.050 20.400 ;
        RECT 682.950 19.950 685.050 20.400 ;
        RECT 10.950 17.400 15.600 18.600 ;
        RECT 16.950 18.600 19.050 19.050 ;
        RECT 22.950 18.600 25.050 19.050 ;
        RECT 16.950 17.400 25.050 18.600 ;
        RECT 10.950 16.950 13.050 17.400 ;
        RECT 16.950 16.950 19.050 17.400 ;
        RECT 22.950 16.950 25.050 17.400 ;
        RECT 25.950 18.600 28.050 19.050 ;
        RECT 34.950 18.600 37.050 19.050 ;
        RECT 25.950 17.400 37.050 18.600 ;
        RECT 25.950 16.950 28.050 17.400 ;
        RECT 34.950 16.950 37.050 17.400 ;
        RECT 124.950 18.600 127.050 19.050 ;
        RECT 133.950 18.600 136.050 19.050 ;
        RECT 139.950 18.600 142.050 19.050 ;
        RECT 124.950 17.400 142.050 18.600 ;
        RECT 124.950 16.950 127.050 17.400 ;
        RECT 133.950 16.950 136.050 17.400 ;
        RECT 139.950 16.950 142.050 17.400 ;
        RECT 142.950 18.600 145.050 19.050 ;
        RECT 154.950 18.600 157.050 19.050 ;
        RECT 223.950 18.600 226.050 19.050 ;
        RECT 142.950 17.400 226.050 18.600 ;
        RECT 142.950 16.950 145.050 17.400 ;
        RECT 154.950 16.950 157.050 17.400 ;
        RECT 223.950 16.950 226.050 17.400 ;
        RECT 289.950 16.950 292.050 19.050 ;
        RECT 295.950 18.600 298.050 19.050 ;
        RECT 310.950 18.600 313.050 19.050 ;
        RECT 295.950 17.400 313.050 18.600 ;
        RECT 295.950 16.950 298.050 17.400 ;
        RECT 310.950 16.950 313.050 17.400 ;
        RECT 319.950 18.600 322.050 19.050 ;
        RECT 358.950 18.600 361.050 19.050 ;
        RECT 370.950 18.600 373.050 19.050 ;
        RECT 319.950 17.400 373.050 18.600 ;
        RECT 319.950 16.950 322.050 17.400 ;
        RECT 358.950 16.950 361.050 17.400 ;
        RECT 370.950 16.950 373.050 17.400 ;
        RECT 439.950 16.950 442.050 19.050 ;
        RECT 448.950 18.600 451.050 19.050 ;
        RECT 460.950 18.600 463.050 19.050 ;
        RECT 448.950 17.400 463.050 18.600 ;
        RECT 448.950 16.950 451.050 17.400 ;
        RECT 460.950 16.950 463.050 17.400 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 598.950 18.600 601.050 19.050 ;
        RECT 613.950 18.600 616.050 19.050 ;
        RECT 598.950 17.400 616.050 18.600 ;
        RECT 598.950 16.950 601.050 17.400 ;
        RECT 613.950 16.950 616.050 17.400 ;
        RECT 658.950 18.600 661.050 19.050 ;
        RECT 676.950 18.600 679.050 19.050 ;
        RECT 658.950 17.400 679.050 18.600 ;
        RECT 658.950 16.950 661.050 17.400 ;
        RECT 676.950 16.950 679.050 17.400 ;
        RECT 685.950 16.950 688.050 19.050 ;
        RECT 689.400 18.600 690.600 20.400 ;
        RECT 691.950 20.400 727.050 21.600 ;
        RECT 691.950 19.950 694.050 20.400 ;
        RECT 724.950 19.950 727.050 20.400 ;
        RECT 748.950 21.600 751.050 22.050 ;
        RECT 754.950 21.600 757.050 22.050 ;
        RECT 784.950 21.600 787.050 22.050 ;
        RECT 748.950 20.400 757.050 21.600 ;
        RECT 748.950 19.950 751.050 20.400 ;
        RECT 754.950 19.950 757.050 20.400 ;
        RECT 758.400 20.400 787.050 21.600 ;
        RECT 758.400 18.600 759.600 20.400 ;
        RECT 784.950 19.950 787.050 20.400 ;
        RECT 802.950 21.600 805.050 22.050 ;
        RECT 823.950 21.600 826.050 22.050 ;
        RECT 802.950 20.400 826.050 21.600 ;
        RECT 802.950 19.950 805.050 20.400 ;
        RECT 823.950 19.950 826.050 20.400 ;
        RECT 838.950 21.600 841.050 22.050 ;
        RECT 847.950 21.600 850.050 22.050 ;
        RECT 838.950 20.400 850.050 21.600 ;
        RECT 838.950 19.950 841.050 20.400 ;
        RECT 847.950 19.950 850.050 20.400 ;
        RECT 689.400 17.400 759.600 18.600 ;
        RECT 787.950 18.600 790.050 19.050 ;
        RECT 805.950 18.600 808.050 19.050 ;
        RECT 787.950 17.400 808.050 18.600 ;
        RECT 787.950 16.950 790.050 17.400 ;
        RECT 805.950 16.950 808.050 17.400 ;
        RECT 814.950 18.600 817.050 19.050 ;
        RECT 850.950 18.600 853.050 19.050 ;
        RECT 814.950 17.400 853.050 18.600 ;
        RECT 814.950 16.950 817.050 17.400 ;
        RECT 850.950 16.950 853.050 17.400 ;
        RECT 28.950 15.600 31.050 16.050 ;
        RECT 118.950 15.600 121.050 16.050 ;
        RECT 28.950 14.400 121.050 15.600 ;
        RECT 28.950 13.950 31.050 14.400 ;
        RECT 118.950 13.950 121.050 14.400 ;
        RECT 277.950 15.600 280.050 16.050 ;
        RECT 290.400 15.600 291.600 16.950 ;
        RECT 313.950 15.600 316.050 16.050 ;
        RECT 277.950 14.400 316.050 15.600 ;
        RECT 277.950 13.950 280.050 14.400 ;
        RECT 313.950 13.950 316.050 14.400 ;
        RECT 415.950 15.600 418.050 16.050 ;
        RECT 433.950 15.600 436.050 16.050 ;
        RECT 472.950 15.600 475.050 16.050 ;
        RECT 415.950 14.400 475.050 15.600 ;
        RECT 415.950 13.950 418.050 14.400 ;
        RECT 433.950 13.950 436.050 14.400 ;
        RECT 472.950 13.950 475.050 14.400 ;
        RECT 544.950 15.600 547.050 16.050 ;
        RECT 679.950 15.600 682.050 16.050 ;
        RECT 544.950 14.400 682.050 15.600 ;
        RECT 686.400 15.600 687.600 16.950 ;
        RECT 694.950 15.600 697.050 16.050 ;
        RECT 686.400 14.400 697.050 15.600 ;
        RECT 544.950 13.950 547.050 14.400 ;
        RECT 679.950 13.950 682.050 14.400 ;
        RECT 694.950 13.950 697.050 14.400 ;
  END
END ALU8_Mult
END LIBRARY

