magic
tech scmos
magscale 1 2
timestamp 1728292262
<< metal1 >>
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 1167 4697 1213 4703
rect 2507 4637 2533 4643
rect 5142 4578 5202 4818
rect 5110 4562 5202 4578
rect 1157 4477 1173 4483
rect 1157 4427 1163 4477
rect 1417 4477 1433 4483
rect 1417 4443 1423 4477
rect 1407 4437 1423 4443
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 867 4217 923 4223
rect 917 4183 923 4217
rect 917 4177 953 4183
rect 1237 4163 1243 4233
rect 1927 4197 1943 4203
rect 1937 4167 1943 4197
rect 4517 4183 4523 4213
rect 4517 4177 4533 4183
rect 1237 4157 1253 4163
rect 5142 4098 5202 4562
rect 5110 4082 5202 4098
rect 2287 3997 2303 4003
rect 2297 3963 2303 3997
rect 2297 3957 2313 3963
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 4067 3777 4083 3783
rect 817 3683 823 3733
rect 2757 3707 2763 3733
rect 817 3677 833 3683
rect 1387 3677 1413 3683
rect 1687 3677 1713 3683
rect 4077 3667 4083 3777
rect 4407 3757 4423 3763
rect 4337 3683 4343 3713
rect 4337 3677 4353 3683
rect 4417 3683 4423 3757
rect 4717 3703 4723 3773
rect 4707 3697 4723 3703
rect 4417 3677 4433 3683
rect 5142 3618 5202 4082
rect 5110 3602 5202 3618
rect 417 3467 423 3513
rect 857 3483 863 3533
rect 857 3477 873 3483
rect 2177 3463 2183 3553
rect 2837 3537 2853 3543
rect 2837 3467 2843 3537
rect 3537 3537 3553 3543
rect 2177 3457 2193 3463
rect 3537 3443 3543 3537
rect 3527 3437 3543 3443
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 397 3223 403 3293
rect 367 3217 403 3223
rect 1837 3203 1843 3293
rect 3847 3277 3863 3283
rect 1837 3197 1873 3203
rect 3857 3203 3863 3277
rect 3997 3277 4013 3283
rect 3857 3197 3873 3203
rect 3997 3203 4003 3277
rect 4067 3277 4083 3283
rect 3987 3197 4003 3203
rect 4077 3203 4083 3277
rect 4537 3277 4553 3283
rect 4067 3197 4083 3203
rect 4537 3203 4543 3277
rect 4617 3237 4633 3243
rect 4617 3207 4623 3237
rect 4527 3197 4543 3203
rect 4817 3203 4823 3273
rect 4817 3197 4833 3203
rect 4897 3203 4903 3233
rect 4887 3197 4903 3203
rect 5142 3138 5202 3602
rect 5110 3122 5202 3138
rect 4497 3077 4513 3083
rect 3647 3037 3673 3043
rect 4497 2987 4503 3077
rect 4597 3017 4613 3023
rect 4597 2963 4603 3017
rect 4877 2983 4883 3053
rect 4867 2977 4883 2983
rect 4587 2957 4603 2963
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 4107 2817 4123 2823
rect 2577 2723 2583 2813
rect 4117 2747 4123 2817
rect 2577 2717 2613 2723
rect 4317 2723 4323 2773
rect 4317 2717 4333 2723
rect 5142 2658 5202 3122
rect 5110 2642 5202 2658
rect 4657 2597 4673 2603
rect 187 2577 203 2583
rect 197 2503 203 2577
rect 4337 2557 4353 2563
rect 4337 2547 4343 2557
rect 4657 2523 4663 2597
rect 4727 2557 4763 2563
rect 4627 2517 4663 2523
rect 197 2497 213 2503
rect 4757 2483 4763 2557
rect 5007 2557 5053 2563
rect 4747 2477 4763 2483
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 3167 2317 3183 2323
rect 3037 2297 3053 2303
rect 3037 2243 3043 2297
rect 3177 2267 3183 2317
rect 3697 2267 3703 2333
rect 3907 2297 3923 2303
rect 3027 2237 3043 2243
rect 3917 2243 3923 2297
rect 4427 2297 4463 2303
rect 4457 2247 4463 2297
rect 3917 2237 3963 2243
rect 3957 2223 3963 2237
rect 3957 2217 3973 2223
rect 4687 2217 4713 2223
rect 5142 2178 5202 2642
rect 5110 2162 5202 2178
rect 3097 2097 3113 2103
rect 3097 2023 3103 2097
rect 3877 2097 3893 2103
rect 3877 2027 3883 2097
rect 4087 2077 4123 2083
rect 4117 2047 4123 2077
rect 3097 2017 3113 2023
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 2287 1857 2303 1863
rect 2297 1783 2303 1857
rect 4867 1857 4883 1863
rect 2367 1837 2383 1843
rect 2267 1777 2303 1783
rect 2377 1763 2383 1837
rect 3517 1783 3523 1833
rect 4437 1817 4453 1823
rect 3507 1777 3523 1783
rect 4437 1783 4443 1817
rect 4427 1777 4443 1783
rect 2367 1757 2383 1763
rect 3107 1757 3153 1763
rect 4617 1747 4623 1833
rect 4877 1743 4883 1857
rect 4877 1737 4893 1743
rect 5142 1698 5202 2162
rect 5110 1682 5202 1698
rect 217 1547 223 1593
rect 1177 1563 1183 1633
rect 3307 1617 3323 1623
rect 1167 1557 1183 1563
rect 3317 1543 3323 1617
rect 3887 1617 3903 1623
rect 3677 1597 3713 1603
rect 3677 1547 3683 1597
rect 3787 1597 3823 1603
rect 3317 1537 3333 1543
rect 3797 1507 3803 1573
rect 3817 1543 3823 1597
rect 3897 1587 3903 1617
rect 4567 1617 4603 1623
rect 3817 1537 3833 1543
rect 4597 1523 4603 1617
rect 4777 1597 4813 1603
rect 4777 1547 4783 1597
rect 4907 1597 4933 1603
rect 4597 1517 4613 1523
rect 4877 1523 4883 1533
rect 4997 1527 5003 1593
rect 4877 1517 4893 1523
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 17 1303 23 1373
rect 2157 1357 2173 1363
rect 907 1337 923 1343
rect 17 1297 33 1303
rect 917 1287 923 1337
rect 1117 1303 1123 1353
rect 1777 1343 1783 1353
rect 1747 1337 1783 1343
rect 2157 1323 2163 1357
rect 2147 1317 2163 1323
rect 2437 1307 2443 1353
rect 2457 1307 2463 1373
rect 2687 1337 2743 1343
rect 1087 1297 1123 1303
rect 2557 1283 2563 1333
rect 2737 1287 2743 1337
rect 2547 1277 2563 1283
rect 2817 1283 2823 1393
rect 3287 1377 3303 1383
rect 3297 1307 3303 1377
rect 3637 1377 3673 1383
rect 3537 1303 3543 1333
rect 3637 1307 3643 1377
rect 4817 1377 4833 1383
rect 3957 1357 3973 1363
rect 3957 1343 3963 1357
rect 4217 1357 4233 1363
rect 3937 1337 3963 1343
rect 3537 1297 3573 1303
rect 2807 1277 2823 1283
rect 3937 1283 3943 1337
rect 4217 1287 4223 1357
rect 4817 1303 4823 1377
rect 4807 1297 4823 1303
rect 3927 1277 3943 1283
rect 5142 1218 5202 1682
rect 5110 1202 5202 1218
rect 1007 1137 1023 1143
rect 1017 1087 1023 1137
rect 3647 1137 3663 1143
rect 2397 1117 2413 1123
rect 2397 1043 2403 1117
rect 3657 1063 3663 1137
rect 3767 1097 3783 1103
rect 3647 1057 3663 1063
rect 2397 1037 2413 1043
rect 3777 1043 3783 1097
rect 3777 1037 3793 1043
rect -62 962 30 978
rect -62 498 -2 962
rect 2207 897 2253 903
rect 3647 897 3663 903
rect 2217 787 2223 873
rect 2897 823 2903 853
rect 2887 817 2903 823
rect 3657 823 3663 897
rect 3647 817 3663 823
rect 5142 738 5202 1202
rect 5110 722 5202 738
rect 4387 657 4403 663
rect 207 637 233 643
rect 2957 637 2973 643
rect 2957 563 2963 637
rect 4397 567 4403 657
rect 2957 557 2973 563
rect -62 482 30 498
rect -62 18 -2 482
rect 17 417 33 423
rect 17 327 23 417
rect 3617 417 3633 423
rect 2577 343 2583 393
rect 2577 337 2613 343
rect 3187 337 3253 343
rect 3617 343 3623 417
rect 3907 397 3923 403
rect 3607 337 3623 343
rect 3917 327 3923 397
rect 5142 258 5202 722
rect 5110 242 5202 258
rect 1747 117 1773 123
rect 4327 97 4353 103
rect -62 2 30 18
rect 5142 2 5202 242
<< m2contact >>
rect 4430 4773 4444 4787
rect 5010 4773 5024 4787
rect 1153 4693 1167 4707
rect 1213 4693 1227 4707
rect 2493 4633 2507 4647
rect 2533 4633 2547 4647
rect 1173 4473 1187 4487
rect 1393 4433 1407 4447
rect 1433 4473 1447 4487
rect 1153 4413 1167 4427
rect 4513 4313 4527 4327
rect 1233 4233 1247 4247
rect 853 4213 867 4227
rect 953 4173 967 4187
rect 4513 4213 4527 4227
rect 1913 4193 1927 4207
rect 4533 4173 4547 4187
rect 1253 4153 1267 4167
rect 1933 4153 1947 4167
rect 2273 3993 2287 4007
rect 2313 3953 2327 3967
rect 4053 3773 4067 3787
rect 813 3733 827 3747
rect 2753 3733 2767 3747
rect 2753 3693 2767 3707
rect 833 3673 847 3687
rect 1373 3673 1387 3687
rect 1413 3673 1427 3687
rect 1673 3673 1687 3687
rect 1713 3673 1727 3687
rect 4713 3773 4727 3787
rect 4393 3753 4407 3767
rect 4333 3713 4347 3727
rect 4353 3673 4367 3687
rect 4693 3693 4707 3707
rect 4433 3673 4447 3687
rect 4073 3653 4087 3667
rect 2173 3553 2187 3567
rect 853 3533 867 3547
rect 413 3513 427 3527
rect 873 3473 887 3487
rect 413 3453 427 3467
rect 2853 3533 2867 3547
rect 2193 3453 2207 3467
rect 2833 3453 2847 3467
rect 3513 3433 3527 3447
rect 3553 3533 3567 3547
rect 393 3293 407 3307
rect 1833 3293 1847 3307
rect 353 3213 367 3227
rect 3833 3273 3847 3287
rect 1873 3193 1887 3207
rect 3873 3193 3887 3207
rect 3973 3193 3987 3207
rect 4013 3273 4027 3287
rect 4053 3273 4067 3287
rect 4053 3193 4067 3207
rect 4513 3193 4527 3207
rect 4553 3273 4567 3287
rect 4813 3273 4827 3287
rect 4633 3233 4647 3247
rect 4613 3193 4627 3207
rect 4893 3233 4907 3247
rect 4833 3193 4847 3207
rect 4873 3193 4887 3207
rect 3633 3033 3647 3047
rect 3673 3033 3687 3047
rect 4513 3073 4527 3087
rect 4873 3053 4887 3067
rect 4493 2973 4507 2987
rect 4573 2953 4587 2967
rect 4613 3013 4627 3027
rect 4853 2973 4867 2987
rect 2573 2813 2587 2827
rect 4093 2813 4107 2827
rect 4313 2773 4327 2787
rect 4113 2733 4127 2747
rect 2613 2713 2627 2727
rect 4333 2713 4347 2727
rect 173 2573 187 2587
rect 4353 2553 4367 2567
rect 4333 2533 4347 2547
rect 4613 2513 4627 2527
rect 4673 2593 4687 2607
rect 4713 2553 4727 2567
rect 213 2493 227 2507
rect 4733 2473 4747 2487
rect 4993 2553 5007 2567
rect 5053 2553 5067 2567
rect 3693 2333 3707 2347
rect 3153 2313 3167 2327
rect 3013 2233 3027 2247
rect 3053 2293 3067 2307
rect 3893 2293 3907 2307
rect 3173 2253 3187 2267
rect 3693 2253 3707 2267
rect 4413 2293 4427 2307
rect 4453 2233 4467 2247
rect 3973 2213 3987 2227
rect 4673 2213 4687 2227
rect 4713 2213 4727 2227
rect 3113 2093 3127 2107
rect 3893 2093 3907 2107
rect 4073 2073 4087 2087
rect 4113 2033 4127 2047
rect 3113 2013 3127 2027
rect 3873 2013 3887 2027
rect 2273 1853 2287 1867
rect 2253 1773 2267 1787
rect 4853 1853 4867 1867
rect 2353 1833 2367 1847
rect 2353 1753 2367 1767
rect 3513 1833 3527 1847
rect 4613 1833 4627 1847
rect 3493 1773 3507 1787
rect 4413 1773 4427 1787
rect 4453 1813 4467 1827
rect 3093 1753 3107 1767
rect 3153 1753 3167 1767
rect 4613 1733 4627 1747
rect 4893 1733 4907 1747
rect 1173 1633 1187 1647
rect 213 1593 227 1607
rect 1153 1553 1167 1567
rect 3293 1613 3307 1627
rect 213 1533 227 1547
rect 3873 1613 3887 1627
rect 3713 1593 3727 1607
rect 3773 1593 3787 1607
rect 3793 1573 3807 1587
rect 3333 1533 3347 1547
rect 3673 1533 3687 1547
rect 4553 1613 4567 1627
rect 3893 1573 3907 1587
rect 3833 1533 3847 1547
rect 4813 1593 4827 1607
rect 4893 1593 4907 1607
rect 4933 1593 4947 1607
rect 4993 1593 5007 1607
rect 4773 1533 4787 1547
rect 4873 1533 4887 1547
rect 4613 1513 4627 1527
rect 4893 1513 4907 1527
rect 4993 1513 5007 1527
rect 3793 1493 3807 1507
rect 2813 1393 2827 1407
rect 13 1373 27 1387
rect 2453 1373 2467 1387
rect 1113 1353 1127 1367
rect 1773 1353 1787 1367
rect 893 1333 907 1347
rect 33 1293 47 1307
rect 1073 1293 1087 1307
rect 1733 1333 1747 1347
rect 2133 1313 2147 1327
rect 2173 1353 2187 1367
rect 2433 1353 2447 1367
rect 2553 1333 2567 1347
rect 2673 1333 2687 1347
rect 2433 1293 2447 1307
rect 2453 1293 2467 1307
rect 913 1273 927 1287
rect 2533 1273 2547 1287
rect 2733 1273 2747 1287
rect 2793 1273 2807 1287
rect 3273 1373 3287 1387
rect 3533 1333 3547 1347
rect 3293 1293 3307 1307
rect 3673 1373 3687 1387
rect 3973 1353 3987 1367
rect 3573 1293 3587 1307
rect 3633 1293 3647 1307
rect 3913 1273 3927 1287
rect 4233 1353 4247 1367
rect 4793 1293 4807 1307
rect 4833 1373 4847 1387
rect 4213 1273 4227 1287
rect 993 1133 1007 1147
rect 3633 1133 3647 1147
rect 1013 1073 1027 1087
rect 2413 1113 2427 1127
rect 3633 1053 3647 1067
rect 3753 1093 3767 1107
rect 2413 1033 2427 1047
rect 3793 1033 3807 1047
rect 2193 893 2207 907
rect 2253 893 2267 907
rect 3633 893 3647 907
rect 2213 873 2227 887
rect 2893 853 2907 867
rect 2873 813 2887 827
rect 3633 813 3647 827
rect 2213 773 2227 787
rect 4373 653 4387 667
rect 193 633 207 647
rect 233 633 247 647
rect 2973 633 2987 647
rect 2973 553 2987 567
rect 4393 553 4407 567
rect 33 413 47 427
rect 2573 393 2587 407
rect 2613 333 2627 347
rect 3173 333 3187 347
rect 3253 333 3267 347
rect 3593 333 3607 347
rect 3633 413 3647 427
rect 3893 393 3907 407
rect 13 313 27 327
rect 3913 313 3927 327
rect 1733 113 1747 127
rect 1773 113 1787 127
rect 4313 93 4327 107
rect 4353 93 4367 107
<< metal2 >>
rect 2276 4856 2303 4863
rect 56 4676 83 4683
rect 116 4676 143 4683
rect 36 4647 43 4663
rect 56 4456 63 4493
rect 76 4487 83 4676
rect 136 4587 143 4676
rect 216 4676 223 4713
rect 176 4667 183 4673
rect 196 4647 203 4663
rect 236 4647 243 4663
rect 316 4643 323 4673
rect 396 4667 403 4683
rect 296 4636 323 4643
rect 336 4587 343 4663
rect 376 4563 383 4663
rect 356 4556 383 4563
rect 36 4427 43 4443
rect 56 4207 63 4413
rect 76 4227 83 4433
rect 96 4427 103 4473
rect 116 4447 123 4493
rect 136 4456 143 4533
rect 196 4476 203 4513
rect 176 4387 183 4463
rect 216 4223 223 4433
rect 256 4227 263 4253
rect 276 4247 283 4453
rect 356 4436 363 4556
rect 376 4456 383 4533
rect 396 4267 403 4653
rect 456 4587 463 4683
rect 616 4676 643 4683
rect 516 4507 523 4663
rect 536 4607 543 4673
rect 636 4667 643 4676
rect 696 4676 703 4753
rect 736 4687 743 4713
rect 647 4656 663 4663
rect 596 4627 603 4643
rect 656 4643 663 4656
rect 716 4647 723 4663
rect 656 4636 673 4643
rect 616 4607 623 4633
rect 476 4443 483 4453
rect 456 4436 483 4443
rect 496 4443 503 4473
rect 576 4447 583 4513
rect 596 4456 603 4533
rect 736 4527 743 4643
rect 776 4627 783 4753
rect 796 4676 823 4683
rect 856 4676 883 4683
rect 796 4607 803 4676
rect 676 4476 683 4513
rect 696 4496 743 4503
rect 736 4447 743 4496
rect 756 4487 763 4593
rect 776 4487 783 4513
rect 796 4476 803 4533
rect 836 4476 843 4493
rect 856 4487 863 4676
rect 996 4676 1003 4713
rect 1336 4696 1363 4703
rect 1396 4696 1423 4703
rect 1036 4656 1063 4663
rect 1016 4647 1023 4653
rect 756 4463 763 4473
rect 756 4456 783 4463
rect 496 4436 523 4443
rect 416 4407 423 4433
rect 196 4216 223 4223
rect 76 4167 83 4183
rect 116 4167 123 4213
rect 196 4187 203 4216
rect 336 4216 363 4223
rect 56 4023 63 4163
rect 36 4016 63 4023
rect 36 3996 43 4016
rect 96 3976 103 4033
rect 136 3927 143 3993
rect 156 3987 163 4183
rect 236 4147 243 4203
rect 276 4027 283 4193
rect 296 3983 303 4193
rect 316 4187 323 4203
rect 356 4027 363 4216
rect 376 4163 383 4213
rect 376 4156 403 4163
rect 156 3967 163 3973
rect 236 3967 243 3983
rect 276 3976 303 3983
rect 336 3963 343 3993
rect 336 3956 363 3963
rect 16 3727 23 3813
rect 36 3747 43 3793
rect 56 3516 63 3753
rect 116 3723 123 3873
rect 416 3787 423 4093
rect 436 4047 443 4413
rect 556 4387 563 4443
rect 756 4427 763 4456
rect 916 4407 923 4453
rect 936 4447 943 4553
rect 496 4216 543 4223
rect 496 4196 503 4216
rect 536 4207 543 4216
rect 436 3976 443 3993
rect 456 3967 463 4013
rect 476 3976 483 3993
rect 116 3716 143 3723
rect 136 3707 143 3716
rect 76 3627 83 3703
rect 156 3687 163 3703
rect 156 3547 163 3673
rect 196 3667 203 3703
rect 256 3567 263 3703
rect 276 3687 283 3723
rect 316 3687 323 3773
rect 356 3716 363 3733
rect 396 3727 403 3753
rect 416 3743 423 3773
rect 416 3736 443 3743
rect 436 3716 443 3736
rect 496 3723 503 3963
rect 516 3767 523 4183
rect 556 4083 563 4253
rect 616 4187 623 4213
rect 636 4167 643 4203
rect 696 4147 703 4183
rect 536 4076 563 4083
rect 536 3907 543 4076
rect 716 4067 723 4233
rect 736 4147 743 4203
rect 816 4183 823 4233
rect 856 4196 863 4213
rect 876 4207 883 4333
rect 896 4196 903 4213
rect 936 4203 943 4253
rect 956 4247 963 4493
rect 976 4487 983 4533
rect 996 4476 1003 4553
rect 1036 4476 1043 4593
rect 1056 4347 1063 4656
rect 1116 4627 1123 4693
rect 1156 4676 1163 4693
rect 1136 4643 1143 4663
rect 1216 4647 1223 4693
rect 1256 4676 1263 4693
rect 1296 4667 1303 4683
rect 1276 4647 1283 4663
rect 1136 4636 1163 4643
rect 1096 4496 1103 4533
rect 1116 4476 1123 4533
rect 1136 4367 1143 4613
rect 1156 4527 1163 4636
rect 1176 4627 1183 4643
rect 1176 4487 1183 4513
rect 1236 4476 1243 4493
rect 1156 4447 1163 4473
rect 1216 4447 1223 4463
rect 1256 4447 1263 4533
rect 1296 4476 1303 4613
rect 1316 4507 1323 4693
rect 1336 4687 1343 4696
rect 1336 4487 1343 4493
rect 1276 4456 1283 4473
rect 1316 4447 1323 4463
rect 1356 4447 1363 4653
rect 1376 4527 1383 4683
rect 1416 4647 1423 4696
rect 1456 4667 1463 4713
rect 1476 4607 1483 4653
rect 1496 4627 1503 4643
rect 1396 4496 1403 4533
rect 1447 4476 1463 4483
rect 1496 4476 1503 4553
rect 1596 4523 1603 4733
rect 1616 4627 1623 4683
rect 1676 4656 1703 4663
rect 1596 4516 1623 4523
rect 1516 4476 1523 4493
rect 1596 4476 1603 4493
rect 936 4196 963 4203
rect 756 4167 763 4183
rect 796 4176 823 4183
rect 596 4016 603 4033
rect 576 3967 583 3983
rect 636 3983 643 4053
rect 776 4016 783 4053
rect 616 3976 643 3983
rect 536 3807 543 3893
rect 596 3847 603 3973
rect 656 3967 663 3983
rect 536 3727 543 3793
rect 596 3727 603 3793
rect 496 3716 523 3723
rect 616 3723 623 3753
rect 616 3716 643 3723
rect 676 3716 683 3973
rect 696 3947 703 3963
rect 736 3927 743 3953
rect 756 3947 763 4013
rect 716 3807 723 3833
rect 756 3827 763 3913
rect 796 3867 803 3983
rect 576 3607 583 3703
rect 616 3687 623 3716
rect 716 3703 723 3793
rect 816 3747 823 4176
rect 916 4167 923 4193
rect 1036 4183 1043 4213
rect 967 4176 983 4183
rect 1016 4176 1043 4183
rect 936 4007 943 4173
rect 1016 4127 1023 4176
rect 836 3996 863 4003
rect 836 3767 843 3996
rect 976 3996 983 4113
rect 836 3747 843 3753
rect 856 3716 863 3733
rect 296 3536 303 3553
rect 96 3516 123 3523
rect 116 3367 123 3516
rect 136 3516 163 3523
rect 136 3307 143 3516
rect 336 3507 343 3533
rect 396 3516 403 3553
rect 427 3516 433 3523
rect 56 3236 63 3253
rect 76 3187 83 3203
rect 96 3047 103 3293
rect 116 3267 123 3273
rect 176 3247 183 3503
rect 216 3447 223 3503
rect 276 3467 283 3503
rect 276 3236 283 3433
rect 196 3187 203 3233
rect 116 3036 123 3073
rect 176 3036 183 3073
rect 216 3043 223 3223
rect 296 3207 303 3493
rect 416 3483 423 3493
rect 496 3487 503 3553
rect 576 3547 583 3593
rect 416 3476 443 3483
rect 316 3256 323 3313
rect 376 3307 383 3473
rect 396 3427 403 3473
rect 416 3447 423 3453
rect 436 3447 443 3476
rect 476 3467 483 3473
rect 416 3327 423 3433
rect 596 3347 603 3653
rect 656 3587 663 3703
rect 696 3696 723 3703
rect 616 3536 673 3543
rect 616 3527 623 3536
rect 676 3516 683 3533
rect 756 3507 763 3703
rect 816 3647 823 3713
rect 836 3687 843 3703
rect 836 3667 843 3673
rect 876 3647 883 3693
rect 916 3663 923 3933
rect 936 3727 943 3813
rect 1016 3787 1023 4113
rect 1056 3976 1063 4203
rect 1076 4147 1083 4183
rect 1116 4147 1123 4183
rect 1136 4087 1143 4273
rect 1156 4247 1163 4413
rect 1356 4267 1363 4433
rect 1396 4407 1403 4433
rect 1416 4387 1423 4473
rect 1476 4447 1483 4463
rect 1536 4407 1543 4463
rect 1227 4236 1233 4243
rect 1236 4216 1263 4223
rect 1296 4216 1323 4223
rect 1156 4127 1163 4173
rect 1176 4147 1183 4183
rect 1216 4167 1223 4183
rect 1236 4167 1243 4216
rect 1316 4207 1323 4216
rect 1256 4027 1263 4153
rect 1276 4147 1283 4203
rect 1376 4196 1383 4253
rect 1416 4207 1423 4233
rect 1456 4227 1463 4373
rect 1496 4216 1503 4233
rect 1316 4167 1323 4193
rect 1336 4187 1343 4193
rect 1096 3996 1123 4003
rect 1156 3996 1183 4003
rect 1096 3967 1103 3996
rect 1176 3983 1183 3996
rect 1176 3976 1203 3983
rect 1036 3847 1043 3963
rect 1076 3947 1083 3963
rect 996 3727 1003 3733
rect 936 3687 943 3713
rect 956 3707 963 3723
rect 976 3667 983 3703
rect 1016 3687 1023 3703
rect 896 3656 923 3663
rect 796 3536 803 3633
rect 856 3547 863 3633
rect 896 3547 903 3656
rect 916 3536 923 3633
rect 836 3516 863 3523
rect 736 3427 743 3483
rect 396 3307 403 3313
rect 396 3243 403 3273
rect 416 3267 423 3293
rect 516 3287 523 3313
rect 456 3267 463 3273
rect 696 3256 703 3293
rect 756 3287 763 3473
rect 776 3467 783 3503
rect 796 3447 803 3473
rect 856 3267 863 3516
rect 876 3507 883 3533
rect 936 3487 943 3653
rect 996 3536 1003 3633
rect 1016 3547 1023 3573
rect 1036 3567 1043 3773
rect 1096 3747 1103 3893
rect 1116 3887 1123 3953
rect 1136 3887 1143 3973
rect 1196 3827 1203 3976
rect 1236 3947 1243 3963
rect 1236 3927 1243 3933
rect 1136 3787 1143 3813
rect 1116 3727 1123 3773
rect 1196 3707 1203 3713
rect 1096 3667 1103 3683
rect 1176 3683 1183 3703
rect 1147 3676 1183 3683
rect 1076 3547 1083 3633
rect 1116 3536 1123 3633
rect 1076 3503 1083 3533
rect 1056 3496 1083 3503
rect 876 3427 883 3473
rect 996 3447 1003 3493
rect 736 3256 763 3263
rect 376 3236 403 3243
rect 316 3183 323 3213
rect 296 3176 323 3183
rect 196 3036 223 3043
rect 236 3036 263 3043
rect 76 2723 83 2813
rect 56 2716 83 2723
rect 116 2707 123 2743
rect 176 2607 183 2873
rect 196 2783 203 3036
rect 256 2867 263 3036
rect 196 2776 223 2783
rect 216 2767 223 2776
rect 276 2763 283 3113
rect 296 2907 303 3176
rect 356 3023 363 3213
rect 376 3067 383 3073
rect 336 3016 363 3023
rect 376 3016 383 3053
rect 436 3027 443 3243
rect 476 3207 483 3243
rect 496 3056 503 3113
rect 416 3007 423 3023
rect 536 3023 543 3193
rect 556 3127 563 3233
rect 576 3207 583 3223
rect 296 2787 303 2893
rect 356 2807 363 2833
rect 436 2807 443 3013
rect 476 2907 483 3023
rect 516 3016 543 3023
rect 516 2827 523 3016
rect 556 2996 563 3113
rect 616 3067 623 3223
rect 636 3167 643 3243
rect 676 3067 683 3253
rect 636 3056 663 3063
rect 536 2807 543 2933
rect 596 2807 603 3003
rect 636 2947 643 3056
rect 716 3047 723 3243
rect 756 3227 763 3256
rect 816 3236 823 3253
rect 896 3236 903 3253
rect 756 3187 763 3213
rect 776 3207 783 3233
rect 836 3187 843 3223
rect 856 3147 863 3233
rect 876 3207 883 3223
rect 876 3087 883 3193
rect 936 3187 943 3243
rect 956 3207 963 3333
rect 996 3283 1003 3433
rect 976 3276 1003 3283
rect 916 3056 923 3133
rect 676 2807 683 3023
rect 716 3003 723 3033
rect 796 3027 803 3053
rect 956 3043 963 3133
rect 976 3067 983 3276
rect 996 3207 1003 3243
rect 1036 3236 1043 3273
rect 996 3167 1003 3193
rect 1016 3127 1023 3223
rect 1076 3123 1083 3373
rect 1116 3287 1123 3493
rect 1176 3327 1183 3653
rect 1216 3523 1223 3753
rect 1236 3687 1243 3853
rect 1256 3736 1263 3873
rect 1276 3847 1283 3873
rect 1296 3823 1303 4153
rect 1336 4087 1343 4173
rect 1356 4147 1363 4183
rect 1396 4127 1403 4183
rect 1436 4127 1443 4183
rect 1316 3967 1323 4073
rect 1396 3996 1403 4053
rect 1416 3996 1423 4113
rect 1456 4027 1463 4213
rect 1476 4167 1483 4183
rect 1276 3816 1303 3823
rect 1276 3767 1283 3816
rect 1296 3736 1303 3793
rect 1316 3707 1323 3773
rect 1196 3516 1223 3523
rect 1196 3467 1203 3516
rect 1236 3387 1243 3503
rect 1276 3496 1283 3693
rect 1296 3287 1303 3693
rect 1336 3687 1343 3703
rect 1376 3687 1383 3703
rect 1316 3447 1323 3633
rect 1356 3567 1363 3683
rect 1396 3667 1403 3953
rect 1436 3947 1443 3983
rect 1476 3803 1483 3973
rect 1516 3927 1523 4233
rect 1536 4227 1543 4253
rect 1536 4167 1543 4183
rect 1556 4147 1563 4413
rect 1616 4307 1623 4516
rect 1636 4407 1643 4493
rect 1676 4483 1683 4656
rect 1756 4647 1763 4693
rect 1776 4676 1803 4683
rect 1856 4676 1863 4713
rect 1916 4683 1923 4813
rect 2296 4727 2303 4856
rect 2436 4827 2443 4863
rect 1896 4676 1923 4683
rect 1776 4667 1783 4676
rect 1656 4476 1683 4483
rect 1656 4427 1663 4476
rect 1696 4456 1703 4493
rect 1716 4467 1723 4633
rect 1816 4567 1823 4643
rect 1916 4607 1923 4676
rect 1936 4567 1943 4663
rect 1976 4627 1983 4663
rect 1996 4627 2003 4713
rect 2056 4676 2063 4713
rect 2016 4656 2043 4663
rect 2016 4563 2023 4656
rect 2116 4643 2123 4653
rect 2116 4636 2143 4643
rect 1996 4556 2023 4563
rect 1996 4547 2003 4556
rect 1576 4216 1583 4293
rect 1656 4247 1663 4413
rect 1676 4407 1683 4443
rect 1756 4407 1763 4493
rect 1776 4427 1783 4443
rect 1816 4427 1823 4443
rect 1836 4387 1843 4513
rect 2016 4487 2023 4533
rect 1616 4227 1623 4233
rect 1696 4196 1703 4233
rect 1756 4207 1763 4353
rect 1796 4267 1803 4353
rect 1796 4196 1803 4253
rect 1576 4007 1583 4173
rect 1556 3976 1563 3993
rect 1516 3867 1523 3913
rect 1476 3796 1503 3803
rect 1476 3736 1483 3773
rect 1496 3703 1503 3796
rect 1516 3787 1523 3853
rect 1536 3747 1543 3953
rect 1576 3927 1583 3963
rect 1556 3716 1563 3833
rect 1596 3747 1603 4113
rect 1616 4107 1623 4173
rect 1676 4147 1683 4183
rect 1636 4003 1643 4093
rect 1696 4067 1703 4153
rect 1716 4147 1723 4183
rect 1736 4127 1743 4183
rect 1616 3996 1643 4003
rect 1676 3996 1683 4053
rect 1616 3967 1623 3996
rect 1716 3983 1723 4013
rect 1696 3976 1723 3983
rect 1616 3883 1623 3953
rect 1636 3903 1643 3953
rect 1656 3927 1663 3973
rect 1716 3907 1723 3976
rect 1636 3896 1663 3903
rect 1616 3876 1643 3883
rect 1616 3716 1623 3773
rect 1636 3747 1643 3876
rect 1656 3716 1663 3896
rect 1736 3887 1743 4033
rect 1756 3967 1763 4153
rect 1776 4147 1783 4183
rect 1816 3967 1823 4183
rect 1836 4147 1843 4233
rect 1856 4227 1863 4253
rect 1916 4207 1923 4413
rect 1956 4387 1963 4443
rect 1836 4007 1843 4053
rect 1876 4003 1883 4203
rect 1936 4183 1943 4233
rect 1976 4196 1983 4293
rect 1996 4187 2003 4433
rect 2036 4367 2043 4633
rect 2076 4567 2083 4633
rect 2076 4456 2083 4473
rect 2096 4467 2103 4593
rect 2116 4456 2123 4513
rect 2136 4507 2143 4636
rect 2176 4627 2183 4673
rect 2196 4667 2203 4713
rect 2236 4667 2243 4693
rect 2136 4447 2143 4493
rect 2236 4476 2243 4653
rect 2276 4627 2283 4693
rect 2296 4676 2303 4713
rect 2356 4696 2383 4703
rect 2336 4667 2343 4673
rect 2376 4647 2383 4696
rect 2276 4476 2283 4533
rect 2316 4476 2323 4493
rect 2216 4447 2223 4473
rect 2056 4407 2063 4443
rect 2156 4423 2163 4443
rect 2156 4416 2183 4423
rect 2076 4227 2083 4413
rect 1936 4176 1963 4183
rect 1916 4047 1923 4173
rect 1856 3996 1883 4003
rect 1756 3947 1763 3953
rect 1476 3696 1503 3703
rect 1427 3676 1443 3683
rect 1336 3516 1343 3533
rect 1376 3516 1383 3573
rect 1116 3263 1123 3273
rect 1116 3256 1143 3263
rect 1136 3247 1143 3256
rect 1196 3236 1223 3243
rect 1096 3227 1103 3233
rect 1116 3207 1123 3223
rect 1056 3116 1083 3123
rect 956 3036 983 3043
rect 716 2996 743 3003
rect 816 2996 823 3033
rect 656 2787 663 2793
rect 316 2776 343 2783
rect 256 2756 283 2763
rect 296 2747 303 2773
rect 236 2727 243 2743
rect 316 2727 323 2776
rect 396 2723 403 2773
rect 456 2747 463 2783
rect 556 2776 583 2783
rect 496 2743 503 2763
rect 476 2736 503 2743
rect 476 2723 483 2736
rect 536 2727 543 2763
rect 576 2727 583 2776
rect 596 2776 623 2783
rect 396 2716 483 2723
rect 596 2707 603 2776
rect 836 2776 863 2783
rect 636 2747 643 2763
rect 716 2707 723 2763
rect 816 2707 823 2763
rect 856 2727 863 2776
rect 896 2743 903 2793
rect 956 2767 963 3013
rect 996 2987 1003 3023
rect 1036 3016 1043 3053
rect 996 2967 1003 2973
rect 1056 2887 1063 3116
rect 1076 2907 1083 3093
rect 1156 3087 1163 3223
rect 1216 3207 1223 3236
rect 1236 3087 1243 3273
rect 1336 3256 1343 3333
rect 1376 3267 1383 3293
rect 1396 3267 1403 3553
rect 1416 3516 1423 3593
rect 1436 3567 1443 3676
rect 1476 3547 1483 3696
rect 1456 3516 1483 3523
rect 1436 3483 1443 3493
rect 1476 3487 1483 3516
rect 1416 3476 1443 3483
rect 1096 3016 1103 3053
rect 1116 3007 1123 3033
rect 1136 2887 1143 2973
rect 1016 2787 1023 2853
rect 1136 2847 1143 2873
rect 1056 2776 1083 2783
rect 1116 2776 1123 2793
rect 1036 2747 1043 2753
rect 876 2727 883 2743
rect 896 2736 943 2743
rect 1016 2727 1023 2743
rect 1056 2727 1063 2776
rect 1136 2743 1143 2813
rect 1156 2807 1163 3003
rect 1176 2947 1183 3053
rect 1256 3036 1263 3223
rect 1296 3167 1303 3193
rect 1196 2987 1203 3033
rect 1296 2927 1303 3013
rect 1356 2983 1363 3233
rect 1396 3187 1403 3213
rect 1416 3087 1423 3476
rect 1476 3427 1483 3433
rect 1436 3047 1443 3153
rect 1476 3107 1483 3413
rect 1496 3387 1503 3673
rect 1516 3516 1523 3573
rect 1536 3536 1543 3593
rect 1556 3567 1563 3673
rect 1576 3587 1583 3703
rect 1556 3516 1563 3553
rect 1596 3547 1603 3693
rect 1636 3667 1643 3703
rect 1676 3687 1683 3703
rect 1696 3667 1703 3833
rect 1716 3747 1723 3873
rect 1856 3847 1863 3996
rect 1896 3987 1903 3993
rect 1916 3956 1923 4033
rect 1936 4007 1943 4153
rect 1936 3976 1943 3993
rect 1956 3987 1963 4176
rect 1976 3976 1983 4013
rect 1996 3996 2003 4133
rect 2016 4067 2023 4203
rect 2096 4183 2103 4293
rect 2076 4176 2103 4183
rect 2076 4043 2083 4176
rect 2136 4147 2143 4163
rect 2156 4107 2163 4313
rect 2176 4247 2183 4416
rect 2196 4387 2203 4433
rect 2216 4216 2243 4223
rect 2196 4167 2203 4203
rect 2236 4163 2243 4216
rect 2256 4196 2263 4293
rect 2296 4167 2303 4433
rect 2316 4407 2323 4433
rect 2336 4243 2343 4633
rect 2396 4623 2403 4733
rect 2476 4687 2483 4753
rect 2636 4703 2643 4863
rect 3176 4827 3183 4863
rect 3216 4856 3263 4863
rect 2616 4696 2643 4703
rect 2556 4676 2563 4693
rect 2416 4643 2423 4663
rect 2416 4636 2463 4643
rect 2396 4616 2423 4623
rect 2356 4487 2363 4513
rect 2376 4476 2383 4593
rect 2416 4487 2423 4616
rect 2456 4456 2463 4636
rect 2496 4607 2503 4633
rect 2516 4607 2523 4673
rect 2536 4647 2543 4663
rect 2496 4443 2503 4493
rect 2536 4487 2543 4613
rect 2576 4587 2583 4663
rect 2616 4647 2623 4696
rect 2616 4496 2623 4593
rect 2476 4436 2503 4443
rect 2516 4476 2533 4483
rect 2436 4287 2443 4433
rect 2416 4247 2423 4273
rect 2336 4236 2363 4243
rect 2316 4196 2323 4213
rect 2336 4167 2343 4183
rect 2236 4156 2263 4163
rect 2176 4107 2183 4153
rect 2056 4036 2083 4043
rect 2056 3996 2063 4036
rect 2096 3996 2123 4003
rect 2116 3987 2123 3996
rect 1756 3736 1763 3833
rect 1736 3683 1743 3723
rect 1727 3676 1743 3683
rect 1616 3567 1623 3653
rect 1756 3643 1763 3693
rect 1776 3667 1783 3773
rect 1796 3703 1803 3733
rect 1836 3727 1843 3833
rect 1796 3696 1823 3703
rect 1756 3636 1783 3643
rect 1576 3536 1593 3543
rect 1576 3516 1583 3536
rect 1536 3467 1543 3493
rect 1596 3487 1603 3503
rect 1556 3236 1563 3473
rect 1596 3447 1603 3473
rect 1636 3467 1643 3503
rect 1676 3467 1683 3553
rect 1716 3496 1723 3513
rect 1756 3483 1763 3513
rect 1696 3467 1703 3483
rect 1736 3476 1763 3483
rect 1636 3447 1643 3453
rect 1496 3107 1503 3223
rect 1576 3187 1583 3223
rect 1616 3203 1623 3393
rect 1636 3227 1643 3253
rect 1616 3196 1643 3203
rect 1387 3036 1403 3043
rect 1396 3016 1403 3036
rect 1456 3036 1463 3053
rect 1496 3043 1503 3073
rect 1496 3036 1523 3043
rect 1416 2983 1423 3003
rect 1436 2987 1443 3013
rect 1516 2987 1523 3036
rect 1576 3036 1603 3043
rect 1616 3036 1623 3053
rect 1356 2976 1423 2983
rect 1296 2827 1303 2913
rect 1156 2747 1163 2763
rect 1116 2736 1143 2743
rect 16 1407 23 2593
rect 296 2587 303 2593
rect 96 2576 123 2583
rect 36 2527 43 2543
rect 116 2523 123 2576
rect 156 2576 173 2583
rect 156 2536 163 2576
rect 196 2523 203 2553
rect 236 2536 243 2573
rect 456 2563 463 2573
rect 436 2556 463 2563
rect 116 2516 143 2523
rect 176 2516 203 2523
rect 116 2287 123 2516
rect 36 2023 43 2233
rect 136 2227 143 2263
rect 156 2127 163 2283
rect 176 2267 183 2516
rect 216 2507 223 2523
rect 416 2483 423 2543
rect 396 2476 423 2483
rect 356 2296 363 2333
rect 76 2096 103 2103
rect 96 2087 103 2096
rect 56 2047 63 2063
rect 36 2016 63 2023
rect 56 1827 63 2016
rect 96 1827 103 2073
rect 136 2056 143 2093
rect 176 1847 183 2033
rect 216 2027 223 2043
rect 236 1987 243 2253
rect 256 2207 263 2263
rect 396 2247 403 2476
rect 456 2427 463 2556
rect 596 2556 603 2573
rect 476 2527 483 2533
rect 516 2487 523 2553
rect 536 2507 543 2543
rect 616 2507 623 2553
rect 636 2547 643 2593
rect 656 2547 663 2573
rect 676 2536 683 2553
rect 776 2536 783 2553
rect 276 2167 283 2243
rect 416 2207 423 2283
rect 256 2056 283 2063
rect 316 2056 323 2073
rect 256 2047 263 2056
rect 356 2043 363 2093
rect 396 2056 403 2153
rect 416 2107 423 2193
rect 436 2167 443 2303
rect 336 2036 363 2043
rect 116 1816 143 1823
rect 176 1816 203 1823
rect 116 1807 123 1816
rect 36 1767 43 1803
rect 96 1767 103 1783
rect 36 1583 43 1733
rect 36 1576 63 1583
rect 76 1567 83 1753
rect 96 1596 103 1753
rect 116 1627 123 1793
rect 136 1583 143 1773
rect 156 1607 163 1773
rect 196 1767 203 1816
rect 116 1576 143 1583
rect 176 1576 183 1613
rect 216 1607 223 1773
rect 236 1747 243 1823
rect 276 1816 283 1993
rect 16 1367 23 1373
rect 56 1347 63 1553
rect 16 1307 23 1333
rect 76 1316 83 1353
rect 36 1287 43 1293
rect 16 1107 23 1233
rect 36 843 43 1173
rect 56 1116 63 1213
rect 76 1136 83 1273
rect 96 1267 103 1303
rect 116 1247 123 1576
rect 216 1563 223 1573
rect 236 1567 243 1583
rect 196 1556 223 1563
rect 216 1347 223 1533
rect 256 1327 263 1773
rect 296 1747 303 1833
rect 316 1747 323 2013
rect 376 2007 383 2033
rect 416 2007 423 2043
rect 336 1816 343 1833
rect 376 1827 383 1853
rect 436 1847 443 2113
rect 476 2087 483 2153
rect 496 2076 503 2413
rect 536 2287 543 2303
rect 576 2296 583 2353
rect 516 2267 523 2283
rect 596 2267 603 2493
rect 636 2276 643 2493
rect 716 2347 723 2533
rect 816 2487 823 2553
rect 716 2287 723 2333
rect 756 2296 763 2313
rect 836 2307 843 2633
rect 876 2576 883 2653
rect 916 2527 923 2613
rect 976 2556 983 2593
rect 996 2576 1003 2673
rect 1016 2607 1023 2713
rect 1036 2543 1043 2593
rect 936 2527 943 2543
rect 1016 2536 1043 2543
rect 616 2227 623 2263
rect 656 2207 663 2263
rect 656 2147 663 2153
rect 536 2087 543 2093
rect 456 2027 463 2073
rect 576 2056 583 2093
rect 656 2076 663 2133
rect 596 2027 603 2043
rect 676 2027 683 2253
rect 396 1787 403 1803
rect 416 1747 423 1823
rect 456 1816 463 1993
rect 276 1596 283 1633
rect 316 1367 323 1693
rect 296 1327 303 1343
rect 336 1336 343 1733
rect 476 1707 483 1853
rect 356 1576 363 1633
rect 416 1596 423 1653
rect 396 1507 403 1583
rect 156 1247 163 1283
rect 116 1136 123 1213
rect 147 1116 163 1123
rect 16 836 43 843
rect 16 547 23 836
rect 76 723 83 1093
rect 156 863 163 1116
rect 236 1107 243 1313
rect 276 1247 283 1323
rect 276 1127 283 1233
rect 356 1227 363 1393
rect 436 1367 443 1673
rect 476 1616 483 1653
rect 496 1607 503 1833
rect 616 1816 623 1833
rect 576 1796 583 1813
rect 516 1767 523 1783
rect 556 1747 563 1763
rect 596 1727 603 1793
rect 456 1567 463 1583
rect 476 1547 483 1573
rect 516 1556 523 1693
rect 636 1627 643 1803
rect 676 1767 683 1973
rect 696 1747 703 1833
rect 716 1807 723 2033
rect 736 1867 743 2293
rect 776 2167 783 2283
rect 796 2187 803 2303
rect 876 2276 903 2283
rect 796 2056 803 2113
rect 836 2107 843 2243
rect 876 2167 883 2276
rect 1076 2263 1083 2493
rect 1096 2287 1103 2673
rect 1036 2256 1083 2263
rect 916 2187 923 2243
rect 836 2087 843 2093
rect 876 2056 883 2153
rect 856 2027 863 2043
rect 896 2036 903 2093
rect 916 2056 923 2173
rect 936 2076 943 2133
rect 716 1763 723 1793
rect 796 1787 803 1813
rect 856 1807 863 1913
rect 916 1796 923 1813
rect 716 1756 743 1763
rect 536 1576 543 1613
rect 556 1547 563 1563
rect 336 1136 343 1153
rect 376 1147 383 1353
rect 556 1347 563 1533
rect 576 1527 583 1593
rect 596 1563 603 1613
rect 676 1563 683 1693
rect 736 1647 743 1756
rect 756 1747 763 1763
rect 776 1747 783 1783
rect 776 1687 783 1733
rect 716 1576 723 1633
rect 776 1616 783 1633
rect 796 1603 803 1773
rect 816 1627 823 1773
rect 836 1767 843 1783
rect 876 1667 883 1783
rect 896 1747 903 1773
rect 936 1707 943 1783
rect 976 1767 983 1783
rect 976 1727 983 1733
rect 836 1607 843 1633
rect 796 1596 823 1603
rect 596 1556 623 1563
rect 656 1556 683 1563
rect 656 1507 663 1533
rect 696 1527 703 1563
rect 596 1336 623 1343
rect 396 1187 403 1293
rect 456 1287 463 1333
rect 616 1327 623 1336
rect 436 1267 443 1283
rect 476 1267 483 1303
rect 396 1116 403 1153
rect 316 1096 363 1103
rect 256 867 263 1083
rect 136 856 163 863
rect 136 807 143 856
rect 176 827 183 843
rect 116 767 123 803
rect 136 723 143 793
rect 76 716 103 723
rect 16 367 23 513
rect 36 427 43 633
rect 76 616 83 653
rect 96 627 103 716
rect 116 716 143 723
rect 116 627 123 716
rect 136 636 143 693
rect 196 667 203 833
rect 216 787 223 843
rect 236 807 243 853
rect 296 836 303 953
rect 316 767 323 823
rect 336 787 343 953
rect 376 887 383 1093
rect 416 1083 423 1103
rect 416 1076 443 1083
rect 376 856 383 873
rect 416 856 423 1053
rect 436 847 443 1076
rect 496 847 503 1253
rect 576 1247 583 1323
rect 616 1307 623 1313
rect 636 1287 643 1353
rect 656 1323 663 1493
rect 656 1316 683 1323
rect 756 1267 763 1533
rect 776 1307 783 1573
rect 816 1547 823 1596
rect 916 1596 923 1653
rect 976 1616 983 1713
rect 996 1627 1003 2213
rect 1056 2076 1063 2233
rect 1116 2227 1123 2736
rect 1176 2543 1183 2733
rect 1196 2707 1203 2763
rect 1236 2607 1243 2793
rect 1276 2727 1283 2763
rect 1276 2576 1303 2583
rect 1276 2547 1283 2576
rect 1156 2536 1183 2543
rect 1276 2263 1283 2533
rect 1296 2287 1303 2533
rect 1096 2096 1103 2133
rect 1116 2047 1123 2063
rect 1016 1783 1023 1833
rect 1076 1807 1083 2033
rect 1136 1907 1143 2213
rect 1156 2107 1163 2233
rect 1156 1947 1163 2093
rect 1176 2076 1183 2253
rect 1216 2247 1223 2263
rect 1256 2256 1283 2263
rect 1216 2096 1223 2133
rect 1236 2127 1243 2243
rect 1256 2107 1263 2256
rect 1296 2076 1303 2173
rect 1316 2163 1323 2243
rect 1336 2227 1343 2893
rect 1396 2723 1403 2773
rect 1436 2756 1443 2773
rect 1396 2716 1423 2723
rect 1416 2556 1423 2716
rect 1456 2687 1463 2743
rect 1496 2723 1503 2853
rect 1536 2756 1543 2813
rect 1556 2787 1563 3013
rect 1596 2907 1603 3036
rect 1636 3027 1643 3196
rect 1656 3107 1663 3243
rect 1696 3236 1703 3253
rect 1736 3223 1743 3453
rect 1756 3267 1763 3476
rect 1776 3407 1783 3636
rect 1796 3407 1803 3473
rect 1836 3463 1843 3653
rect 1856 3587 1863 3703
rect 1876 3627 1883 3653
rect 1876 3487 1883 3553
rect 1896 3496 1903 3833
rect 1916 3727 1923 3893
rect 1956 3787 1963 3953
rect 2016 3947 2023 3983
rect 2136 3947 2143 4013
rect 1976 3787 1983 3933
rect 2156 3927 2163 4053
rect 2196 4027 2203 4033
rect 2216 3996 2223 4053
rect 2256 3996 2263 4156
rect 2356 4127 2363 4236
rect 2416 4183 2423 4213
rect 2276 3976 2283 3993
rect 2296 3947 2303 4013
rect 2356 3987 2363 4113
rect 1956 3736 1963 3773
rect 1976 3703 1983 3773
rect 2036 3747 2043 3833
rect 2056 3716 2063 3853
rect 2076 3747 2083 3813
rect 2156 3723 2163 3733
rect 2136 3716 2163 3723
rect 1976 3696 2003 3703
rect 1976 3516 1983 3533
rect 2016 3516 2023 3553
rect 2036 3547 2043 3693
rect 2116 3627 2123 3703
rect 1936 3487 1943 3503
rect 1996 3483 2003 3503
rect 1996 3476 2023 3483
rect 1816 3456 1843 3463
rect 1776 3267 1783 3353
rect 1816 3327 1823 3456
rect 1836 3307 1843 3353
rect 1836 3223 1843 3273
rect 1676 3187 1683 3223
rect 1716 3216 1743 3223
rect 1696 3187 1703 3193
rect 1656 3047 1663 3073
rect 1596 2887 1603 2893
rect 1616 2843 1623 2933
rect 1696 2927 1703 3173
rect 1716 2947 1723 3216
rect 1776 3107 1783 3223
rect 1816 3216 1843 3223
rect 1796 3127 1803 3203
rect 1776 3036 1783 3073
rect 1816 3036 1823 3053
rect 1856 3047 1863 3333
rect 1956 3307 1963 3473
rect 1976 3307 1983 3453
rect 2016 3427 2023 3476
rect 2036 3447 2043 3503
rect 2016 3387 2023 3413
rect 2016 3236 2023 3353
rect 1916 3207 1923 3223
rect 1887 3196 1903 3203
rect 1936 3167 1943 3213
rect 1596 2836 1623 2843
rect 1496 2716 1523 2723
rect 1436 2607 1443 2673
rect 1396 2287 1403 2543
rect 1436 2536 1443 2593
rect 1456 2563 1463 2573
rect 1456 2556 1483 2563
rect 1516 2556 1523 2716
rect 1576 2667 1583 2763
rect 1596 2643 1603 2836
rect 1696 2787 1703 2893
rect 1736 2776 1743 2853
rect 1616 2747 1623 2773
rect 1656 2756 1683 2763
rect 1676 2727 1683 2756
rect 1576 2636 1603 2643
rect 1456 2387 1463 2556
rect 1436 2247 1443 2263
rect 1476 2227 1483 2253
rect 1496 2247 1503 2543
rect 1536 2536 1543 2593
rect 1516 2243 1523 2373
rect 1556 2276 1563 2553
rect 1576 2487 1583 2636
rect 1596 2527 1603 2573
rect 1636 2447 1643 2543
rect 1596 2276 1603 2433
rect 1636 2276 1663 2283
rect 1636 2263 1643 2276
rect 1616 2256 1643 2263
rect 1516 2236 1543 2243
rect 1316 2156 1343 2163
rect 1236 2047 1243 2063
rect 1096 1796 1103 1893
rect 1016 1776 1043 1783
rect 1076 1747 1083 1763
rect 1156 1747 1163 1783
rect 856 1567 863 1583
rect 856 1307 863 1553
rect 896 1547 903 1583
rect 936 1567 943 1613
rect 956 1596 963 1613
rect 896 1347 903 1473
rect 1016 1347 1023 1653
rect 1036 1507 1043 1613
rect 1056 1567 1063 1633
rect 1096 1616 1103 1733
rect 1176 1727 1183 1813
rect 1256 1783 1263 1913
rect 1276 1807 1283 2053
rect 1336 1887 1343 2156
rect 1416 2076 1443 2083
rect 1356 2027 1363 2043
rect 1356 1823 1363 2013
rect 1396 1847 1403 2033
rect 1416 2027 1423 2076
rect 1516 2076 1523 2113
rect 1456 2047 1463 2053
rect 1496 2047 1503 2063
rect 1536 1987 1543 2236
rect 1556 2207 1563 2233
rect 1556 2067 1563 2093
rect 1576 2027 1583 2063
rect 1616 2047 1623 2063
rect 1336 1816 1363 1823
rect 1356 1783 1363 1816
rect 1416 1816 1423 1873
rect 1076 1367 1083 1573
rect 1116 1367 1123 1713
rect 1176 1647 1183 1693
rect 1196 1667 1203 1783
rect 1236 1776 1263 1783
rect 1336 1776 1363 1783
rect 1216 1643 1223 1673
rect 1196 1636 1223 1643
rect 1156 1627 1163 1633
rect 1136 1567 1143 1583
rect 1156 1567 1163 1573
rect 916 1307 923 1333
rect 516 887 523 1103
rect 536 1047 543 1213
rect 556 1127 563 1173
rect 576 1136 583 1213
rect 576 1083 583 1093
rect 656 1083 663 1213
rect 736 1096 743 1113
rect 576 1076 603 1083
rect 636 1076 663 1083
rect 596 823 603 893
rect 516 807 523 823
rect 536 807 543 823
rect 576 816 603 823
rect 616 856 643 863
rect 316 707 323 753
rect 327 696 343 703
rect 196 647 203 653
rect 216 623 223 633
rect 56 583 63 603
rect 56 576 83 583
rect 56 527 63 553
rect 36 376 43 393
rect 76 387 83 576
rect 156 547 163 623
rect 196 616 223 623
rect 236 616 243 633
rect 216 527 223 616
rect 276 616 283 633
rect 256 596 263 613
rect 16 327 23 333
rect 76 156 83 253
rect 96 167 103 413
rect 116 376 123 393
rect 276 387 283 493
rect 296 383 303 413
rect 316 407 323 673
rect 336 636 343 696
rect 556 687 563 803
rect 356 547 363 623
rect 396 616 423 623
rect 416 587 423 616
rect 436 567 443 633
rect 456 507 463 613
rect 496 567 503 633
rect 536 596 543 633
rect 576 487 583 603
rect 596 587 603 633
rect 616 627 623 856
rect 716 863 723 1083
rect 796 907 803 1293
rect 836 1287 843 1303
rect 816 1187 823 1283
rect 896 1276 913 1283
rect 856 1136 863 1173
rect 816 887 823 1113
rect 776 867 783 873
rect 716 856 743 863
rect 716 843 723 856
rect 796 856 823 863
rect 656 767 663 843
rect 696 836 723 843
rect 756 687 763 833
rect 796 767 803 856
rect 836 667 843 843
rect 876 727 883 1133
rect 896 1067 903 1103
rect 936 967 943 1303
rect 956 1267 963 1293
rect 976 1287 983 1313
rect 1056 1267 1063 1303
rect 1076 1287 1083 1293
rect 976 1096 983 1153
rect 996 1147 1003 1153
rect 1016 1107 1023 1173
rect 956 1047 963 1083
rect 996 1067 1003 1083
rect 916 836 923 853
rect 936 807 943 933
rect 956 867 963 1033
rect 996 856 1003 913
rect 976 703 983 843
rect 956 696 983 703
rect 296 376 323 383
rect 356 376 363 393
rect 136 347 143 363
rect 276 347 283 373
rect 116 123 123 253
rect 176 187 183 333
rect 196 327 203 343
rect 216 156 223 173
rect 276 136 283 313
rect 336 307 343 353
rect 396 347 403 393
rect 396 267 403 333
rect 476 307 483 383
rect 516 376 543 383
rect 336 156 343 173
rect 396 163 403 233
rect 396 156 423 163
rect 376 127 383 153
rect 116 116 143 123
rect 356 116 373 123
rect 416 123 423 156
rect 456 136 463 273
rect 536 247 543 376
rect 556 327 563 433
rect 496 156 503 233
rect 536 156 543 213
rect 616 167 623 613
rect 696 607 703 623
rect 736 616 763 623
rect 736 607 743 616
rect 776 607 783 653
rect 816 636 843 643
rect 696 367 703 513
rect 716 367 723 453
rect 736 387 743 593
rect 756 327 763 593
rect 816 527 823 636
rect 796 356 803 373
rect 856 363 863 613
rect 916 487 923 693
rect 836 356 863 363
rect 656 307 663 323
rect 676 187 683 313
rect 516 127 523 143
rect 616 136 623 153
rect 656 136 663 173
rect 696 147 703 313
rect 816 187 823 343
rect 836 287 843 356
rect 876 307 883 413
rect 896 387 903 473
rect 956 447 963 696
rect 976 667 983 673
rect 996 656 1003 753
rect 1016 707 1023 1073
rect 1036 1067 1043 1233
rect 1076 1136 1083 1193
rect 1096 1167 1103 1353
rect 1176 1347 1183 1613
rect 1196 1596 1203 1636
rect 1236 1623 1243 1733
rect 1216 1616 1243 1623
rect 1256 1607 1263 1693
rect 1276 1576 1283 1673
rect 1256 1507 1263 1563
rect 1276 1347 1283 1493
rect 1296 1487 1303 1553
rect 1116 1143 1123 1333
rect 1256 1316 1263 1333
rect 1176 1296 1203 1303
rect 1156 1223 1163 1283
rect 1136 1216 1163 1223
rect 1136 1187 1143 1216
rect 1107 1136 1123 1143
rect 1096 1116 1103 1133
rect 1056 1087 1063 1103
rect 1156 1096 1163 1193
rect 1176 1087 1183 1273
rect 1196 1247 1203 1296
rect 1036 856 1063 863
rect 1096 856 1123 863
rect 1036 687 1043 856
rect 1076 767 1083 843
rect 1116 807 1123 856
rect 1076 656 1083 673
rect 976 647 983 653
rect 1016 636 1043 643
rect 1016 467 1023 636
rect 1116 627 1123 793
rect 1096 616 1113 623
rect 936 387 943 393
rect 1016 376 1023 433
rect 916 347 923 363
rect 996 327 1003 363
rect 716 156 743 163
rect 416 116 443 123
rect 636 116 643 133
rect 716 87 723 156
rect 796 127 803 143
rect 816 136 823 173
rect 856 147 863 153
rect 936 147 943 273
rect 956 156 963 313
rect 996 156 1003 193
rect 1016 156 1023 213
rect 1056 156 1063 233
rect 1076 183 1083 513
rect 1096 376 1103 573
rect 1136 447 1143 1073
rect 1196 1067 1203 1173
rect 1216 1167 1223 1253
rect 1236 1227 1243 1303
rect 1276 1287 1283 1303
rect 1256 1207 1263 1273
rect 1216 1096 1223 1133
rect 1276 1116 1283 1213
rect 1296 1187 1303 1453
rect 1316 1367 1323 1673
rect 1336 1527 1343 1776
rect 1436 1767 1443 1813
rect 1356 1627 1363 1753
rect 1356 1596 1363 1613
rect 1436 1596 1443 1633
rect 1376 1547 1383 1583
rect 1356 1336 1363 1533
rect 1376 1303 1383 1513
rect 1396 1347 1403 1513
rect 1416 1407 1423 1583
rect 1456 1467 1463 1833
rect 1476 1827 1483 1853
rect 1556 1827 1563 1873
rect 1516 1816 1543 1823
rect 1496 1727 1503 1803
rect 1536 1787 1543 1816
rect 1596 1816 1603 1833
rect 1516 1727 1523 1773
rect 1616 1707 1623 1993
rect 1676 1867 1683 2193
rect 1696 2107 1703 2733
rect 1716 2536 1723 2763
rect 1756 2647 1763 2893
rect 1796 2827 1803 3033
rect 1876 2887 1883 3113
rect 1896 2947 1903 3153
rect 1916 3056 1923 3133
rect 1956 3127 1963 3223
rect 1976 3067 1983 3193
rect 2016 3127 2023 3193
rect 2036 3167 2043 3223
rect 2056 3187 2063 3473
rect 2076 3447 2083 3553
rect 2096 3467 2103 3573
rect 2136 3567 2143 3693
rect 2176 3567 2183 3913
rect 2216 3703 2223 3933
rect 2316 3867 2323 3953
rect 2336 3947 2343 3983
rect 2376 3887 2383 4013
rect 2396 3987 2403 4183
rect 2416 4176 2443 4183
rect 2416 4087 2423 4176
rect 2436 4016 2443 4053
rect 2456 4016 2463 4413
rect 2516 4307 2523 4476
rect 2696 4483 2703 4673
rect 2716 4643 2723 4713
rect 2756 4676 2783 4683
rect 2716 4636 2743 4643
rect 2576 4476 2603 4483
rect 2596 4467 2603 4476
rect 2676 4476 2703 4483
rect 2676 4447 2683 4476
rect 2716 4456 2723 4513
rect 2756 4503 2763 4633
rect 2776 4627 2783 4676
rect 2876 4647 2883 4663
rect 2756 4496 2783 4503
rect 2556 4147 2563 4373
rect 2656 4327 2663 4413
rect 2676 4307 2683 4433
rect 2696 4423 2703 4443
rect 2696 4416 2723 4423
rect 2716 4327 2723 4416
rect 2616 4196 2623 4213
rect 2496 4007 2503 4073
rect 2596 3996 2603 4183
rect 2676 4167 2683 4293
rect 2696 4147 2703 4183
rect 2716 4067 2723 4313
rect 2756 4267 2763 4496
rect 2736 4127 2743 4183
rect 2776 4176 2783 4233
rect 2816 4187 2823 4613
rect 2836 4587 2843 4633
rect 2836 4367 2843 4573
rect 2916 4567 2923 4663
rect 2916 4496 2923 4553
rect 2876 4456 2883 4493
rect 2856 4227 2863 4433
rect 2896 4423 2903 4443
rect 2876 4416 2903 4423
rect 2856 4167 2863 4183
rect 2416 3927 2423 3983
rect 2456 3927 2463 3973
rect 2196 3696 2223 3703
rect 2236 3696 2263 3703
rect 2156 3527 2163 3553
rect 2136 3496 2143 3513
rect 2156 3467 2163 3483
rect 2176 3467 2183 3533
rect 2196 3516 2203 3533
rect 2076 3227 2083 3253
rect 2116 3143 2123 3433
rect 2136 3223 2143 3433
rect 2156 3367 2163 3453
rect 2136 3216 2163 3223
rect 2096 3136 2123 3143
rect 1796 2756 1803 2813
rect 1776 2727 1783 2743
rect 1776 2556 1783 2693
rect 1836 2667 1843 2763
rect 1856 2727 1863 2853
rect 1856 2707 1863 2713
rect 1816 2556 1823 2613
rect 1856 2556 1863 2613
rect 1876 2607 1883 2833
rect 1896 2807 1903 2933
rect 1916 2756 1923 2873
rect 1956 2787 1963 3013
rect 1976 2967 1983 3003
rect 2016 2967 2023 3003
rect 2016 2867 2023 2953
rect 2036 2847 2043 3073
rect 2056 3056 2063 3113
rect 2056 2867 2063 2973
rect 1896 2587 1903 2743
rect 1936 2703 1943 2723
rect 1976 2707 1983 2733
rect 1916 2696 1943 2703
rect 1916 2587 1923 2696
rect 1996 2687 2003 2813
rect 2036 2787 2043 2833
rect 2056 2756 2063 2833
rect 2076 2727 2083 2743
rect 1936 2576 1983 2583
rect 1716 2207 1723 2473
rect 1756 2467 1763 2543
rect 1876 2487 1883 2543
rect 1916 2527 1923 2573
rect 1936 2567 1943 2576
rect 1876 2447 1883 2473
rect 1836 2263 1843 2313
rect 1816 2256 1843 2263
rect 1716 2076 1723 2153
rect 1776 2083 1783 2173
rect 1756 2076 1783 2083
rect 1816 2076 1823 2213
rect 1836 2087 1843 2133
rect 1856 2096 1883 2103
rect 1696 2056 1703 2073
rect 1636 1796 1643 1853
rect 1476 1607 1483 1633
rect 1476 1447 1483 1553
rect 1496 1527 1503 1613
rect 1556 1596 1603 1603
rect 1516 1547 1523 1563
rect 1436 1336 1443 1393
rect 1476 1336 1483 1433
rect 1516 1336 1523 1473
rect 1356 1296 1383 1303
rect 1316 1143 1323 1193
rect 1296 1136 1323 1143
rect 1296 1107 1303 1136
rect 1356 1083 1363 1296
rect 1416 1247 1423 1323
rect 1376 1136 1383 1213
rect 1456 1187 1463 1333
rect 1496 1287 1503 1323
rect 1416 1147 1423 1173
rect 1416 1103 1423 1133
rect 1496 1116 1523 1123
rect 1416 1096 1443 1103
rect 1336 1076 1363 1083
rect 1156 867 1163 1013
rect 1236 883 1243 1073
rect 1216 876 1243 883
rect 1196 856 1203 873
rect 1156 647 1163 693
rect 1176 616 1183 653
rect 1196 596 1203 673
rect 1216 643 1223 876
rect 1236 663 1243 833
rect 1256 787 1263 823
rect 1296 707 1303 823
rect 1316 767 1323 1053
rect 1276 683 1283 693
rect 1276 676 1303 683
rect 1236 656 1253 663
rect 1216 636 1243 643
rect 1256 636 1263 653
rect 1296 636 1303 676
rect 1316 647 1323 693
rect 1236 427 1243 636
rect 1116 347 1123 363
rect 1156 287 1163 363
rect 1076 176 1103 183
rect 796 107 803 113
rect 976 87 983 143
rect 1076 136 1083 153
rect 1096 147 1103 176
rect 1136 156 1143 213
rect 1176 156 1183 353
rect 1236 287 1243 383
rect 1276 363 1283 593
rect 1336 587 1343 1076
rect 1516 1067 1523 1116
rect 1376 863 1383 973
rect 1376 856 1403 863
rect 1396 743 1403 856
rect 1436 827 1443 1053
rect 1496 856 1503 1033
rect 1416 747 1423 823
rect 1476 807 1483 843
rect 1516 807 1523 993
rect 1536 927 1543 1453
rect 1556 1347 1563 1596
rect 1596 1576 1603 1596
rect 1636 1547 1643 1753
rect 1656 1667 1663 1783
rect 1676 1643 1683 1813
rect 1696 1687 1703 1853
rect 1716 1783 1723 1973
rect 1736 1967 1743 2063
rect 1796 1967 1803 2063
rect 1856 2047 1863 2096
rect 1756 1807 1763 1933
rect 1796 1796 1803 1813
rect 1716 1776 1743 1783
rect 1656 1636 1683 1643
rect 1576 1316 1583 1393
rect 1596 1347 1603 1433
rect 1616 1316 1623 1533
rect 1656 1347 1663 1636
rect 1736 1596 1743 1653
rect 1796 1627 1803 1693
rect 1836 1667 1843 1973
rect 1856 1947 1863 2033
rect 1876 1767 1883 2053
rect 1916 2027 1923 2433
rect 1956 2227 1963 2353
rect 1996 2287 2003 2593
rect 1976 2167 1983 2263
rect 2016 2147 2023 2553
rect 2056 2443 2063 2673
rect 2076 2556 2083 2613
rect 2096 2447 2103 3136
rect 2156 3036 2163 3193
rect 2176 3107 2183 3453
rect 2196 3287 2203 3453
rect 2216 3387 2223 3673
rect 2256 3587 2263 3696
rect 2236 3563 2243 3573
rect 2236 3556 2263 3563
rect 2256 3516 2263 3556
rect 2316 3547 2323 3773
rect 2356 3747 2363 3813
rect 2416 3703 2423 3733
rect 2356 3696 2383 3703
rect 2396 3696 2423 3703
rect 2336 3667 2343 3693
rect 2236 3476 2263 3483
rect 2256 3427 2263 3476
rect 2196 3207 2203 3223
rect 2216 3087 2223 3373
rect 2256 3087 2263 3413
rect 2276 3307 2283 3533
rect 2336 3516 2343 3553
rect 2316 3367 2323 3503
rect 2376 3447 2383 3696
rect 2456 3667 2463 3913
rect 2476 3727 2483 3773
rect 2496 3727 2503 3793
rect 2396 3427 2403 3613
rect 2416 3516 2423 3593
rect 2456 3527 2463 3613
rect 2316 3223 2323 3313
rect 2376 3256 2383 3313
rect 2416 3256 2423 3473
rect 2436 3347 2443 3493
rect 2296 3203 2303 3223
rect 2316 3216 2343 3223
rect 2436 3207 2443 3293
rect 2296 3196 2323 3203
rect 2296 3036 2303 3053
rect 2136 2887 2143 3023
rect 2176 2987 2183 3023
rect 2136 2807 2143 2873
rect 2116 2707 2123 2763
rect 2136 2727 2143 2743
rect 2176 2723 2183 2743
rect 2196 2727 2203 2993
rect 2216 2987 2223 3033
rect 2236 2967 2243 3023
rect 2276 3007 2283 3023
rect 2316 2987 2323 3196
rect 2456 3147 2463 3453
rect 2476 3327 2483 3593
rect 2496 3287 2503 3653
rect 2536 3627 2543 3813
rect 2596 3627 2603 3703
rect 2616 3667 2623 3693
rect 2636 3627 2643 3733
rect 2656 3647 2663 4033
rect 2856 4007 2863 4153
rect 2876 4107 2883 4416
rect 2896 4407 2903 4416
rect 2936 4387 2943 4463
rect 2676 3736 2683 3953
rect 2716 3927 2723 4003
rect 2716 3736 2723 3873
rect 2736 3747 2743 3973
rect 2756 3747 2763 3933
rect 2776 3927 2783 4003
rect 2876 3963 2883 4093
rect 2856 3956 2883 3963
rect 2747 3716 2783 3723
rect 2816 3716 2823 3873
rect 2516 3496 2523 3533
rect 2536 3516 2543 3553
rect 2596 3547 2603 3593
rect 2556 3307 2563 3503
rect 2616 3496 2623 3593
rect 2656 3547 2663 3613
rect 2676 3607 2683 3693
rect 2656 3483 2663 3513
rect 2396 3056 2403 3113
rect 2236 2887 2243 2953
rect 2256 2756 2263 2793
rect 2276 2787 2283 2973
rect 2356 2887 2363 2993
rect 2296 2776 2303 2853
rect 2336 2787 2343 2873
rect 2156 2716 2183 2723
rect 2116 2556 2123 2593
rect 2156 2447 2163 2716
rect 2216 2527 2223 2733
rect 2236 2667 2243 2743
rect 2276 2736 2303 2743
rect 2256 2687 2263 2713
rect 2296 2707 2303 2736
rect 2316 2727 2323 2763
rect 2256 2587 2263 2653
rect 2336 2587 2343 2733
rect 2356 2707 2363 2873
rect 2376 2807 2383 3023
rect 2396 2783 2403 2833
rect 2376 2776 2403 2783
rect 2376 2647 2383 2776
rect 2416 2756 2423 2793
rect 2436 2767 2443 3053
rect 2456 2987 2463 3043
rect 2496 3027 2503 3223
rect 2516 2867 2523 3093
rect 2536 3067 2543 3193
rect 2556 3107 2563 3273
rect 2576 3243 2583 3373
rect 2596 3347 2603 3483
rect 2636 3476 2663 3483
rect 2616 3267 2623 3373
rect 2676 3307 2683 3533
rect 2696 3467 2703 3633
rect 2756 3627 2763 3693
rect 2716 3496 2723 3553
rect 2776 3543 2783 3673
rect 2796 3647 2803 3703
rect 2856 3687 2863 3956
rect 2916 3787 2923 4333
rect 2956 4167 2963 4653
rect 2896 3716 2903 3733
rect 2776 3536 2803 3543
rect 2756 3427 2763 3503
rect 2836 3483 2843 3553
rect 2856 3547 2863 3593
rect 2876 3496 2883 3533
rect 2816 3476 2843 3483
rect 2716 3267 2723 3273
rect 2576 3236 2603 3243
rect 2636 3236 2643 3253
rect 2536 3036 2563 3043
rect 2576 3036 2583 3133
rect 2556 3007 2563 3036
rect 2236 2556 2263 2563
rect 2036 2436 2063 2443
rect 2036 2267 2043 2436
rect 2176 2276 2183 2333
rect 2216 2276 2223 2473
rect 2236 2347 2243 2556
rect 1936 1927 1943 2093
rect 1976 2056 1983 2093
rect 1996 2036 2003 2113
rect 1916 1903 1923 1913
rect 1916 1896 1943 1903
rect 1896 1767 1903 1783
rect 1916 1767 1923 1873
rect 1936 1803 1943 1896
rect 1936 1796 1963 1803
rect 1976 1796 1983 1893
rect 1996 1807 2003 1913
rect 2036 1887 2043 2253
rect 2056 2227 2063 2253
rect 2076 2227 2083 2263
rect 2116 2127 2123 2263
rect 2136 2243 2143 2273
rect 2136 2236 2163 2243
rect 2056 2076 2063 2113
rect 2116 2107 2123 2113
rect 2156 2076 2163 2236
rect 2256 2227 2263 2513
rect 2276 2487 2283 2543
rect 2316 2527 2323 2543
rect 2336 2507 2343 2553
rect 2296 2207 2303 2243
rect 2296 2147 2303 2173
rect 2216 2076 2223 2133
rect 2236 2076 2263 2083
rect 2176 2056 2203 2063
rect 2076 1907 2083 2053
rect 2196 2047 2203 2056
rect 1856 1627 1863 1713
rect 1856 1596 1863 1613
rect 1676 1576 1683 1593
rect 1716 1527 1723 1583
rect 1556 1227 1563 1293
rect 1596 1207 1603 1303
rect 1636 1267 1643 1293
rect 1656 1247 1663 1313
rect 1576 1087 1583 1133
rect 1596 1096 1603 1173
rect 1616 1127 1623 1193
rect 1596 1007 1603 1053
rect 1536 867 1543 893
rect 1536 836 1543 853
rect 1576 803 1583 913
rect 1616 836 1623 953
rect 1636 887 1643 1173
rect 1676 1147 1683 1373
rect 1696 1367 1703 1473
rect 1736 1427 1743 1493
rect 1736 1327 1743 1333
rect 1756 1327 1763 1593
rect 1776 1367 1783 1593
rect 1836 1567 1843 1583
rect 1876 1507 1883 1653
rect 1916 1607 1923 1653
rect 1936 1603 1943 1693
rect 1956 1623 1963 1796
rect 2016 1707 2023 1783
rect 1956 1616 1983 1623
rect 1936 1596 1963 1603
rect 1916 1547 1923 1563
rect 1836 1407 1843 1453
rect 1796 1336 1803 1373
rect 1876 1347 1883 1493
rect 1916 1347 1923 1353
rect 1696 1127 1703 1303
rect 1756 1247 1763 1273
rect 1776 1207 1783 1333
rect 1836 1327 1843 1343
rect 1816 1307 1823 1323
rect 1856 1307 1863 1323
rect 1896 1307 1903 1323
rect 1856 1287 1863 1293
rect 1656 967 1663 1113
rect 1716 1103 1723 1133
rect 1696 1096 1723 1103
rect 1736 1096 1743 1133
rect 1796 1116 1803 1233
rect 1656 836 1663 913
rect 1676 887 1683 1083
rect 1776 927 1783 1093
rect 1816 967 1823 1213
rect 1836 1103 1843 1213
rect 1876 1167 1883 1273
rect 1876 1136 1883 1153
rect 1836 1096 1863 1103
rect 1836 947 1843 1096
rect 1556 796 1583 803
rect 1376 736 1403 743
rect 1376 667 1383 736
rect 1396 447 1403 713
rect 1476 603 1483 733
rect 1496 616 1503 633
rect 1416 567 1423 603
rect 1456 596 1483 603
rect 1516 596 1523 613
rect 1576 607 1583 753
rect 1376 376 1403 383
rect 1256 356 1283 363
rect 1296 356 1323 363
rect 1256 323 1263 356
rect 1256 316 1283 323
rect 1316 207 1323 356
rect 1396 363 1403 376
rect 1476 376 1483 573
rect 1516 376 1523 453
rect 1556 383 1563 603
rect 1596 587 1603 793
rect 1636 747 1643 813
rect 1676 807 1683 823
rect 1616 727 1623 733
rect 1616 636 1623 713
rect 1636 656 1643 693
rect 1656 647 1663 653
rect 1676 467 1683 773
rect 1696 687 1703 873
rect 1756 856 1763 873
rect 1736 767 1743 843
rect 1776 807 1783 853
rect 1796 836 1803 893
rect 1856 863 1863 993
rect 1836 856 1863 863
rect 1836 836 1843 856
rect 1756 707 1763 713
rect 1696 667 1703 673
rect 1756 656 1763 693
rect 1716 567 1723 633
rect 1776 627 1783 733
rect 1816 616 1823 733
rect 1856 727 1863 753
rect 1856 683 1863 713
rect 1876 707 1883 1093
rect 1896 1047 1903 1233
rect 1936 1207 1943 1573
rect 1976 1467 1983 1616
rect 1996 1596 2003 1633
rect 2016 1627 2023 1693
rect 2036 1647 2043 1793
rect 2056 1627 2063 1833
rect 2076 1667 2083 1783
rect 2116 1767 2123 1783
rect 2136 1743 2143 2013
rect 2176 1807 2183 1893
rect 2116 1736 2143 1743
rect 2016 1547 2023 1573
rect 2056 1507 2063 1583
rect 1956 1187 1963 1353
rect 1936 1096 1943 1153
rect 1996 1147 2003 1323
rect 2036 1267 2043 1413
rect 2056 1407 2063 1473
rect 2076 1427 2083 1553
rect 2096 1403 2103 1613
rect 2116 1567 2123 1736
rect 2156 1667 2163 1773
rect 2196 1767 2203 2033
rect 2236 1847 2243 2076
rect 2276 1867 2283 2113
rect 2296 2067 2303 2133
rect 2316 2127 2323 2433
rect 2356 2387 2363 2593
rect 2396 2587 2403 2743
rect 2436 2667 2443 2723
rect 2416 2556 2423 2613
rect 2436 2507 2443 2543
rect 2436 2487 2443 2493
rect 2416 2327 2423 2373
rect 2376 2263 2383 2293
rect 2416 2263 2423 2313
rect 2376 2256 2403 2263
rect 2416 2256 2443 2263
rect 2456 2187 2463 2473
rect 2476 2123 2483 2853
rect 2496 2707 2503 2763
rect 2536 2756 2543 2853
rect 2576 2827 2583 2973
rect 2596 2847 2603 3236
rect 2676 3223 2683 3233
rect 2676 3216 2703 3223
rect 2736 3127 2743 3313
rect 2816 3307 2823 3476
rect 2896 3467 2903 3483
rect 2576 2687 2583 2793
rect 2596 2747 2603 2773
rect 2616 2756 2623 2773
rect 2536 2507 2543 2673
rect 2556 2263 2563 2313
rect 2516 2256 2543 2263
rect 2556 2256 2583 2263
rect 2536 2207 2543 2256
rect 2576 2227 2583 2256
rect 2456 2116 2483 2123
rect 2336 2056 2343 2073
rect 2376 2043 2383 2073
rect 2416 2056 2423 2073
rect 2256 1807 2263 1813
rect 2247 1776 2253 1783
rect 2276 1727 2283 1803
rect 2296 1707 2303 2013
rect 2316 1847 2323 2033
rect 2356 2027 2363 2043
rect 2376 2036 2403 2043
rect 2356 1847 2363 1953
rect 2376 1823 2383 1873
rect 2396 1867 2403 1953
rect 2456 1927 2463 2116
rect 2496 1967 2503 2113
rect 2536 2076 2543 2173
rect 2516 1887 2523 2043
rect 2536 1967 2543 1993
rect 2356 1816 2383 1823
rect 2336 1763 2343 1803
rect 2336 1756 2353 1763
rect 2136 1596 2143 1633
rect 2156 1607 2163 1653
rect 2176 1596 2183 1613
rect 2196 1596 2203 1653
rect 2276 1647 2283 1693
rect 2136 1523 2143 1533
rect 2127 1516 2143 1523
rect 2096 1396 2123 1403
rect 2056 1347 2063 1393
rect 2056 1287 2063 1303
rect 2076 1227 2083 1393
rect 2096 1336 2103 1373
rect 2116 1347 2123 1396
rect 2136 1347 2143 1413
rect 2136 1307 2143 1313
rect 2016 1136 2023 1193
rect 1996 1116 2003 1133
rect 2056 1107 2063 1193
rect 2096 1143 2103 1293
rect 2116 1147 2123 1173
rect 2076 1136 2103 1143
rect 2036 1087 2043 1103
rect 1896 867 1903 1033
rect 2016 847 2023 1053
rect 2076 907 2083 1136
rect 2136 1127 2143 1273
rect 2156 1227 2163 1493
rect 2216 1387 2223 1633
rect 2256 1596 2283 1603
rect 2236 1527 2243 1563
rect 2176 1336 2183 1353
rect 2216 1336 2223 1353
rect 2196 1167 2203 1323
rect 2156 1107 2163 1133
rect 2196 1123 2203 1153
rect 2236 1127 2243 1253
rect 2256 1147 2263 1433
rect 2276 1367 2283 1596
rect 2296 1507 2303 1693
rect 2336 1447 2343 1673
rect 2356 1627 2363 1733
rect 2376 1727 2383 1816
rect 2396 1647 2403 1813
rect 2476 1807 2483 1873
rect 2496 1816 2503 1853
rect 2536 1816 2543 1893
rect 2556 1783 2563 2213
rect 2576 2167 2583 2213
rect 2576 2027 2583 2153
rect 2596 2107 2603 2553
rect 2616 2487 2623 2713
rect 2636 2667 2643 3113
rect 2656 2987 2663 3053
rect 2676 2967 2683 3073
rect 2736 3063 2743 3113
rect 2756 3087 2763 3213
rect 2776 3067 2783 3293
rect 2836 3247 2843 3453
rect 2856 3223 2863 3373
rect 2896 3267 2903 3453
rect 2916 3347 2923 3653
rect 2936 3287 2943 3673
rect 2956 3547 2963 4053
rect 2976 4047 2983 4813
rect 3196 4667 3203 4673
rect 3016 4456 3023 4493
rect 3036 4476 3043 4663
rect 3156 4656 3183 4663
rect 3076 4476 3103 4483
rect 3096 4467 3103 4476
rect 3056 4447 3063 4463
rect 3056 4267 3063 4433
rect 3116 4427 3123 4483
rect 3176 4407 3183 4656
rect 3196 4476 3203 4653
rect 3236 4476 3243 4513
rect 3256 4447 3263 4856
rect 4016 4727 4023 4863
rect 3296 4467 3303 4673
rect 3116 4216 3123 4233
rect 3076 4196 3083 4213
rect 3096 4027 3103 4183
rect 3116 4087 3123 4173
rect 3196 4143 3203 4433
rect 3196 4136 3223 4143
rect 3176 4016 3183 4033
rect 3156 4007 3163 4013
rect 3107 3996 3123 4003
rect 3196 3967 3203 3983
rect 2996 3927 3003 3963
rect 3036 3887 3043 3963
rect 3216 3947 3223 4136
rect 3256 4007 3263 4253
rect 3296 4047 3303 4183
rect 3316 3963 3323 4713
rect 3376 4676 3383 4713
rect 3536 4696 3563 4703
rect 3476 4667 3483 4683
rect 3416 4627 3423 4663
rect 3456 4647 3463 4663
rect 3376 4476 3383 4513
rect 3356 4227 3363 4453
rect 3436 4427 3443 4443
rect 3496 4407 3503 4693
rect 3536 4687 3543 4696
rect 3576 4667 3583 4683
rect 3636 4656 3643 4693
rect 3876 4676 3883 4713
rect 4436 4683 4443 4773
rect 4476 4696 4503 4703
rect 4016 4676 4043 4683
rect 3756 4647 3763 4663
rect 3516 4507 3523 4613
rect 3556 4476 3583 4483
rect 3556 4463 3563 4476
rect 3536 4456 3563 4463
rect 3336 4167 3343 4183
rect 3356 4143 3363 4213
rect 3336 4136 3363 4143
rect 3336 3996 3343 4136
rect 3376 4003 3383 4093
rect 3356 3996 3383 4003
rect 3316 3956 3343 3963
rect 3036 3747 3043 3833
rect 2987 3736 3003 3743
rect 2976 3647 2983 3733
rect 3076 3516 3083 3553
rect 2976 3487 2983 3503
rect 2976 3467 2983 3473
rect 2996 3467 3003 3493
rect 3016 3447 3023 3503
rect 2796 3127 2803 3223
rect 2836 3216 2863 3223
rect 2836 3207 2843 3216
rect 2856 3143 2863 3173
rect 2856 3136 2883 3143
rect 2736 3056 2763 3063
rect 2696 3036 2723 3043
rect 2796 3036 2803 3093
rect 2656 2756 2663 2833
rect 2676 2743 2683 2813
rect 2696 2783 2703 3036
rect 2736 2987 2743 3023
rect 2856 3016 2863 3053
rect 2736 2807 2743 2973
rect 2696 2776 2723 2783
rect 2716 2756 2723 2776
rect 2756 2756 2763 2793
rect 2836 2747 2843 2893
rect 2876 2887 2883 3136
rect 2896 3107 2903 3253
rect 2916 3187 2923 3273
rect 2956 3247 2963 3433
rect 3036 3403 3043 3453
rect 3056 3427 3063 3493
rect 3036 3396 3063 3403
rect 2956 3223 2963 3233
rect 2996 3223 3003 3293
rect 2936 3216 2963 3223
rect 2976 3216 3003 3223
rect 2676 2736 2703 2743
rect 2636 2556 2643 2593
rect 2616 2083 2623 2193
rect 2636 2167 2643 2263
rect 2656 2187 2663 2693
rect 2676 2556 2683 2613
rect 2736 2587 2743 2743
rect 2856 2727 2863 2743
rect 2836 2567 2843 2713
rect 2676 2163 2683 2513
rect 2696 2287 2703 2333
rect 2716 2307 2723 2433
rect 2756 2296 2763 2313
rect 2656 2156 2683 2163
rect 2596 2076 2623 2083
rect 2616 1983 2623 2053
rect 2616 1976 2643 1983
rect 2556 1776 2583 1783
rect 2356 1596 2363 1613
rect 2276 1307 2283 1323
rect 2316 1316 2323 1393
rect 2336 1347 2343 1413
rect 2376 1387 2383 1633
rect 2396 1596 2403 1633
rect 2436 1596 2443 1653
rect 2436 1367 2443 1553
rect 2456 1507 2463 1753
rect 2496 1687 2503 1773
rect 2496 1596 2503 1613
rect 2456 1387 2463 1433
rect 2476 1427 2483 1563
rect 2516 1547 2523 1633
rect 2496 1387 2503 1453
rect 2416 1336 2443 1343
rect 2436 1327 2443 1336
rect 2296 1287 2303 1303
rect 2336 1267 2343 1293
rect 2356 1243 2363 1323
rect 2376 1316 2403 1323
rect 2376 1287 2383 1316
rect 2456 1323 2463 1353
rect 2496 1347 2503 1373
rect 2516 1347 2523 1533
rect 2536 1487 2543 1553
rect 2576 1487 2583 1753
rect 2596 1747 2603 1913
rect 2616 1663 2623 1753
rect 2636 1687 2643 1976
rect 2656 1967 2663 2156
rect 2736 2147 2743 2193
rect 2776 2167 2783 2313
rect 2856 2307 2863 2673
rect 2876 2667 2883 2853
rect 2896 2787 2903 3093
rect 2916 3007 2923 3023
rect 2876 2556 2883 2593
rect 2896 2487 2903 2713
rect 2916 2607 2923 2993
rect 2936 2687 2943 2893
rect 2956 2787 2963 3133
rect 2976 2927 2983 3193
rect 2996 3027 3003 3113
rect 3016 2963 3023 3053
rect 3036 2987 3043 3333
rect 3056 3147 3063 3396
rect 3076 3307 3083 3473
rect 3116 3363 3123 3933
rect 3216 3707 3223 3733
rect 3176 3687 3183 3703
rect 3136 3527 3143 3633
rect 3136 3387 3143 3483
rect 3156 3407 3163 3453
rect 3176 3427 3183 3483
rect 3196 3447 3203 3553
rect 3216 3447 3223 3693
rect 3236 3487 3243 3523
rect 3276 3467 3283 3913
rect 3296 3703 3303 3833
rect 3296 3696 3323 3703
rect 3296 3523 3303 3673
rect 3296 3516 3323 3523
rect 3116 3356 3143 3363
rect 3016 2956 3043 2963
rect 2956 2647 2963 2743
rect 2916 2556 2923 2573
rect 2936 2443 2943 2633
rect 2936 2436 2963 2443
rect 2936 2347 2943 2413
rect 2676 2076 2683 2093
rect 2716 2076 2723 2113
rect 2696 1867 2703 2073
rect 2736 2047 2743 2133
rect 2756 2087 2763 2133
rect 2776 2056 2783 2153
rect 2796 2107 2803 2293
rect 2936 2283 2943 2333
rect 2956 2287 2963 2436
rect 2976 2347 2983 2853
rect 2996 2727 3003 2743
rect 2996 2447 3003 2673
rect 3016 2527 3023 2933
rect 3036 2847 3043 2956
rect 3076 2947 3083 3273
rect 3096 3087 3103 3133
rect 3096 2967 3103 3033
rect 3036 2536 3043 2833
rect 3056 2776 3063 2813
rect 3096 2807 3103 2953
rect 3076 2667 3083 2763
rect 3116 2687 3123 3253
rect 3136 3067 3143 3356
rect 3156 3047 3163 3293
rect 3196 3247 3203 3393
rect 3236 3243 3243 3413
rect 3216 3236 3243 3243
rect 3216 3127 3223 3236
rect 3256 3207 3263 3293
rect 3176 2967 3183 3003
rect 3196 2847 3203 3093
rect 3216 2987 3223 3003
rect 3276 2887 3283 3433
rect 3296 3407 3303 3516
rect 3336 3467 3343 3956
rect 3356 3847 3363 3996
rect 3356 3647 3363 3703
rect 3356 3516 3363 3533
rect 3376 3487 3383 3953
rect 3396 3767 3403 4393
rect 3416 4187 3423 4233
rect 3416 3967 3423 4173
rect 3436 4107 3443 4183
rect 3456 4107 3463 4273
rect 3536 4263 3543 4456
rect 3596 4447 3603 4463
rect 3516 4256 3543 4263
rect 3436 4087 3443 4093
rect 3516 4027 3523 4256
rect 3536 4216 3553 4223
rect 3536 4187 3543 4216
rect 3596 4216 3603 4233
rect 3696 4227 3703 4433
rect 3736 4327 3743 4433
rect 3676 4196 3683 4213
rect 3656 4167 3663 4183
rect 3576 3996 3583 4013
rect 3596 4003 3603 4113
rect 3696 4047 3703 4183
rect 3676 4027 3683 4033
rect 3596 3996 3623 4003
rect 3436 3887 3443 3953
rect 3396 3647 3403 3753
rect 3436 3703 3443 3873
rect 3476 3867 3483 3963
rect 3496 3927 3503 3993
rect 3556 3967 3563 3983
rect 3416 3696 3443 3703
rect 3456 3687 3463 3703
rect 3476 3567 3483 3853
rect 3516 3703 3523 3893
rect 3496 3696 3523 3703
rect 3516 3587 3523 3613
rect 3336 3427 3343 3453
rect 3356 3427 3363 3473
rect 3296 3067 3303 3243
rect 3316 3167 3323 3223
rect 3356 3016 3363 3193
rect 3376 3067 3383 3433
rect 3416 3287 3423 3513
rect 3436 3256 3443 3553
rect 3496 3516 3503 3533
rect 3536 3487 3543 3633
rect 3556 3547 3563 3933
rect 3576 3707 3583 3713
rect 3616 3543 3623 3996
rect 3656 3827 3663 3853
rect 3676 3703 3683 4013
rect 3696 3996 3703 4013
rect 3716 3947 3723 4273
rect 3776 4227 3783 4593
rect 3816 4343 3823 4673
rect 4036 4667 4043 4676
rect 4056 4676 4083 4683
rect 4056 4643 4063 4676
rect 4156 4667 4163 4683
rect 4436 4676 4463 4683
rect 4056 4636 4083 4643
rect 3876 4476 3883 4633
rect 3796 4336 3823 4343
rect 3716 3827 3723 3913
rect 3756 3883 3763 4093
rect 3796 3887 3803 4336
rect 3836 4067 3843 4183
rect 3756 3876 3783 3883
rect 3656 3696 3683 3703
rect 3616 3536 3643 3543
rect 3636 3523 3643 3536
rect 3636 3516 3663 3523
rect 3676 3516 3683 3553
rect 3696 3547 3703 3703
rect 3716 3687 3723 3813
rect 3756 3627 3763 3693
rect 3776 3687 3783 3876
rect 3816 3703 3823 3753
rect 3816 3696 3843 3703
rect 3756 3547 3763 3613
rect 3696 3516 3723 3523
rect 3616 3507 3623 3513
rect 3616 3483 3623 3493
rect 3476 3387 3483 3473
rect 3476 3267 3483 3373
rect 3436 3203 3443 3213
rect 3416 3196 3443 3203
rect 3396 3043 3403 3073
rect 3416 3047 3423 3196
rect 3456 3147 3463 3243
rect 3496 3107 3503 3473
rect 3516 3267 3523 3433
rect 3556 3427 3563 3483
rect 3596 3476 3623 3483
rect 3656 3447 3663 3516
rect 3536 3327 3543 3393
rect 3576 3367 3583 3413
rect 3556 3247 3563 3313
rect 3596 3247 3603 3353
rect 3696 3347 3703 3516
rect 3736 3427 3743 3503
rect 3776 3496 3783 3633
rect 3756 3363 3763 3473
rect 3796 3463 3803 3613
rect 3836 3587 3843 3673
rect 3856 3627 3863 4113
rect 3896 4087 3903 4183
rect 3916 4127 3923 4633
rect 3956 4447 3963 4483
rect 3996 4436 4023 4443
rect 3956 4207 3963 4373
rect 3996 4247 4003 4436
rect 4036 4243 4043 4413
rect 4056 4387 4063 4443
rect 4036 4236 4063 4243
rect 3996 4207 4003 4233
rect 4056 4203 4063 4236
rect 4036 4196 4063 4203
rect 3956 4183 3963 4193
rect 3956 4176 3983 4183
rect 3896 3987 3903 4033
rect 3916 3996 3923 4053
rect 3956 4003 3963 4013
rect 3956 3996 3983 4003
rect 3876 3687 3883 3873
rect 3836 3487 3843 3513
rect 3736 3356 3763 3363
rect 3776 3456 3803 3463
rect 3636 3256 3643 3273
rect 3716 3267 3723 3313
rect 3516 3127 3523 3233
rect 3616 3223 3623 3253
rect 3676 3227 3683 3253
rect 3736 3247 3743 3356
rect 3756 3287 3763 3313
rect 3536 3207 3543 3223
rect 3616 3216 3643 3223
rect 3596 3147 3603 3193
rect 3376 3036 3403 3043
rect 3336 2987 3343 3003
rect 3376 2996 3383 3036
rect 3416 2967 3423 3003
rect 3136 2756 3143 2813
rect 3176 2723 3183 2813
rect 3156 2716 3183 2723
rect 3016 2296 3023 2393
rect 3076 2387 3083 2543
rect 3047 2296 3053 2303
rect 3096 2287 3103 2473
rect 3116 2327 3123 2633
rect 3176 2607 3183 2716
rect 3256 2687 3263 2743
rect 3276 2607 3283 2793
rect 3296 2707 3303 2933
rect 3316 2756 3323 2813
rect 3336 2683 3343 2873
rect 3416 2787 3423 2953
rect 3376 2756 3383 2773
rect 3316 2676 3343 2683
rect 3196 2536 3223 2543
rect 3196 2367 3203 2536
rect 3236 2527 3243 2573
rect 3256 2547 3263 2593
rect 3296 2523 3303 2573
rect 3276 2516 3303 2523
rect 3156 2307 3163 2313
rect 3176 2287 3183 2313
rect 3216 2287 3223 2473
rect 3236 2307 3243 2373
rect 2916 2276 2943 2283
rect 3056 2276 3083 2283
rect 2816 2107 2823 2233
rect 2856 2203 2863 2263
rect 2836 2196 2863 2203
rect 2836 2087 2843 2196
rect 2756 1947 2763 2053
rect 2696 1816 2703 1833
rect 2676 1727 2683 1783
rect 2616 1656 2643 1663
rect 2616 1596 2623 1633
rect 2636 1587 2643 1656
rect 2676 1576 2683 1673
rect 2696 1607 2703 1673
rect 2576 1427 2583 1453
rect 2556 1347 2563 1353
rect 2456 1316 2483 1323
rect 2516 1316 2523 1333
rect 2596 1327 2603 1353
rect 2336 1236 2363 1243
rect 2276 1207 2283 1233
rect 2336 1187 2343 1236
rect 2316 1136 2323 1153
rect 2176 1116 2203 1123
rect 2176 1096 2183 1116
rect 2196 963 2203 1083
rect 2216 1047 2223 1113
rect 2176 956 2203 963
rect 2096 887 2103 953
rect 2176 887 2183 956
rect 2196 907 2203 933
rect 2216 887 2223 933
rect 2236 927 2243 1093
rect 2256 1067 2263 1083
rect 2267 896 2273 903
rect 1896 767 1903 833
rect 1916 787 1923 843
rect 1936 747 1943 823
rect 1976 807 1983 823
rect 2016 767 2023 803
rect 2036 767 2043 823
rect 2056 767 2063 873
rect 2096 856 2103 873
rect 2196 856 2223 863
rect 2076 827 2083 853
rect 1856 676 1883 683
rect 1836 667 1843 673
rect 1556 376 1583 383
rect 1636 376 1643 453
rect 1396 356 1423 363
rect 1236 136 1243 173
rect 1276 147 1283 173
rect 1316 143 1323 193
rect 1316 136 1343 143
rect 1356 116 1363 233
rect 1416 123 1423 356
rect 1456 327 1463 363
rect 1476 136 1483 253
rect 1536 207 1543 363
rect 1576 343 1583 376
rect 1576 336 1603 343
rect 1536 156 1543 193
rect 1556 147 1563 273
rect 1596 187 1603 233
rect 1616 176 1623 213
rect 1576 156 1583 173
rect 1656 167 1663 343
rect 1676 267 1683 413
rect 1696 287 1703 453
rect 1736 376 1743 573
rect 1756 467 1763 613
rect 1796 427 1803 603
rect 1836 596 1843 653
rect 1856 627 1863 653
rect 1876 387 1883 676
rect 1896 627 1903 733
rect 2096 683 2103 813
rect 2116 787 2123 843
rect 2116 747 2123 773
rect 2176 727 2183 843
rect 2216 827 2223 856
rect 2216 787 2223 793
rect 2076 676 2103 683
rect 1956 656 1963 673
rect 1996 623 2003 653
rect 1976 616 2003 623
rect 2016 596 2023 673
rect 1676 187 1683 253
rect 1756 227 1763 363
rect 1796 343 1803 373
rect 1796 336 1823 343
rect 1836 247 1843 323
rect 1676 143 1683 173
rect 1716 163 1723 213
rect 1716 156 1743 163
rect 1816 156 1823 213
rect 1656 136 1683 143
rect 1696 136 1703 153
rect 1736 143 1743 156
rect 1836 147 1843 233
rect 1856 156 1863 273
rect 1896 247 1903 473
rect 1916 376 1923 593
rect 1996 347 2003 573
rect 2056 487 2063 603
rect 2036 387 2043 453
rect 2076 427 2083 676
rect 2096 407 2103 653
rect 2116 616 2123 713
rect 2176 647 2183 693
rect 2236 667 2243 893
rect 2256 687 2263 873
rect 2296 847 2303 1073
rect 2316 867 2323 1093
rect 2356 887 2363 1213
rect 2376 1007 2383 1153
rect 2336 856 2343 873
rect 2396 863 2403 1293
rect 2436 1247 2443 1293
rect 2456 1187 2463 1293
rect 2536 1287 2543 1303
rect 2556 1287 2563 1313
rect 2636 1287 2643 1533
rect 2656 1447 2663 1563
rect 2696 1547 2703 1563
rect 2716 1543 2723 1933
rect 2816 1867 2823 2053
rect 2756 1807 2763 1833
rect 2736 1707 2743 1783
rect 2776 1667 2783 1773
rect 2796 1687 2803 1853
rect 2856 1787 2863 2173
rect 2896 2083 2903 2263
rect 2956 2147 2963 2173
rect 2956 2107 2963 2113
rect 2976 2103 2983 2213
rect 3016 2207 3023 2233
rect 3036 2227 3043 2273
rect 3056 2243 3063 2276
rect 3056 2236 3083 2243
rect 3076 2203 3083 2236
rect 3096 2227 3103 2243
rect 3076 2196 3103 2203
rect 2996 2147 3003 2193
rect 3096 2167 3103 2196
rect 2976 2096 3003 2103
rect 2876 2076 2903 2083
rect 2876 2067 2883 2076
rect 2916 2056 2923 2093
rect 2976 2047 2983 2063
rect 2876 1827 2883 2033
rect 2896 2003 2903 2043
rect 2896 1996 2923 2003
rect 2836 1747 2843 1783
rect 2736 1567 2743 1653
rect 2756 1587 2763 1613
rect 2816 1596 2823 1713
rect 2876 1687 2883 1783
rect 2796 1567 2803 1583
rect 2856 1576 2863 1653
rect 2716 1536 2743 1543
rect 2676 1407 2683 1433
rect 2696 1363 2703 1393
rect 2716 1387 2723 1493
rect 2687 1356 2703 1363
rect 2676 1316 2683 1333
rect 2716 1316 2723 1373
rect 2736 1307 2743 1536
rect 2756 1367 2763 1513
rect 2776 1367 2783 1553
rect 2796 1407 2803 1493
rect 2816 1407 2823 1473
rect 2776 1327 2783 1353
rect 2416 1127 2423 1153
rect 2476 1116 2483 1133
rect 2516 1123 2523 1273
rect 2536 1227 2543 1273
rect 2596 1183 2603 1283
rect 2576 1176 2603 1183
rect 2576 1167 2583 1176
rect 2496 1116 2523 1123
rect 2416 987 2423 1033
rect 2456 927 2463 1103
rect 2476 1007 2483 1073
rect 2496 1067 2503 1116
rect 2596 1116 2603 1153
rect 2616 1116 2623 1153
rect 2536 1087 2543 1103
rect 2516 907 2523 1073
rect 2576 1067 2583 1103
rect 2376 856 2403 863
rect 2276 787 2283 813
rect 2296 707 2303 803
rect 2196 636 2223 643
rect 2156 607 2163 623
rect 2016 283 2023 353
rect 2096 343 2103 373
rect 2116 356 2123 473
rect 2136 367 2143 593
rect 2196 587 2203 636
rect 2296 627 2303 633
rect 2276 616 2293 623
rect 2316 607 2323 693
rect 2376 627 2383 673
rect 2396 643 2403 856
rect 2416 856 2443 863
rect 2416 787 2423 856
rect 2536 856 2543 953
rect 2456 667 2463 843
rect 2516 807 2523 843
rect 2556 747 2563 973
rect 2576 827 2583 1053
rect 2636 1027 2643 1233
rect 2676 1116 2683 1193
rect 2696 1187 2703 1283
rect 2756 1283 2763 1303
rect 2747 1276 2763 1283
rect 2776 1276 2793 1283
rect 2656 947 2663 1033
rect 2696 987 2703 1173
rect 2616 867 2623 933
rect 2716 927 2723 1273
rect 2736 967 2743 1273
rect 2776 1136 2783 1153
rect 2816 1143 2823 1373
rect 2836 1307 2843 1333
rect 2836 1147 2843 1253
rect 2856 1187 2863 1303
rect 2876 1267 2883 1373
rect 2896 1347 2903 1973
rect 2916 1967 2923 1996
rect 2936 1927 2943 2043
rect 2956 1827 2963 1833
rect 2916 1727 2923 1813
rect 2936 1747 2943 1783
rect 2916 1387 2923 1693
rect 2976 1667 2983 1933
rect 2996 1927 3003 2096
rect 3076 2087 3083 2153
rect 3116 2107 3123 2253
rect 3156 2087 3163 2253
rect 3176 2227 3183 2253
rect 3196 2203 3203 2263
rect 3216 2227 3223 2243
rect 3236 2203 3243 2263
rect 3256 2223 3263 2333
rect 3276 2243 3283 2493
rect 3296 2447 3303 2516
rect 3316 2423 3323 2676
rect 3376 2627 3383 2713
rect 3356 2587 3363 2613
rect 3296 2416 3323 2423
rect 3296 2267 3303 2416
rect 3316 2296 3323 2393
rect 3336 2327 3343 2513
rect 3356 2387 3363 2543
rect 3376 2507 3383 2593
rect 3396 2587 3403 2753
rect 3416 2687 3423 2733
rect 3436 2707 3443 3053
rect 3456 2987 3463 3073
rect 3536 3016 3543 3033
rect 3416 2556 3423 2633
rect 3276 2236 3303 2243
rect 3256 2216 3283 2223
rect 3176 2196 3203 2203
rect 3216 2196 3243 2203
rect 3176 2167 3183 2196
rect 3216 2183 3223 2196
rect 3196 2176 3223 2183
rect 3096 2076 3143 2083
rect 3096 2067 3103 2076
rect 3136 2056 3143 2076
rect 3016 1827 3023 1913
rect 3076 1887 3083 2043
rect 2936 1587 2943 1633
rect 2996 1623 3003 1753
rect 3016 1687 3023 1773
rect 3036 1767 3043 1853
rect 3056 1816 3063 1833
rect 3096 1807 3103 2013
rect 3116 1867 3123 2013
rect 3116 1847 3123 1853
rect 3076 1767 3083 1783
rect 3096 1767 3103 1793
rect 3116 1727 3123 1833
rect 2996 1616 3023 1623
rect 2956 1596 2963 1613
rect 3016 1587 3023 1616
rect 2856 1167 2863 1173
rect 2796 1136 2823 1143
rect 2796 1083 2803 1136
rect 2856 1116 2863 1133
rect 2876 1127 2883 1213
rect 2916 1163 2923 1333
rect 2956 1316 2963 1433
rect 2976 1347 2983 1573
rect 3016 1303 3023 1533
rect 3036 1467 3043 1713
rect 3076 1576 3083 1613
rect 3116 1576 3123 1673
rect 3136 1607 3143 1953
rect 3156 1827 3163 2043
rect 3176 1967 3183 2153
rect 3196 2107 3203 2176
rect 3216 2083 3223 2113
rect 3236 2087 3243 2173
rect 3196 2076 3223 2083
rect 3196 2056 3203 2076
rect 3216 2036 3223 2053
rect 3196 2007 3203 2013
rect 3176 1796 3183 1913
rect 3196 1847 3203 1993
rect 3256 1887 3263 2013
rect 3276 1887 3283 2216
rect 3296 2167 3303 2236
rect 3316 2207 3323 2233
rect 3336 2123 3343 2253
rect 3356 2187 3363 2213
rect 3376 2207 3383 2283
rect 3336 2116 3363 2123
rect 3356 2107 3363 2116
rect 3336 2056 3343 2093
rect 3296 2023 3303 2053
rect 3356 2027 3363 2043
rect 3296 2016 3323 2023
rect 3216 1796 3223 1833
rect 3296 1816 3303 1833
rect 3156 1767 3163 1783
rect 3156 1576 3163 1673
rect 3176 1603 3183 1733
rect 3196 1627 3203 1783
rect 3256 1767 3263 1793
rect 3236 1747 3243 1753
rect 3176 1596 3203 1603
rect 3036 1363 3043 1453
rect 3056 1427 3063 1563
rect 3136 1387 3143 1553
rect 3176 1547 3183 1563
rect 3196 1467 3203 1596
rect 3216 1547 3223 1653
rect 3236 1576 3243 1733
rect 3256 1596 3263 1713
rect 3276 1667 3283 1783
rect 3316 1727 3323 2016
rect 3336 1827 3343 1853
rect 3376 1843 3383 2033
rect 3396 1987 3403 2553
rect 3436 2527 3443 2673
rect 3456 2567 3463 2773
rect 3476 2743 3483 2913
rect 3556 2787 3563 3073
rect 3616 3056 3623 3133
rect 3636 3067 3643 3216
rect 3576 2967 3583 2993
rect 3596 2867 3603 2993
rect 3476 2736 3503 2743
rect 3476 2556 3483 2653
rect 3496 2447 3503 2736
rect 3556 2663 3563 2743
rect 3576 2687 3583 2723
rect 3616 2687 3623 3013
rect 3636 2987 3643 3033
rect 3656 3023 3663 3093
rect 3696 3087 3703 3213
rect 3716 3207 3723 3223
rect 3716 3187 3723 3193
rect 3736 3163 3743 3203
rect 3756 3167 3763 3213
rect 3716 3156 3743 3163
rect 3716 3127 3723 3156
rect 3776 3147 3783 3456
rect 3796 3387 3803 3433
rect 3816 3387 3823 3453
rect 3836 3287 3843 3453
rect 3876 3363 3883 3553
rect 3896 3543 3903 3873
rect 3936 3747 3943 3973
rect 3976 3887 3983 3996
rect 4036 3907 4043 4003
rect 4056 3943 4063 4133
rect 4076 3967 4083 4636
rect 4176 4607 4183 4653
rect 4096 4147 4103 4463
rect 4136 4307 4143 4553
rect 4176 4467 4183 4593
rect 4336 4563 4343 4643
rect 4336 4556 4363 4563
rect 4356 4527 4363 4556
rect 4356 4496 4383 4503
rect 4376 4467 4383 4496
rect 4136 4063 4143 4293
rect 4216 4183 4223 4453
rect 4196 4176 4223 4183
rect 4176 4147 4183 4153
rect 4116 4056 4143 4063
rect 4116 4016 4123 4056
rect 4056 3936 4083 3943
rect 4056 3787 4063 3793
rect 3916 3567 3923 3693
rect 3936 3647 3943 3703
rect 3976 3696 4003 3703
rect 3996 3687 4003 3696
rect 4056 3683 4063 3753
rect 4076 3727 4083 3936
rect 4136 3787 4143 4033
rect 4156 3767 4163 4073
rect 4176 3996 4183 4133
rect 4236 4067 4243 4313
rect 4276 4187 4283 4373
rect 4196 3996 4223 4003
rect 4196 3987 4203 3996
rect 4196 3827 4203 3973
rect 4216 3716 4223 3733
rect 4076 3687 4083 3713
rect 4156 3707 4163 3713
rect 3896 3536 3923 3543
rect 3916 3516 3923 3536
rect 3856 3356 3883 3363
rect 3796 3256 3803 3273
rect 3836 3256 3843 3273
rect 3816 3227 3823 3243
rect 3856 3223 3863 3356
rect 3896 3247 3903 3513
rect 3916 3267 3923 3473
rect 3936 3267 3943 3613
rect 3956 3516 3963 3573
rect 3976 3487 3983 3673
rect 4016 3667 4023 3683
rect 4036 3676 4063 3683
rect 4016 3547 4023 3653
rect 4016 3487 4023 3513
rect 4036 3467 4043 3676
rect 3976 3227 3983 3253
rect 3856 3216 3883 3223
rect 3736 3087 3743 3133
rect 3687 3036 3703 3043
rect 3736 3036 3743 3073
rect 3656 3016 3683 3023
rect 3656 2767 3663 3016
rect 3716 3003 3723 3023
rect 3776 3003 3783 3023
rect 3716 2996 3783 3003
rect 3696 2967 3703 2993
rect 3636 2707 3643 2743
rect 3676 2727 3683 2743
rect 3556 2656 3583 2663
rect 3516 2543 3523 2613
rect 3516 2536 3543 2543
rect 3436 2307 3443 2433
rect 3456 2276 3463 2393
rect 3516 2276 3523 2393
rect 3536 2307 3543 2513
rect 3556 2323 3563 2533
rect 3576 2427 3583 2656
rect 3616 2536 3623 2553
rect 3656 2547 3663 2573
rect 3596 2487 3603 2523
rect 3676 2507 3683 2713
rect 3696 2547 3703 2773
rect 3716 2727 3723 2853
rect 3736 2607 3743 2953
rect 3796 2907 3803 3193
rect 3836 3127 3843 3213
rect 3916 3207 3923 3223
rect 3876 3167 3883 3193
rect 3956 3167 3963 3223
rect 3976 3167 3983 3193
rect 3996 3147 4003 3313
rect 4016 3307 4023 3413
rect 4056 3407 4063 3653
rect 4076 3647 4083 3653
rect 4096 3607 4103 3703
rect 4136 3683 4143 3703
rect 4176 3683 4183 3693
rect 4136 3676 4183 3683
rect 4136 3587 4143 3613
rect 4076 3516 4083 3553
rect 4116 3516 4123 3573
rect 4136 3496 4143 3513
rect 4056 3287 4063 3353
rect 4016 3256 4023 3273
rect 3816 3036 3823 3093
rect 3736 2536 3743 2553
rect 3556 2316 3583 2323
rect 3416 2227 3423 2273
rect 3436 2247 3443 2263
rect 3416 2087 3423 2173
rect 3436 2076 3443 2173
rect 3456 2047 3463 2153
rect 3416 2027 3423 2043
rect 3476 2007 3483 2233
rect 3496 2227 3503 2263
rect 3516 2127 3523 2213
rect 3536 2127 3543 2263
rect 3516 2056 3523 2073
rect 3356 1836 3383 1843
rect 3356 1816 3363 1836
rect 3416 1783 3423 1953
rect 3456 1823 3463 1993
rect 3516 1847 3523 1993
rect 3556 1947 3563 2253
rect 3576 2167 3583 2316
rect 3596 2276 3603 2373
rect 3696 2347 3703 2453
rect 3716 2367 3723 2523
rect 3756 2516 3763 2613
rect 3776 2536 3783 2713
rect 3816 2687 3823 2763
rect 3796 2503 3803 2593
rect 3816 2536 3823 2633
rect 3836 2607 3843 2973
rect 3876 2867 3883 2893
rect 3876 2763 3883 2773
rect 3896 2763 3903 3033
rect 3916 2927 3923 3113
rect 3936 2983 3943 3133
rect 4016 3127 4023 3213
rect 4036 3203 4043 3243
rect 4036 3196 4053 3203
rect 3956 3047 3963 3113
rect 3976 3016 3983 3033
rect 3996 2996 4003 3073
rect 4016 3027 4023 3093
rect 4076 3067 4083 3453
rect 4096 3407 4103 3473
rect 4116 3287 4123 3433
rect 4116 3247 4123 3273
rect 4096 3207 4103 3213
rect 4116 3167 4123 3203
rect 4136 3127 4143 3223
rect 4156 3083 4163 3633
rect 4236 3607 4243 3953
rect 4256 3516 4263 3813
rect 4276 3667 4283 3933
rect 4296 3907 4303 4213
rect 4356 4203 4363 4453
rect 4396 4207 4403 4333
rect 4456 4227 4463 4653
rect 4476 4547 4483 4696
rect 4616 4676 4643 4683
rect 4476 4456 4483 4533
rect 4336 4196 4363 4203
rect 4316 4107 4323 4173
rect 4356 4047 4363 4173
rect 4376 4107 4383 4183
rect 4416 4087 4423 4213
rect 4476 4207 4483 4393
rect 4516 4327 4523 4443
rect 4556 4327 4563 4663
rect 4576 4307 4583 4443
rect 4636 4427 4643 4676
rect 4676 4463 4683 4813
rect 4736 4607 4743 4683
rect 4656 4456 4683 4463
rect 4516 4227 4523 4293
rect 4656 4267 4663 4456
rect 4576 4207 4583 4253
rect 4376 4007 4383 4073
rect 4416 4027 4423 4033
rect 4436 4027 4443 4203
rect 4456 4167 4463 4183
rect 4516 4127 4523 4193
rect 4616 4183 4623 4233
rect 4676 4223 4683 4253
rect 4656 4216 4683 4223
rect 4736 4223 4743 4433
rect 4756 4247 4763 4863
rect 4796 4827 4803 4863
rect 4936 4856 4963 4863
rect 4776 4476 4803 4483
rect 4836 4476 4843 4493
rect 4916 4487 4923 4643
rect 4936 4507 4943 4856
rect 5016 4683 5023 4773
rect 5056 4727 5063 4863
rect 5056 4696 5083 4703
rect 5016 4676 5043 4683
rect 5036 4496 5043 4653
rect 5056 4547 5063 4696
rect 4776 4407 4783 4476
rect 4776 4227 4783 4293
rect 4736 4216 4763 4223
rect 4656 4196 4663 4216
rect 4756 4196 4763 4216
rect 4536 4167 4543 4173
rect 4456 4007 4463 4113
rect 4316 3727 4323 3753
rect 4336 3727 4343 3753
rect 4356 3747 4363 3973
rect 4396 3947 4403 3983
rect 4416 3947 4423 3973
rect 4396 3767 4403 3893
rect 4456 3727 4463 3953
rect 4476 3747 4483 4053
rect 4496 3996 4503 4033
rect 4556 3976 4563 4113
rect 4336 3683 4343 3693
rect 4316 3676 4343 3683
rect 4356 3647 4363 3673
rect 4196 3496 4203 3513
rect 4236 3507 4243 3513
rect 4236 3483 4243 3493
rect 4176 3467 4183 3483
rect 4216 3476 4243 3483
rect 4176 3447 4183 3453
rect 4136 3076 4163 3083
rect 4096 3056 4103 3073
rect 4056 3036 4063 3053
rect 4036 2987 4043 3033
rect 3936 2976 3963 2983
rect 3956 2847 3963 2976
rect 4056 2967 4063 2993
rect 3936 2807 3943 2833
rect 3876 2756 3903 2763
rect 3856 2707 3863 2743
rect 3896 2707 3903 2723
rect 3896 2687 3903 2693
rect 3876 2556 3883 2613
rect 3796 2496 3823 2503
rect 3716 2347 3723 2353
rect 3676 2327 3683 2333
rect 3716 2323 3723 2333
rect 3696 2316 3723 2323
rect 3636 2307 3643 2313
rect 3636 2276 3643 2293
rect 3676 2287 3683 2313
rect 3696 2283 3703 2316
rect 3696 2276 3723 2283
rect 3756 2276 3763 2353
rect 3616 2207 3623 2233
rect 3576 2076 3583 2133
rect 3616 2096 3623 2133
rect 3636 2127 3643 2193
rect 3656 2127 3663 2263
rect 3596 2047 3603 2063
rect 3636 2007 3643 2063
rect 3656 2047 3663 2093
rect 3696 2056 3703 2253
rect 3736 2247 3743 2263
rect 3796 2227 3803 2473
rect 3816 2387 3823 2496
rect 3816 2267 3823 2353
rect 3836 2276 3843 2293
rect 3816 2207 3823 2253
rect 3856 2247 3863 2453
rect 3896 2307 3903 2593
rect 3916 2556 3923 2613
rect 3936 2607 3943 2793
rect 4056 2767 4063 2913
rect 4096 2827 4103 3013
rect 4116 2987 4123 3023
rect 4136 3007 4143 3076
rect 4176 3067 4183 3313
rect 4196 3236 4203 3253
rect 4336 3243 4343 3493
rect 4356 3467 4363 3483
rect 4316 3236 4343 3243
rect 4196 3107 4203 3153
rect 4236 3127 4243 3233
rect 4296 3147 4303 3223
rect 4336 3207 4343 3236
rect 4356 3147 4363 3393
rect 4396 3267 4403 3473
rect 4416 3467 4423 3713
rect 4436 3527 4443 3673
rect 4456 3647 4463 3683
rect 4476 3667 4483 3703
rect 4496 3507 4503 3873
rect 4516 3847 4523 3973
rect 4576 3787 4583 4153
rect 4596 4067 4603 4183
rect 4616 4176 4643 4183
rect 4636 4087 4643 4176
rect 4636 4027 4643 4053
rect 4656 4047 4663 4153
rect 4676 4107 4683 4183
rect 4716 4107 4723 4183
rect 4596 3967 4603 4013
rect 4656 3996 4663 4033
rect 4676 4016 4683 4073
rect 4736 4067 4743 4163
rect 4776 4127 4783 4213
rect 4736 4016 4743 4033
rect 4776 4007 4783 4113
rect 4616 3803 4623 3983
rect 4656 3807 4663 3953
rect 4596 3796 4623 3803
rect 4596 3743 4603 3796
rect 4576 3736 4603 3743
rect 4576 3727 4583 3736
rect 4516 3627 4523 3703
rect 4556 3683 4563 3703
rect 4616 3687 4623 3773
rect 4656 3716 4663 3793
rect 4716 3787 4723 3973
rect 4676 3747 4683 3773
rect 4736 3763 4743 3913
rect 4756 3787 4763 3983
rect 4796 3767 4803 4413
rect 4816 4367 4823 4453
rect 4836 4247 4843 4253
rect 4836 4196 4843 4233
rect 4856 4227 4863 4433
rect 4876 4347 4883 4443
rect 4816 4027 4823 4153
rect 4836 4107 4843 4153
rect 4836 4016 4843 4093
rect 4856 4027 4863 4183
rect 4916 4047 4923 4313
rect 4956 4287 4963 4433
rect 4996 4307 5003 4463
rect 5016 4243 5023 4473
rect 5076 4463 5083 4533
rect 5116 4507 5123 4613
rect 5136 4587 5143 4673
rect 5056 4456 5083 4463
rect 4996 4236 5023 4243
rect 4936 4147 4943 4163
rect 4816 3996 4823 4013
rect 4716 3756 4743 3763
rect 4696 3707 4703 3723
rect 4556 3676 4573 3683
rect 4636 3667 4643 3703
rect 4416 3307 4423 3453
rect 4436 3447 4443 3483
rect 4476 3407 4483 3483
rect 4516 3347 4523 3613
rect 4376 3207 4383 3223
rect 4156 3036 4163 3053
rect 4176 3007 4183 3023
rect 4136 2907 4143 2953
rect 4116 2767 4123 2813
rect 4156 2783 4163 2893
rect 4176 2807 4183 2993
rect 4216 2887 4223 3023
rect 4256 2883 4263 3053
rect 4296 3016 4303 3093
rect 4396 3067 4403 3193
rect 4416 3167 4423 3223
rect 4456 3216 4483 3223
rect 4456 3167 4463 3216
rect 4496 3163 4503 3203
rect 4476 3156 4503 3163
rect 4316 3056 4343 3063
rect 4316 3047 4323 3056
rect 4376 3036 4403 3043
rect 4436 3036 4443 3053
rect 4376 3023 4383 3036
rect 4356 3016 4383 3023
rect 4316 2967 4323 2993
rect 4336 2907 4343 3013
rect 4416 2947 4423 3023
rect 4456 3016 4463 3153
rect 4476 3127 4483 3156
rect 4436 2947 4443 2993
rect 4476 2983 4483 3033
rect 4496 3007 4503 3133
rect 4516 3087 4523 3193
rect 4536 3167 4543 3473
rect 4556 3287 4563 3653
rect 4596 3256 4603 3273
rect 4616 3223 4623 3633
rect 4636 3527 4643 3593
rect 4656 3587 4663 3673
rect 4656 3283 4663 3553
rect 4676 3387 4683 3503
rect 4696 3467 4703 3533
rect 4636 3276 4663 3283
rect 4636 3247 4643 3276
rect 4716 3267 4723 3756
rect 4836 3743 4843 3973
rect 4876 3887 4883 4033
rect 4936 3996 4943 4013
rect 4976 3987 4983 4193
rect 4996 4027 5003 4236
rect 5036 4047 5043 4183
rect 5076 4176 5103 4183
rect 5056 4007 5063 4153
rect 4916 3947 4923 3983
rect 4816 3736 4843 3743
rect 4736 3547 4743 3693
rect 4756 3667 4763 3733
rect 4776 3543 4783 3713
rect 4816 3667 4823 3736
rect 4876 3727 4883 3853
rect 4836 3716 4863 3723
rect 4836 3627 4843 3716
rect 4756 3536 4803 3543
rect 4816 3516 4823 3613
rect 4736 3427 4743 3493
rect 4836 3483 4843 3513
rect 4876 3496 4883 3533
rect 4916 3507 4923 3793
rect 4936 3747 4943 3953
rect 4996 3927 5003 3983
rect 4936 3667 4943 3703
rect 4836 3476 4863 3483
rect 4816 3287 4823 3473
rect 4896 3467 4903 3483
rect 4756 3247 4763 3273
rect 4836 3263 4843 3413
rect 4816 3256 4843 3263
rect 4596 3216 4623 3223
rect 4536 3047 4543 3113
rect 4556 3087 4563 3173
rect 4596 3167 4603 3216
rect 4576 3067 4583 3073
rect 4576 3016 4583 3053
rect 4516 2987 4523 3003
rect 4556 2996 4563 3013
rect 4456 2976 4483 2983
rect 4456 2923 4463 2976
rect 4436 2916 4463 2923
rect 4256 2876 4283 2883
rect 4256 2827 4263 2853
rect 4136 2776 4163 2783
rect 3956 2747 3963 2763
rect 4096 2756 4113 2763
rect 3956 2723 3963 2733
rect 4036 2723 4043 2743
rect 3956 2716 4043 2723
rect 3996 2583 4003 2633
rect 4036 2583 4043 2593
rect 3996 2576 4023 2583
rect 4036 2576 4063 2583
rect 3956 2556 3963 2573
rect 3996 2567 4003 2576
rect 3936 2427 3943 2533
rect 3916 2263 3923 2333
rect 3916 2260 3943 2263
rect 3916 2256 3947 2260
rect 3933 2247 3947 2256
rect 3736 2167 3743 2193
rect 3716 2083 3723 2153
rect 3756 2147 3763 2193
rect 3796 2183 3803 2193
rect 3896 2183 3903 2233
rect 3796 2176 3823 2183
rect 3716 2076 3743 2083
rect 3456 1816 3473 1823
rect 3516 1816 3543 1823
rect 3576 1816 3583 1953
rect 3616 1887 3623 1913
rect 3416 1776 3443 1783
rect 3476 1776 3493 1783
rect 3336 1767 3343 1773
rect 3287 1616 3293 1623
rect 3036 1356 3063 1363
rect 3056 1336 3063 1356
rect 3096 1336 3103 1373
rect 2996 1296 3023 1303
rect 2896 1156 2923 1163
rect 2796 1076 2823 1083
rect 2616 847 2623 853
rect 2636 847 2643 913
rect 2656 836 2663 893
rect 2756 847 2763 893
rect 2396 636 2423 643
rect 2496 636 2503 653
rect 2376 603 2383 613
rect 2356 596 2383 603
rect 2236 467 2243 533
rect 2316 467 2323 593
rect 2236 376 2243 453
rect 2196 347 2203 373
rect 2036 327 2043 343
rect 2076 336 2103 343
rect 2036 283 2043 293
rect 2016 276 2043 283
rect 1916 207 1923 273
rect 1736 136 1763 143
rect 1756 127 1763 136
rect 1916 136 1923 193
rect 1956 147 1963 173
rect 1396 116 1423 123
rect 1716 116 1733 123
rect 1787 116 1793 123
rect 1976 116 1983 153
rect 1996 147 2003 193
rect 2036 123 2043 276
rect 2016 116 2043 123
rect 2076 47 2083 233
rect 2096 156 2103 313
rect 2156 287 2163 313
rect 2176 247 2183 343
rect 2276 307 2283 383
rect 2296 287 2303 363
rect 2176 127 2183 233
rect 2196 147 2203 153
rect 2216 116 2223 173
rect 2236 136 2243 173
rect 2276 123 2283 253
rect 2316 203 2323 413
rect 2336 347 2343 363
rect 2356 307 2363 383
rect 2396 376 2403 573
rect 2516 427 2523 633
rect 2536 627 2543 733
rect 2596 707 2603 823
rect 2676 807 2683 843
rect 2556 596 2563 653
rect 2376 283 2383 353
rect 2256 116 2283 123
rect 2296 196 2323 203
rect 2336 276 2383 283
rect 2296 27 2303 196
rect 2316 136 2323 173
rect 2336 156 2343 276
rect 2376 167 2383 213
rect 2396 156 2403 233
rect 2416 227 2423 393
rect 2556 376 2563 473
rect 2576 407 2583 413
rect 2596 407 2603 603
rect 2616 487 2623 673
rect 2636 603 2643 733
rect 2656 647 2663 733
rect 2696 683 2703 833
rect 2716 727 2723 833
rect 2776 723 2783 953
rect 2816 856 2823 1076
rect 2896 923 2903 1156
rect 2956 1107 2963 1133
rect 2996 1083 3003 1296
rect 3116 1287 3123 1313
rect 3136 1307 3143 1343
rect 3176 1336 3183 1393
rect 3196 1347 3203 1453
rect 3216 1447 3223 1533
rect 3236 1367 3243 1473
rect 3276 1387 3283 1583
rect 3316 1563 3323 1653
rect 3376 1607 3383 1773
rect 3436 1763 3443 1776
rect 3436 1756 3473 1763
rect 3516 1747 3523 1816
rect 3556 1787 3563 1793
rect 3396 1616 3403 1673
rect 3436 1623 3443 1733
rect 3536 1687 3543 1773
rect 3596 1747 3603 1873
rect 3636 1807 3643 1833
rect 3696 1803 3703 2013
rect 3716 1967 3723 2043
rect 3736 1807 3743 2076
rect 3776 2056 3783 2153
rect 3796 2067 3803 2133
rect 3816 2063 3823 2176
rect 3876 2176 3903 2183
rect 3876 2163 3883 2176
rect 3856 2156 3883 2163
rect 3856 2147 3863 2156
rect 3816 2056 3843 2063
rect 3776 1827 3783 2013
rect 3836 1987 3843 2056
rect 3876 2043 3883 2133
rect 3896 2107 3903 2153
rect 3956 2147 3963 2353
rect 3976 2287 3983 2373
rect 3996 2347 4003 2553
rect 4036 2447 4043 2473
rect 3996 2223 4003 2233
rect 3987 2216 4003 2223
rect 4016 2167 4023 2433
rect 4056 2407 4063 2576
rect 4036 2263 4043 2393
rect 4076 2387 4083 2743
rect 4096 2627 4103 2713
rect 4116 2667 4123 2733
rect 4136 2707 4143 2776
rect 4156 2647 4163 2713
rect 4196 2707 4203 2783
rect 4256 2767 4263 2813
rect 4276 2787 4283 2876
rect 4296 2787 4303 2893
rect 4316 2787 4323 2873
rect 4216 2756 4243 2763
rect 4216 2687 4223 2756
rect 4276 2756 4283 2773
rect 4356 2756 4363 2773
rect 4256 2707 4263 2723
rect 4116 2536 4123 2573
rect 4156 2536 4163 2553
rect 4216 2547 4223 2573
rect 4076 2287 4083 2293
rect 4096 2287 4103 2493
rect 4216 2407 4223 2453
rect 4036 2256 4063 2263
rect 4016 2087 4023 2093
rect 3976 2076 4003 2083
rect 3856 2036 3883 2043
rect 3676 1796 3703 1803
rect 3436 1616 3463 1623
rect 3456 1596 3463 1616
rect 3536 1596 3543 1613
rect 3436 1563 3443 1593
rect 3316 1556 3343 1563
rect 3296 1387 3303 1553
rect 3236 1316 3243 1353
rect 3296 1327 3303 1373
rect 3316 1347 3323 1556
rect 3336 1347 3343 1533
rect 3376 1467 3383 1563
rect 3416 1556 3443 1563
rect 3336 1316 3343 1333
rect 3016 1116 3023 1133
rect 2996 1076 3023 1083
rect 2936 1067 2943 1073
rect 2916 987 2923 1053
rect 2896 916 2923 923
rect 2896 867 2903 893
rect 2796 747 2803 853
rect 2836 827 2843 843
rect 2776 716 2803 723
rect 2696 676 2723 683
rect 2636 596 2663 603
rect 2696 596 2703 653
rect 2716 647 2723 676
rect 2756 667 2763 673
rect 2796 636 2803 716
rect 2716 616 2743 623
rect 2436 156 2443 373
rect 2516 356 2543 363
rect 2496 347 2503 353
rect 2476 287 2483 323
rect 2516 307 2523 356
rect 2576 327 2583 373
rect 2616 367 2623 383
rect 2656 376 2663 553
rect 2736 547 2743 616
rect 2476 247 2483 273
rect 2516 267 2523 293
rect 2356 127 2363 143
rect 2456 136 2463 193
rect 2496 163 2503 173
rect 2496 156 2523 163
rect 2536 143 2543 313
rect 2596 247 2603 363
rect 2616 327 2623 333
rect 2636 307 2643 363
rect 2616 183 2623 253
rect 2596 176 2623 183
rect 2596 163 2603 176
rect 2576 156 2603 163
rect 2536 136 2563 143
rect 2556 127 2563 136
rect 2596 -24 2603 13
rect 2636 -24 2643 213
rect 2656 -17 2663 213
rect 2676 27 2683 433
rect 2696 227 2703 473
rect 2736 387 2743 453
rect 2756 387 2763 593
rect 2776 547 2783 613
rect 2796 487 2803 593
rect 2816 507 2823 813
rect 2856 707 2863 863
rect 2876 807 2883 813
rect 2896 747 2903 833
rect 2916 667 2923 916
rect 2936 727 2943 843
rect 2996 807 3003 823
rect 2836 636 2863 643
rect 2836 567 2843 636
rect 2936 636 2943 673
rect 2956 627 2963 693
rect 3016 647 3023 1076
rect 3036 867 3043 933
rect 3076 887 3083 1273
rect 3176 1267 3183 1293
rect 3196 1283 3203 1313
rect 3256 1283 3263 1303
rect 3196 1276 3263 1283
rect 3116 1096 3123 1113
rect 3156 1087 3163 1173
rect 3136 987 3143 1083
rect 3176 947 3183 1133
rect 3196 1116 3203 1173
rect 3236 1116 3243 1133
rect 3276 1123 3283 1253
rect 3296 1183 3303 1293
rect 3316 1287 3323 1303
rect 3296 1176 3323 1183
rect 3316 1127 3323 1176
rect 3276 1116 3303 1123
rect 3296 1107 3303 1116
rect 3336 1107 3343 1193
rect 3356 1187 3363 1303
rect 3396 1143 3403 1433
rect 3416 1307 3423 1556
rect 3476 1467 3483 1583
rect 3496 1527 3503 1553
rect 3516 1527 3523 1573
rect 3556 1447 3563 1733
rect 3656 1687 3663 1783
rect 3596 1596 3603 1673
rect 3696 1627 3703 1773
rect 3716 1767 3723 1783
rect 3736 1667 3743 1763
rect 3636 1607 3643 1613
rect 3576 1407 3583 1593
rect 3456 1316 3463 1333
rect 3396 1136 3423 1143
rect 3216 1067 3223 1103
rect 3256 1087 3263 1103
rect 3256 987 3263 1073
rect 3276 987 3283 1013
rect 3096 836 3123 843
rect 3036 807 3043 823
rect 3056 783 3063 793
rect 3036 776 3063 783
rect 3036 667 3043 776
rect 3076 667 3083 803
rect 3116 687 3123 836
rect 3176 836 3183 933
rect 3256 856 3263 873
rect 3296 856 3303 993
rect 3336 867 3343 993
rect 3356 907 3363 1083
rect 3376 947 3383 1133
rect 3356 863 3363 893
rect 3396 887 3403 1136
rect 3436 867 3443 1093
rect 3456 1067 3463 1193
rect 3476 947 3483 1393
rect 3596 1367 3603 1493
rect 3616 1487 3623 1583
rect 3656 1576 3663 1613
rect 3696 1576 3703 1593
rect 3716 1556 3723 1593
rect 3736 1576 3743 1633
rect 3756 1607 3763 1783
rect 3776 1607 3783 1793
rect 3816 1783 3823 1973
rect 3836 1863 3843 1933
rect 3856 1927 3863 2036
rect 3876 2007 3883 2013
rect 3896 1947 3903 2073
rect 3836 1856 3863 1863
rect 3796 1776 3823 1783
rect 3796 1587 3803 1753
rect 3836 1747 3843 1783
rect 3816 1587 3823 1733
rect 3856 1607 3863 1856
rect 3876 1627 3883 1853
rect 3916 1843 3923 2013
rect 3936 1907 3943 2033
rect 3956 1987 3963 2033
rect 3996 1987 4003 2076
rect 4056 2076 4063 2093
rect 4076 2087 4083 2233
rect 4136 2227 4143 2393
rect 4236 2363 4243 2523
rect 4256 2363 4263 2613
rect 4276 2467 4283 2573
rect 4296 2563 4303 2743
rect 4316 2587 4323 2753
rect 4336 2567 4343 2713
rect 4356 2567 4363 2573
rect 4296 2556 4323 2563
rect 4316 2536 4323 2556
rect 4376 2543 4383 2713
rect 4396 2587 4403 2673
rect 4416 2576 4423 2653
rect 4436 2587 4443 2916
rect 4456 2707 4463 2813
rect 4476 2776 4483 2953
rect 4496 2807 4503 2973
rect 4567 2956 4573 2963
rect 4596 2947 4603 3133
rect 4616 3027 4623 3193
rect 4636 3067 4643 3213
rect 4656 3207 4663 3233
rect 4656 3056 4663 3193
rect 4676 3187 4683 3223
rect 4716 3187 4723 3223
rect 4736 3207 4743 3223
rect 4696 3056 4703 3073
rect 4736 3067 4743 3113
rect 4516 2787 4523 2893
rect 4356 2536 4383 2543
rect 4296 2487 4303 2523
rect 4336 2516 4343 2533
rect 4236 2356 4263 2363
rect 4216 2296 4223 2313
rect 4156 2247 4163 2283
rect 4036 1987 4043 2063
rect 4016 1847 4023 1853
rect 3916 1836 3943 1843
rect 3896 1816 3903 1833
rect 3936 1827 3943 1836
rect 3976 1807 3983 1833
rect 3916 1727 3923 1803
rect 4016 1796 4023 1833
rect 4056 1783 4063 1813
rect 4036 1776 4063 1783
rect 3896 1627 3903 1693
rect 3916 1627 3923 1713
rect 3936 1616 3943 1693
rect 3896 1603 3903 1613
rect 3896 1596 3923 1603
rect 3956 1596 3963 1613
rect 3776 1543 3783 1573
rect 3816 1556 3843 1563
rect 3756 1536 3783 1543
rect 3676 1527 3683 1533
rect 3516 1336 3533 1343
rect 3516 1316 3523 1336
rect 3536 1287 3543 1313
rect 3576 1307 3583 1343
rect 3616 1336 3623 1353
rect 3636 1327 3643 1373
rect 3516 1096 3523 1113
rect 3556 1087 3563 1293
rect 3536 1007 3543 1083
rect 3576 1027 3583 1173
rect 3636 1147 3643 1293
rect 3656 1147 3663 1393
rect 3676 1387 3683 1393
rect 3696 1363 3703 1413
rect 3676 1356 3703 1363
rect 3676 1347 3683 1356
rect 3596 1067 3603 1083
rect 3636 1047 3643 1053
rect 3356 856 3383 863
rect 3136 807 3143 833
rect 3156 787 3163 823
rect 2876 587 2883 623
rect 2976 616 2983 633
rect 2736 356 2743 373
rect 2796 363 2803 453
rect 2836 407 2843 413
rect 2776 356 2803 363
rect 2816 356 2823 373
rect 2836 367 2843 393
rect 2856 356 2863 453
rect 2936 407 2943 593
rect 2956 567 2963 593
rect 3056 587 3063 653
rect 3076 607 3083 633
rect 2976 567 2983 573
rect 3156 567 3163 623
rect 3176 567 3183 793
rect 3196 787 3203 803
rect 3256 707 3263 733
rect 3216 667 3223 673
rect 3216 547 3223 613
rect 3236 603 3243 693
rect 3276 687 3283 843
rect 3376 843 3383 856
rect 3456 863 3463 933
rect 3456 856 3483 863
rect 3376 836 3403 843
rect 3356 807 3363 833
rect 3476 827 3483 856
rect 3416 767 3423 823
rect 3456 816 3473 823
rect 3496 787 3503 843
rect 3536 836 3543 953
rect 3596 836 3603 953
rect 3636 907 3643 1013
rect 3656 887 3663 1113
rect 3716 1087 3723 1213
rect 3736 1096 3743 1153
rect 3756 1107 3763 1536
rect 3796 1523 3803 1553
rect 3776 1516 3803 1523
rect 3776 1347 3783 1516
rect 3796 1387 3803 1493
rect 3816 1347 3823 1556
rect 3836 1407 3843 1533
rect 3876 1387 3883 1553
rect 3896 1467 3903 1573
rect 3936 1507 3943 1573
rect 3976 1567 3983 1673
rect 3956 1427 3963 1553
rect 3996 1543 4003 1753
rect 4016 1607 4023 1753
rect 4036 1747 4043 1776
rect 4056 1623 4063 1673
rect 4076 1647 4083 1933
rect 4096 1767 4103 2213
rect 4156 2127 4163 2233
rect 4196 2147 4203 2273
rect 4236 2263 4243 2333
rect 4256 2307 4263 2356
rect 4276 2287 4283 2413
rect 4316 2327 4323 2493
rect 4356 2447 4363 2493
rect 4376 2347 4383 2536
rect 4396 2527 4403 2543
rect 4336 2283 4343 2313
rect 4316 2276 4343 2283
rect 4236 2256 4263 2263
rect 4116 2067 4123 2113
rect 4156 2107 4163 2113
rect 4216 2103 4223 2253
rect 4216 2096 4243 2103
rect 4116 2007 4123 2033
rect 4136 1967 4143 2093
rect 4136 1807 4143 1933
rect 4196 1867 4203 2053
rect 4216 1967 4223 2053
rect 4236 2027 4243 2096
rect 4256 2027 4263 2153
rect 4296 2147 4303 2263
rect 4276 2087 4283 2133
rect 4316 2107 4323 2276
rect 4356 2243 4363 2293
rect 4396 2287 4403 2373
rect 4416 2367 4423 2533
rect 4436 2343 4443 2553
rect 4456 2536 4463 2653
rect 4476 2627 4483 2733
rect 4496 2667 4503 2763
rect 4516 2687 4523 2733
rect 4516 2627 4523 2633
rect 4476 2556 4483 2593
rect 4516 2556 4523 2613
rect 4416 2336 4443 2343
rect 4416 2307 4423 2336
rect 4436 2276 4443 2293
rect 4456 2263 4463 2453
rect 4496 2447 4503 2543
rect 4536 2507 4543 2833
rect 4556 2807 4563 2913
rect 4576 2787 4583 2893
rect 4576 2756 4583 2773
rect 4596 2767 4603 2913
rect 4616 2887 4623 2993
rect 4636 2987 4643 3013
rect 4656 2907 4663 3013
rect 4676 2987 4683 3023
rect 4676 2847 4683 2953
rect 4696 2887 4703 3013
rect 4756 2967 4763 3153
rect 4776 3027 4783 3173
rect 4796 3147 4803 3233
rect 4816 3167 4823 3256
rect 4896 3247 4903 3433
rect 4936 3283 4943 3573
rect 4956 3567 4963 3873
rect 4976 3736 4983 3753
rect 4996 3747 5003 3893
rect 4916 3276 4943 3283
rect 4836 3207 4843 3223
rect 4876 3216 4893 3223
rect 4836 3187 4843 3193
rect 4796 3087 4803 3093
rect 4796 3036 4803 3073
rect 4816 3056 4823 3093
rect 4836 3036 4843 3053
rect 4856 3043 4863 3153
rect 4876 3067 4883 3193
rect 4896 3087 4903 3213
rect 4916 3167 4923 3276
rect 4956 3263 4963 3493
rect 5016 3487 5023 3973
rect 5036 3947 5043 3983
rect 5076 3963 5083 4153
rect 5096 4143 5103 4176
rect 5116 4167 5123 4453
rect 5096 4136 5123 4143
rect 5056 3956 5083 3963
rect 5036 3587 5043 3913
rect 4936 3256 4963 3263
rect 4896 3056 4903 3073
rect 4856 3036 4883 3043
rect 4916 3036 4923 3113
rect 4856 3003 4863 3013
rect 4836 2996 4863 3003
rect 4696 2776 4703 2853
rect 4636 2723 4643 2763
rect 4596 2716 4643 2723
rect 4476 2296 4483 2313
rect 4456 2256 4483 2263
rect 4476 2247 4483 2256
rect 4356 2236 4383 2243
rect 4296 2083 4303 2093
rect 4296 2076 4323 2083
rect 4316 2036 4323 2076
rect 4336 2056 4343 2113
rect 4216 1816 4223 1833
rect 4116 1727 4123 1783
rect 4156 1747 4163 1783
rect 4136 1707 4143 1733
rect 4056 1616 4083 1623
rect 4096 1607 4103 1653
rect 3996 1536 4023 1543
rect 3976 1487 3983 1513
rect 3796 1247 3803 1303
rect 3816 1207 3823 1333
rect 3856 1316 3863 1333
rect 3896 1316 3903 1333
rect 3836 1267 3843 1303
rect 3876 1287 3883 1303
rect 3676 1047 3683 1083
rect 3776 1007 3783 1173
rect 3876 1123 3883 1273
rect 3916 1187 3923 1273
rect 3936 1207 3943 1353
rect 3956 1303 3963 1393
rect 3996 1387 4003 1393
rect 3976 1347 3983 1353
rect 3996 1307 4003 1373
rect 4016 1347 4023 1536
rect 4076 1527 4083 1573
rect 4036 1347 4043 1413
rect 3956 1296 3983 1303
rect 3956 1267 3963 1296
rect 4036 1267 4043 1303
rect 3856 1116 3883 1123
rect 3836 1087 3843 1103
rect 3796 907 3803 1033
rect 3656 843 3663 873
rect 3647 836 3663 843
rect 3676 827 3683 843
rect 3516 747 3523 823
rect 3616 767 3623 823
rect 3276 616 3283 653
rect 3316 616 3343 623
rect 3236 596 3263 603
rect 3336 567 3343 616
rect 3076 376 3083 513
rect 2716 183 2723 333
rect 2756 307 2763 343
rect 2896 267 2903 373
rect 3036 367 3043 373
rect 2916 327 2923 343
rect 2756 227 2763 253
rect 2707 176 2723 183
rect 2696 156 2703 173
rect 2736 156 2743 173
rect 2716 127 2723 143
rect 2756 136 2763 213
rect 2936 163 2943 273
rect 2956 207 2963 343
rect 2996 227 3003 333
rect 3016 187 3023 363
rect 2916 156 2943 163
rect 2916 143 2923 156
rect 3016 147 3023 173
rect 3036 163 3043 353
rect 3056 287 3063 363
rect 3096 347 3103 473
rect 3116 367 3123 453
rect 3216 387 3223 413
rect 3356 387 3363 673
rect 3376 616 3383 653
rect 3436 636 3443 673
rect 3636 663 3643 813
rect 3656 687 3663 813
rect 3676 807 3683 813
rect 3696 807 3703 863
rect 3756 847 3763 893
rect 3696 787 3703 793
rect 3776 787 3783 853
rect 3796 827 3803 843
rect 3636 656 3663 663
rect 3456 603 3463 653
rect 3516 607 3523 653
rect 3536 616 3563 623
rect 3556 607 3563 616
rect 3456 596 3483 603
rect 3436 527 3443 593
rect 3556 387 3563 593
rect 3596 447 3603 613
rect 3636 607 3643 623
rect 3156 336 3173 343
rect 3156 307 3163 336
rect 3176 307 3183 313
rect 3036 156 3063 163
rect 3096 156 3103 273
rect 3136 156 3143 173
rect 2896 136 2923 143
rect 3176 136 3183 293
rect 3196 267 3203 363
rect 3236 267 3243 363
rect 3276 347 3283 363
rect 3316 347 3323 373
rect 3336 356 3343 373
rect 3256 327 3263 333
rect 3396 267 3403 343
rect 3416 227 3423 373
rect 3436 307 3443 353
rect 3456 327 3463 383
rect 3476 347 3483 363
rect 3516 267 3523 353
rect 3616 347 3623 513
rect 3636 427 3643 573
rect 3656 427 3663 656
rect 3676 636 3683 693
rect 3816 667 3823 853
rect 3876 847 3883 1093
rect 3896 967 3903 1083
rect 3936 1076 3943 1173
rect 3956 1103 3963 1153
rect 3996 1136 4003 1173
rect 4016 1147 4023 1213
rect 4056 1107 4063 1353
rect 4076 1347 4083 1433
rect 4096 1343 4103 1353
rect 4116 1343 4123 1693
rect 4176 1667 4183 1773
rect 4196 1747 4203 1803
rect 4236 1783 4243 1973
rect 4216 1776 4243 1783
rect 4136 1627 4143 1653
rect 4136 1367 4143 1553
rect 4096 1336 4123 1343
rect 4096 1316 4103 1336
rect 4076 1287 4083 1303
rect 4076 1116 4083 1273
rect 4116 1227 4123 1303
rect 4136 1187 4143 1313
rect 4116 1116 4123 1153
rect 3956 1096 3983 1103
rect 4136 1096 4143 1133
rect 3896 823 3903 933
rect 3936 907 3943 933
rect 3956 907 3963 1033
rect 3976 967 3983 1033
rect 3996 1007 4003 1093
rect 3936 836 3943 853
rect 3976 836 3983 953
rect 4056 887 4063 993
rect 4096 987 4103 1073
rect 3876 816 3903 823
rect 3756 616 3763 633
rect 3736 387 3743 613
rect 3776 607 3783 653
rect 3756 387 3763 573
rect 3816 507 3823 603
rect 3656 347 3663 383
rect 3536 307 3543 343
rect 3576 336 3593 343
rect 3676 327 3683 363
rect 3816 363 3823 433
rect 3796 356 3823 363
rect 3536 287 3543 293
rect 3676 287 3683 313
rect 3716 267 3723 353
rect 3736 307 3743 343
rect 3116 127 3123 133
rect 3216 127 3223 173
rect 3256 136 3263 213
rect 3316 156 3323 173
rect 3396 123 3403 193
rect 3456 147 3463 173
rect 3516 156 3523 193
rect 3536 156 3543 213
rect 3576 156 3583 233
rect 3656 176 3663 213
rect 3596 136 3603 173
rect 3736 163 3743 173
rect 3756 163 3763 313
rect 3796 247 3803 356
rect 3836 347 3843 673
rect 3876 667 3883 816
rect 3896 623 3903 793
rect 3916 747 3923 823
rect 3956 687 3963 823
rect 3876 616 3903 623
rect 3916 656 3943 663
rect 3916 567 3923 656
rect 3976 607 3983 633
rect 3996 587 4003 653
rect 3916 447 3923 553
rect 3896 407 3903 413
rect 3896 376 3903 393
rect 3816 307 3823 333
rect 3876 327 3883 363
rect 3916 343 3923 393
rect 3916 336 3943 343
rect 3976 327 3983 343
rect 3876 207 3883 293
rect 3736 156 3763 163
rect 3876 156 3883 193
rect 3916 183 3923 313
rect 3956 307 3963 323
rect 4016 307 4023 813
rect 4036 747 4043 863
rect 4056 807 4063 843
rect 4076 707 4083 813
rect 4096 663 4103 933
rect 4116 887 4123 1073
rect 4156 887 4163 1633
rect 4176 1387 4183 1613
rect 4196 1547 4203 1713
rect 4216 1596 4223 1776
rect 4256 1667 4263 1953
rect 4276 1747 4283 1973
rect 4296 1947 4303 2013
rect 4356 1927 4363 2213
rect 4376 2087 4383 2236
rect 4396 2056 4403 2153
rect 4456 2107 4463 2233
rect 4516 2227 4523 2293
rect 4536 2267 4543 2273
rect 4416 2036 4423 2073
rect 4436 2067 4443 2093
rect 4476 2076 4483 2193
rect 4296 1887 4303 1893
rect 4296 1816 4303 1873
rect 4316 1843 4323 1913
rect 4436 1907 4443 1993
rect 4316 1836 4343 1843
rect 4336 1827 4343 1836
rect 4356 1827 4363 1853
rect 4376 1807 4383 1873
rect 4456 1863 4463 2073
rect 4536 2047 4543 2063
rect 4476 2007 4483 2033
rect 4436 1856 4463 1863
rect 4296 1727 4303 1773
rect 4316 1767 4323 1803
rect 4256 1616 4263 1633
rect 4216 1403 4223 1513
rect 4236 1507 4243 1583
rect 4256 1487 4263 1533
rect 4276 1487 4283 1583
rect 4216 1396 4243 1403
rect 4216 1303 4223 1373
rect 4236 1367 4243 1396
rect 4256 1367 4263 1473
rect 4276 1363 4283 1393
rect 4296 1387 4303 1633
rect 4336 1627 4343 1773
rect 4356 1707 4363 1783
rect 4396 1703 4403 1783
rect 4416 1747 4423 1773
rect 4376 1696 4403 1703
rect 4376 1627 4383 1696
rect 4396 1563 4403 1673
rect 4436 1663 4443 1856
rect 4456 1827 4463 1833
rect 4476 1727 4483 1753
rect 4476 1687 4483 1713
rect 4496 1687 4503 1913
rect 4416 1656 4443 1663
rect 4416 1607 4423 1656
rect 4516 1647 4523 2013
rect 4536 1967 4543 2033
rect 4556 1987 4563 2573
rect 4576 2556 4583 2633
rect 4596 2587 4603 2693
rect 4636 2607 4643 2716
rect 4656 2683 4663 2713
rect 4676 2707 4683 2753
rect 4656 2676 4683 2683
rect 4576 2207 4583 2493
rect 4596 2447 4603 2543
rect 4636 2527 4643 2543
rect 4616 2467 4623 2513
rect 4636 2507 4643 2513
rect 4656 2327 4663 2633
rect 4676 2607 4683 2676
rect 4696 2583 4703 2713
rect 4716 2707 4723 2933
rect 4796 2927 4803 2973
rect 4756 2783 4763 2893
rect 4776 2787 4783 2873
rect 4736 2776 4763 2783
rect 4736 2643 4743 2776
rect 4776 2756 4783 2773
rect 4796 2767 4803 2833
rect 4816 2767 4823 2833
rect 4836 2807 4843 2996
rect 4856 2887 4863 2973
rect 4876 2927 4883 3036
rect 4896 2907 4903 3013
rect 4936 2923 4943 3256
rect 4916 2916 4943 2923
rect 4896 2776 4903 2813
rect 4756 2663 4763 2743
rect 4836 2723 4843 2763
rect 4796 2716 4843 2723
rect 4756 2656 4783 2663
rect 4776 2647 4783 2656
rect 4736 2636 4763 2643
rect 4736 2587 4743 2593
rect 4696 2576 4723 2583
rect 4716 2567 4723 2576
rect 4696 2536 4703 2553
rect 4736 2547 4743 2573
rect 4616 2187 4623 2283
rect 4636 2267 4643 2303
rect 4576 2043 4583 2113
rect 4616 2067 4623 2133
rect 4636 2107 4643 2253
rect 4676 2227 4683 2453
rect 4736 2347 4743 2473
rect 4756 2427 4763 2636
rect 4776 2587 4783 2613
rect 4776 2556 4783 2573
rect 4816 2556 4823 2716
rect 4836 2563 4843 2693
rect 4856 2627 4863 2753
rect 4876 2747 4883 2763
rect 4836 2556 4863 2563
rect 4796 2467 4803 2543
rect 4796 2447 4803 2453
rect 4696 2167 4703 2313
rect 4716 2296 4723 2333
rect 4756 2287 4763 2293
rect 4796 2287 4803 2393
rect 4736 2267 4743 2283
rect 4776 2276 4793 2283
rect 4727 2216 4743 2223
rect 4656 2067 4663 2073
rect 4696 2056 4703 2133
rect 4716 2087 4723 2113
rect 4576 2036 4603 2043
rect 4556 1807 4563 1813
rect 4596 1796 4603 1853
rect 4616 1847 4623 1993
rect 4436 1636 4503 1643
rect 4436 1596 4443 1636
rect 4496 1627 4503 1636
rect 4536 1623 4543 1783
rect 4616 1763 4623 1813
rect 4636 1796 4643 1853
rect 4676 1847 4683 2033
rect 4716 1967 4723 2043
rect 4736 1967 4743 2216
rect 4776 2083 4783 2093
rect 4756 2076 4783 2083
rect 4756 2023 4763 2076
rect 4796 2067 4803 2153
rect 4816 2127 4823 2333
rect 4856 2303 4863 2556
rect 4876 2327 4883 2713
rect 4916 2707 4923 2916
rect 4936 2807 4943 2893
rect 4956 2827 4963 3023
rect 4976 2807 4983 3473
rect 5016 3247 5023 3453
rect 5056 3427 5063 3956
rect 5076 3907 5083 3933
rect 5076 3527 5083 3833
rect 5096 3447 5103 4013
rect 5116 3647 5123 4136
rect 5136 4087 5143 4233
rect 5136 3927 5143 4033
rect 5136 3467 5143 3893
rect 5056 3256 5083 3263
rect 5056 3227 5063 3256
rect 5016 3187 5023 3203
rect 5036 3187 5043 3223
rect 5116 3223 5123 3273
rect 5096 3216 5123 3223
rect 5056 3043 5063 3153
rect 5076 3067 5083 3213
rect 5056 3036 5083 3043
rect 4996 2907 5003 2993
rect 5016 2987 5023 3023
rect 4896 2607 4903 2673
rect 4936 2667 4943 2763
rect 4956 2687 4963 2783
rect 4996 2776 5003 2833
rect 4916 2587 4923 2593
rect 4936 2556 4943 2653
rect 4976 2567 4983 2613
rect 4996 2567 5003 2733
rect 5016 2667 5023 2873
rect 5016 2547 5023 2573
rect 4896 2527 4903 2543
rect 4896 2307 4903 2493
rect 4916 2487 4923 2533
rect 4956 2527 4963 2543
rect 4996 2536 5013 2543
rect 4936 2307 4943 2513
rect 4856 2296 4883 2303
rect 4876 2287 4883 2296
rect 4856 2227 4863 2263
rect 4896 2256 4923 2263
rect 4836 2056 4843 2093
rect 4916 2087 4923 2256
rect 4956 2247 4963 2263
rect 4936 2067 4943 2093
rect 4816 2036 4823 2053
rect 4756 2016 4783 2023
rect 4716 1827 4723 1953
rect 4676 1763 4683 1773
rect 4616 1756 4643 1763
rect 4607 1736 4613 1743
rect 4536 1616 4553 1623
rect 4356 1527 4363 1563
rect 4376 1556 4403 1563
rect 4316 1367 4323 1453
rect 4276 1356 4303 1363
rect 4296 1323 4303 1356
rect 4376 1336 4383 1556
rect 4416 1527 4423 1563
rect 4436 1507 4443 1553
rect 4216 1296 4243 1303
rect 4176 1067 4183 1253
rect 4196 1147 4203 1273
rect 4216 1147 4223 1273
rect 4196 967 4203 1093
rect 4236 1007 4243 1296
rect 4256 1287 4263 1323
rect 4296 1316 4323 1323
rect 4296 1247 4303 1273
rect 4316 1247 4323 1293
rect 4336 1207 4343 1313
rect 4356 1267 4363 1323
rect 4136 787 4143 863
rect 4176 856 4203 863
rect 4156 767 4163 833
rect 4176 667 4183 813
rect 4196 747 4203 856
rect 4236 863 4243 973
rect 4256 867 4263 1193
rect 4296 1116 4303 1173
rect 4316 1067 4323 1103
rect 4227 856 4243 863
rect 4236 843 4243 856
rect 4236 836 4263 843
rect 4236 787 4243 803
rect 4096 656 4123 663
rect 4076 587 4083 603
rect 3896 176 3923 183
rect 3916 167 3923 176
rect 3376 116 3403 123
rect 3736 116 3743 156
rect 3956 136 3963 253
rect 3936 107 3943 123
rect 3996 123 4003 293
rect 4036 267 4043 433
rect 4116 347 4123 656
rect 4196 647 4203 673
rect 4256 656 4263 693
rect 4276 667 4283 823
rect 4156 636 4183 643
rect 4176 607 4183 636
rect 4216 636 4223 653
rect 4136 587 4143 603
rect 4196 587 4203 613
rect 4256 487 4263 613
rect 4276 607 4283 623
rect 4216 376 4243 383
rect 4276 376 4283 393
rect 4176 367 4183 373
rect 4096 336 4113 343
rect 4096 327 4103 336
rect 4076 267 4083 323
rect 4136 307 4143 363
rect 4076 123 4083 253
rect 4116 167 4123 173
rect 4156 163 4163 343
rect 4216 267 4223 376
rect 4256 187 4263 363
rect 4136 156 4163 163
rect 4116 136 4123 153
rect 4136 127 4143 156
rect 4176 136 4183 153
rect 4216 136 4223 173
rect 4296 167 4303 873
rect 4316 787 4323 913
rect 4336 867 4343 1073
rect 4356 987 4363 1233
rect 4376 1227 4383 1293
rect 4396 1187 4403 1453
rect 4416 1163 4423 1473
rect 4436 1327 4443 1353
rect 4456 1327 4463 1613
rect 4476 1596 4483 1613
rect 4476 1327 4483 1393
rect 4496 1347 4503 1433
rect 4516 1307 4523 1513
rect 4536 1487 4543 1583
rect 4556 1527 4563 1553
rect 4576 1507 4583 1733
rect 4596 1467 4603 1653
rect 4616 1627 4623 1653
rect 4636 1627 4643 1756
rect 4656 1756 4683 1763
rect 4656 1707 4663 1756
rect 4676 1647 4683 1733
rect 4716 1687 4723 1783
rect 4736 1767 4743 1803
rect 4736 1687 4743 1713
rect 4616 1576 4623 1613
rect 4676 1603 4683 1633
rect 4676 1596 4703 1603
rect 4736 1596 4743 1613
rect 4756 1607 4763 1973
rect 4776 1847 4783 2016
rect 4836 1843 4843 1973
rect 4856 1927 4863 2053
rect 4896 2047 4903 2063
rect 4956 2027 4963 2193
rect 4976 2187 4983 2283
rect 4996 2263 5003 2413
rect 5036 2407 5043 2953
rect 5076 2947 5083 3036
rect 5056 2627 5063 2913
rect 5076 2767 5083 2813
rect 5056 2447 5063 2553
rect 5076 2547 5083 2753
rect 5076 2347 5083 2513
rect 5096 2467 5103 3093
rect 5116 3047 5123 3193
rect 5116 2827 5123 3013
rect 5116 2727 5123 2793
rect 4996 2256 5023 2263
rect 5016 2247 5023 2256
rect 4996 2203 5003 2233
rect 5036 2227 5043 2303
rect 5076 2296 5083 2313
rect 4996 2196 5023 2203
rect 4996 2096 5003 2173
rect 5016 2107 5023 2196
rect 4856 1867 4863 1893
rect 4836 1836 4863 1843
rect 4836 1787 4843 1803
rect 4656 1547 4663 1583
rect 4616 1407 4623 1513
rect 4676 1447 4683 1513
rect 4436 1247 4443 1273
rect 4456 1227 4463 1283
rect 4396 1156 4423 1163
rect 4376 1096 4383 1133
rect 4396 1116 4403 1156
rect 4476 1103 4483 1253
rect 4516 1207 4523 1253
rect 4536 1227 4543 1323
rect 4556 1187 4563 1313
rect 4576 1287 4583 1323
rect 4596 1227 4603 1293
rect 4616 1283 4623 1373
rect 4636 1347 4643 1373
rect 4636 1316 4643 1333
rect 4656 1327 4663 1413
rect 4676 1316 4683 1433
rect 4696 1343 4703 1553
rect 4716 1547 4723 1583
rect 4776 1567 4783 1713
rect 4796 1667 4803 1693
rect 4816 1667 4823 1783
rect 4796 1576 4803 1633
rect 4816 1607 4823 1613
rect 4836 1576 4843 1693
rect 4856 1627 4863 1836
rect 4876 1747 4883 2013
rect 4976 1947 4983 2013
rect 4916 1847 4923 1873
rect 4996 1867 5003 2053
rect 5016 2047 5023 2063
rect 4896 1816 4903 1833
rect 4716 1427 4723 1533
rect 4736 1367 4743 1553
rect 4696 1336 4723 1343
rect 4716 1303 4723 1336
rect 4756 1316 4763 1413
rect 4776 1347 4783 1533
rect 4836 1387 4843 1533
rect 4856 1507 4863 1563
rect 4876 1547 4883 1693
rect 4896 1663 4903 1733
rect 4916 1687 4923 1793
rect 4936 1787 4943 1813
rect 4956 1796 4983 1803
rect 4976 1767 4983 1796
rect 4996 1787 5003 1823
rect 5036 1816 5043 2033
rect 5056 1987 5063 2233
rect 5076 2047 5083 2253
rect 5096 2227 5103 2433
rect 4896 1656 4923 1663
rect 4896 1607 4903 1633
rect 4916 1627 4923 1656
rect 4987 1596 4993 1603
rect 4896 1543 4903 1593
rect 4936 1556 4943 1593
rect 4896 1536 4923 1543
rect 4916 1523 4923 1536
rect 4916 1516 4943 1523
rect 4896 1423 4903 1513
rect 4876 1416 4903 1423
rect 4796 1307 4803 1323
rect 4616 1276 4643 1283
rect 4396 847 4403 1073
rect 4416 1067 4423 1103
rect 4456 1096 4483 1103
rect 4436 1047 4443 1073
rect 4456 1047 4463 1096
rect 4496 1087 4503 1133
rect 4516 1107 4523 1153
rect 4556 1083 4563 1153
rect 4536 1076 4563 1083
rect 4416 843 4423 953
rect 4476 887 4483 1013
rect 4416 836 4443 843
rect 4336 767 4343 833
rect 4316 616 4323 733
rect 4356 727 4363 823
rect 4456 807 4463 863
rect 4496 856 4503 1013
rect 4516 883 4523 973
rect 4536 907 4543 933
rect 4516 876 4543 883
rect 4516 827 4523 853
rect 4536 727 4543 876
rect 4556 856 4563 993
rect 4576 927 4583 1213
rect 4636 1147 4643 1276
rect 4656 1247 4663 1283
rect 4656 1207 4663 1233
rect 4696 1203 4703 1303
rect 4716 1296 4743 1303
rect 4756 1247 4763 1273
rect 4676 1196 4703 1203
rect 4656 1127 4663 1133
rect 4616 1027 4623 1093
rect 4636 1047 4643 1103
rect 4656 867 4663 1053
rect 4676 887 4683 1196
rect 4696 1116 4703 1173
rect 4716 1147 4723 1233
rect 4756 1096 4763 1153
rect 4596 807 4603 853
rect 4616 827 4623 843
rect 4656 836 4663 853
rect 4696 827 4703 833
rect 4676 787 4683 823
rect 4336 656 4373 663
rect 4336 636 4343 656
rect 4376 636 4403 643
rect 4416 636 4423 673
rect 4456 636 4463 653
rect 4396 587 4403 636
rect 4396 467 4403 553
rect 4336 367 4343 393
rect 4496 387 4503 653
rect 4516 636 4523 673
rect 4556 636 4563 673
rect 4636 627 4643 733
rect 4576 616 4623 623
rect 4596 587 4603 616
rect 4656 616 4663 693
rect 4636 596 4643 613
rect 4676 487 4683 603
rect 4696 567 4703 713
rect 4396 356 4403 373
rect 4616 356 4623 393
rect 4636 367 4643 473
rect 4716 407 4723 873
rect 4776 867 4783 1303
rect 4816 1287 4823 1373
rect 4876 1367 4883 1416
rect 4796 947 4803 1273
rect 4816 1147 4823 1253
rect 4836 1187 4843 1323
rect 4856 1167 4863 1343
rect 4896 1336 4903 1393
rect 4876 1287 4883 1313
rect 4876 1187 4883 1253
rect 4896 1143 4903 1293
rect 4876 1136 4903 1143
rect 4916 1143 4923 1413
rect 4936 1367 4943 1516
rect 4956 1387 4963 1533
rect 4976 1487 4983 1563
rect 4996 1547 5003 1573
rect 4976 1407 4983 1453
rect 4996 1447 5003 1513
rect 5016 1467 5023 1733
rect 5036 1443 5043 1773
rect 5056 1727 5063 1933
rect 5076 1727 5083 1953
rect 5096 1923 5103 2213
rect 5116 1947 5123 2693
rect 5136 2647 5143 3313
rect 5096 1916 5123 1923
rect 5096 1767 5103 1833
rect 5076 1607 5083 1613
rect 5076 1576 5083 1593
rect 5096 1587 5103 1733
rect 5116 1667 5123 1916
rect 5136 1787 5143 2613
rect 5096 1556 5103 1573
rect 5056 1507 5063 1513
rect 5016 1436 5043 1443
rect 4976 1367 4983 1393
rect 4956 1327 4963 1343
rect 4996 1336 5003 1413
rect 4936 1167 4943 1323
rect 4916 1136 4943 1143
rect 4816 887 4823 1113
rect 4856 1067 4863 1103
rect 4876 907 4883 1093
rect 4896 1087 4903 1103
rect 4916 927 4923 1113
rect 4736 823 4743 853
rect 4776 836 4783 853
rect 4856 847 4863 863
rect 4896 856 4923 863
rect 4736 816 4763 823
rect 4836 807 4843 843
rect 4756 596 4763 693
rect 4776 616 4783 633
rect 4736 376 4763 383
rect 4656 356 4663 373
rect 4316 307 4323 323
rect 4336 147 4343 313
rect 4416 207 4423 343
rect 4496 287 4503 343
rect 4536 307 4543 313
rect 4416 143 4423 193
rect 4396 136 4423 143
rect 4556 136 4563 153
rect 4576 143 4583 193
rect 4596 187 4603 333
rect 4676 327 4683 353
rect 4756 347 4763 376
rect 4776 287 4783 573
rect 4816 403 4823 633
rect 4836 407 4843 793
rect 4856 667 4863 833
rect 4916 827 4923 856
rect 4936 827 4943 1136
rect 4956 1127 4963 1273
rect 4976 1267 4983 1323
rect 4976 1207 4983 1253
rect 4996 1163 5003 1293
rect 5016 1207 5023 1436
rect 5036 1287 5043 1373
rect 5056 1363 5063 1493
rect 5076 1427 5083 1533
rect 5096 1367 5103 1433
rect 5056 1356 5083 1363
rect 5076 1343 5083 1356
rect 5116 1347 5123 1533
rect 5136 1507 5143 1713
rect 5076 1336 5103 1343
rect 5056 1267 5063 1323
rect 5096 1316 5103 1336
rect 5076 1283 5083 1303
rect 5076 1276 5103 1283
rect 5076 1223 5083 1253
rect 5096 1227 5103 1276
rect 5116 1247 5123 1303
rect 5056 1216 5083 1223
rect 4996 1156 5023 1163
rect 4996 1076 5003 1133
rect 5016 1096 5023 1156
rect 5036 1087 5043 1173
rect 5056 1027 5063 1216
rect 4936 647 4943 653
rect 4876 607 4883 623
rect 4936 616 4943 633
rect 4956 607 4963 873
rect 4996 836 5003 1013
rect 5036 836 5043 913
rect 5056 807 5063 973
rect 4976 627 4983 673
rect 4996 583 5003 603
rect 4976 576 5003 583
rect 4976 407 4983 576
rect 4796 396 4823 403
rect 4736 167 4743 193
rect 4776 156 4783 233
rect 4796 167 4803 396
rect 4576 136 4603 143
rect 4676 136 4683 153
rect 4836 147 4843 353
rect 4856 347 4863 383
rect 4876 307 4883 363
rect 4856 136 4863 193
rect 4876 156 4883 273
rect 4896 207 4903 363
rect 4916 347 4923 383
rect 4996 363 5003 553
rect 5016 367 5023 753
rect 5076 387 5083 1193
rect 5096 1107 5103 1213
rect 5116 1067 5123 1213
rect 5136 987 5143 1413
rect 4976 356 5003 363
rect 4976 156 4983 356
rect 5076 327 5083 373
rect 5096 367 5103 893
rect 4996 136 5003 293
rect 3996 116 4023 123
rect 4056 116 4083 123
rect 4096 107 4103 123
rect 4236 116 4283 123
rect 4316 107 4323 123
rect 4376 103 4383 123
rect 4367 96 4383 103
rect 4096 87 4103 93
rect 4656 87 4663 123
rect 2656 -24 2683 -17
rect 2716 -24 2723 33
rect 5116 27 5123 933
rect 2876 -24 2883 13
rect 5036 -24 5043 13
<< m3contact >>
rect 1913 4813 1927 4827
rect 693 4753 707 4767
rect 773 4753 787 4767
rect 213 4713 227 4727
rect 33 4633 47 4647
rect 53 4493 67 4507
rect 93 4653 107 4667
rect 173 4673 187 4687
rect 273 4673 287 4687
rect 313 4673 327 4687
rect 353 4673 367 4687
rect 173 4653 187 4667
rect 193 4633 207 4647
rect 233 4633 247 4647
rect 133 4573 147 4587
rect 333 4573 347 4587
rect 393 4653 407 4667
rect 133 4533 147 4547
rect 113 4493 127 4507
rect 73 4473 87 4487
rect 93 4473 107 4487
rect 73 4433 87 4447
rect 33 4413 47 4427
rect 53 4413 67 4427
rect 193 4513 207 4527
rect 153 4473 167 4487
rect 113 4433 127 4447
rect 93 4413 107 4427
rect 233 4453 247 4467
rect 273 4453 287 4467
rect 333 4453 347 4467
rect 213 4433 227 4447
rect 253 4433 267 4447
rect 173 4373 187 4387
rect 73 4213 87 4227
rect 113 4213 127 4227
rect 133 4213 147 4227
rect 253 4253 267 4267
rect 313 4433 327 4447
rect 373 4533 387 4547
rect 493 4673 507 4687
rect 533 4673 547 4687
rect 573 4673 587 4687
rect 473 4653 487 4667
rect 453 4573 467 4587
rect 653 4673 667 4687
rect 733 4713 747 4727
rect 733 4673 747 4687
rect 753 4673 767 4687
rect 553 4653 567 4667
rect 633 4653 647 4667
rect 613 4633 627 4647
rect 673 4653 687 4667
rect 673 4633 687 4647
rect 713 4633 727 4647
rect 593 4613 607 4627
rect 533 4593 547 4607
rect 613 4593 627 4607
rect 593 4533 607 4547
rect 573 4513 587 4527
rect 513 4493 527 4507
rect 493 4473 507 4487
rect 433 4453 447 4467
rect 473 4453 487 4467
rect 413 4433 427 4447
rect 533 4453 547 4467
rect 1593 4733 1607 4747
rect 993 4713 1007 4727
rect 1453 4713 1467 4727
rect 773 4613 787 4627
rect 833 4653 847 4667
rect 753 4593 767 4607
rect 793 4593 807 4607
rect 673 4513 687 4527
rect 733 4513 747 4527
rect 613 4473 627 4487
rect 653 4473 667 4487
rect 713 4473 727 4487
rect 633 4453 647 4467
rect 793 4533 807 4547
rect 773 4513 787 4527
rect 753 4473 767 4487
rect 773 4473 787 4487
rect 833 4493 847 4507
rect 953 4673 967 4687
rect 1113 4693 1127 4707
rect 1253 4693 1267 4707
rect 1313 4693 1327 4707
rect 893 4653 907 4667
rect 973 4653 987 4667
rect 1013 4653 1027 4667
rect 1013 4633 1027 4647
rect 1033 4593 1047 4607
rect 933 4553 947 4567
rect 993 4553 1007 4567
rect 853 4473 867 4487
rect 433 4413 447 4427
rect 413 4393 427 4407
rect 393 4253 407 4267
rect 273 4233 287 4247
rect 53 4193 67 4207
rect 33 4173 47 4187
rect 93 4173 107 4187
rect 253 4213 267 4227
rect 293 4213 307 4227
rect 73 4153 87 4167
rect 113 4153 127 4167
rect 93 4033 107 4047
rect 73 3993 87 4007
rect 53 3973 67 3987
rect 133 3993 147 4007
rect 193 4173 207 4187
rect 273 4193 287 4207
rect 293 4193 307 4207
rect 233 4133 247 4147
rect 193 4013 207 4027
rect 273 4013 287 4027
rect 213 3993 227 4007
rect 253 3993 267 4007
rect 153 3973 167 3987
rect 173 3973 187 3987
rect 313 4173 327 4187
rect 373 4213 387 4227
rect 413 4193 427 4207
rect 413 4093 427 4107
rect 353 4013 367 4027
rect 333 3993 347 4007
rect 153 3953 167 3967
rect 233 3953 247 3967
rect 373 3973 387 3987
rect 393 3953 407 3967
rect 133 3913 147 3927
rect 113 3873 127 3887
rect 13 3813 27 3827
rect 33 3793 47 3807
rect 53 3753 67 3767
rect 33 3733 47 3747
rect 13 3713 27 3727
rect 33 3693 47 3707
rect 573 4433 587 4447
rect 733 4433 747 4447
rect 813 4453 827 4467
rect 873 4453 887 4467
rect 913 4453 927 4467
rect 853 4433 867 4447
rect 893 4433 907 4447
rect 753 4413 767 4427
rect 973 4533 987 4547
rect 953 4493 967 4507
rect 933 4433 947 4447
rect 913 4393 927 4407
rect 553 4373 567 4387
rect 873 4333 887 4347
rect 553 4253 567 4267
rect 453 4193 467 4207
rect 533 4193 547 4207
rect 473 4153 487 4167
rect 433 4033 447 4047
rect 453 4013 467 4027
rect 433 3993 447 4007
rect 473 3993 487 4007
rect 453 3953 467 3967
rect 313 3773 327 3787
rect 413 3773 427 3787
rect 173 3713 187 3727
rect 233 3713 247 3727
rect 133 3693 147 3707
rect 153 3673 167 3687
rect 73 3613 87 3627
rect 213 3693 227 3707
rect 193 3653 207 3667
rect 393 3753 407 3767
rect 353 3733 367 3747
rect 393 3713 407 3727
rect 473 3713 487 3727
rect 713 4233 727 4247
rect 813 4233 827 4247
rect 613 4213 627 4227
rect 573 4193 587 4207
rect 613 4173 627 4187
rect 673 4193 687 4207
rect 653 4173 667 4187
rect 593 4153 607 4167
rect 633 4153 647 4167
rect 693 4133 707 4147
rect 773 4193 787 4207
rect 933 4253 947 4267
rect 893 4213 907 4227
rect 873 4193 887 4207
rect 913 4193 927 4207
rect 973 4473 987 4487
rect 973 4453 987 4467
rect 1013 4453 1027 4467
rect 1073 4653 1087 4667
rect 1193 4673 1207 4687
rect 1233 4653 1247 4667
rect 1293 4653 1307 4667
rect 1113 4613 1127 4627
rect 1133 4613 1147 4627
rect 1093 4533 1107 4547
rect 1113 4533 1127 4547
rect 1073 4473 1087 4487
rect 1213 4633 1227 4647
rect 1273 4633 1287 4647
rect 1173 4613 1187 4627
rect 1293 4613 1307 4627
rect 1253 4533 1267 4547
rect 1153 4513 1167 4527
rect 1173 4513 1187 4527
rect 1233 4493 1247 4507
rect 1153 4473 1167 4487
rect 1193 4473 1207 4487
rect 1173 4453 1187 4467
rect 1273 4473 1287 4487
rect 1333 4673 1347 4687
rect 1353 4653 1367 4667
rect 1313 4493 1327 4507
rect 1333 4493 1347 4507
rect 1333 4473 1347 4487
rect 1433 4673 1447 4687
rect 1533 4673 1547 4687
rect 1453 4653 1467 4667
rect 1473 4653 1487 4667
rect 1413 4633 1427 4647
rect 1553 4633 1567 4647
rect 1493 4613 1507 4627
rect 1473 4593 1487 4607
rect 1493 4553 1507 4567
rect 1393 4533 1407 4547
rect 1373 4513 1387 4527
rect 1413 4473 1427 4487
rect 1853 4713 1867 4727
rect 1753 4693 1767 4707
rect 1653 4673 1667 4687
rect 1633 4653 1647 4667
rect 1613 4613 1627 4627
rect 1513 4493 1527 4507
rect 1593 4493 1607 4507
rect 1553 4473 1567 4487
rect 1373 4453 1387 4467
rect 1153 4433 1167 4447
rect 1213 4433 1227 4447
rect 1253 4433 1267 4447
rect 1313 4433 1327 4447
rect 1353 4433 1367 4447
rect 1133 4353 1147 4367
rect 1053 4333 1067 4347
rect 1133 4273 1147 4287
rect 953 4233 967 4247
rect 1033 4213 1047 4227
rect 993 4193 1007 4207
rect 753 4153 767 4167
rect 733 4133 747 4147
rect 633 4053 647 4067
rect 713 4053 727 4067
rect 773 4053 787 4067
rect 593 4033 607 4047
rect 553 3993 567 4007
rect 593 3973 607 3987
rect 673 4013 687 4027
rect 753 4013 767 4027
rect 573 3953 587 3967
rect 533 3893 547 3907
rect 673 3973 687 3987
rect 713 3973 727 3987
rect 653 3953 667 3967
rect 593 3833 607 3847
rect 533 3793 547 3807
rect 593 3793 607 3807
rect 513 3753 527 3767
rect 613 3753 627 3767
rect 533 3713 547 3727
rect 553 3713 567 3727
rect 593 3713 607 3727
rect 733 3953 747 3967
rect 693 3933 707 3947
rect 753 3933 767 3947
rect 733 3913 747 3927
rect 753 3913 767 3927
rect 713 3833 727 3847
rect 793 3853 807 3867
rect 753 3813 767 3827
rect 713 3793 727 3807
rect 333 3693 347 3707
rect 413 3693 427 3707
rect 453 3693 467 3707
rect 273 3673 287 3687
rect 313 3673 327 3687
rect 373 3673 387 3687
rect 533 3673 547 3687
rect 833 4173 847 4187
rect 933 4173 947 4187
rect 873 4153 887 4167
rect 913 4153 927 4167
rect 973 4113 987 4127
rect 1013 4113 1027 4127
rect 893 3993 907 4007
rect 933 3993 947 4007
rect 913 3933 927 3947
rect 833 3753 847 3767
rect 833 3733 847 3747
rect 853 3733 867 3747
rect 733 3713 747 3727
rect 773 3713 787 3727
rect 813 3713 827 3727
rect 893 3713 907 3727
rect 613 3673 627 3687
rect 593 3653 607 3667
rect 573 3593 587 3607
rect 253 3553 267 3567
rect 293 3553 307 3567
rect 393 3553 407 3567
rect 493 3553 507 3567
rect 153 3533 167 3547
rect 193 3533 207 3547
rect 333 3533 347 3547
rect 113 3353 127 3367
rect 353 3513 367 3527
rect 433 3513 447 3527
rect 93 3293 107 3307
rect 133 3293 147 3307
rect 53 3253 67 3267
rect 73 3173 87 3187
rect 53 3053 67 3067
rect 113 3273 127 3287
rect 113 3253 127 3267
rect 153 3253 167 3267
rect 293 3493 307 3507
rect 333 3493 347 3507
rect 373 3493 387 3507
rect 413 3493 427 3507
rect 453 3493 467 3507
rect 273 3453 287 3467
rect 213 3433 227 3447
rect 273 3433 287 3447
rect 133 3233 147 3247
rect 173 3233 187 3247
rect 193 3233 207 3247
rect 233 3233 247 3247
rect 193 3173 207 3187
rect 113 3073 127 3087
rect 173 3073 187 3087
rect 93 3033 107 3047
rect 153 3033 167 3047
rect 373 3473 387 3487
rect 393 3473 407 3487
rect 573 3533 587 3547
rect 533 3513 547 3527
rect 573 3513 587 3527
rect 513 3493 527 3507
rect 553 3493 567 3507
rect 313 3313 327 3327
rect 473 3473 487 3487
rect 493 3473 507 3487
rect 473 3453 487 3467
rect 413 3433 427 3447
rect 433 3433 447 3447
rect 393 3413 407 3427
rect 653 3573 667 3587
rect 673 3533 687 3547
rect 613 3513 627 3527
rect 633 3513 647 3527
rect 793 3693 807 3707
rect 873 3693 887 3707
rect 833 3653 847 3667
rect 933 3813 947 3827
rect 1093 4193 1107 4207
rect 1073 4133 1087 4147
rect 1113 4133 1127 4147
rect 1393 4393 1407 4407
rect 1433 4453 1447 4467
rect 1473 4433 1487 4447
rect 1573 4453 1587 4467
rect 1553 4413 1567 4427
rect 1533 4393 1547 4407
rect 1413 4373 1427 4387
rect 1453 4373 1467 4387
rect 1353 4253 1367 4267
rect 1373 4253 1387 4267
rect 1153 4233 1167 4247
rect 1213 4233 1227 4247
rect 1153 4193 1167 4207
rect 1193 4193 1207 4207
rect 1153 4173 1167 4187
rect 1213 4153 1227 4167
rect 1233 4153 1247 4167
rect 1173 4133 1187 4147
rect 1153 4113 1167 4127
rect 1133 4073 1147 4087
rect 1313 4193 1327 4207
rect 1333 4193 1347 4207
rect 1413 4233 1427 4247
rect 1533 4253 1547 4267
rect 1493 4233 1507 4247
rect 1513 4233 1527 4247
rect 1453 4213 1467 4227
rect 1413 4193 1427 4207
rect 1333 4173 1347 4187
rect 1293 4153 1307 4167
rect 1313 4153 1327 4167
rect 1273 4133 1287 4147
rect 1133 4013 1147 4027
rect 1213 4013 1227 4027
rect 1253 4013 1267 4027
rect 1133 3973 1147 3987
rect 1093 3953 1107 3967
rect 1113 3953 1127 3967
rect 1073 3933 1087 3947
rect 1093 3893 1107 3907
rect 1033 3833 1047 3847
rect 1013 3773 1027 3787
rect 1033 3773 1047 3787
rect 993 3733 1007 3747
rect 933 3713 947 3727
rect 993 3713 1007 3727
rect 953 3693 967 3707
rect 933 3673 947 3687
rect 1013 3673 1027 3687
rect 793 3633 807 3647
rect 813 3633 827 3647
rect 853 3633 867 3647
rect 873 3633 887 3647
rect 933 3653 947 3667
rect 973 3653 987 3667
rect 913 3633 927 3647
rect 873 3533 887 3547
rect 893 3533 907 3547
rect 613 3493 627 3507
rect 653 3493 667 3507
rect 713 3493 727 3507
rect 753 3493 767 3507
rect 693 3473 707 3487
rect 753 3473 767 3487
rect 733 3413 747 3427
rect 593 3333 607 3347
rect 393 3313 407 3327
rect 413 3313 427 3327
rect 513 3313 527 3327
rect 373 3293 387 3307
rect 413 3293 427 3307
rect 393 3273 407 3287
rect 353 3253 367 3267
rect 333 3233 347 3247
rect 693 3293 707 3307
rect 453 3273 467 3287
rect 513 3273 527 3287
rect 413 3253 427 3267
rect 453 3253 467 3267
rect 493 3253 507 3267
rect 533 3253 547 3267
rect 673 3253 687 3267
rect 813 3493 827 3507
rect 793 3473 807 3487
rect 773 3453 787 3467
rect 793 3433 807 3447
rect 753 3273 767 3287
rect 873 3493 887 3507
rect 893 3493 907 3507
rect 993 3633 1007 3647
rect 1013 3573 1027 3587
rect 1113 3873 1127 3887
rect 1133 3873 1147 3887
rect 1253 3973 1267 3987
rect 1273 3953 1287 3967
rect 1233 3933 1247 3947
rect 1233 3913 1247 3927
rect 1253 3873 1267 3887
rect 1273 3873 1287 3887
rect 1233 3853 1247 3867
rect 1133 3813 1147 3827
rect 1193 3813 1207 3827
rect 1113 3773 1127 3787
rect 1133 3773 1147 3787
rect 1093 3733 1107 3747
rect 1213 3753 1227 3767
rect 1073 3713 1087 3727
rect 1113 3713 1127 3727
rect 1153 3713 1167 3727
rect 1193 3713 1207 3727
rect 1053 3693 1067 3707
rect 1133 3693 1147 3707
rect 1133 3673 1147 3687
rect 1193 3693 1207 3707
rect 1093 3653 1107 3667
rect 1173 3653 1187 3667
rect 1073 3633 1087 3647
rect 1113 3633 1127 3647
rect 1033 3553 1047 3567
rect 1013 3533 1027 3547
rect 1033 3533 1047 3547
rect 1073 3533 1087 3547
rect 953 3513 967 3527
rect 973 3493 987 3507
rect 993 3493 1007 3507
rect 1013 3493 1027 3507
rect 1153 3513 1167 3527
rect 1093 3493 1107 3507
rect 1113 3493 1127 3507
rect 1133 3493 1147 3507
rect 933 3473 947 3487
rect 993 3433 1007 3447
rect 873 3413 887 3427
rect 953 3333 967 3347
rect 313 3213 327 3227
rect 253 3193 267 3207
rect 293 3193 307 3207
rect 273 3113 287 3127
rect 33 3013 47 3027
rect 93 3013 107 3027
rect 133 3013 147 3027
rect 173 2873 187 2887
rect 73 2813 87 2827
rect 33 2753 47 2767
rect 93 2753 107 2767
rect 133 2753 147 2767
rect 153 2733 167 2747
rect 113 2693 127 2707
rect 213 2993 227 3007
rect 253 2853 267 2867
rect 213 2753 227 2767
rect 373 3073 387 3087
rect 373 3053 387 3067
rect 393 3053 407 3067
rect 513 3233 527 3247
rect 553 3233 567 3247
rect 593 3233 607 3247
rect 473 3193 487 3207
rect 533 3193 547 3207
rect 493 3113 507 3127
rect 433 3013 447 3027
rect 573 3193 587 3207
rect 553 3113 567 3127
rect 313 2993 327 3007
rect 353 2993 367 3007
rect 413 2993 427 3007
rect 293 2893 307 2907
rect 353 2833 367 2847
rect 473 2893 487 2907
rect 633 3153 647 3167
rect 613 3053 627 3067
rect 573 3013 587 3027
rect 533 2933 547 2947
rect 513 2813 527 2827
rect 673 3053 687 3067
rect 813 3253 827 3267
rect 853 3253 867 3267
rect 893 3253 907 3267
rect 773 3233 787 3247
rect 853 3233 867 3247
rect 753 3213 767 3227
rect 793 3213 807 3227
rect 773 3193 787 3207
rect 753 3173 767 3187
rect 833 3173 847 3187
rect 913 3213 927 3227
rect 873 3193 887 3207
rect 853 3133 867 3147
rect 1073 3373 1087 3387
rect 953 3193 967 3207
rect 933 3173 947 3187
rect 913 3133 927 3147
rect 953 3133 967 3147
rect 873 3073 887 3087
rect 793 3053 807 3067
rect 713 3033 727 3047
rect 633 2933 647 2947
rect 813 3033 827 3047
rect 1033 3273 1047 3287
rect 993 3193 1007 3207
rect 993 3153 1007 3167
rect 1053 3213 1067 3227
rect 1013 3113 1027 3127
rect 1273 3833 1287 3847
rect 1353 4133 1367 4147
rect 1393 4113 1407 4127
rect 1413 4113 1427 4127
rect 1433 4113 1447 4127
rect 1313 4073 1327 4087
rect 1333 4073 1347 4087
rect 1393 4053 1407 4067
rect 1353 3993 1367 4007
rect 1473 4153 1487 4167
rect 1453 4013 1467 4027
rect 1453 3993 1467 4007
rect 1493 3993 1507 4007
rect 1333 3973 1347 3987
rect 1373 3973 1387 3987
rect 1313 3953 1327 3967
rect 1393 3953 1407 3967
rect 1293 3793 1307 3807
rect 1273 3753 1287 3767
rect 1313 3773 1327 3787
rect 1273 3713 1287 3727
rect 1273 3693 1287 3707
rect 1293 3693 1307 3707
rect 1313 3693 1327 3707
rect 1233 3673 1247 3687
rect 1253 3513 1267 3527
rect 1193 3453 1207 3467
rect 1233 3373 1247 3387
rect 1173 3313 1187 3327
rect 1333 3673 1347 3687
rect 1313 3633 1327 3647
rect 1473 3973 1487 3987
rect 1433 3933 1447 3947
rect 1533 4213 1547 4227
rect 1533 4153 1547 4167
rect 1633 4493 1647 4507
rect 1733 4653 1747 4667
rect 2433 4813 2447 4827
rect 2473 4753 2487 4767
rect 2393 4733 2407 4747
rect 1993 4713 2007 4727
rect 2053 4713 2067 4727
rect 2193 4713 2207 4727
rect 2293 4713 2307 4727
rect 1773 4653 1787 4667
rect 1833 4653 1847 4667
rect 1873 4653 1887 4667
rect 1713 4633 1727 4647
rect 1753 4633 1767 4647
rect 1693 4493 1707 4507
rect 1913 4593 1927 4607
rect 1953 4633 1967 4647
rect 2093 4673 2107 4687
rect 2133 4673 2147 4687
rect 2173 4673 2187 4687
rect 1973 4613 1987 4627
rect 1993 4613 2007 4627
rect 1813 4553 1827 4567
rect 1933 4553 1947 4567
rect 2113 4653 2127 4667
rect 2153 4653 2167 4667
rect 2033 4633 2047 4647
rect 2073 4633 2087 4647
rect 1993 4533 2007 4547
rect 2013 4533 2027 4547
rect 1833 4513 1847 4527
rect 1753 4493 1767 4507
rect 1713 4453 1727 4467
rect 1733 4453 1747 4467
rect 1653 4413 1667 4427
rect 1633 4393 1647 4407
rect 1573 4293 1587 4307
rect 1613 4293 1627 4307
rect 1713 4433 1727 4447
rect 1793 4453 1807 4467
rect 1773 4413 1787 4427
rect 1813 4413 1827 4427
rect 1673 4393 1687 4407
rect 1753 4393 1767 4407
rect 1893 4473 1907 4487
rect 1933 4473 1947 4487
rect 2013 4473 2027 4487
rect 1873 4453 1887 4467
rect 1913 4453 1927 4467
rect 1973 4453 1987 4467
rect 1913 4413 1927 4427
rect 1833 4373 1847 4387
rect 1753 4353 1767 4367
rect 1793 4353 1807 4367
rect 1613 4233 1627 4247
rect 1653 4233 1667 4247
rect 1693 4233 1707 4247
rect 1613 4213 1627 4227
rect 1593 4193 1607 4207
rect 1653 4193 1667 4207
rect 1793 4253 1807 4267
rect 1853 4253 1867 4267
rect 1753 4193 1767 4207
rect 1833 4233 1847 4247
rect 1573 4173 1587 4187
rect 1613 4173 1627 4187
rect 1553 4133 1567 4147
rect 1593 4113 1607 4127
rect 1553 3993 1567 4007
rect 1573 3993 1587 4007
rect 1533 3953 1547 3967
rect 1513 3913 1527 3927
rect 1513 3853 1527 3867
rect 1473 3773 1487 3787
rect 1433 3733 1447 3747
rect 1453 3713 1467 3727
rect 1513 3773 1527 3787
rect 1573 3913 1587 3927
rect 1553 3833 1567 3847
rect 1533 3733 1547 3747
rect 1513 3713 1527 3727
rect 1693 4153 1707 4167
rect 1673 4133 1687 4147
rect 1613 4093 1627 4107
rect 1633 4093 1647 4107
rect 1713 4133 1727 4147
rect 1753 4153 1767 4167
rect 1733 4113 1747 4127
rect 1673 4053 1687 4067
rect 1693 4053 1707 4067
rect 1733 4033 1747 4047
rect 1713 4013 1727 4027
rect 1653 3973 1667 3987
rect 1613 3953 1627 3967
rect 1633 3953 1647 3967
rect 1653 3913 1667 3927
rect 1613 3773 1627 3787
rect 1593 3733 1607 3747
rect 1633 3733 1647 3747
rect 1713 3893 1727 3907
rect 1773 4133 1787 4147
rect 1773 3993 1787 4007
rect 1853 4213 1867 4227
rect 1893 4213 1907 4227
rect 1993 4433 2007 4447
rect 1953 4373 1967 4387
rect 1973 4293 1987 4307
rect 1933 4233 1947 4247
rect 1833 4133 1847 4147
rect 1833 4053 1847 4067
rect 1833 3993 1847 4007
rect 1913 4173 1927 4187
rect 2093 4593 2107 4607
rect 2073 4553 2087 4567
rect 2073 4473 2087 4487
rect 2113 4513 2127 4527
rect 2093 4453 2107 4467
rect 2233 4693 2247 4707
rect 2273 4693 2287 4707
rect 2253 4673 2267 4687
rect 2193 4653 2207 4667
rect 2233 4653 2247 4667
rect 2173 4613 2187 4627
rect 2133 4493 2147 4507
rect 2213 4473 2227 4487
rect 2313 4693 2327 4707
rect 2333 4673 2347 4687
rect 2333 4653 2347 4667
rect 2333 4633 2347 4647
rect 2373 4633 2387 4647
rect 2273 4613 2287 4627
rect 2273 4533 2287 4547
rect 2313 4493 2327 4507
rect 2173 4453 2187 4467
rect 2253 4453 2267 4467
rect 2293 4453 2307 4467
rect 2093 4433 2107 4447
rect 2133 4433 2147 4447
rect 2073 4413 2087 4427
rect 2193 4433 2207 4447
rect 2213 4433 2227 4447
rect 2293 4433 2307 4447
rect 2313 4433 2327 4447
rect 2053 4393 2067 4407
rect 2033 4353 2047 4367
rect 2153 4313 2167 4327
rect 2093 4293 2107 4307
rect 2073 4213 2087 4227
rect 1913 4033 1927 4047
rect 1753 3953 1767 3967
rect 1793 3953 1807 3967
rect 1813 3953 1827 3967
rect 1753 3933 1767 3947
rect 1713 3873 1727 3887
rect 1733 3873 1747 3887
rect 1693 3833 1707 3847
rect 1393 3653 1407 3667
rect 1413 3593 1427 3607
rect 1373 3573 1387 3587
rect 1353 3553 1367 3567
rect 1333 3533 1347 3547
rect 1353 3533 1367 3547
rect 1393 3553 1407 3567
rect 1313 3433 1327 3447
rect 1333 3333 1347 3347
rect 1113 3273 1127 3287
rect 1233 3273 1247 3287
rect 1293 3273 1307 3287
rect 1093 3233 1107 3247
rect 1133 3233 1147 3247
rect 1093 3213 1107 3227
rect 1113 3193 1127 3207
rect 973 3053 987 3067
rect 1033 3053 1047 3067
rect 1013 3033 1027 3047
rect 753 3013 767 3027
rect 793 3013 807 3027
rect 773 2993 787 3007
rect 833 3013 847 3027
rect 933 3013 947 3027
rect 953 3013 967 3027
rect 853 2993 867 3007
rect 353 2793 367 2807
rect 433 2793 447 2807
rect 533 2793 547 2807
rect 593 2793 607 2807
rect 653 2793 667 2807
rect 673 2793 687 2807
rect 893 2793 907 2807
rect 293 2773 307 2787
rect 193 2733 207 2747
rect 293 2733 307 2747
rect 373 2773 387 2787
rect 393 2773 407 2787
rect 413 2773 427 2787
rect 353 2753 367 2767
rect 233 2713 247 2727
rect 313 2713 327 2727
rect 433 2753 447 2767
rect 513 2773 527 2787
rect 473 2753 487 2767
rect 453 2733 467 2747
rect 533 2713 547 2727
rect 573 2713 587 2727
rect 653 2773 667 2787
rect 693 2773 707 2787
rect 733 2773 747 2787
rect 793 2773 807 2787
rect 673 2753 687 2767
rect 633 2733 647 2747
rect 913 2773 927 2787
rect 993 2973 1007 2987
rect 993 2953 1007 2967
rect 1073 3093 1087 3107
rect 1173 3193 1187 3207
rect 1213 3193 1227 3207
rect 1373 3293 1387 3307
rect 1433 3553 1447 3567
rect 1533 3693 1547 3707
rect 1493 3673 1507 3687
rect 1553 3673 1567 3687
rect 1433 3533 1447 3547
rect 1473 3533 1487 3547
rect 1433 3493 1447 3507
rect 1373 3253 1387 3267
rect 1393 3253 1407 3267
rect 1273 3233 1287 3247
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1153 3073 1167 3087
rect 1233 3073 1247 3087
rect 1093 3053 1107 3067
rect 1173 3053 1187 3067
rect 1233 3053 1247 3067
rect 1113 3033 1127 3047
rect 1133 3013 1147 3027
rect 1113 2993 1127 3007
rect 1133 2973 1147 2987
rect 1073 2893 1087 2907
rect 1053 2873 1067 2887
rect 1133 2873 1147 2887
rect 1013 2853 1027 2867
rect 1133 2833 1147 2847
rect 1133 2813 1147 2827
rect 1113 2793 1127 2807
rect 1013 2773 1027 2787
rect 953 2753 967 2767
rect 993 2753 1007 2767
rect 1033 2753 1047 2767
rect 973 2733 987 2747
rect 1033 2733 1047 2747
rect 1093 2753 1107 2767
rect 1193 3033 1207 3047
rect 1213 3033 1227 3047
rect 1293 3193 1307 3207
rect 1293 3153 1307 3167
rect 1293 3053 1307 3067
rect 1273 3033 1287 3047
rect 1313 3033 1327 3047
rect 1293 3013 1307 3027
rect 1193 2973 1207 2987
rect 1173 2933 1187 2947
rect 1393 3213 1407 3227
rect 1393 3173 1407 3187
rect 1473 3473 1487 3487
rect 1473 3433 1487 3447
rect 1473 3413 1487 3427
rect 1453 3233 1467 3247
rect 1433 3193 1447 3207
rect 1433 3153 1447 3167
rect 1413 3073 1427 3087
rect 1533 3593 1547 3607
rect 1513 3573 1527 3587
rect 1593 3693 1607 3707
rect 1573 3573 1587 3587
rect 1553 3553 1567 3567
rect 1893 3993 1907 4007
rect 1893 3973 1907 3987
rect 1873 3953 1887 3967
rect 1933 3993 1947 4007
rect 1993 4173 2007 4187
rect 1993 4133 2007 4147
rect 1973 4013 1987 4027
rect 1953 3973 1967 3987
rect 2053 4193 2067 4207
rect 2033 4173 2047 4187
rect 2113 4193 2127 4207
rect 2013 4053 2027 4067
rect 2133 4133 2147 4147
rect 2193 4373 2207 4387
rect 2253 4293 2267 4307
rect 2173 4233 2187 4247
rect 2173 4213 2187 4227
rect 2173 4153 2187 4167
rect 2193 4153 2207 4167
rect 2273 4173 2287 4187
rect 2313 4393 2327 4407
rect 2553 4693 2567 4707
rect 2973 4813 2987 4827
rect 3173 4813 3187 4827
rect 2713 4713 2727 4727
rect 2433 4673 2447 4687
rect 2473 4673 2487 4687
rect 2513 4673 2527 4687
rect 2593 4673 2607 4687
rect 2453 4653 2467 4667
rect 2493 4653 2507 4667
rect 2373 4593 2387 4607
rect 2353 4513 2367 4527
rect 2353 4473 2367 4487
rect 2413 4473 2427 4487
rect 2353 4453 2367 4467
rect 2393 4453 2407 4467
rect 2533 4613 2547 4627
rect 2493 4593 2507 4607
rect 2513 4593 2527 4607
rect 2493 4493 2507 4507
rect 2433 4433 2447 4447
rect 2673 4693 2687 4707
rect 2653 4673 2667 4687
rect 2693 4673 2707 4687
rect 2613 4633 2627 4647
rect 2613 4593 2627 4607
rect 2573 4573 2587 4587
rect 2553 4493 2567 4507
rect 2453 4413 2467 4427
rect 2413 4273 2427 4287
rect 2433 4273 2447 4287
rect 2313 4213 2327 4227
rect 2153 4093 2167 4107
rect 2173 4093 2187 4107
rect 2153 4053 2167 4067
rect 2213 4053 2227 4067
rect 2033 3993 2047 4007
rect 2073 4013 2087 4027
rect 2133 4013 2147 4027
rect 1953 3953 1967 3967
rect 1913 3893 1927 3907
rect 1753 3833 1767 3847
rect 1833 3833 1847 3847
rect 1853 3833 1867 3847
rect 1893 3833 1907 3847
rect 1713 3733 1727 3747
rect 1773 3773 1787 3787
rect 1753 3693 1767 3707
rect 1613 3653 1627 3667
rect 1633 3653 1647 3667
rect 1693 3653 1707 3667
rect 1793 3733 1807 3747
rect 1833 3713 1847 3727
rect 1873 3713 1887 3727
rect 1773 3653 1787 3667
rect 1833 3653 1847 3667
rect 1613 3553 1627 3567
rect 1673 3553 1687 3567
rect 1593 3533 1607 3547
rect 1613 3513 1627 3527
rect 1653 3513 1667 3527
rect 1533 3493 1547 3507
rect 1553 3473 1567 3487
rect 1593 3473 1607 3487
rect 1533 3453 1547 3467
rect 1493 3373 1507 3387
rect 1513 3233 1527 3247
rect 1713 3513 1727 3527
rect 1753 3513 1767 3527
rect 1633 3453 1647 3467
rect 1673 3453 1687 3467
rect 1693 3453 1707 3467
rect 1733 3453 1747 3467
rect 1593 3433 1607 3447
rect 1633 3433 1647 3447
rect 1613 3393 1627 3407
rect 1533 3213 1547 3227
rect 1633 3253 1647 3267
rect 1693 3253 1707 3267
rect 1633 3213 1647 3227
rect 1573 3173 1587 3187
rect 1473 3093 1487 3107
rect 1493 3093 1507 3107
rect 1493 3073 1507 3087
rect 1453 3053 1467 3067
rect 1473 3053 1487 3067
rect 1373 3033 1387 3047
rect 1433 3033 1447 3047
rect 1553 3053 1567 3067
rect 1613 3053 1627 3067
rect 1433 3013 1447 3027
rect 1373 2993 1387 3007
rect 1533 3033 1547 3047
rect 1553 3013 1567 3027
rect 1433 2973 1447 2987
rect 1513 2973 1527 2987
rect 1293 2913 1307 2927
rect 1333 2893 1347 2907
rect 1293 2813 1307 2827
rect 1153 2793 1167 2807
rect 1233 2793 1247 2807
rect 1173 2773 1187 2787
rect 1213 2773 1227 2787
rect 853 2713 867 2727
rect 873 2713 887 2727
rect 1013 2713 1027 2727
rect 1053 2713 1067 2727
rect 593 2693 607 2707
rect 713 2693 727 2707
rect 813 2693 827 2707
rect 993 2673 1007 2687
rect 873 2653 887 2667
rect 833 2633 847 2647
rect 13 2593 27 2607
rect 173 2593 187 2607
rect 293 2593 307 2607
rect 633 2593 647 2607
rect 73 2553 87 2567
rect 33 2513 47 2527
rect 233 2573 247 2587
rect 293 2573 307 2587
rect 453 2573 467 2587
rect 493 2573 507 2587
rect 553 2573 567 2587
rect 593 2573 607 2587
rect 193 2553 207 2567
rect 393 2553 407 2567
rect 313 2533 327 2547
rect 373 2533 387 2547
rect 53 2273 67 2287
rect 113 2273 127 2287
rect 93 2253 107 2267
rect 33 2233 47 2247
rect 73 2233 87 2247
rect 133 2213 147 2227
rect 253 2513 267 2527
rect 353 2333 367 2347
rect 213 2273 227 2287
rect 173 2253 187 2267
rect 233 2253 247 2267
rect 153 2113 167 2127
rect 133 2093 147 2107
rect 93 2073 107 2087
rect 53 2033 67 2047
rect 193 2053 207 2067
rect 113 2033 127 2047
rect 153 2033 167 2047
rect 173 2033 187 2047
rect 213 2013 227 2027
rect 313 2253 327 2267
rect 373 2253 387 2267
rect 513 2553 527 2567
rect 613 2553 627 2567
rect 473 2533 487 2547
rect 473 2513 487 2527
rect 573 2533 587 2547
rect 653 2573 667 2587
rect 673 2553 687 2567
rect 773 2553 787 2567
rect 813 2553 827 2567
rect 633 2533 647 2547
rect 653 2533 667 2547
rect 713 2533 727 2547
rect 733 2533 747 2547
rect 653 2513 667 2527
rect 693 2513 707 2527
rect 533 2493 547 2507
rect 593 2493 607 2507
rect 613 2493 627 2507
rect 633 2493 647 2507
rect 513 2473 527 2487
rect 453 2413 467 2427
rect 493 2413 507 2427
rect 253 2193 267 2207
rect 393 2233 407 2247
rect 413 2193 427 2207
rect 273 2153 287 2167
rect 393 2153 407 2167
rect 353 2093 367 2107
rect 313 2073 327 2087
rect 253 2033 267 2047
rect 293 2033 307 2047
rect 473 2293 487 2307
rect 453 2273 467 2287
rect 433 2153 447 2167
rect 473 2153 487 2167
rect 433 2113 447 2127
rect 413 2093 427 2107
rect 373 2033 387 2047
rect 313 2013 327 2027
rect 273 1993 287 2007
rect 233 1973 247 1987
rect 173 1833 187 1847
rect 53 1813 67 1827
rect 93 1813 107 1827
rect 73 1793 87 1807
rect 113 1793 127 1807
rect 153 1793 167 1807
rect 53 1773 67 1787
rect 33 1753 47 1767
rect 73 1753 87 1767
rect 93 1753 107 1767
rect 33 1733 47 1747
rect 133 1773 147 1787
rect 153 1773 167 1787
rect 113 1613 127 1627
rect 213 1793 227 1807
rect 213 1773 227 1787
rect 193 1753 207 1767
rect 173 1613 187 1627
rect 153 1593 167 1607
rect 293 1833 307 1847
rect 253 1793 267 1807
rect 253 1773 267 1787
rect 233 1733 247 1747
rect 53 1553 67 1567
rect 73 1553 87 1567
rect 13 1393 27 1407
rect 13 1353 27 1367
rect 73 1353 87 1367
rect 13 1333 27 1347
rect 53 1333 67 1347
rect 33 1313 47 1327
rect 13 1293 27 1307
rect 53 1293 67 1307
rect 33 1273 47 1287
rect 73 1273 87 1287
rect 13 1233 27 1247
rect 53 1213 67 1227
rect 33 1173 47 1187
rect 13 1093 27 1107
rect 93 1253 107 1267
rect 213 1573 227 1587
rect 153 1553 167 1567
rect 233 1553 247 1567
rect 213 1333 227 1347
rect 373 1993 387 2007
rect 413 1993 427 2007
rect 373 1853 387 1867
rect 333 1833 347 1847
rect 453 2073 467 2087
rect 473 2073 487 2087
rect 573 2353 587 2367
rect 533 2273 547 2287
rect 553 2273 567 2287
rect 753 2513 767 2527
rect 793 2513 807 2527
rect 813 2473 827 2487
rect 713 2333 727 2347
rect 753 2313 767 2327
rect 733 2293 747 2307
rect 913 2613 927 2627
rect 853 2533 867 2547
rect 973 2593 987 2607
rect 1093 2673 1107 2687
rect 1013 2593 1027 2607
rect 1033 2593 1047 2607
rect 1053 2533 1067 2547
rect 913 2513 927 2527
rect 933 2513 947 2527
rect 1033 2513 1047 2527
rect 1073 2513 1087 2527
rect 1073 2493 1087 2507
rect 673 2273 687 2287
rect 713 2273 727 2287
rect 513 2253 527 2267
rect 593 2253 607 2267
rect 613 2213 627 2227
rect 673 2253 687 2267
rect 653 2193 667 2207
rect 653 2153 667 2167
rect 653 2133 667 2147
rect 533 2093 547 2107
rect 573 2093 587 2107
rect 633 2093 647 2107
rect 533 2073 547 2087
rect 473 2053 487 2067
rect 513 2053 527 2067
rect 553 2033 567 2047
rect 693 2053 707 2067
rect 713 2033 727 2047
rect 453 2013 467 2027
rect 593 2013 607 2027
rect 673 2013 687 2027
rect 453 1993 467 2007
rect 433 1833 447 1847
rect 373 1813 387 1827
rect 353 1793 367 1807
rect 393 1773 407 1787
rect 673 1973 687 1987
rect 473 1853 487 1867
rect 433 1793 447 1807
rect 293 1733 307 1747
rect 313 1733 327 1747
rect 333 1733 347 1747
rect 413 1733 427 1747
rect 313 1693 327 1707
rect 273 1633 287 1647
rect 293 1613 307 1627
rect 313 1353 327 1367
rect 493 1833 507 1847
rect 613 1833 627 1847
rect 473 1693 487 1707
rect 433 1673 447 1687
rect 413 1653 427 1667
rect 353 1633 367 1647
rect 373 1593 387 1607
rect 393 1493 407 1507
rect 353 1393 367 1407
rect 133 1313 147 1327
rect 193 1313 207 1327
rect 233 1313 247 1327
rect 253 1313 267 1327
rect 173 1293 187 1307
rect 213 1293 227 1307
rect 113 1233 127 1247
rect 153 1233 167 1247
rect 113 1213 127 1227
rect 93 1113 107 1127
rect 133 1113 147 1127
rect 73 1093 87 1107
rect 53 793 67 807
rect 293 1313 307 1327
rect 313 1313 327 1327
rect 273 1233 287 1247
rect 473 1653 487 1667
rect 573 1813 587 1827
rect 653 1813 667 1827
rect 533 1793 547 1807
rect 593 1793 607 1807
rect 513 1753 527 1767
rect 553 1733 567 1747
rect 593 1713 607 1727
rect 513 1693 527 1707
rect 493 1593 507 1607
rect 473 1573 487 1587
rect 493 1573 507 1587
rect 453 1553 467 1567
rect 693 1833 707 1847
rect 673 1753 687 1767
rect 833 2293 847 2307
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 793 2173 807 2187
rect 773 2153 787 2167
rect 793 2113 807 2127
rect 933 2273 947 2287
rect 1013 2273 1027 2287
rect 1053 2273 1067 2287
rect 953 2253 967 2267
rect 993 2253 1007 2267
rect 1093 2273 1107 2287
rect 1053 2233 1067 2247
rect 993 2213 1007 2227
rect 913 2173 927 2187
rect 873 2153 887 2167
rect 833 2093 847 2107
rect 833 2073 847 2087
rect 893 2093 907 2107
rect 773 2033 787 2047
rect 813 2033 827 2047
rect 933 2133 947 2147
rect 953 2093 967 2107
rect 973 2073 987 2087
rect 853 2013 867 2027
rect 853 1913 867 1927
rect 733 1853 747 1867
rect 793 1813 807 1827
rect 713 1793 727 1807
rect 913 1813 927 1827
rect 813 1793 827 1807
rect 853 1793 867 1807
rect 953 1793 967 1807
rect 733 1773 747 1787
rect 693 1733 707 1747
rect 673 1693 687 1707
rect 533 1613 547 1627
rect 593 1613 607 1627
rect 633 1613 647 1627
rect 573 1593 587 1607
rect 473 1533 487 1547
rect 553 1533 567 1547
rect 373 1353 387 1367
rect 433 1353 447 1367
rect 353 1213 367 1227
rect 333 1153 347 1167
rect 633 1573 647 1587
rect 793 1773 807 1787
rect 813 1773 827 1787
rect 753 1733 767 1747
rect 773 1733 787 1747
rect 773 1673 787 1687
rect 713 1633 727 1647
rect 733 1633 747 1647
rect 773 1633 787 1647
rect 753 1593 767 1607
rect 833 1753 847 1767
rect 893 1773 907 1787
rect 893 1733 907 1747
rect 973 1753 987 1767
rect 973 1733 987 1747
rect 973 1713 987 1727
rect 933 1693 947 1707
rect 873 1653 887 1667
rect 913 1653 927 1667
rect 833 1633 847 1647
rect 813 1613 827 1627
rect 773 1573 787 1587
rect 653 1533 667 1547
rect 573 1513 587 1527
rect 733 1553 747 1567
rect 753 1533 767 1547
rect 693 1513 707 1527
rect 653 1493 667 1507
rect 633 1353 647 1367
rect 453 1333 467 1347
rect 553 1333 567 1347
rect 413 1313 427 1327
rect 393 1293 407 1307
rect 493 1313 507 1327
rect 533 1313 547 1327
rect 453 1273 467 1287
rect 513 1273 527 1287
rect 433 1253 447 1267
rect 473 1253 487 1267
rect 493 1253 507 1267
rect 393 1173 407 1187
rect 393 1153 407 1167
rect 373 1133 387 1147
rect 273 1113 287 1127
rect 433 1113 447 1127
rect 173 1093 187 1107
rect 233 1093 247 1107
rect 273 1093 287 1107
rect 373 1093 387 1107
rect 293 1073 307 1087
rect 293 953 307 967
rect 333 953 347 967
rect 93 833 107 847
rect 193 853 207 867
rect 233 853 247 867
rect 253 853 267 867
rect 193 833 207 847
rect 173 813 187 827
rect 133 793 147 807
rect 113 753 127 767
rect 73 653 87 667
rect 33 633 47 647
rect 13 533 27 547
rect 13 513 27 527
rect 133 693 147 707
rect 253 833 267 847
rect 233 793 247 807
rect 273 793 287 807
rect 213 773 227 787
rect 453 1093 467 1107
rect 413 1053 427 1067
rect 373 873 387 887
rect 613 1313 627 1327
rect 613 1293 627 1307
rect 713 1313 727 1327
rect 693 1293 707 1307
rect 733 1293 747 1307
rect 633 1273 647 1287
rect 833 1593 847 1607
rect 873 1593 887 1607
rect 933 1613 947 1627
rect 953 1613 967 1627
rect 1153 2733 1167 2747
rect 1173 2733 1187 2747
rect 1193 2693 1207 2707
rect 1253 2773 1267 2787
rect 1293 2773 1307 2787
rect 1273 2713 1287 2727
rect 1233 2593 1247 2607
rect 1193 2553 1207 2567
rect 1253 2553 1267 2567
rect 1213 2533 1227 2547
rect 1273 2533 1287 2547
rect 1293 2533 1307 2547
rect 1313 2533 1327 2547
rect 1133 2273 1147 2287
rect 1173 2253 1187 2267
rect 1293 2273 1307 2287
rect 1153 2233 1167 2247
rect 1113 2213 1127 2227
rect 1133 2213 1147 2227
rect 1093 2133 1107 2147
rect 1073 2053 1087 2067
rect 1073 2033 1087 2047
rect 1113 2033 1127 2047
rect 1013 1833 1027 1847
rect 1153 2093 1167 2107
rect 1213 2233 1227 2247
rect 1213 2133 1227 2147
rect 1233 2113 1247 2127
rect 1293 2173 1307 2187
rect 1253 2093 1267 2107
rect 1253 2073 1267 2087
rect 1493 2853 1507 2867
rect 1393 2773 1407 2787
rect 1433 2773 1447 2787
rect 1373 2753 1387 2767
rect 1353 2713 1367 2727
rect 1473 2753 1487 2767
rect 1413 2733 1427 2747
rect 1373 2553 1387 2567
rect 1533 2813 1547 2827
rect 1793 3513 1807 3527
rect 1793 3473 1807 3487
rect 1813 3473 1827 3487
rect 1873 3653 1887 3667
rect 1873 3613 1887 3627
rect 1853 3573 1867 3587
rect 1873 3553 1887 3567
rect 1853 3513 1867 3527
rect 2113 3973 2127 3987
rect 1973 3933 1987 3947
rect 2013 3933 2027 3947
rect 2133 3933 2147 3947
rect 2193 4033 2207 4047
rect 2193 4013 2207 4027
rect 2293 4153 2307 4167
rect 2333 4153 2347 4167
rect 2413 4233 2427 4247
rect 2413 4213 2427 4227
rect 2353 4113 2367 4127
rect 2293 4013 2307 4027
rect 2313 4013 2327 4027
rect 2173 3973 2187 3987
rect 2233 3973 2247 3987
rect 2373 4013 2387 4027
rect 2213 3933 2227 3947
rect 2293 3933 2307 3947
rect 2153 3913 2167 3927
rect 2173 3913 2187 3927
rect 2053 3853 2067 3867
rect 2033 3833 2047 3847
rect 1953 3773 1967 3787
rect 1973 3773 1987 3787
rect 1913 3713 1927 3727
rect 1933 3693 1947 3707
rect 2033 3733 2047 3747
rect 2073 3813 2087 3827
rect 2073 3733 2087 3747
rect 2153 3733 2167 3747
rect 2093 3713 2107 3727
rect 2033 3693 2047 3707
rect 2073 3693 2087 3707
rect 2013 3553 2027 3567
rect 1973 3533 1987 3547
rect 1913 3513 1927 3527
rect 1953 3513 1967 3527
rect 2133 3693 2147 3707
rect 2113 3613 2127 3627
rect 2093 3573 2107 3587
rect 2073 3553 2087 3567
rect 2033 3533 2047 3547
rect 2053 3513 2067 3527
rect 1873 3473 1887 3487
rect 1933 3473 1947 3487
rect 1953 3473 1967 3487
rect 1773 3393 1787 3407
rect 1793 3393 1807 3407
rect 1773 3353 1787 3367
rect 1833 3353 1847 3367
rect 1813 3313 1827 3327
rect 1853 3333 1867 3347
rect 1833 3273 1847 3287
rect 1753 3253 1767 3267
rect 1773 3253 1787 3267
rect 1693 3193 1707 3207
rect 1673 3173 1687 3187
rect 1693 3173 1707 3187
rect 1653 3093 1667 3107
rect 1653 3073 1667 3087
rect 1653 3033 1667 3047
rect 1673 3033 1687 3047
rect 1633 3013 1647 3027
rect 1653 2993 1667 3007
rect 1613 2933 1627 2947
rect 1593 2893 1607 2907
rect 1593 2873 1607 2887
rect 1793 3113 1807 3127
rect 1773 3093 1787 3107
rect 1773 3073 1787 3087
rect 1753 3053 1767 3067
rect 1733 3033 1747 3047
rect 1813 3053 1827 3067
rect 1833 3053 1847 3067
rect 1793 3033 1807 3047
rect 1973 3453 1987 3467
rect 2053 3473 2067 3487
rect 2033 3433 2047 3447
rect 2013 3413 2027 3427
rect 2013 3373 2027 3387
rect 2013 3353 2027 3367
rect 1953 3293 1967 3307
rect 1973 3293 1987 3307
rect 1973 3233 1987 3247
rect 1873 3213 1887 3227
rect 1933 3213 1947 3227
rect 1913 3193 1927 3207
rect 1893 3153 1907 3167
rect 1933 3153 1947 3167
rect 1873 3113 1887 3127
rect 1853 3033 1867 3047
rect 1713 2933 1727 2947
rect 1693 2913 1707 2927
rect 1693 2893 1707 2907
rect 1753 2893 1767 2907
rect 1553 2773 1567 2787
rect 1513 2733 1527 2747
rect 1553 2733 1567 2747
rect 1433 2673 1447 2687
rect 1453 2673 1467 2687
rect 1433 2593 1447 2607
rect 1453 2573 1467 2587
rect 1573 2653 1587 2667
rect 1733 2853 1747 2867
rect 1613 2773 1627 2787
rect 1693 2773 1707 2787
rect 1613 2733 1627 2747
rect 1693 2733 1707 2747
rect 1633 2713 1647 2727
rect 1673 2713 1687 2727
rect 1533 2593 1547 2607
rect 1453 2373 1467 2387
rect 1373 2273 1387 2287
rect 1393 2273 1407 2287
rect 1413 2273 1427 2287
rect 1353 2253 1367 2267
rect 1473 2253 1487 2267
rect 1393 2233 1407 2247
rect 1433 2233 1447 2247
rect 1453 2233 1467 2247
rect 1553 2553 1567 2567
rect 1513 2373 1527 2387
rect 1493 2233 1507 2247
rect 1593 2573 1607 2587
rect 1653 2573 1667 2587
rect 1613 2553 1627 2567
rect 1593 2513 1607 2527
rect 1573 2473 1587 2487
rect 1673 2533 1687 2547
rect 1593 2433 1607 2447
rect 1633 2433 1647 2447
rect 1533 2253 1547 2267
rect 1573 2253 1587 2267
rect 1333 2213 1347 2227
rect 1473 2213 1487 2227
rect 1193 2053 1207 2067
rect 1273 2053 1287 2067
rect 1313 2053 1327 2067
rect 1233 2033 1247 2047
rect 1153 1933 1167 1947
rect 1253 1913 1267 1927
rect 1093 1893 1107 1907
rect 1133 1893 1147 1907
rect 1053 1793 1067 1807
rect 1073 1793 1087 1807
rect 1173 1813 1187 1827
rect 1113 1773 1127 1787
rect 1133 1753 1147 1767
rect 1073 1733 1087 1747
rect 1093 1733 1107 1747
rect 1153 1733 1167 1747
rect 1013 1653 1027 1667
rect 993 1613 1007 1627
rect 853 1553 867 1567
rect 813 1533 827 1547
rect 993 1593 1007 1607
rect 933 1553 947 1567
rect 893 1533 907 1547
rect 893 1473 907 1487
rect 1053 1633 1067 1647
rect 1033 1613 1047 1627
rect 1513 2113 1527 2127
rect 1373 2053 1387 2067
rect 1393 2033 1407 2047
rect 1353 2013 1367 2027
rect 1333 1873 1347 1887
rect 1293 1813 1307 1827
rect 1473 2073 1487 2087
rect 1453 2053 1467 2067
rect 1453 2033 1467 2047
rect 1493 2033 1507 2047
rect 1413 2013 1427 2027
rect 1553 2233 1567 2247
rect 1673 2233 1687 2247
rect 1553 2193 1567 2207
rect 1673 2193 1687 2207
rect 1553 2093 1567 2107
rect 1593 2093 1607 2107
rect 1633 2073 1647 2087
rect 1553 2053 1567 2067
rect 1613 2033 1627 2047
rect 1573 2013 1587 2027
rect 1613 1993 1627 2007
rect 1533 1973 1547 1987
rect 1413 1873 1427 1887
rect 1553 1873 1567 1887
rect 1393 1833 1407 1847
rect 1273 1793 1287 1807
rect 1313 1793 1327 1807
rect 1373 1813 1387 1827
rect 1473 1853 1487 1867
rect 1453 1833 1467 1847
rect 1433 1813 1447 1827
rect 1393 1793 1407 1807
rect 1113 1713 1127 1727
rect 1173 1713 1187 1727
rect 1073 1573 1087 1587
rect 1053 1553 1067 1567
rect 1033 1493 1047 1507
rect 1173 1693 1187 1707
rect 1213 1753 1227 1767
rect 1233 1733 1247 1747
rect 1213 1673 1227 1687
rect 1193 1653 1207 1667
rect 1153 1633 1167 1647
rect 1153 1613 1167 1627
rect 1173 1613 1187 1627
rect 1153 1573 1167 1587
rect 1133 1553 1147 1567
rect 1073 1353 1087 1367
rect 1093 1353 1107 1367
rect 913 1333 927 1347
rect 953 1333 967 1347
rect 1013 1333 1027 1347
rect 873 1313 887 1327
rect 973 1313 987 1327
rect 1033 1313 1047 1327
rect 1073 1313 1087 1327
rect 773 1293 787 1307
rect 793 1293 807 1307
rect 753 1253 767 1267
rect 573 1233 587 1247
rect 533 1213 547 1227
rect 573 1213 587 1227
rect 653 1213 667 1227
rect 553 1173 567 1187
rect 553 1113 567 1127
rect 573 1093 587 1107
rect 613 1093 627 1107
rect 733 1113 747 1127
rect 773 1093 787 1107
rect 533 1033 547 1047
rect 593 893 607 907
rect 513 873 527 887
rect 393 833 407 847
rect 433 833 447 847
rect 453 833 467 847
rect 493 833 507 847
rect 473 813 487 827
rect 513 793 527 807
rect 533 793 547 807
rect 333 773 347 787
rect 313 753 327 767
rect 313 693 327 707
rect 313 673 327 687
rect 193 653 207 667
rect 173 633 187 647
rect 213 633 227 647
rect 273 633 287 647
rect 93 613 107 627
rect 113 613 127 627
rect 93 593 107 607
rect 53 553 67 567
rect 53 513 67 527
rect 33 393 47 407
rect 153 533 167 547
rect 253 613 267 627
rect 293 593 307 607
rect 213 513 227 527
rect 273 493 287 507
rect 93 413 107 427
rect 73 373 87 387
rect 13 353 27 367
rect 53 353 67 367
rect 13 333 27 347
rect 73 253 87 267
rect 53 173 67 187
rect 33 153 47 167
rect 113 393 127 407
rect 293 413 307 427
rect 153 373 167 387
rect 273 373 287 387
rect 553 673 567 687
rect 453 653 467 667
rect 373 633 387 647
rect 433 633 447 647
rect 493 633 507 647
rect 533 633 547 647
rect 593 633 607 647
rect 413 573 427 587
rect 453 613 467 627
rect 473 613 487 627
rect 433 553 447 567
rect 353 533 367 547
rect 513 613 527 627
rect 553 613 567 627
rect 493 553 507 567
rect 453 493 467 507
rect 673 853 687 867
rect 753 1073 767 1087
rect 853 1293 867 1307
rect 913 1293 927 1307
rect 833 1273 847 1287
rect 813 1173 827 1187
rect 853 1173 867 1187
rect 873 1133 887 1147
rect 913 1133 927 1147
rect 813 1113 827 1127
rect 793 893 807 907
rect 833 1093 847 1107
rect 773 873 787 887
rect 813 873 827 887
rect 773 853 787 867
rect 753 833 767 847
rect 653 753 667 767
rect 853 853 867 867
rect 793 753 807 767
rect 753 673 767 687
rect 893 1053 907 1067
rect 953 1293 967 1307
rect 993 1293 1007 1307
rect 1013 1293 1027 1307
rect 973 1273 987 1287
rect 1073 1273 1087 1287
rect 953 1253 967 1267
rect 1053 1253 1067 1267
rect 1033 1233 1047 1247
rect 1013 1173 1027 1187
rect 973 1153 987 1167
rect 993 1153 1007 1167
rect 1013 1093 1027 1107
rect 993 1053 1007 1067
rect 953 1033 967 1047
rect 933 953 947 967
rect 933 933 947 947
rect 913 853 927 867
rect 893 813 907 827
rect 993 913 1007 927
rect 953 853 967 867
rect 933 793 947 807
rect 873 713 887 727
rect 913 693 927 707
rect 993 753 1007 767
rect 733 653 747 667
rect 773 653 787 667
rect 833 653 847 667
rect 873 653 887 667
rect 673 633 687 647
rect 713 633 727 647
rect 613 613 627 627
rect 653 613 667 627
rect 593 573 607 587
rect 573 473 587 487
rect 553 433 567 447
rect 313 393 327 407
rect 353 393 367 407
rect 393 393 407 407
rect 173 353 187 367
rect 213 353 227 367
rect 253 353 267 367
rect 333 353 347 367
rect 133 333 147 347
rect 173 333 187 347
rect 113 253 127 267
rect 93 153 107 167
rect 233 333 247 347
rect 273 333 287 347
rect 193 313 207 327
rect 273 313 287 327
rect 173 173 187 187
rect 213 173 227 187
rect 153 153 167 167
rect 253 153 267 167
rect 233 133 247 147
rect 413 353 427 367
rect 453 353 467 367
rect 393 333 407 347
rect 333 293 347 307
rect 433 313 447 327
rect 493 353 507 367
rect 473 293 487 307
rect 453 273 467 287
rect 393 253 407 267
rect 393 233 407 247
rect 333 173 347 187
rect 373 153 387 167
rect 373 113 387 127
rect 593 353 607 367
rect 553 313 567 327
rect 493 233 507 247
rect 533 233 547 247
rect 533 213 547 227
rect 693 593 707 607
rect 733 593 747 607
rect 753 593 767 607
rect 773 593 787 607
rect 693 513 707 527
rect 713 453 727 467
rect 733 373 747 387
rect 673 353 687 367
rect 693 353 707 367
rect 713 353 727 367
rect 633 333 647 347
rect 733 333 747 347
rect 853 613 867 627
rect 893 613 907 627
rect 813 513 827 527
rect 793 373 807 387
rect 933 613 947 627
rect 893 473 907 487
rect 913 473 927 487
rect 873 413 887 427
rect 773 333 787 347
rect 673 313 687 327
rect 693 313 707 327
rect 753 313 767 327
rect 653 293 667 307
rect 653 173 667 187
rect 673 173 687 187
rect 573 153 587 167
rect 613 153 627 167
rect 553 133 567 147
rect 633 133 647 147
rect 973 673 987 687
rect 973 653 987 667
rect 1073 1193 1087 1207
rect 1253 1693 1267 1707
rect 1273 1673 1287 1687
rect 1313 1673 1327 1687
rect 1233 1593 1247 1607
rect 1253 1593 1267 1607
rect 1293 1553 1307 1567
rect 1253 1493 1267 1507
rect 1273 1493 1287 1507
rect 1293 1473 1307 1487
rect 1293 1453 1307 1467
rect 1113 1333 1127 1347
rect 1173 1333 1187 1347
rect 1253 1333 1267 1347
rect 1273 1333 1287 1347
rect 1093 1153 1107 1167
rect 1093 1133 1107 1147
rect 1213 1313 1227 1327
rect 1133 1293 1147 1307
rect 1173 1273 1187 1287
rect 1153 1193 1167 1207
rect 1133 1173 1147 1187
rect 1133 1113 1147 1127
rect 1113 1093 1127 1107
rect 1213 1253 1227 1267
rect 1193 1233 1207 1247
rect 1193 1173 1207 1187
rect 1053 1073 1067 1087
rect 1133 1073 1147 1087
rect 1173 1073 1187 1087
rect 1033 1053 1047 1067
rect 1013 693 1027 707
rect 1113 793 1127 807
rect 1073 753 1087 767
rect 1033 673 1047 687
rect 1073 673 1087 687
rect 973 633 987 647
rect 1053 613 1067 627
rect 1113 613 1127 627
rect 1093 573 1107 587
rect 1073 513 1087 527
rect 1013 453 1027 467
rect 953 433 967 447
rect 1013 433 1027 447
rect 933 393 947 407
rect 893 373 907 387
rect 933 373 947 387
rect 973 373 987 387
rect 953 353 967 367
rect 913 333 927 347
rect 953 313 967 327
rect 993 313 1007 327
rect 873 293 887 307
rect 833 273 847 287
rect 933 273 947 287
rect 773 173 787 187
rect 813 173 827 187
rect 693 133 707 147
rect 473 113 487 127
rect 513 113 527 127
rect 673 113 687 127
rect 753 133 767 147
rect 853 153 867 167
rect 1053 233 1067 247
rect 1013 213 1027 227
rect 993 193 1007 207
rect 1253 1273 1267 1287
rect 1273 1273 1287 1287
rect 1233 1213 1247 1227
rect 1273 1213 1287 1227
rect 1253 1193 1267 1207
rect 1213 1153 1227 1167
rect 1213 1133 1227 1147
rect 1233 1113 1247 1127
rect 1353 1753 1367 1767
rect 1433 1753 1447 1767
rect 1433 1633 1447 1647
rect 1353 1613 1367 1627
rect 1393 1593 1407 1607
rect 1353 1533 1367 1547
rect 1373 1533 1387 1547
rect 1333 1513 1347 1527
rect 1313 1353 1327 1367
rect 1313 1333 1327 1347
rect 1373 1513 1387 1527
rect 1393 1513 1407 1527
rect 1333 1313 1347 1327
rect 1593 1833 1607 1847
rect 1473 1813 1487 1827
rect 1553 1813 1567 1827
rect 1573 1793 1587 1807
rect 1513 1773 1527 1787
rect 1533 1773 1547 1787
rect 1493 1713 1507 1727
rect 1513 1713 1527 1727
rect 1913 3133 1927 3147
rect 1993 3213 2007 3227
rect 1973 3193 1987 3207
rect 2013 3193 2027 3207
rect 1953 3113 1967 3127
rect 2353 3973 2367 3987
rect 2333 3933 2347 3947
rect 2413 4073 2427 4087
rect 2433 4053 2447 4067
rect 2533 4473 2547 4487
rect 2753 4633 2767 4647
rect 2713 4513 2727 4527
rect 2593 4453 2607 4467
rect 2633 4453 2647 4467
rect 2853 4673 2867 4687
rect 2833 4653 2847 4667
rect 2833 4633 2847 4647
rect 2873 4633 2887 4647
rect 2773 4613 2787 4627
rect 2813 4613 2827 4627
rect 2673 4433 2687 4447
rect 2653 4413 2667 4427
rect 2553 4373 2567 4387
rect 2513 4293 2527 4307
rect 2473 4213 2487 4227
rect 2513 4213 2527 4227
rect 2493 4193 2507 4207
rect 2653 4313 2667 4327
rect 2733 4433 2747 4447
rect 2713 4313 2727 4327
rect 2673 4293 2687 4307
rect 2613 4213 2627 4227
rect 2573 4193 2587 4207
rect 2553 4133 2567 4147
rect 2493 4073 2507 4087
rect 2493 3993 2507 4007
rect 2633 4173 2647 4187
rect 2673 4153 2687 4167
rect 2693 4133 2707 4147
rect 2793 4453 2807 4467
rect 2753 4253 2767 4267
rect 2773 4233 2787 4247
rect 2833 4573 2847 4587
rect 2953 4653 2967 4667
rect 2913 4553 2927 4567
rect 2873 4493 2887 4507
rect 2853 4433 2867 4447
rect 2833 4353 2847 4367
rect 2853 4213 2867 4227
rect 2813 4173 2827 4187
rect 2853 4153 2867 4167
rect 2733 4113 2747 4127
rect 2713 4053 2727 4067
rect 2653 4033 2667 4047
rect 2633 3993 2647 4007
rect 2393 3973 2407 3987
rect 2453 3973 2467 3987
rect 2473 3973 2487 3987
rect 2413 3913 2427 3927
rect 2453 3913 2467 3927
rect 2373 3873 2387 3887
rect 2313 3853 2327 3867
rect 2353 3813 2367 3827
rect 2313 3773 2327 3787
rect 2213 3673 2227 3687
rect 2133 3553 2147 3567
rect 2153 3553 2167 3567
rect 2173 3533 2187 3547
rect 2193 3533 2207 3547
rect 2133 3513 2147 3527
rect 2153 3513 2167 3527
rect 2113 3473 2127 3487
rect 2093 3453 2107 3467
rect 2153 3453 2167 3467
rect 2173 3453 2187 3467
rect 2073 3433 2087 3447
rect 2113 3433 2127 3447
rect 2133 3433 2147 3447
rect 2073 3253 2087 3267
rect 2073 3213 2087 3227
rect 2053 3173 2067 3187
rect 2033 3153 2047 3167
rect 2153 3353 2167 3367
rect 2153 3193 2167 3207
rect 2013 3113 2027 3127
rect 2053 3113 2067 3127
rect 2033 3073 2047 3087
rect 1973 3053 1987 3067
rect 1933 3013 1947 3027
rect 1953 3013 1967 3027
rect 1993 3013 2007 3027
rect 1893 2933 1907 2947
rect 1873 2873 1887 2887
rect 1853 2853 1867 2867
rect 1793 2813 1807 2827
rect 1813 2733 1827 2747
rect 1773 2713 1787 2727
rect 1773 2693 1787 2707
rect 1753 2633 1767 2647
rect 1733 2553 1747 2567
rect 1873 2833 1887 2847
rect 1853 2713 1867 2727
rect 1853 2693 1867 2707
rect 1833 2653 1847 2667
rect 1813 2613 1827 2627
rect 1853 2613 1867 2627
rect 1913 2873 1927 2887
rect 1893 2793 1907 2807
rect 1973 2953 1987 2967
rect 2013 2953 2027 2967
rect 2013 2853 2027 2867
rect 2073 3013 2087 3027
rect 2053 2973 2067 2987
rect 2053 2853 2067 2867
rect 2033 2833 2047 2847
rect 2053 2833 2067 2847
rect 1993 2813 2007 2827
rect 1953 2773 1967 2787
rect 1953 2753 1967 2767
rect 1873 2593 1887 2607
rect 1973 2733 1987 2747
rect 1973 2693 1987 2707
rect 2033 2773 2047 2787
rect 2013 2753 2027 2767
rect 2033 2733 2047 2747
rect 2073 2713 2087 2727
rect 1993 2673 2007 2687
rect 2053 2673 2067 2687
rect 1993 2593 2007 2607
rect 1893 2573 1907 2587
rect 1913 2573 1927 2587
rect 1893 2553 1907 2567
rect 1713 2473 1727 2487
rect 1833 2533 1847 2547
rect 1933 2553 1947 2567
rect 1953 2533 1967 2547
rect 1913 2513 1927 2527
rect 1873 2473 1887 2487
rect 1753 2453 1767 2467
rect 1873 2433 1887 2447
rect 1913 2433 1927 2447
rect 1833 2313 1847 2327
rect 1773 2253 1787 2267
rect 1893 2253 1907 2267
rect 1813 2213 1827 2227
rect 1713 2193 1727 2207
rect 1773 2173 1787 2187
rect 1713 2153 1727 2167
rect 1693 2093 1707 2107
rect 1693 2073 1707 2087
rect 1833 2133 1847 2147
rect 1833 2073 1847 2087
rect 1713 1973 1727 1987
rect 1633 1853 1647 1867
rect 1673 1853 1687 1867
rect 1693 1853 1707 1867
rect 1673 1813 1687 1827
rect 1633 1753 1647 1767
rect 1613 1693 1627 1707
rect 1473 1633 1487 1647
rect 1493 1613 1507 1627
rect 1473 1593 1487 1607
rect 1473 1553 1487 1567
rect 1453 1453 1467 1467
rect 1533 1593 1547 1607
rect 1513 1533 1527 1547
rect 1493 1513 1507 1527
rect 1513 1473 1527 1487
rect 1473 1433 1487 1447
rect 1413 1393 1427 1407
rect 1433 1393 1447 1407
rect 1393 1333 1407 1347
rect 1453 1333 1467 1347
rect 1533 1453 1547 1467
rect 1313 1193 1327 1207
rect 1293 1173 1307 1187
rect 1253 1093 1267 1107
rect 1293 1093 1307 1107
rect 1333 1093 1347 1107
rect 1233 1073 1247 1087
rect 1413 1233 1427 1247
rect 1373 1213 1387 1227
rect 1493 1273 1507 1287
rect 1413 1173 1427 1187
rect 1453 1173 1467 1187
rect 1413 1133 1427 1147
rect 1453 1133 1467 1147
rect 1393 1093 1407 1107
rect 1473 1093 1487 1107
rect 1193 1053 1207 1067
rect 1153 1013 1167 1027
rect 1193 873 1207 887
rect 1313 1053 1327 1067
rect 1153 853 1167 867
rect 1173 833 1187 847
rect 1153 693 1167 707
rect 1193 673 1207 687
rect 1173 653 1187 667
rect 1153 633 1167 647
rect 1153 593 1167 607
rect 1233 833 1247 847
rect 1273 833 1287 847
rect 1253 773 1267 787
rect 1313 753 1327 767
rect 1273 693 1287 707
rect 1293 693 1307 707
rect 1313 693 1327 707
rect 1253 653 1267 667
rect 1213 613 1227 627
rect 1133 433 1147 447
rect 1313 633 1327 647
rect 1273 613 1287 627
rect 1313 613 1327 627
rect 1273 593 1287 607
rect 1233 413 1247 427
rect 1133 373 1147 387
rect 1193 373 1207 387
rect 1113 333 1127 347
rect 1173 353 1187 367
rect 1213 353 1227 367
rect 1153 273 1167 287
rect 1133 213 1147 227
rect 1073 153 1087 167
rect 853 133 867 147
rect 933 133 947 147
rect 793 113 807 127
rect 833 113 847 127
rect 873 113 887 127
rect 793 93 807 107
rect 1033 133 1047 147
rect 1433 1053 1447 1067
rect 1513 1053 1527 1067
rect 1373 973 1387 987
rect 1353 813 1367 827
rect 1493 1033 1507 1047
rect 1453 853 1467 867
rect 1513 993 1527 1007
rect 1433 813 1447 827
rect 1573 1553 1587 1567
rect 1613 1553 1627 1567
rect 1653 1653 1667 1667
rect 1833 2053 1847 2067
rect 1873 2053 1887 2067
rect 1893 2053 1907 2067
rect 1853 2033 1867 2047
rect 1833 1973 1847 1987
rect 1733 1953 1747 1967
rect 1793 1953 1807 1967
rect 1753 1933 1767 1947
rect 1793 1813 1807 1827
rect 1753 1793 1767 1807
rect 1773 1753 1787 1767
rect 1793 1693 1807 1707
rect 1693 1673 1707 1687
rect 1733 1653 1747 1667
rect 1613 1533 1627 1547
rect 1633 1533 1647 1547
rect 1593 1433 1607 1447
rect 1573 1393 1587 1407
rect 1553 1333 1567 1347
rect 1593 1333 1607 1347
rect 1673 1593 1687 1607
rect 1693 1593 1707 1607
rect 1853 1933 1867 1947
rect 1853 1773 1867 1787
rect 1953 2353 1967 2367
rect 1933 2253 1947 2267
rect 2013 2553 2027 2567
rect 1993 2273 2007 2287
rect 1953 2213 1967 2227
rect 1973 2153 1987 2167
rect 2073 2613 2087 2627
rect 2113 3033 2127 3047
rect 2273 3693 2287 3707
rect 2233 3573 2247 3587
rect 2253 3573 2267 3587
rect 2353 3733 2367 3747
rect 2413 3733 2427 3747
rect 2333 3693 2347 3707
rect 2333 3653 2347 3667
rect 2333 3553 2347 3567
rect 2273 3533 2287 3547
rect 2313 3533 2327 3547
rect 2253 3413 2267 3427
rect 2213 3373 2227 3387
rect 2193 3273 2207 3287
rect 2193 3193 2207 3207
rect 2173 3093 2187 3107
rect 2293 3513 2307 3527
rect 2353 3493 2367 3507
rect 2533 3813 2547 3827
rect 2493 3793 2507 3807
rect 2473 3773 2487 3787
rect 2473 3713 2487 3727
rect 2493 3713 2507 3727
rect 2513 3713 2527 3727
rect 2493 3673 2507 3687
rect 2453 3653 2467 3667
rect 2493 3653 2507 3667
rect 2393 3613 2407 3627
rect 2453 3613 2467 3627
rect 2373 3433 2387 3447
rect 2413 3593 2427 3607
rect 2433 3533 2447 3547
rect 2473 3593 2487 3607
rect 2453 3513 2467 3527
rect 2433 3493 2447 3507
rect 2413 3473 2427 3487
rect 2393 3413 2407 3427
rect 2313 3353 2327 3367
rect 2313 3313 2327 3327
rect 2373 3313 2387 3327
rect 2273 3293 2287 3307
rect 2453 3453 2467 3467
rect 2433 3333 2447 3347
rect 2433 3293 2447 3307
rect 2393 3233 2407 3247
rect 2213 3073 2227 3087
rect 2253 3073 2267 3087
rect 2253 3053 2267 3067
rect 2293 3053 2307 3067
rect 2193 3033 2207 3047
rect 2213 3033 2227 3047
rect 2193 2993 2207 3007
rect 2173 2973 2187 2987
rect 2133 2873 2147 2887
rect 2133 2793 2147 2807
rect 2153 2753 2167 2767
rect 2133 2713 2147 2727
rect 2213 2973 2227 2987
rect 2273 2993 2287 3007
rect 2433 3193 2447 3207
rect 2473 3313 2487 3327
rect 2633 3733 2647 3747
rect 2573 3713 2587 3727
rect 2613 3713 2627 3727
rect 2553 3693 2567 3707
rect 2613 3693 2627 3707
rect 2613 3653 2627 3667
rect 2893 4393 2907 4407
rect 2933 4373 2947 4387
rect 2913 4333 2927 4347
rect 2893 4173 2907 4187
rect 2873 4093 2887 4107
rect 2673 3953 2687 3967
rect 2733 3973 2747 3987
rect 2713 3913 2727 3927
rect 2713 3873 2727 3887
rect 2753 3933 2767 3947
rect 2853 3993 2867 4007
rect 2893 3993 2907 4007
rect 2773 3913 2787 3927
rect 2813 3873 2827 3887
rect 2733 3733 2747 3747
rect 2693 3713 2707 3727
rect 2733 3713 2747 3727
rect 2673 3693 2687 3707
rect 2653 3633 2667 3647
rect 2533 3613 2547 3627
rect 2593 3613 2607 3627
rect 2633 3613 2647 3627
rect 2653 3613 2667 3627
rect 2593 3593 2607 3607
rect 2613 3593 2627 3607
rect 2533 3553 2547 3567
rect 2513 3533 2527 3547
rect 2593 3533 2607 3547
rect 2573 3513 2587 3527
rect 2693 3633 2707 3647
rect 2673 3593 2687 3607
rect 2653 3533 2667 3547
rect 2673 3533 2687 3547
rect 2653 3513 2667 3527
rect 2573 3373 2587 3387
rect 2553 3293 2567 3307
rect 2493 3273 2507 3287
rect 2553 3273 2567 3287
rect 2473 3233 2487 3247
rect 2513 3233 2527 3247
rect 2453 3133 2467 3147
rect 2393 3113 2407 3127
rect 2433 3053 2447 3067
rect 2353 3033 2367 3047
rect 2353 2993 2367 3007
rect 2273 2973 2287 2987
rect 2313 2973 2327 2987
rect 2233 2953 2247 2967
rect 2233 2873 2247 2887
rect 2253 2793 2267 2807
rect 2213 2753 2227 2767
rect 2333 2873 2347 2887
rect 2353 2873 2367 2887
rect 2293 2853 2307 2867
rect 2273 2773 2287 2787
rect 2333 2773 2347 2787
rect 2213 2733 2227 2747
rect 2113 2693 2127 2707
rect 2113 2593 2127 2607
rect 2193 2713 2207 2727
rect 2193 2553 2207 2567
rect 2253 2713 2267 2727
rect 2333 2733 2347 2747
rect 2313 2713 2327 2727
rect 2293 2693 2307 2707
rect 2253 2673 2267 2687
rect 2233 2653 2247 2667
rect 2253 2653 2267 2667
rect 2413 3013 2427 3027
rect 2393 2833 2407 2847
rect 2373 2793 2387 2807
rect 2413 2793 2427 2807
rect 2353 2693 2367 2707
rect 2533 3213 2547 3227
rect 2533 3193 2547 3207
rect 2513 3093 2527 3107
rect 2493 3013 2507 3027
rect 2453 2973 2467 2987
rect 2613 3373 2627 3387
rect 2593 3333 2607 3347
rect 2773 3673 2787 3687
rect 2753 3613 2767 3627
rect 2713 3553 2727 3567
rect 2833 3693 2847 3707
rect 2953 4153 2967 4167
rect 2953 4053 2967 4067
rect 2913 3773 2927 3787
rect 2893 3733 2907 3747
rect 2933 3713 2947 3727
rect 2873 3693 2887 3707
rect 2913 3693 2927 3707
rect 2853 3673 2867 3687
rect 2933 3673 2947 3687
rect 2913 3653 2927 3667
rect 2793 3633 2807 3647
rect 2853 3593 2867 3607
rect 2833 3553 2847 3567
rect 2733 3513 2747 3527
rect 2773 3513 2787 3527
rect 2693 3453 2707 3467
rect 2813 3493 2827 3507
rect 2873 3533 2887 3547
rect 2753 3413 2767 3427
rect 2733 3313 2747 3327
rect 2673 3293 2687 3307
rect 2713 3273 2727 3287
rect 2613 3253 2627 3267
rect 2633 3253 2647 3267
rect 2713 3253 2727 3267
rect 2573 3133 2587 3147
rect 2553 3093 2567 3107
rect 2533 3053 2547 3067
rect 2553 2993 2567 3007
rect 2573 2973 2587 2987
rect 2473 2853 2487 2867
rect 2513 2853 2527 2867
rect 2533 2853 2547 2867
rect 2433 2753 2447 2767
rect 2453 2753 2467 2767
rect 2373 2633 2387 2647
rect 2353 2593 2367 2607
rect 2253 2573 2267 2587
rect 2293 2573 2307 2587
rect 2333 2573 2347 2587
rect 2213 2513 2227 2527
rect 2213 2473 2227 2487
rect 2093 2433 2107 2447
rect 2153 2433 2167 2447
rect 2173 2333 2187 2347
rect 2053 2273 2067 2287
rect 2093 2273 2107 2287
rect 2133 2273 2147 2287
rect 2333 2553 2347 2567
rect 2253 2513 2267 2527
rect 2233 2333 2247 2347
rect 2033 2253 2047 2267
rect 2053 2253 2067 2267
rect 2013 2133 2027 2147
rect 1993 2113 2007 2127
rect 1933 2093 1947 2107
rect 1973 2093 1987 2107
rect 1913 2013 1927 2027
rect 1953 2033 1967 2047
rect 2013 2053 2027 2067
rect 1913 1913 1927 1927
rect 1933 1913 1947 1927
rect 1993 1913 2007 1927
rect 1913 1873 1927 1887
rect 1973 1893 1987 1907
rect 2053 2213 2067 2227
rect 2073 2213 2087 2227
rect 2153 2253 2167 2267
rect 2193 2253 2207 2267
rect 2233 2253 2247 2267
rect 2053 2113 2067 2127
rect 2113 2113 2127 2127
rect 2073 2093 2087 2107
rect 2113 2093 2127 2107
rect 2093 2073 2107 2087
rect 2113 2073 2127 2087
rect 2313 2513 2327 2527
rect 2333 2493 2347 2507
rect 2273 2473 2287 2487
rect 2313 2433 2327 2447
rect 2273 2273 2287 2287
rect 2253 2213 2267 2227
rect 2293 2193 2307 2207
rect 2293 2173 2307 2187
rect 2213 2133 2227 2147
rect 2293 2133 2307 2147
rect 2273 2113 2287 2127
rect 2073 2053 2087 2067
rect 2133 2053 2147 2067
rect 2193 2033 2207 2047
rect 2133 2013 2147 2027
rect 2073 1893 2087 1907
rect 2033 1873 2047 1887
rect 2053 1833 2067 1847
rect 1873 1753 1887 1767
rect 1893 1753 1907 1767
rect 1913 1753 1927 1767
rect 1853 1713 1867 1727
rect 1833 1653 1847 1667
rect 1933 1693 1947 1707
rect 1873 1653 1887 1667
rect 1913 1653 1927 1667
rect 1793 1613 1807 1627
rect 1853 1613 1867 1627
rect 1753 1593 1767 1607
rect 1773 1593 1787 1607
rect 1813 1593 1827 1607
rect 1713 1513 1727 1527
rect 1733 1493 1747 1507
rect 1693 1473 1707 1487
rect 1673 1373 1687 1387
rect 1653 1333 1667 1347
rect 1653 1313 1667 1327
rect 1553 1293 1567 1307
rect 1553 1213 1567 1227
rect 1633 1293 1647 1307
rect 1633 1253 1647 1267
rect 1653 1233 1667 1247
rect 1593 1193 1607 1207
rect 1613 1193 1627 1207
rect 1593 1173 1607 1187
rect 1573 1133 1587 1147
rect 1553 1093 1567 1107
rect 1633 1173 1647 1187
rect 1613 1113 1627 1127
rect 1573 1073 1587 1087
rect 1613 1073 1627 1087
rect 1593 1053 1607 1067
rect 1593 993 1607 1007
rect 1613 953 1627 967
rect 1533 913 1547 927
rect 1573 913 1587 927
rect 1533 893 1547 907
rect 1533 853 1547 867
rect 1473 793 1487 807
rect 1513 793 1527 807
rect 1733 1413 1747 1427
rect 1693 1353 1707 1367
rect 1793 1573 1807 1587
rect 1833 1553 1847 1567
rect 1893 1593 1907 1607
rect 1913 1593 1927 1607
rect 1993 1793 2007 1807
rect 2033 1793 2047 1807
rect 2013 1693 2027 1707
rect 1993 1633 2007 1647
rect 1933 1573 1947 1587
rect 1913 1533 1927 1547
rect 1873 1493 1887 1507
rect 1833 1453 1847 1467
rect 1833 1393 1847 1407
rect 1793 1373 1807 1387
rect 1773 1333 1787 1347
rect 1913 1353 1927 1367
rect 1713 1313 1727 1327
rect 1733 1313 1747 1327
rect 1753 1313 1767 1327
rect 1673 1133 1687 1147
rect 1733 1273 1747 1287
rect 1753 1273 1767 1287
rect 1753 1233 1767 1247
rect 1873 1333 1887 1347
rect 1913 1333 1927 1347
rect 1833 1313 1847 1327
rect 1813 1293 1827 1307
rect 1853 1293 1867 1307
rect 1893 1293 1907 1307
rect 1853 1273 1867 1287
rect 1873 1273 1887 1287
rect 1793 1233 1807 1247
rect 1773 1193 1787 1207
rect 1713 1133 1727 1147
rect 1733 1133 1747 1147
rect 1773 1133 1787 1147
rect 1653 1113 1667 1127
rect 1693 1113 1707 1127
rect 1753 1113 1767 1127
rect 1813 1213 1827 1227
rect 1833 1213 1847 1227
rect 1773 1093 1787 1107
rect 1653 953 1667 967
rect 1653 913 1667 927
rect 1633 873 1647 887
rect 1713 1073 1727 1087
rect 1893 1233 1907 1247
rect 1873 1153 1887 1167
rect 1813 953 1827 967
rect 1873 1093 1887 1107
rect 1853 993 1867 1007
rect 1833 933 1847 947
rect 1773 913 1787 927
rect 1793 893 1807 907
rect 1673 873 1687 887
rect 1693 873 1707 887
rect 1753 873 1767 887
rect 1593 813 1607 827
rect 1633 813 1647 827
rect 1593 793 1607 807
rect 1573 753 1587 767
rect 1413 733 1427 747
rect 1473 733 1487 747
rect 1393 713 1407 727
rect 1353 653 1367 667
rect 1373 653 1387 667
rect 1373 613 1387 627
rect 1333 573 1347 587
rect 1433 613 1447 627
rect 1493 633 1507 647
rect 1513 613 1527 627
rect 1533 613 1547 627
rect 1473 573 1487 587
rect 1413 553 1427 567
rect 1393 433 1407 447
rect 1333 373 1347 387
rect 1233 273 1247 287
rect 1353 353 1367 367
rect 1433 373 1447 387
rect 1513 453 1527 467
rect 1573 593 1587 607
rect 1673 793 1687 807
rect 1673 773 1687 787
rect 1613 733 1627 747
rect 1633 733 1647 747
rect 1613 713 1627 727
rect 1633 693 1647 707
rect 1653 653 1667 667
rect 1653 633 1667 647
rect 1593 573 1607 587
rect 1713 853 1727 867
rect 1773 853 1787 867
rect 1853 813 1867 827
rect 1773 793 1787 807
rect 1813 793 1827 807
rect 1733 753 1747 767
rect 1853 753 1867 767
rect 1773 733 1787 747
rect 1813 733 1827 747
rect 1753 713 1767 727
rect 1753 693 1767 707
rect 1693 673 1707 687
rect 1693 653 1707 667
rect 1713 633 1727 647
rect 1733 633 1747 647
rect 1693 613 1707 627
rect 1753 613 1767 627
rect 1773 613 1787 627
rect 1853 713 1867 727
rect 1833 673 1847 687
rect 2033 1633 2047 1647
rect 2093 1793 2107 1807
rect 2113 1753 2127 1767
rect 2173 1893 2187 1907
rect 2173 1793 2187 1807
rect 2153 1773 2167 1787
rect 2073 1653 2087 1667
rect 2013 1613 2027 1627
rect 2053 1613 2067 1627
rect 2093 1613 2107 1627
rect 2033 1593 2047 1607
rect 2073 1593 2087 1607
rect 2013 1573 2027 1587
rect 2013 1533 2027 1547
rect 2073 1553 2087 1567
rect 2053 1493 2067 1507
rect 2053 1473 2067 1487
rect 1973 1453 1987 1467
rect 2033 1413 2047 1427
rect 1953 1353 1967 1367
rect 1933 1193 1947 1207
rect 1973 1333 1987 1347
rect 2013 1333 2027 1347
rect 1953 1173 1967 1187
rect 1933 1153 1947 1167
rect 2073 1413 2087 1427
rect 2053 1393 2067 1407
rect 2073 1393 2087 1407
rect 2433 2653 2447 2667
rect 2413 2613 2427 2627
rect 2393 2573 2407 2587
rect 2373 2553 2387 2567
rect 2453 2553 2467 2567
rect 2393 2533 2407 2547
rect 2433 2493 2447 2507
rect 2433 2473 2447 2487
rect 2453 2473 2467 2487
rect 2353 2373 2367 2387
rect 2413 2373 2427 2387
rect 2413 2313 2427 2327
rect 2373 2293 2387 2307
rect 2453 2173 2467 2187
rect 2313 2113 2327 2127
rect 2673 3233 2687 3247
rect 2613 3213 2627 3227
rect 2653 3213 2667 3227
rect 2853 3473 2867 3487
rect 2893 3453 2907 3467
rect 2773 3293 2787 3307
rect 2813 3293 2827 3307
rect 2753 3213 2767 3227
rect 2633 3113 2647 3127
rect 2733 3113 2747 3127
rect 2593 2833 2607 2847
rect 2573 2793 2587 2807
rect 2513 2733 2527 2747
rect 2553 2733 2567 2747
rect 2493 2693 2507 2707
rect 2593 2773 2607 2787
rect 2613 2773 2627 2787
rect 2593 2733 2607 2747
rect 2533 2673 2547 2687
rect 2573 2673 2587 2687
rect 2513 2573 2527 2587
rect 2493 2533 2507 2547
rect 2553 2553 2567 2567
rect 2593 2553 2607 2567
rect 2533 2493 2547 2507
rect 2553 2313 2567 2327
rect 2553 2213 2567 2227
rect 2573 2213 2587 2227
rect 2533 2193 2547 2207
rect 2533 2173 2547 2187
rect 2333 2073 2347 2087
rect 2373 2073 2387 2087
rect 2413 2073 2427 2087
rect 2293 2053 2307 2067
rect 2313 2033 2327 2047
rect 2293 2013 2307 2027
rect 2233 1833 2247 1847
rect 2213 1813 2227 1827
rect 2253 1813 2267 1827
rect 2233 1793 2247 1807
rect 2253 1793 2267 1807
rect 2233 1773 2247 1787
rect 2193 1753 2207 1767
rect 2273 1713 2287 1727
rect 2433 2033 2447 2047
rect 2353 2013 2367 2027
rect 2353 1953 2367 1967
rect 2393 1953 2407 1967
rect 2373 1873 2387 1887
rect 2313 1833 2327 1847
rect 2313 1813 2327 1827
rect 2493 2113 2507 2127
rect 2473 2073 2487 2087
rect 2493 1953 2507 1967
rect 2453 1913 2467 1927
rect 2533 1993 2547 2007
rect 2533 1953 2547 1967
rect 2533 1893 2547 1907
rect 2473 1873 2487 1887
rect 2513 1873 2527 1887
rect 2393 1853 2407 1867
rect 2353 1733 2367 1747
rect 2273 1693 2287 1707
rect 2293 1693 2307 1707
rect 2153 1653 2167 1667
rect 2193 1653 2207 1667
rect 2133 1633 2147 1647
rect 2173 1613 2187 1627
rect 2153 1593 2167 1607
rect 2213 1633 2227 1647
rect 2273 1633 2287 1647
rect 2113 1553 2127 1567
rect 2133 1533 2147 1547
rect 2113 1513 2127 1527
rect 2153 1493 2167 1507
rect 2133 1413 2147 1427
rect 2053 1333 2067 1347
rect 2053 1273 2067 1287
rect 2033 1253 2047 1267
rect 2093 1373 2107 1387
rect 2113 1333 2127 1347
rect 2133 1333 2147 1347
rect 2093 1293 2107 1307
rect 2113 1293 2127 1307
rect 2133 1293 2147 1307
rect 2073 1213 2087 1227
rect 2013 1193 2027 1207
rect 2053 1193 2067 1207
rect 1993 1133 2007 1147
rect 1953 1113 1967 1127
rect 2133 1273 2147 1287
rect 2113 1173 2127 1187
rect 1973 1093 1987 1107
rect 2053 1093 2067 1107
rect 2033 1073 2047 1087
rect 2013 1053 2027 1067
rect 1893 1033 1907 1047
rect 1893 853 1907 867
rect 2113 1133 2127 1147
rect 2233 1513 2247 1527
rect 2253 1433 2267 1447
rect 2213 1373 2227 1387
rect 2213 1353 2227 1367
rect 2153 1213 2167 1227
rect 2233 1253 2247 1267
rect 2193 1153 2207 1167
rect 2153 1133 2167 1147
rect 2133 1113 2147 1127
rect 2333 1673 2347 1687
rect 2313 1593 2327 1607
rect 2293 1493 2307 1507
rect 2393 1813 2407 1827
rect 2373 1713 2387 1727
rect 2493 1853 2507 1867
rect 2433 1793 2447 1807
rect 2473 1793 2487 1807
rect 2513 1793 2527 1807
rect 2413 1773 2427 1787
rect 2493 1773 2507 1787
rect 2573 2153 2587 2167
rect 2673 3073 2687 3087
rect 2653 3053 2667 3067
rect 2653 2973 2667 2987
rect 2753 3073 2767 3087
rect 2853 3373 2867 3387
rect 2813 3233 2827 3247
rect 2833 3233 2847 3247
rect 2913 3333 2927 3347
rect 3193 4673 3207 4687
rect 3233 4673 3247 4687
rect 3013 4493 3027 4507
rect 3073 4653 3087 4667
rect 3093 4453 3107 4467
rect 3053 4433 3067 4447
rect 3113 4413 3127 4427
rect 3193 4653 3207 4667
rect 3233 4513 3247 4527
rect 4673 4813 4687 4827
rect 3313 4713 3327 4727
rect 3373 4713 3387 4727
rect 3873 4713 3887 4727
rect 4013 4713 4027 4727
rect 3293 4673 3307 4687
rect 3293 4453 3307 4467
rect 3193 4433 3207 4447
rect 3253 4433 3267 4447
rect 3173 4393 3187 4407
rect 3053 4253 3067 4267
rect 3113 4233 3127 4247
rect 3073 4213 3087 4227
rect 3153 4213 3167 4227
rect 3033 4193 3047 4207
rect 3133 4193 3147 4207
rect 3053 4173 3067 4187
rect 2973 4033 2987 4047
rect 3113 4173 3127 4187
rect 3253 4253 3267 4267
rect 3213 4173 3227 4187
rect 3113 4073 3127 4087
rect 3173 4033 3187 4047
rect 3093 4013 3107 4027
rect 3153 4013 3167 4027
rect 3093 3993 3107 4007
rect 3153 3993 3167 4007
rect 3013 3973 3027 3987
rect 3093 3973 3107 3987
rect 3133 3973 3147 3987
rect 2993 3913 3007 3927
rect 3193 3953 3207 3967
rect 3293 4033 3307 4047
rect 3253 3993 3267 4007
rect 3293 3993 3307 4007
rect 3493 4693 3507 4707
rect 3433 4673 3447 4687
rect 3473 4653 3487 4667
rect 3453 4633 3467 4647
rect 3413 4613 3427 4627
rect 3373 4513 3387 4527
rect 3333 4473 3347 4487
rect 3353 4453 3367 4467
rect 3393 4453 3407 4467
rect 3453 4453 3467 4467
rect 3473 4433 3487 4447
rect 3433 4413 3447 4427
rect 3593 4693 3607 4707
rect 3633 4693 3647 4707
rect 3533 4673 3547 4687
rect 3573 4653 3587 4667
rect 3813 4673 3827 4687
rect 3713 4653 3727 4667
rect 3753 4633 3767 4647
rect 3513 4613 3527 4627
rect 3773 4593 3787 4607
rect 3513 4493 3527 4507
rect 3613 4473 3627 4487
rect 3393 4393 3407 4407
rect 3493 4393 3507 4407
rect 3353 4213 3367 4227
rect 3333 4153 3347 4167
rect 3373 4093 3387 4107
rect 3113 3933 3127 3947
rect 3213 3933 3227 3947
rect 3033 3873 3047 3887
rect 3033 3833 3047 3847
rect 2973 3733 2987 3747
rect 3033 3733 3047 3747
rect 3013 3713 3027 3727
rect 2973 3633 2987 3647
rect 3073 3553 3087 3567
rect 2953 3533 2967 3547
rect 2993 3533 3007 3547
rect 2953 3513 2967 3527
rect 3033 3513 3047 3527
rect 2993 3493 3007 3507
rect 2973 3473 2987 3487
rect 2973 3453 2987 3467
rect 2993 3453 3007 3467
rect 3053 3493 3067 3507
rect 3093 3493 3107 3507
rect 3033 3453 3047 3467
rect 2953 3433 2967 3447
rect 3013 3433 3027 3447
rect 2913 3273 2927 3287
rect 2933 3273 2947 3287
rect 2893 3253 2907 3267
rect 2833 3193 2847 3207
rect 2853 3173 2867 3187
rect 2793 3113 2807 3127
rect 2793 3093 2807 3107
rect 2773 3053 2787 3067
rect 2853 3053 2867 3067
rect 2673 2953 2687 2967
rect 2653 2833 2667 2847
rect 2673 2813 2687 2827
rect 2833 3033 2847 3047
rect 2773 3013 2787 3027
rect 2813 3013 2827 3027
rect 2733 2973 2747 2987
rect 2833 2893 2847 2907
rect 2733 2793 2747 2807
rect 2753 2793 2767 2807
rect 2813 2753 2827 2767
rect 3073 3473 3087 3487
rect 3053 3413 3067 3427
rect 3033 3333 3047 3347
rect 2993 3293 3007 3307
rect 2953 3233 2967 3247
rect 2973 3193 2987 3207
rect 2913 3173 2927 3187
rect 2953 3133 2967 3147
rect 2893 3093 2907 3107
rect 2873 2873 2887 2887
rect 2873 2853 2887 2867
rect 2653 2693 2667 2707
rect 2633 2653 2647 2667
rect 2633 2593 2647 2607
rect 2613 2473 2627 2487
rect 2613 2293 2627 2307
rect 2613 2193 2627 2207
rect 2593 2093 2607 2107
rect 2673 2613 2687 2627
rect 2773 2733 2787 2747
rect 2833 2733 2847 2747
rect 2793 2713 2807 2727
rect 2833 2713 2847 2727
rect 2853 2713 2867 2727
rect 2733 2573 2747 2587
rect 2853 2673 2867 2687
rect 2793 2553 2807 2567
rect 2833 2553 2847 2567
rect 2673 2513 2687 2527
rect 2653 2173 2667 2187
rect 2633 2153 2647 2167
rect 2713 2433 2727 2447
rect 2693 2333 2707 2347
rect 2753 2313 2767 2327
rect 2773 2313 2787 2327
rect 2713 2293 2727 2307
rect 2693 2273 2707 2287
rect 2733 2273 2747 2287
rect 2733 2193 2747 2207
rect 2633 2073 2647 2087
rect 2613 2053 2627 2067
rect 2573 2013 2587 2027
rect 2593 1913 2607 1927
rect 2453 1753 2467 1767
rect 2433 1653 2447 1667
rect 2373 1633 2387 1647
rect 2393 1633 2407 1647
rect 2353 1613 2367 1627
rect 2333 1433 2347 1447
rect 2333 1413 2347 1427
rect 2313 1393 2327 1407
rect 2273 1353 2287 1367
rect 2413 1573 2427 1587
rect 2433 1553 2447 1567
rect 2373 1373 2387 1387
rect 2573 1753 2587 1767
rect 2493 1673 2507 1687
rect 2513 1633 2527 1647
rect 2493 1613 2507 1627
rect 2453 1493 2467 1507
rect 2453 1433 2467 1447
rect 2553 1593 2567 1607
rect 2533 1553 2547 1567
rect 2513 1533 2527 1547
rect 2493 1453 2507 1467
rect 2473 1413 2487 1427
rect 2493 1373 2507 1387
rect 2453 1353 2467 1367
rect 2333 1333 2347 1347
rect 2373 1333 2387 1347
rect 2273 1293 2287 1307
rect 2333 1293 2347 1307
rect 2293 1273 2307 1287
rect 2333 1253 2347 1267
rect 2273 1233 2287 1247
rect 2433 1313 2447 1327
rect 2613 1773 2627 1787
rect 2613 1753 2627 1767
rect 2593 1733 2607 1747
rect 2913 2993 2927 3007
rect 2893 2773 2907 2787
rect 2893 2733 2907 2747
rect 2893 2713 2907 2727
rect 2873 2653 2887 2667
rect 2873 2593 2887 2607
rect 2933 2893 2947 2907
rect 2993 3113 3007 3127
rect 3013 3053 3027 3067
rect 2993 3013 3007 3027
rect 3273 3913 3287 3927
rect 3213 3733 3227 3747
rect 3133 3693 3147 3707
rect 3213 3693 3227 3707
rect 3253 3693 3267 3707
rect 3173 3673 3187 3687
rect 3133 3633 3147 3647
rect 3193 3553 3207 3567
rect 3133 3513 3147 3527
rect 3153 3493 3167 3507
rect 3153 3453 3167 3467
rect 3233 3473 3247 3487
rect 3293 3833 3307 3847
rect 3293 3673 3307 3687
rect 3273 3453 3287 3467
rect 3193 3433 3207 3447
rect 3213 3433 3227 3447
rect 3273 3433 3287 3447
rect 3173 3413 3187 3427
rect 3233 3413 3247 3427
rect 3153 3393 3167 3407
rect 3193 3393 3207 3407
rect 3133 3373 3147 3387
rect 3073 3293 3087 3307
rect 3073 3273 3087 3287
rect 3053 3133 3067 3147
rect 3053 3013 3067 3027
rect 3033 2973 3047 2987
rect 3013 2933 3027 2947
rect 2973 2913 2987 2927
rect 2973 2853 2987 2867
rect 2953 2773 2967 2787
rect 2933 2673 2947 2687
rect 2933 2633 2947 2647
rect 2953 2633 2967 2647
rect 2913 2593 2927 2607
rect 2913 2573 2927 2587
rect 2893 2473 2907 2487
rect 2933 2413 2947 2427
rect 2933 2333 2947 2347
rect 2793 2293 2807 2307
rect 2853 2293 2867 2307
rect 2773 2153 2787 2167
rect 2733 2133 2747 2147
rect 2753 2133 2767 2147
rect 2713 2113 2727 2127
rect 2673 2093 2687 2107
rect 2693 2073 2707 2087
rect 2653 1953 2667 1967
rect 2753 2073 2767 2087
rect 2753 2053 2767 2067
rect 2813 2273 2827 2287
rect 2873 2273 2887 2287
rect 2993 2713 3007 2727
rect 2993 2673 3007 2687
rect 3113 3253 3127 3267
rect 3093 3233 3107 3247
rect 3093 3133 3107 3147
rect 3093 3073 3107 3087
rect 3093 3033 3107 3047
rect 3093 2953 3107 2967
rect 3073 2933 3087 2947
rect 3033 2833 3047 2847
rect 3053 2813 3067 2827
rect 3093 2793 3107 2807
rect 3093 2773 3107 2787
rect 3153 3293 3167 3307
rect 3133 3053 3147 3067
rect 3193 3233 3207 3247
rect 3253 3293 3267 3307
rect 3253 3193 3267 3207
rect 3213 3113 3227 3127
rect 3193 3093 3207 3107
rect 3153 3033 3167 3047
rect 3153 3013 3167 3027
rect 3133 2993 3147 3007
rect 3173 2953 3187 2967
rect 3233 3013 3247 3027
rect 3253 2993 3267 3007
rect 3213 2973 3227 2987
rect 3373 3953 3387 3967
rect 3353 3833 3367 3847
rect 3353 3633 3367 3647
rect 3353 3533 3367 3547
rect 3453 4273 3467 4287
rect 3413 4233 3427 4247
rect 3413 4173 3427 4187
rect 3633 4453 3647 4467
rect 3713 4453 3727 4467
rect 3593 4433 3607 4447
rect 3693 4433 3707 4447
rect 3733 4433 3747 4447
rect 3473 4173 3487 4187
rect 3433 4093 3447 4107
rect 3453 4093 3467 4107
rect 3433 4073 3447 4087
rect 3593 4233 3607 4247
rect 3553 4213 3567 4227
rect 3733 4313 3747 4327
rect 3713 4273 3727 4287
rect 3673 4213 3687 4227
rect 3693 4213 3707 4227
rect 3573 4193 3587 4207
rect 3633 4193 3647 4207
rect 3533 4173 3547 4187
rect 3653 4153 3667 4167
rect 3593 4113 3607 4127
rect 3513 4013 3527 4027
rect 3573 4013 3587 4027
rect 3493 3993 3507 4007
rect 3533 3993 3547 4007
rect 3673 4033 3687 4047
rect 3693 4033 3707 4047
rect 3673 4013 3687 4027
rect 3693 4013 3707 4027
rect 3453 3973 3467 3987
rect 3413 3953 3427 3967
rect 3433 3953 3447 3967
rect 3433 3873 3447 3887
rect 3393 3753 3407 3767
rect 3513 3973 3527 3987
rect 3553 3953 3567 3967
rect 3553 3933 3567 3947
rect 3493 3913 3507 3927
rect 3513 3893 3527 3907
rect 3473 3853 3487 3867
rect 3453 3673 3467 3687
rect 3393 3633 3407 3647
rect 3533 3693 3547 3707
rect 3533 3633 3547 3647
rect 3513 3613 3527 3627
rect 3513 3573 3527 3587
rect 3433 3553 3447 3567
rect 3473 3553 3487 3567
rect 3413 3513 3427 3527
rect 3353 3473 3367 3487
rect 3373 3473 3387 3487
rect 3333 3453 3347 3467
rect 3373 3433 3387 3447
rect 3333 3413 3347 3427
rect 3353 3413 3367 3427
rect 3293 3393 3307 3407
rect 3333 3233 3347 3247
rect 3353 3213 3367 3227
rect 3353 3193 3367 3207
rect 3313 3153 3327 3167
rect 3293 3053 3307 3067
rect 3313 3013 3327 3027
rect 3413 3273 3427 3287
rect 3493 3533 3507 3547
rect 3453 3513 3467 3527
rect 3473 3493 3487 3507
rect 3513 3493 3527 3507
rect 3573 3713 3587 3727
rect 3573 3693 3587 3707
rect 3653 3853 3667 3867
rect 3653 3813 3667 3827
rect 4033 4653 4047 4667
rect 3873 4633 3887 4647
rect 3913 4633 3927 4647
rect 4153 4653 4167 4667
rect 4173 4653 4187 4667
rect 4453 4653 4467 4667
rect 3833 4473 3847 4487
rect 3733 4213 3747 4227
rect 3773 4213 3787 4227
rect 3753 4193 3767 4207
rect 3753 4093 3767 4107
rect 3733 3993 3747 4007
rect 3713 3933 3727 3947
rect 3713 3913 3727 3927
rect 3813 4193 3827 4207
rect 3853 4193 3867 4207
rect 3873 4173 3887 4187
rect 3853 4113 3867 4127
rect 3833 4053 3847 4067
rect 3713 3813 3727 3827
rect 3673 3553 3687 3567
rect 3613 3513 3627 3527
rect 3753 3693 3767 3707
rect 3713 3673 3727 3687
rect 3793 3873 3807 3887
rect 3813 3753 3827 3767
rect 3793 3693 3807 3707
rect 3773 3673 3787 3687
rect 3833 3673 3847 3687
rect 3773 3633 3787 3647
rect 3753 3613 3767 3627
rect 3693 3533 3707 3547
rect 3753 3533 3767 3547
rect 3573 3493 3587 3507
rect 3613 3493 3627 3507
rect 3473 3473 3487 3487
rect 3493 3473 3507 3487
rect 3533 3473 3547 3487
rect 3473 3373 3487 3387
rect 3473 3253 3487 3267
rect 3393 3233 3407 3247
rect 3433 3213 3447 3227
rect 3393 3073 3407 3087
rect 3373 3053 3387 3067
rect 3453 3133 3467 3147
rect 3653 3433 3667 3447
rect 3553 3413 3567 3427
rect 3573 3413 3587 3427
rect 3533 3393 3547 3407
rect 3573 3353 3587 3367
rect 3593 3353 3607 3367
rect 3533 3313 3547 3327
rect 3553 3313 3567 3327
rect 3513 3253 3527 3267
rect 3753 3513 3767 3527
rect 3793 3613 3807 3627
rect 3753 3473 3767 3487
rect 3733 3413 3747 3427
rect 4033 4453 4047 4467
rect 3953 4433 3967 4447
rect 3953 4373 3967 4387
rect 4033 4413 4047 4427
rect 3993 4233 4007 4247
rect 4053 4373 4067 4387
rect 3953 4193 3967 4207
rect 3993 4193 4007 4207
rect 3933 4173 3947 4187
rect 4013 4173 4027 4187
rect 4053 4133 4067 4147
rect 3913 4113 3927 4127
rect 3893 4073 3907 4087
rect 3913 4053 3927 4067
rect 3893 4033 3907 4047
rect 3953 4013 3967 4027
rect 3893 3973 3907 3987
rect 3933 3973 3947 3987
rect 3873 3873 3887 3887
rect 3893 3873 3907 3887
rect 3873 3673 3887 3687
rect 3853 3613 3867 3627
rect 3833 3573 3847 3587
rect 3873 3553 3887 3567
rect 3833 3513 3847 3527
rect 3833 3473 3847 3487
rect 3693 3333 3707 3347
rect 3713 3313 3727 3327
rect 3633 3273 3647 3287
rect 3613 3253 3627 3267
rect 3673 3253 3687 3267
rect 3713 3253 3727 3267
rect 3513 3233 3527 3247
rect 3553 3233 3567 3247
rect 3593 3233 3607 3247
rect 3653 3233 3667 3247
rect 3753 3313 3767 3327
rect 3753 3273 3767 3287
rect 3693 3233 3707 3247
rect 3733 3233 3747 3247
rect 3533 3193 3547 3207
rect 3573 3193 3587 3207
rect 3593 3193 3607 3207
rect 3593 3133 3607 3147
rect 3613 3133 3627 3147
rect 3513 3113 3527 3127
rect 3493 3093 3507 3107
rect 3453 3073 3467 3087
rect 3553 3073 3567 3087
rect 3433 3053 3447 3067
rect 3293 2993 3307 3007
rect 3413 3033 3427 3047
rect 3393 3013 3407 3027
rect 3333 2973 3347 2987
rect 3413 2953 3427 2967
rect 3293 2933 3307 2947
rect 3273 2873 3287 2887
rect 3193 2833 3207 2847
rect 3133 2813 3147 2827
rect 3173 2813 3187 2827
rect 3273 2793 3287 2807
rect 3193 2753 3207 2767
rect 3233 2753 3247 2767
rect 3213 2733 3227 2747
rect 3113 2673 3127 2687
rect 3073 2653 3087 2667
rect 3113 2633 3127 2647
rect 3053 2553 3067 2567
rect 3093 2553 3107 2567
rect 3013 2513 3027 2527
rect 2993 2433 3007 2447
rect 3013 2393 3027 2407
rect 2973 2333 2987 2347
rect 2973 2293 2987 2307
rect 3093 2473 3107 2487
rect 3073 2373 3087 2387
rect 3033 2293 3047 2307
rect 3253 2673 3267 2687
rect 3333 2873 3347 2887
rect 3313 2813 3327 2827
rect 3293 2693 3307 2707
rect 3373 2773 3387 2787
rect 3413 2773 3427 2787
rect 3393 2753 3407 2767
rect 3353 2733 3367 2747
rect 3373 2713 3387 2727
rect 3173 2593 3187 2607
rect 3253 2593 3267 2607
rect 3273 2593 3287 2607
rect 3173 2573 3187 2587
rect 3233 2573 3247 2587
rect 3133 2553 3147 2567
rect 3153 2533 3167 2547
rect 3293 2573 3307 2587
rect 3253 2533 3267 2547
rect 3233 2513 3247 2527
rect 3273 2493 3287 2507
rect 3213 2473 3227 2487
rect 3193 2353 3207 2367
rect 3113 2313 3127 2327
rect 3173 2313 3187 2327
rect 3113 2293 3127 2307
rect 3153 2293 3167 2307
rect 3233 2373 3247 2387
rect 3253 2333 3267 2347
rect 3233 2293 3247 2307
rect 2953 2273 2967 2287
rect 2993 2273 3007 2287
rect 3033 2273 3047 2287
rect 2813 2233 2827 2247
rect 2833 2233 2847 2247
rect 2793 2093 2807 2107
rect 2813 2093 2827 2107
rect 2853 2173 2867 2187
rect 2793 2073 2807 2087
rect 2833 2073 2847 2087
rect 2813 2053 2827 2067
rect 2733 2033 2747 2047
rect 2713 1933 2727 1947
rect 2753 1933 2767 1947
rect 2693 1853 2707 1867
rect 2693 1833 2707 1847
rect 2673 1713 2687 1727
rect 2633 1673 2647 1687
rect 2673 1673 2687 1687
rect 2693 1673 2707 1687
rect 2613 1633 2627 1647
rect 2633 1573 2647 1587
rect 2693 1593 2707 1607
rect 2593 1553 2607 1567
rect 2633 1533 2647 1547
rect 2533 1473 2547 1487
rect 2573 1473 2587 1487
rect 2573 1453 2587 1467
rect 2573 1413 2587 1427
rect 2553 1353 2567 1367
rect 2593 1353 2607 1367
rect 2493 1333 2507 1347
rect 2513 1333 2527 1347
rect 2553 1313 2567 1327
rect 2593 1313 2607 1327
rect 2393 1293 2407 1307
rect 2493 1293 2507 1307
rect 2373 1273 2387 1287
rect 2273 1193 2287 1207
rect 2353 1213 2367 1227
rect 2333 1173 2347 1187
rect 2313 1153 2327 1167
rect 2253 1133 2267 1147
rect 2093 1093 2107 1107
rect 2133 1093 2147 1107
rect 2153 1093 2167 1107
rect 2213 1113 2227 1127
rect 2233 1113 2247 1127
rect 2153 1073 2167 1087
rect 2093 953 2107 967
rect 2233 1093 2247 1107
rect 2273 1093 2287 1107
rect 2313 1093 2327 1107
rect 2333 1093 2347 1107
rect 2213 1033 2227 1047
rect 2073 893 2087 907
rect 2193 933 2207 947
rect 2213 933 2227 947
rect 2293 1073 2307 1087
rect 2253 1053 2267 1067
rect 2233 913 2247 927
rect 2233 893 2247 907
rect 2273 893 2287 907
rect 2053 873 2067 887
rect 2093 873 2107 887
rect 2173 873 2187 887
rect 1893 833 1907 847
rect 1953 833 1967 847
rect 2013 833 2027 847
rect 1913 773 1927 787
rect 1893 753 1907 767
rect 1993 813 2007 827
rect 1973 793 1987 807
rect 2073 853 2087 867
rect 2133 853 2147 867
rect 2153 853 2167 867
rect 2073 813 2087 827
rect 2093 813 2107 827
rect 2013 753 2027 767
rect 2033 753 2047 767
rect 2053 753 2067 767
rect 1893 733 1907 747
rect 1933 733 1947 747
rect 1873 693 1887 707
rect 1833 653 1847 667
rect 1853 653 1867 667
rect 1733 573 1747 587
rect 1713 553 1727 567
rect 1633 453 1647 467
rect 1673 453 1687 467
rect 1693 453 1707 467
rect 1673 413 1687 427
rect 1353 233 1367 247
rect 1313 193 1327 207
rect 1233 173 1247 187
rect 1273 173 1287 187
rect 1093 133 1107 147
rect 1153 133 1167 147
rect 1193 133 1207 147
rect 1273 133 1287 147
rect 1253 113 1267 127
rect 1293 113 1307 127
rect 1373 133 1387 147
rect 1453 313 1467 327
rect 1473 253 1487 267
rect 1553 273 1567 287
rect 1533 193 1547 207
rect 1493 153 1507 167
rect 1593 233 1607 247
rect 1613 213 1627 227
rect 1573 173 1587 187
rect 1593 173 1607 187
rect 1753 453 1767 467
rect 1853 613 1867 627
rect 1793 413 1807 427
rect 1953 673 1967 687
rect 2013 673 2027 687
rect 2113 773 2127 787
rect 2113 733 2127 747
rect 2213 813 2227 827
rect 2213 793 2227 807
rect 2113 713 2127 727
rect 2173 713 2187 727
rect 1993 653 2007 667
rect 1913 633 1927 647
rect 1893 613 1907 627
rect 1933 613 1947 627
rect 1913 593 1927 607
rect 2033 613 2047 627
rect 1893 473 1907 487
rect 1773 373 1787 387
rect 1793 373 1807 387
rect 1873 373 1887 387
rect 1693 273 1707 287
rect 1673 253 1687 267
rect 1853 333 1867 347
rect 1853 273 1867 287
rect 1833 233 1847 247
rect 1713 213 1727 227
rect 1753 213 1767 227
rect 1813 213 1827 227
rect 1673 173 1687 187
rect 1653 153 1667 167
rect 1513 133 1527 147
rect 1553 133 1567 147
rect 1593 133 1607 147
rect 1633 133 1647 147
rect 1693 153 1707 167
rect 1773 173 1787 187
rect 1993 573 2007 587
rect 1953 373 1967 387
rect 1933 353 1947 367
rect 1973 353 1987 367
rect 2053 473 2067 487
rect 2033 453 2047 467
rect 2093 653 2107 667
rect 2073 413 2087 427
rect 2173 693 2187 707
rect 2253 873 2267 887
rect 2373 1153 2387 1167
rect 2373 993 2387 1007
rect 2333 873 2347 887
rect 2353 873 2367 887
rect 2313 853 2327 867
rect 2433 1233 2447 1247
rect 2573 1293 2587 1307
rect 2613 1293 2627 1307
rect 2693 1533 2707 1547
rect 2793 1853 2807 1867
rect 2813 1853 2827 1867
rect 2753 1833 2767 1847
rect 2753 1793 2767 1807
rect 2773 1773 2787 1787
rect 2733 1693 2747 1707
rect 2973 2213 2987 2227
rect 2953 2173 2967 2187
rect 2953 2133 2967 2147
rect 2953 2113 2967 2127
rect 2913 2093 2927 2107
rect 2953 2093 2967 2107
rect 3093 2273 3107 2287
rect 3133 2273 3147 2287
rect 3173 2273 3187 2287
rect 3213 2273 3227 2287
rect 3113 2253 3127 2267
rect 3153 2253 3167 2267
rect 3033 2213 3047 2227
rect 2993 2193 3007 2207
rect 3013 2193 3027 2207
rect 3093 2213 3107 2227
rect 3073 2153 3087 2167
rect 3093 2153 3107 2167
rect 2993 2133 3007 2147
rect 2873 2053 2887 2067
rect 2873 2033 2887 2047
rect 2893 1973 2907 1987
rect 2873 1813 2887 1827
rect 2853 1773 2867 1787
rect 2833 1733 2847 1747
rect 2813 1713 2827 1727
rect 2793 1673 2807 1687
rect 2733 1653 2747 1667
rect 2773 1653 2787 1667
rect 2753 1613 2767 1627
rect 2773 1593 2787 1607
rect 2873 1673 2887 1687
rect 2853 1653 2867 1667
rect 2753 1573 2767 1587
rect 2733 1553 2747 1567
rect 2773 1553 2787 1567
rect 2793 1553 2807 1567
rect 2833 1553 2847 1567
rect 2873 1553 2887 1567
rect 2713 1493 2727 1507
rect 2653 1433 2667 1447
rect 2673 1433 2687 1447
rect 2673 1393 2687 1407
rect 2693 1393 2707 1407
rect 2673 1353 2687 1367
rect 2713 1373 2727 1387
rect 2753 1513 2767 1527
rect 2793 1493 2807 1507
rect 2813 1473 2827 1487
rect 2793 1393 2807 1407
rect 2813 1373 2827 1387
rect 2873 1373 2887 1387
rect 2753 1353 2767 1367
rect 2773 1353 2787 1367
rect 2773 1313 2787 1327
rect 2653 1293 2667 1307
rect 2733 1293 2747 1307
rect 2513 1273 2527 1287
rect 2553 1273 2567 1287
rect 2453 1173 2467 1187
rect 2413 1153 2427 1167
rect 2473 1133 2487 1147
rect 2433 1113 2447 1127
rect 2533 1213 2547 1227
rect 2633 1273 2647 1287
rect 2633 1233 2647 1247
rect 2573 1153 2587 1167
rect 2593 1153 2607 1167
rect 2613 1153 2627 1167
rect 2413 1093 2427 1107
rect 2413 973 2427 987
rect 2473 1073 2487 1087
rect 2553 1113 2567 1127
rect 2513 1073 2527 1087
rect 2533 1073 2547 1087
rect 2493 1053 2507 1067
rect 2473 993 2487 1007
rect 2453 913 2467 927
rect 2573 1053 2587 1067
rect 2553 973 2567 987
rect 2533 953 2547 967
rect 2513 893 2527 907
rect 2293 833 2307 847
rect 2353 833 2367 847
rect 2273 813 2287 827
rect 2313 813 2327 827
rect 2273 773 2287 787
rect 2293 693 2307 707
rect 2313 693 2327 707
rect 2253 673 2267 687
rect 2233 653 2247 667
rect 2253 653 2267 667
rect 2133 633 2147 647
rect 2173 633 2187 647
rect 2133 593 2147 607
rect 2153 593 2167 607
rect 2113 473 2127 487
rect 2093 393 2107 407
rect 2033 373 2047 387
rect 2093 373 2107 387
rect 2013 353 2027 367
rect 2053 353 2067 367
rect 1993 333 2007 347
rect 1913 273 1927 287
rect 2293 633 2307 647
rect 2233 613 2247 627
rect 2293 613 2307 627
rect 2373 673 2387 687
rect 2333 633 2347 647
rect 2473 853 2487 867
rect 2493 853 2507 867
rect 2413 773 2427 787
rect 2513 793 2527 807
rect 2673 1193 2687 1207
rect 2713 1273 2727 1287
rect 2793 1293 2807 1307
rect 2693 1173 2707 1187
rect 2653 1073 2667 1087
rect 2653 1033 2667 1047
rect 2633 1013 2647 1027
rect 2693 973 2707 987
rect 2613 933 2627 947
rect 2653 933 2667 947
rect 2773 1153 2787 1167
rect 2833 1333 2847 1347
rect 2833 1293 2847 1307
rect 2833 1253 2847 1267
rect 2913 1953 2927 1967
rect 2973 2033 2987 2047
rect 2973 1933 2987 1947
rect 2933 1913 2947 1927
rect 2953 1833 2967 1847
rect 2913 1813 2927 1827
rect 2953 1813 2967 1827
rect 2933 1733 2947 1747
rect 2913 1713 2927 1727
rect 2913 1693 2927 1707
rect 3173 2213 3187 2227
rect 3213 2213 3227 2227
rect 3293 2433 3307 2447
rect 3353 2613 3367 2627
rect 3373 2613 3387 2627
rect 3373 2593 3387 2607
rect 3333 2573 3347 2587
rect 3353 2573 3367 2587
rect 3333 2513 3347 2527
rect 3313 2393 3327 2407
rect 3413 2733 3427 2747
rect 3533 3033 3547 3047
rect 3493 3013 3507 3027
rect 3473 2993 3487 3007
rect 3513 2993 3527 3007
rect 3453 2973 3467 2987
rect 3473 2913 3487 2927
rect 3453 2773 3467 2787
rect 3433 2693 3447 2707
rect 3413 2673 3427 2687
rect 3433 2673 3447 2687
rect 3413 2633 3427 2647
rect 3393 2573 3407 2587
rect 3393 2553 3407 2567
rect 3373 2493 3387 2507
rect 3353 2373 3367 2387
rect 3333 2313 3347 2327
rect 3353 2293 3367 2307
rect 3333 2273 3347 2287
rect 3293 2253 3307 2267
rect 3333 2253 3347 2267
rect 3173 2153 3187 2167
rect 3073 2073 3087 2087
rect 3013 2053 3027 2067
rect 3053 2053 3067 2067
rect 3093 2053 3107 2067
rect 3153 2073 3167 2087
rect 3033 2033 3047 2047
rect 2993 1913 3007 1927
rect 3013 1913 3027 1927
rect 3113 2033 3127 2047
rect 3093 2013 3107 2027
rect 3073 1873 3087 1887
rect 3033 1853 3047 1867
rect 3013 1813 3027 1827
rect 2993 1773 3007 1787
rect 3013 1773 3027 1787
rect 2993 1753 3007 1767
rect 2973 1653 2987 1667
rect 2933 1633 2947 1647
rect 2953 1613 2967 1627
rect 3053 1833 3067 1847
rect 3133 1953 3147 1967
rect 3113 1853 3127 1867
rect 3113 1833 3127 1847
rect 3093 1793 3107 1807
rect 3033 1753 3047 1767
rect 3073 1753 3087 1767
rect 3033 1713 3047 1727
rect 3113 1713 3127 1727
rect 3013 1673 3027 1687
rect 2993 1593 3007 1607
rect 2933 1573 2947 1587
rect 2973 1573 2987 1587
rect 3013 1573 3027 1587
rect 2953 1433 2967 1447
rect 2913 1373 2927 1387
rect 2893 1333 2907 1347
rect 2913 1333 2927 1347
rect 2893 1293 2907 1307
rect 2873 1253 2887 1267
rect 2873 1213 2887 1227
rect 2853 1173 2867 1187
rect 2853 1153 2867 1167
rect 2753 1093 2767 1107
rect 2833 1133 2847 1147
rect 2853 1133 2867 1147
rect 2813 1113 2827 1127
rect 3013 1533 3027 1547
rect 2973 1333 2987 1347
rect 2993 1313 3007 1327
rect 2933 1293 2947 1307
rect 2973 1293 2987 1307
rect 3113 1673 3127 1687
rect 3073 1613 3087 1627
rect 3233 2173 3247 2187
rect 3213 2113 3227 2127
rect 3193 2093 3207 2107
rect 3233 2073 3247 2087
rect 3213 2053 3227 2067
rect 3233 2053 3247 2067
rect 3253 2033 3267 2047
rect 3193 2013 3207 2027
rect 3253 2013 3267 2027
rect 3193 1993 3207 2007
rect 3173 1953 3187 1967
rect 3173 1913 3187 1927
rect 3153 1813 3167 1827
rect 3313 2233 3327 2247
rect 3313 2193 3327 2207
rect 3293 2153 3307 2167
rect 3353 2213 3367 2227
rect 3373 2193 3387 2207
rect 3353 2173 3367 2187
rect 3333 2093 3347 2107
rect 3353 2093 3367 2107
rect 3293 2053 3307 2067
rect 3373 2073 3387 2087
rect 3313 2033 3327 2047
rect 3373 2033 3387 2047
rect 3253 1873 3267 1887
rect 3273 1873 3287 1887
rect 3193 1833 3207 1847
rect 3213 1833 3227 1847
rect 3293 1833 3307 1847
rect 3253 1793 3267 1807
rect 3173 1733 3187 1747
rect 3153 1673 3167 1687
rect 3133 1593 3147 1607
rect 3233 1773 3247 1787
rect 3233 1753 3247 1767
rect 3253 1753 3267 1767
rect 3233 1733 3247 1747
rect 3213 1653 3227 1667
rect 3193 1613 3207 1627
rect 3033 1453 3047 1467
rect 3093 1553 3107 1567
rect 3133 1553 3147 1567
rect 3053 1413 3067 1427
rect 3173 1533 3187 1547
rect 3253 1713 3267 1727
rect 3353 2013 3367 2027
rect 3333 1853 3347 1867
rect 3673 3213 3687 3227
rect 3693 3213 3707 3227
rect 3653 3093 3667 3107
rect 3633 3053 3647 3067
rect 3593 3013 3607 3027
rect 3613 3013 3627 3027
rect 3573 2993 3587 3007
rect 3593 2993 3607 3007
rect 3573 2953 3587 2967
rect 3593 2853 3607 2867
rect 3553 2773 3567 2787
rect 3493 2753 3507 2767
rect 3533 2753 3547 2767
rect 3593 2753 3607 2767
rect 3473 2653 3487 2667
rect 3453 2553 3467 2567
rect 3433 2513 3447 2527
rect 3453 2513 3467 2527
rect 3513 2733 3527 2747
rect 3753 3213 3767 3227
rect 3713 3193 3727 3207
rect 3713 3173 3727 3187
rect 3753 3153 3767 3167
rect 3813 3453 3827 3467
rect 3833 3453 3847 3467
rect 3793 3433 3807 3447
rect 3793 3373 3807 3387
rect 3813 3373 3827 3387
rect 4173 4593 4187 4607
rect 4133 4553 4147 4567
rect 4353 4513 4367 4527
rect 4173 4453 4187 4467
rect 4213 4453 4227 4467
rect 4353 4453 4367 4467
rect 4373 4453 4387 4467
rect 4133 4293 4147 4307
rect 4093 4133 4107 4147
rect 4153 4173 4167 4187
rect 4273 4373 4287 4387
rect 4233 4313 4247 4327
rect 4173 4153 4187 4167
rect 4173 4133 4187 4147
rect 4153 4073 4167 4087
rect 4133 4033 4147 4047
rect 4093 3973 4107 3987
rect 4073 3953 4087 3967
rect 4033 3893 4047 3907
rect 3973 3873 3987 3887
rect 4053 3793 4067 3807
rect 4053 3753 4067 3767
rect 3933 3733 3947 3747
rect 3913 3713 3927 3727
rect 3953 3713 3967 3727
rect 3913 3693 3927 3707
rect 4033 3693 4047 3707
rect 3973 3673 3987 3687
rect 3993 3673 4007 3687
rect 4133 3773 4147 3787
rect 4293 4213 4307 4227
rect 4273 4173 4287 4187
rect 4233 4053 4247 4067
rect 4193 3973 4207 3987
rect 4253 3973 4267 3987
rect 4233 3953 4247 3967
rect 4273 3953 4287 3967
rect 4193 3813 4207 3827
rect 4153 3753 4167 3767
rect 4213 3733 4227 3747
rect 4073 3713 4087 3727
rect 4113 3713 4127 3727
rect 4153 3713 4167 3727
rect 3933 3633 3947 3647
rect 3933 3613 3947 3627
rect 3913 3553 3927 3567
rect 3893 3513 3907 3527
rect 3793 3273 3807 3287
rect 3813 3213 3827 3227
rect 3833 3213 3847 3227
rect 3913 3473 3927 3487
rect 3953 3573 3967 3587
rect 4013 3653 4027 3667
rect 4013 3533 4027 3547
rect 4013 3513 4027 3527
rect 3973 3473 3987 3487
rect 4013 3473 4027 3487
rect 4073 3673 4087 3687
rect 4053 3653 4067 3667
rect 4033 3453 4047 3467
rect 4013 3413 4027 3427
rect 3993 3313 4007 3327
rect 3913 3253 3927 3267
rect 3933 3253 3947 3267
rect 3973 3253 3987 3267
rect 3893 3233 3907 3247
rect 3933 3233 3947 3247
rect 3793 3193 3807 3207
rect 3733 3133 3747 3147
rect 3773 3133 3787 3147
rect 3713 3113 3727 3127
rect 3693 3073 3707 3087
rect 3733 3073 3747 3087
rect 3753 3053 3767 3067
rect 3633 2973 3647 2987
rect 3693 2993 3707 3007
rect 3693 2953 3707 2967
rect 3733 2953 3747 2967
rect 3713 2853 3727 2867
rect 3693 2773 3707 2787
rect 3653 2753 3667 2767
rect 3673 2713 3687 2727
rect 3633 2693 3647 2707
rect 3573 2673 3587 2687
rect 3613 2673 3627 2687
rect 3513 2613 3527 2627
rect 3553 2573 3567 2587
rect 3553 2533 3567 2547
rect 3533 2513 3547 2527
rect 3433 2433 3447 2447
rect 3493 2433 3507 2447
rect 3453 2393 3467 2407
rect 3513 2393 3527 2407
rect 3433 2293 3447 2307
rect 3413 2273 3427 2287
rect 3653 2573 3667 2587
rect 3613 2553 3627 2567
rect 3653 2533 3667 2547
rect 3633 2513 3647 2527
rect 3713 2713 3727 2727
rect 3913 3193 3927 3207
rect 3973 3213 3987 3227
rect 3873 3153 3887 3167
rect 3953 3153 3967 3167
rect 3973 3153 3987 3167
rect 4073 3633 4087 3647
rect 4153 3693 4167 3707
rect 4173 3693 4187 3707
rect 4193 3673 4207 3687
rect 4153 3633 4167 3647
rect 4133 3613 4147 3627
rect 4093 3593 4107 3607
rect 4113 3573 4127 3587
rect 4133 3573 4147 3587
rect 4073 3553 4087 3567
rect 4133 3513 4147 3527
rect 4093 3493 4107 3507
rect 4093 3473 4107 3487
rect 4073 3453 4087 3467
rect 4053 3393 4067 3407
rect 4053 3353 4067 3367
rect 4013 3293 4027 3307
rect 4053 3253 4067 3267
rect 4013 3213 4027 3227
rect 3933 3133 3947 3147
rect 3993 3133 4007 3147
rect 3833 3113 3847 3127
rect 3913 3113 3927 3127
rect 3813 3093 3827 3107
rect 3853 3033 3867 3047
rect 3893 3033 3907 3047
rect 3833 3013 3847 3027
rect 3873 3013 3887 3027
rect 3833 2973 3847 2987
rect 3793 2893 3807 2907
rect 3753 2773 3767 2787
rect 3793 2773 3807 2787
rect 3773 2753 3787 2767
rect 3773 2713 3787 2727
rect 3753 2613 3767 2627
rect 3733 2593 3747 2607
rect 3733 2553 3747 2567
rect 3693 2533 3707 2547
rect 3673 2493 3687 2507
rect 3593 2473 3607 2487
rect 3693 2453 3707 2467
rect 3573 2413 3587 2427
rect 3593 2373 3607 2387
rect 3533 2293 3547 2307
rect 3553 2273 3567 2287
rect 3473 2253 3487 2267
rect 3433 2233 3447 2247
rect 3473 2233 3487 2247
rect 3413 2213 3427 2227
rect 3413 2173 3427 2187
rect 3433 2173 3447 2187
rect 3413 2073 3427 2087
rect 3453 2153 3467 2167
rect 3453 2033 3467 2047
rect 3413 2013 3427 2027
rect 3493 2213 3507 2227
rect 3513 2213 3527 2227
rect 3553 2253 3567 2267
rect 3513 2113 3527 2127
rect 3533 2113 3547 2127
rect 3513 2073 3527 2087
rect 3493 2033 3507 2047
rect 3533 2033 3547 2047
rect 3453 1993 3467 2007
rect 3473 1993 3487 2007
rect 3513 1993 3527 2007
rect 3393 1973 3407 1987
rect 3413 1953 3427 1967
rect 3333 1813 3347 1827
rect 3393 1813 3407 1827
rect 3373 1793 3387 1807
rect 3333 1773 3347 1787
rect 3373 1773 3387 1787
rect 3813 2673 3827 2687
rect 3813 2633 3827 2647
rect 3793 2593 3807 2607
rect 3873 2893 3887 2907
rect 3873 2853 3887 2867
rect 3873 2773 3887 2787
rect 3953 3113 3967 3127
rect 4013 3113 4027 3127
rect 4013 3093 4027 3107
rect 3993 3073 4007 3087
rect 3953 3033 3967 3047
rect 3973 3033 3987 3047
rect 3953 2993 3967 3007
rect 4113 3433 4127 3447
rect 4093 3393 4107 3407
rect 4113 3273 4127 3287
rect 4113 3233 4127 3247
rect 4093 3213 4107 3227
rect 4093 3193 4107 3207
rect 4113 3153 4127 3167
rect 4133 3113 4147 3127
rect 4093 3073 4107 3087
rect 4273 3933 4287 3947
rect 4253 3813 4267 3827
rect 4233 3593 4247 3607
rect 4193 3513 4207 3527
rect 4233 3513 4247 3527
rect 4393 4333 4407 4347
rect 4573 4673 4587 4687
rect 4473 4533 4487 4547
rect 4473 4393 4487 4407
rect 4413 4213 4427 4227
rect 4453 4213 4467 4227
rect 4393 4193 4407 4207
rect 4313 4173 4327 4187
rect 4353 4173 4367 4187
rect 4313 4093 4327 4107
rect 4393 4153 4407 4167
rect 4373 4093 4387 4107
rect 4593 4633 4607 4647
rect 4593 4453 4607 4467
rect 4553 4313 4567 4327
rect 4613 4433 4627 4447
rect 4653 4673 4667 4687
rect 4733 4593 4747 4607
rect 4693 4473 4707 4487
rect 4733 4473 4747 4487
rect 4633 4413 4647 4427
rect 4513 4293 4527 4307
rect 4573 4293 4587 4307
rect 4713 4453 4727 4467
rect 4733 4433 4747 4447
rect 4573 4253 4587 4267
rect 4653 4253 4667 4267
rect 4673 4253 4687 4267
rect 4613 4233 4627 4247
rect 4373 4073 4387 4087
rect 4413 4073 4427 4087
rect 4353 4033 4367 4047
rect 4353 4013 4367 4027
rect 4413 4033 4427 4047
rect 4473 4193 4487 4207
rect 4513 4193 4527 4207
rect 4533 4193 4547 4207
rect 4573 4193 4587 4207
rect 4493 4173 4507 4187
rect 4453 4153 4467 4167
rect 4553 4173 4567 4187
rect 4793 4813 4807 4827
rect 4813 4493 4827 4507
rect 4833 4493 4847 4507
rect 5053 4713 5067 4727
rect 5033 4653 5047 4667
rect 4933 4493 4947 4507
rect 4973 4493 4987 4507
rect 5133 4673 5147 4687
rect 5113 4613 5127 4627
rect 5053 4533 5067 4547
rect 5073 4533 5087 4547
rect 4913 4473 4927 4487
rect 5013 4473 5027 4487
rect 4813 4453 4827 4467
rect 4893 4453 4907 4467
rect 4933 4453 4947 4467
rect 4793 4413 4807 4427
rect 4773 4393 4787 4407
rect 4773 4293 4787 4307
rect 4753 4233 4767 4247
rect 4693 4193 4707 4207
rect 4773 4213 4787 4227
rect 4533 4153 4547 4167
rect 4573 4153 4587 4167
rect 4453 4113 4467 4127
rect 4513 4113 4527 4127
rect 4553 4113 4567 4127
rect 4413 4013 4427 4027
rect 4433 4013 4447 4027
rect 4473 4053 4487 4067
rect 4333 3993 4347 4007
rect 4373 3993 4387 4007
rect 4453 3993 4467 4007
rect 4353 3973 4367 3987
rect 4293 3893 4307 3907
rect 4313 3753 4327 3767
rect 4333 3753 4347 3767
rect 4413 3973 4427 3987
rect 4433 3973 4447 3987
rect 4453 3953 4467 3967
rect 4393 3933 4407 3947
rect 4413 3933 4427 3947
rect 4393 3893 4407 3907
rect 4353 3733 4367 3747
rect 4393 3733 4407 3747
rect 4493 4033 4507 4047
rect 4533 3993 4547 4007
rect 4513 3973 4527 3987
rect 4493 3873 4507 3887
rect 4473 3733 4487 3747
rect 4293 3713 4307 3727
rect 4313 3713 4327 3727
rect 4373 3713 4387 3727
rect 4413 3713 4427 3727
rect 4453 3713 4467 3727
rect 4333 3693 4347 3707
rect 4273 3653 4287 3667
rect 4353 3633 4367 3647
rect 4293 3513 4307 3527
rect 4233 3493 4247 3507
rect 4333 3493 4347 3507
rect 4373 3493 4387 3507
rect 4173 3453 4187 3467
rect 4173 3433 4187 3447
rect 4173 3313 4187 3327
rect 4053 3053 4067 3067
rect 4073 3053 4087 3067
rect 4033 3033 4047 3047
rect 4013 3013 4027 3027
rect 4073 3013 4087 3027
rect 4093 3013 4107 3027
rect 4053 2993 4067 3007
rect 3913 2913 3927 2927
rect 4033 2973 4047 2987
rect 4053 2953 4067 2967
rect 4053 2913 4067 2927
rect 3933 2833 3947 2847
rect 3953 2833 3967 2847
rect 3933 2793 3947 2807
rect 3913 2753 3927 2767
rect 3853 2693 3867 2707
rect 3893 2693 3907 2707
rect 3893 2673 3907 2687
rect 3873 2613 3887 2627
rect 3913 2613 3927 2627
rect 3833 2593 3847 2607
rect 3833 2553 3847 2567
rect 3893 2593 3907 2607
rect 3853 2533 3867 2547
rect 3793 2473 3807 2487
rect 3713 2353 3727 2367
rect 3753 2353 3767 2367
rect 3673 2333 3687 2347
rect 3713 2333 3727 2347
rect 3633 2313 3647 2327
rect 3673 2313 3687 2327
rect 3633 2293 3647 2307
rect 3673 2273 3687 2287
rect 3613 2233 3627 2247
rect 3613 2193 3627 2207
rect 3633 2193 3647 2207
rect 3573 2153 3587 2167
rect 3573 2133 3587 2147
rect 3613 2133 3627 2147
rect 3633 2113 3647 2127
rect 3653 2113 3667 2127
rect 3653 2093 3667 2107
rect 3593 2033 3607 2047
rect 3773 2253 3787 2267
rect 3733 2233 3747 2247
rect 3853 2453 3867 2467
rect 3813 2373 3827 2387
rect 3813 2353 3827 2367
rect 3833 2293 3847 2307
rect 3813 2253 3827 2267
rect 3793 2213 3807 2227
rect 4193 3253 4207 3267
rect 4233 3233 4247 3247
rect 4273 3233 4287 3247
rect 4393 3473 4407 3487
rect 4353 3453 4367 3467
rect 4353 3393 4367 3407
rect 4213 3193 4227 3207
rect 4193 3153 4207 3167
rect 4253 3213 4267 3227
rect 4333 3193 4347 3207
rect 4433 3693 4447 3707
rect 4473 3653 4487 3667
rect 4453 3633 4467 3647
rect 4433 3513 4447 3527
rect 4513 3833 4527 3847
rect 4653 4153 4667 4167
rect 4633 4073 4647 4087
rect 4593 4053 4607 4067
rect 4633 4053 4647 4067
rect 4673 4093 4687 4107
rect 4713 4093 4727 4107
rect 4673 4073 4687 4087
rect 4653 4033 4667 4047
rect 4593 4013 4607 4027
rect 4633 4013 4647 4027
rect 4773 4113 4787 4127
rect 4733 4053 4747 4067
rect 4733 4033 4747 4047
rect 4693 3993 4707 4007
rect 4773 3993 4787 4007
rect 4593 3953 4607 3967
rect 4713 3973 4727 3987
rect 4653 3953 4667 3967
rect 4573 3773 4587 3787
rect 4653 3793 4667 3807
rect 4613 3773 4627 3787
rect 4533 3713 4547 3727
rect 4573 3713 4587 3727
rect 4593 3693 4607 3707
rect 4733 3913 4747 3927
rect 4673 3773 4687 3787
rect 4753 3773 4767 3787
rect 4853 4433 4867 4447
rect 4813 4353 4827 4367
rect 4833 4253 4847 4267
rect 4833 4233 4847 4247
rect 4913 4433 4927 4447
rect 4953 4433 4967 4447
rect 4873 4333 4887 4347
rect 4913 4313 4927 4327
rect 4853 4213 4867 4227
rect 4873 4193 4887 4207
rect 4813 4173 4827 4187
rect 4813 4153 4827 4167
rect 4833 4153 4847 4167
rect 4833 4093 4847 4107
rect 4813 4013 4827 4027
rect 4893 4173 4907 4187
rect 4993 4293 5007 4307
rect 4953 4273 4967 4287
rect 5133 4573 5147 4587
rect 5113 4493 5127 4507
rect 5113 4453 5127 4467
rect 4953 4193 4967 4207
rect 4973 4193 4987 4207
rect 4933 4133 4947 4147
rect 4873 4033 4887 4047
rect 4913 4033 4927 4047
rect 4853 4013 4867 4027
rect 4853 3993 4867 4007
rect 4833 3973 4847 3987
rect 4673 3733 4687 3747
rect 4573 3673 4587 3687
rect 4613 3673 4627 3687
rect 4673 3693 4687 3707
rect 4653 3673 4667 3687
rect 4553 3653 4567 3667
rect 4633 3653 4647 3667
rect 4513 3613 4527 3627
rect 4453 3493 4467 3507
rect 4493 3493 4507 3507
rect 4413 3453 4427 3467
rect 4433 3433 4447 3447
rect 4473 3393 4487 3407
rect 4533 3493 4547 3507
rect 4533 3473 4547 3487
rect 4513 3333 4527 3347
rect 4413 3293 4427 3307
rect 4393 3253 4407 3267
rect 4393 3233 4407 3247
rect 4433 3233 4447 3247
rect 4373 3193 4387 3207
rect 4393 3193 4407 3207
rect 4293 3133 4307 3147
rect 4353 3133 4367 3147
rect 4233 3113 4247 3127
rect 4193 3093 4207 3107
rect 4293 3093 4307 3107
rect 4153 3053 4167 3067
rect 4173 3053 4187 3067
rect 4253 3053 4267 3067
rect 4193 3033 4207 3047
rect 4233 3033 4247 3047
rect 4133 2993 4147 3007
rect 4173 2993 4187 3007
rect 4113 2973 4127 2987
rect 4133 2953 4147 2967
rect 4133 2893 4147 2907
rect 4153 2893 4167 2907
rect 4113 2813 4127 2827
rect 4213 2873 4227 2887
rect 4513 3213 4527 3227
rect 4413 3153 4427 3167
rect 4453 3153 4467 3167
rect 4393 3053 4407 3067
rect 4433 3053 4447 3067
rect 4313 3033 4327 3047
rect 4333 3013 4347 3027
rect 4273 2993 4287 3007
rect 4313 2993 4327 3007
rect 4313 2953 4327 2967
rect 4493 3133 4507 3147
rect 4473 3113 4487 3127
rect 4473 3033 4487 3047
rect 4433 2993 4447 3007
rect 4613 3633 4627 3647
rect 4593 3273 4607 3287
rect 4553 3253 4567 3267
rect 4573 3233 4587 3247
rect 4633 3593 4647 3607
rect 4653 3573 4667 3587
rect 4653 3553 4667 3567
rect 4633 3513 4647 3527
rect 4693 3533 4707 3547
rect 4693 3453 4707 3467
rect 4673 3373 4687 3387
rect 4793 3753 4807 3767
rect 4753 3733 4767 3747
rect 4793 3733 4807 3747
rect 4933 4013 4947 4027
rect 4893 3993 4907 4007
rect 5013 4193 5027 4207
rect 5053 4193 5067 4207
rect 5053 4153 5067 4167
rect 5073 4153 5087 4167
rect 5033 4033 5047 4047
rect 4993 4013 5007 4027
rect 5013 4013 5027 4027
rect 5053 3993 5067 4007
rect 4953 3973 4967 3987
rect 4973 3973 4987 3987
rect 4933 3953 4947 3967
rect 4913 3933 4927 3947
rect 4873 3873 4887 3887
rect 4873 3853 4887 3867
rect 4733 3713 4747 3727
rect 4733 3693 4747 3707
rect 4773 3713 4787 3727
rect 4753 3653 4767 3667
rect 4733 3533 4747 3547
rect 4913 3793 4927 3807
rect 4813 3653 4827 3667
rect 4873 3713 4887 3727
rect 4893 3713 4907 3727
rect 4813 3613 4827 3627
rect 4833 3613 4847 3627
rect 4773 3513 4787 3527
rect 4873 3533 4887 3547
rect 4833 3513 4847 3527
rect 4733 3493 4747 3507
rect 4813 3473 4827 3487
rect 5013 3973 5027 3987
rect 4993 3913 5007 3927
rect 4993 3893 5007 3907
rect 4953 3873 4967 3887
rect 4933 3733 4947 3747
rect 4933 3653 4947 3667
rect 4933 3573 4947 3587
rect 4913 3493 4927 3507
rect 4733 3413 4747 3427
rect 4893 3453 4907 3467
rect 4893 3433 4907 3447
rect 4833 3413 4847 3427
rect 4753 3273 4767 3287
rect 4713 3253 4727 3267
rect 4653 3233 4667 3247
rect 4693 3233 4707 3247
rect 4753 3233 4767 3247
rect 4793 3233 4807 3247
rect 4553 3173 4567 3187
rect 4533 3153 4547 3167
rect 4533 3113 4547 3127
rect 4633 3213 4647 3227
rect 4593 3153 4607 3167
rect 4593 3133 4607 3147
rect 4553 3073 4567 3087
rect 4573 3073 4587 3087
rect 4573 3053 4587 3067
rect 4533 3033 4547 3047
rect 4533 3013 4547 3027
rect 4553 3013 4567 3027
rect 4493 2993 4507 3007
rect 4413 2933 4427 2947
rect 4433 2933 4447 2947
rect 4513 2973 4527 2987
rect 4473 2953 4487 2967
rect 4293 2893 4307 2907
rect 4333 2893 4347 2907
rect 4253 2853 4267 2867
rect 4253 2813 4267 2827
rect 4173 2793 4187 2807
rect 3993 2753 4007 2767
rect 4053 2753 4067 2767
rect 4113 2753 4127 2767
rect 3953 2733 3967 2747
rect 3973 2733 3987 2747
rect 4013 2733 4027 2747
rect 3993 2633 4007 2647
rect 3933 2593 3947 2607
rect 3953 2573 3967 2587
rect 4033 2593 4047 2607
rect 3993 2553 4007 2567
rect 3933 2533 3947 2547
rect 3973 2533 3987 2547
rect 3933 2413 3947 2427
rect 3973 2373 3987 2387
rect 3953 2353 3967 2367
rect 3913 2333 3927 2347
rect 3893 2273 3907 2287
rect 3873 2253 3887 2267
rect 3853 2233 3867 2247
rect 3893 2233 3907 2247
rect 3933 2233 3947 2247
rect 3733 2193 3747 2207
rect 3753 2193 3767 2207
rect 3793 2193 3807 2207
rect 3813 2193 3827 2207
rect 3713 2153 3727 2167
rect 3733 2153 3747 2167
rect 3773 2153 3787 2167
rect 3753 2133 3767 2147
rect 3653 2033 3667 2047
rect 3673 2033 3687 2047
rect 3693 2013 3707 2027
rect 3633 1993 3647 2007
rect 3573 1953 3587 1967
rect 3553 1933 3567 1947
rect 3473 1813 3487 1827
rect 3613 1913 3627 1927
rect 3593 1873 3607 1887
rect 3613 1873 3627 1887
rect 3453 1793 3467 1807
rect 3493 1793 3507 1807
rect 3333 1753 3347 1767
rect 3313 1713 3327 1727
rect 3273 1653 3287 1667
rect 3313 1653 3327 1667
rect 3273 1613 3287 1627
rect 3293 1593 3307 1607
rect 3213 1533 3227 1547
rect 3193 1453 3207 1467
rect 3173 1393 3187 1407
rect 3093 1373 3107 1387
rect 3133 1373 3147 1387
rect 3073 1313 3087 1327
rect 3113 1313 3127 1327
rect 2873 1113 2887 1127
rect 2833 1093 2847 1107
rect 2873 1093 2887 1107
rect 2733 953 2747 967
rect 2773 953 2787 967
rect 2633 913 2647 927
rect 2713 913 2727 927
rect 2613 853 2627 867
rect 2653 893 2667 907
rect 2753 893 2767 907
rect 2613 833 2627 847
rect 2633 833 2647 847
rect 2693 853 2707 867
rect 2733 853 2747 867
rect 2573 813 2587 827
rect 2533 733 2547 747
rect 2553 733 2567 747
rect 2453 653 2467 667
rect 2493 653 2507 667
rect 2453 633 2467 647
rect 2513 633 2527 647
rect 2373 613 2387 627
rect 2433 613 2447 627
rect 2473 613 2487 627
rect 2313 593 2327 607
rect 2193 573 2207 587
rect 2233 533 2247 547
rect 2393 573 2407 587
rect 2233 453 2247 467
rect 2313 453 2327 467
rect 2193 373 2207 387
rect 2313 413 2327 427
rect 2133 353 2147 367
rect 2153 353 2167 367
rect 2253 353 2267 367
rect 2033 313 2047 327
rect 2093 313 2107 327
rect 2133 313 2147 327
rect 2153 313 2167 327
rect 2033 293 2047 307
rect 1893 233 1907 247
rect 1913 193 1927 207
rect 1993 193 2007 207
rect 1893 153 1907 167
rect 1793 133 1807 147
rect 1833 133 1847 147
rect 1873 133 1887 147
rect 1953 173 1967 187
rect 1973 153 1987 167
rect 1953 133 1967 147
rect 1673 113 1687 127
rect 1753 113 1767 127
rect 1793 113 1807 127
rect 1993 133 2007 147
rect 2073 233 2087 247
rect 713 73 727 87
rect 973 73 987 87
rect 2153 273 2167 287
rect 2193 333 2207 347
rect 2273 293 2287 307
rect 2293 273 2307 287
rect 2273 253 2287 267
rect 2173 233 2187 247
rect 2133 173 2147 187
rect 2113 133 2127 147
rect 2153 133 2167 147
rect 2213 173 2227 187
rect 2233 173 2247 187
rect 2193 153 2207 167
rect 2193 133 2207 147
rect 2173 113 2187 127
rect 2333 333 2347 347
rect 2693 833 2707 847
rect 2713 833 2727 847
rect 2753 833 2767 847
rect 2633 793 2647 807
rect 2673 793 2687 807
rect 2633 733 2647 747
rect 2653 733 2667 747
rect 2593 693 2607 707
rect 2613 673 2627 687
rect 2553 653 2567 667
rect 2533 613 2547 627
rect 2573 613 2587 627
rect 2553 473 2567 487
rect 2513 413 2527 427
rect 2413 393 2427 407
rect 2373 353 2387 367
rect 2353 293 2367 307
rect 2073 33 2087 47
rect 2313 173 2327 187
rect 2393 233 2407 247
rect 2373 213 2387 227
rect 2373 153 2387 167
rect 2433 373 2447 387
rect 2513 373 2527 387
rect 2573 413 2587 427
rect 2713 713 2727 727
rect 2793 853 2807 867
rect 2953 1133 2967 1147
rect 2953 1093 2967 1107
rect 2933 1073 2947 1087
rect 2973 1073 2987 1087
rect 3233 1473 3247 1487
rect 3213 1433 3227 1447
rect 3293 1553 3307 1567
rect 3473 1753 3487 1767
rect 3553 1793 3567 1807
rect 3533 1773 3547 1787
rect 3553 1773 3567 1787
rect 3433 1733 3447 1747
rect 3513 1733 3527 1747
rect 3393 1673 3407 1687
rect 3633 1833 3647 1847
rect 3633 1793 3647 1807
rect 3713 1953 3727 1967
rect 3793 2133 3807 2147
rect 3793 2053 3807 2067
rect 3893 2153 3907 2167
rect 3853 2133 3867 2147
rect 3873 2133 3887 2147
rect 3833 2093 3847 2107
rect 3753 2033 3767 2047
rect 3793 2033 3807 2047
rect 3773 2013 3787 2027
rect 3853 2053 3867 2067
rect 4033 2533 4047 2547
rect 4033 2473 4047 2487
rect 4013 2433 4027 2447
rect 4033 2433 4047 2447
rect 3993 2333 4007 2347
rect 3973 2273 3987 2287
rect 3993 2273 4007 2287
rect 3973 2233 3987 2247
rect 3993 2233 4007 2247
rect 4033 2393 4047 2407
rect 4053 2393 4067 2407
rect 4093 2713 4107 2727
rect 4173 2753 4187 2767
rect 4153 2713 4167 2727
rect 4133 2693 4147 2707
rect 4113 2653 4127 2667
rect 4313 2873 4327 2887
rect 4273 2773 4287 2787
rect 4293 2773 4307 2787
rect 4353 2773 4367 2787
rect 4193 2693 4207 2707
rect 4253 2753 4267 2767
rect 4313 2753 4327 2767
rect 4393 2753 4407 2767
rect 4253 2693 4267 2707
rect 4213 2673 4227 2687
rect 4153 2633 4167 2647
rect 4093 2613 4107 2627
rect 4253 2613 4267 2627
rect 4113 2573 4127 2587
rect 4213 2573 4227 2587
rect 4153 2553 4167 2567
rect 4173 2533 4187 2547
rect 4213 2533 4227 2547
rect 4093 2513 4107 2527
rect 4133 2513 4147 2527
rect 4193 2513 4207 2527
rect 4093 2493 4107 2507
rect 4073 2373 4087 2387
rect 4073 2293 4087 2307
rect 4213 2453 4227 2467
rect 4133 2393 4147 2407
rect 4213 2393 4227 2407
rect 4073 2273 4087 2287
rect 4093 2273 4107 2287
rect 4113 2273 4127 2287
rect 4073 2233 4087 2247
rect 4093 2233 4107 2247
rect 4013 2153 4027 2167
rect 3953 2133 3967 2147
rect 4013 2093 4027 2107
rect 4053 2093 4067 2107
rect 3893 2073 3907 2087
rect 3933 2073 3947 2087
rect 3813 1973 3827 1987
rect 3833 1973 3847 1987
rect 3773 1813 3787 1827
rect 3733 1793 3747 1807
rect 3773 1793 3787 1807
rect 3613 1773 3627 1787
rect 3553 1733 3567 1747
rect 3593 1733 3607 1747
rect 3533 1673 3547 1687
rect 3373 1593 3387 1607
rect 3433 1593 3447 1607
rect 3533 1613 3547 1627
rect 3493 1593 3507 1607
rect 3353 1573 3367 1587
rect 3413 1573 3427 1587
rect 3293 1373 3307 1387
rect 3233 1353 3247 1367
rect 3193 1333 3207 1347
rect 3153 1313 3167 1327
rect 3193 1313 3207 1327
rect 3373 1453 3387 1467
rect 3393 1433 3407 1447
rect 3313 1333 3327 1347
rect 3333 1333 3347 1347
rect 3273 1313 3287 1327
rect 3293 1313 3307 1327
rect 3373 1313 3387 1327
rect 3133 1293 3147 1307
rect 3173 1293 3187 1307
rect 3073 1273 3087 1287
rect 3113 1273 3127 1287
rect 3013 1133 3027 1147
rect 3033 1133 3047 1147
rect 3053 1113 3067 1127
rect 2913 1053 2927 1067
rect 2933 1053 2947 1067
rect 2913 973 2927 987
rect 2893 893 2907 907
rect 2813 813 2827 827
rect 2833 813 2847 827
rect 2793 733 2807 747
rect 2693 653 2707 667
rect 2653 633 2667 647
rect 2673 613 2687 627
rect 2753 673 2767 687
rect 2753 653 2767 667
rect 2713 633 2727 647
rect 2653 553 2667 567
rect 2613 473 2627 487
rect 2593 393 2607 407
rect 2573 373 2587 387
rect 2413 213 2427 227
rect 2453 353 2467 367
rect 2493 353 2507 367
rect 2493 333 2507 347
rect 2773 613 2787 627
rect 2753 593 2767 607
rect 2733 533 2747 547
rect 2693 473 2707 487
rect 2673 433 2687 447
rect 2533 313 2547 327
rect 2573 313 2587 327
rect 2513 293 2527 307
rect 2473 273 2487 287
rect 2513 253 2527 267
rect 2473 233 2487 247
rect 2453 193 2467 207
rect 2413 133 2427 147
rect 2493 173 2507 187
rect 2613 353 2627 367
rect 2613 313 2627 327
rect 2633 293 2647 307
rect 2613 253 2627 267
rect 2593 233 2607 247
rect 2633 213 2647 227
rect 2653 213 2667 227
rect 2613 133 2627 147
rect 2353 113 2367 127
rect 2553 113 2567 127
rect 2293 13 2307 27
rect 2593 13 2607 27
rect 2733 453 2747 467
rect 2793 593 2807 607
rect 2773 533 2787 547
rect 2873 833 2887 847
rect 2893 833 2907 847
rect 2873 793 2887 807
rect 2893 733 2907 747
rect 2853 693 2867 707
rect 2973 833 2987 847
rect 2953 813 2967 827
rect 2993 793 3007 807
rect 2933 713 2947 727
rect 2953 693 2967 707
rect 2933 673 2947 687
rect 2913 653 2927 667
rect 2893 633 2907 647
rect 3033 933 3047 947
rect 3213 1293 3227 1307
rect 3173 1253 3187 1267
rect 3273 1253 3287 1267
rect 3153 1173 3167 1187
rect 3193 1173 3207 1187
rect 3113 1113 3127 1127
rect 3173 1133 3187 1147
rect 3093 1073 3107 1087
rect 3153 1073 3167 1087
rect 3133 973 3147 987
rect 3233 1133 3247 1147
rect 3313 1273 3327 1287
rect 3333 1193 3347 1207
rect 3313 1113 3327 1127
rect 3353 1173 3367 1187
rect 3373 1133 3387 1147
rect 3513 1573 3527 1587
rect 3493 1553 3507 1567
rect 3493 1513 3507 1527
rect 3513 1513 3527 1527
rect 3473 1453 3487 1467
rect 3693 1773 3707 1787
rect 3593 1673 3607 1687
rect 3653 1673 3667 1687
rect 3573 1593 3587 1607
rect 3713 1753 3727 1767
rect 3733 1653 3747 1667
rect 3733 1633 3747 1647
rect 3633 1613 3647 1627
rect 3653 1613 3667 1627
rect 3693 1613 3707 1627
rect 3633 1593 3647 1607
rect 3553 1433 3567 1447
rect 3593 1493 3607 1507
rect 3473 1393 3487 1407
rect 3573 1393 3587 1407
rect 3453 1333 3467 1347
rect 3413 1293 3427 1307
rect 3433 1273 3447 1287
rect 3453 1193 3467 1207
rect 3293 1093 3307 1107
rect 3333 1093 3347 1107
rect 3253 1073 3267 1087
rect 3313 1073 3327 1087
rect 3213 1053 3227 1067
rect 3273 1013 3287 1027
rect 3293 993 3307 1007
rect 3333 993 3347 1007
rect 3253 973 3267 987
rect 3273 973 3287 987
rect 3173 933 3187 947
rect 3073 873 3087 887
rect 3033 853 3047 867
rect 3053 833 3067 847
rect 3033 793 3047 807
rect 3053 793 3067 807
rect 3133 833 3147 847
rect 3253 873 3267 887
rect 3373 933 3387 947
rect 3353 893 3367 907
rect 3333 853 3347 867
rect 3433 1093 3447 1107
rect 3393 873 3407 887
rect 3453 1053 3467 1067
rect 3693 1593 3707 1607
rect 3833 1933 3847 1947
rect 3873 1993 3887 2007
rect 3913 2053 3927 2067
rect 3953 2053 3967 2067
rect 3933 2033 3947 2047
rect 3953 2033 3967 2047
rect 3913 2013 3927 2027
rect 3893 1933 3907 1947
rect 3853 1913 3867 1927
rect 3793 1753 3807 1767
rect 3753 1593 3767 1607
rect 3813 1733 3827 1747
rect 3833 1733 3847 1747
rect 3873 1853 3887 1867
rect 3893 1833 3907 1847
rect 4013 2073 4027 2087
rect 4273 2573 4287 2587
rect 4333 2733 4347 2747
rect 4373 2733 4387 2747
rect 4413 2733 4427 2747
rect 4373 2713 4387 2727
rect 4313 2573 4327 2587
rect 4353 2573 4367 2587
rect 4333 2553 4347 2567
rect 4393 2673 4407 2687
rect 4413 2653 4427 2667
rect 4393 2573 4407 2587
rect 4453 2813 4467 2827
rect 4553 2953 4567 2967
rect 4653 3193 4667 3207
rect 4633 3053 4647 3067
rect 4773 3213 4787 3227
rect 4733 3193 4747 3207
rect 4673 3173 4687 3187
rect 4713 3173 4727 3187
rect 4773 3173 4787 3187
rect 4753 3153 4767 3167
rect 4733 3113 4747 3127
rect 4693 3073 4707 3087
rect 4733 3053 4747 3067
rect 4733 3033 4747 3047
rect 4633 3013 4647 3027
rect 4653 3013 4667 3027
rect 4613 2993 4627 3007
rect 4593 2933 4607 2947
rect 4553 2913 4567 2927
rect 4593 2913 4607 2927
rect 4513 2893 4527 2907
rect 4493 2793 4507 2807
rect 4533 2833 4547 2847
rect 4513 2773 4527 2787
rect 4473 2733 4487 2747
rect 4453 2693 4467 2707
rect 4453 2653 4467 2667
rect 4433 2573 4447 2587
rect 4433 2553 4447 2567
rect 4313 2493 4327 2507
rect 4353 2493 4367 2507
rect 4293 2473 4307 2487
rect 4273 2453 4287 2467
rect 4273 2413 4287 2427
rect 4233 2333 4247 2347
rect 4213 2313 4227 2327
rect 4173 2293 4187 2307
rect 4193 2273 4207 2287
rect 4153 2233 4167 2247
rect 4093 2213 4107 2227
rect 4133 2213 4147 2227
rect 4073 2053 4087 2067
rect 3953 1973 3967 1987
rect 3993 1973 4007 1987
rect 4033 1973 4047 1987
rect 4073 1933 4087 1947
rect 3933 1893 3947 1907
rect 4013 1853 4027 1867
rect 3973 1833 3987 1847
rect 4013 1833 4027 1847
rect 3933 1813 3947 1827
rect 3973 1793 3987 1807
rect 4053 1813 4067 1827
rect 3953 1773 3967 1787
rect 3993 1773 4007 1787
rect 3993 1753 4007 1767
rect 4013 1753 4027 1767
rect 3913 1713 3927 1727
rect 3893 1693 3907 1707
rect 3933 1693 3947 1707
rect 3893 1613 3907 1627
rect 3913 1613 3927 1627
rect 3973 1673 3987 1687
rect 3953 1613 3967 1627
rect 3853 1593 3867 1607
rect 3773 1573 3787 1587
rect 3813 1573 3827 1587
rect 3853 1573 3867 1587
rect 3933 1573 3947 1587
rect 3753 1553 3767 1567
rect 3793 1553 3807 1567
rect 3673 1513 3687 1527
rect 3613 1473 3627 1487
rect 3693 1413 3707 1427
rect 3653 1393 3667 1407
rect 3673 1393 3687 1407
rect 3633 1373 3647 1387
rect 3593 1353 3607 1367
rect 3613 1353 3627 1367
rect 3533 1313 3547 1327
rect 3553 1313 3567 1327
rect 3593 1313 3607 1327
rect 3633 1313 3647 1327
rect 3553 1293 3567 1307
rect 3493 1273 3507 1287
rect 3533 1273 3547 1287
rect 3513 1113 3527 1127
rect 3573 1173 3587 1187
rect 3493 1073 3507 1087
rect 3553 1073 3567 1087
rect 3673 1333 3687 1347
rect 3713 1333 3727 1347
rect 3693 1313 3707 1327
rect 3733 1293 3747 1307
rect 3713 1213 3727 1227
rect 3653 1133 3667 1147
rect 3653 1113 3667 1127
rect 3613 1093 3627 1107
rect 3633 1073 3647 1087
rect 3593 1053 3607 1067
rect 3633 1033 3647 1047
rect 3573 1013 3587 1027
rect 3633 1013 3647 1027
rect 3533 993 3547 1007
rect 3533 953 3547 967
rect 3593 953 3607 967
rect 3453 933 3467 947
rect 3473 933 3487 947
rect 3213 833 3227 847
rect 3133 793 3147 807
rect 3173 793 3187 807
rect 3153 773 3167 787
rect 3113 673 3127 687
rect 3033 653 3047 667
rect 3053 653 3067 667
rect 3073 653 3087 667
rect 3133 653 3147 667
rect 3013 633 3027 647
rect 2913 613 2927 627
rect 2953 613 2967 627
rect 3013 613 3027 627
rect 2933 593 2947 607
rect 2953 593 2967 607
rect 2993 593 3007 607
rect 3033 593 3047 607
rect 2873 573 2887 587
rect 2833 553 2847 567
rect 2813 493 2827 507
rect 2793 473 2807 487
rect 2793 453 2807 467
rect 2853 453 2867 467
rect 2733 373 2747 387
rect 2753 373 2767 387
rect 2833 413 2847 427
rect 2833 393 2847 407
rect 2813 373 2827 387
rect 2833 353 2847 367
rect 3073 633 3087 647
rect 3093 633 3107 647
rect 3113 613 3127 627
rect 3073 593 3087 607
rect 2973 573 2987 587
rect 3053 573 3067 587
rect 3193 773 3207 787
rect 3253 733 3267 747
rect 3233 693 3247 707
rect 3253 693 3267 707
rect 3213 673 3227 687
rect 3213 653 3227 667
rect 3193 613 3207 627
rect 3213 613 3227 627
rect 2953 553 2967 567
rect 3153 553 3167 567
rect 3173 553 3187 567
rect 3333 833 3347 847
rect 3353 833 3367 847
rect 3433 853 3447 867
rect 3433 833 3447 847
rect 3313 793 3327 807
rect 3353 793 3367 807
rect 3473 813 3487 827
rect 3693 1093 3707 1107
rect 3733 1153 3747 1167
rect 3793 1373 3807 1387
rect 3873 1553 3887 1567
rect 3833 1393 3847 1407
rect 3953 1553 3967 1567
rect 3973 1553 3987 1567
rect 3933 1493 3947 1507
rect 3893 1453 3907 1467
rect 4033 1733 4047 1747
rect 4053 1673 4067 1687
rect 4213 2253 4227 2267
rect 4253 2293 4267 2307
rect 4353 2433 4367 2447
rect 4413 2533 4427 2547
rect 4393 2513 4407 2527
rect 4393 2373 4407 2387
rect 4373 2333 4387 2347
rect 4313 2313 4327 2327
rect 4333 2313 4347 2327
rect 4273 2273 4287 2287
rect 4353 2293 4367 2307
rect 4193 2133 4207 2147
rect 4113 2113 4127 2127
rect 4153 2113 4167 2127
rect 4133 2093 4147 2107
rect 4153 2093 4167 2107
rect 4193 2093 4207 2107
rect 4253 2153 4267 2167
rect 4113 2053 4127 2067
rect 4113 1993 4127 2007
rect 4153 2073 4167 2087
rect 4173 2053 4187 2067
rect 4193 2053 4207 2067
rect 4213 2053 4227 2067
rect 4133 1953 4147 1967
rect 4133 1933 4147 1947
rect 4273 2133 4287 2147
rect 4293 2133 4307 2147
rect 4413 2353 4427 2367
rect 4513 2733 4527 2747
rect 4513 2673 4527 2687
rect 4493 2653 4507 2667
rect 4513 2633 4527 2647
rect 4473 2613 4487 2627
rect 4513 2613 4527 2627
rect 4473 2593 4487 2607
rect 4453 2453 4467 2467
rect 4433 2293 4447 2307
rect 4393 2273 4407 2287
rect 4373 2253 4387 2267
rect 4573 2893 4587 2907
rect 4553 2793 4567 2807
rect 4573 2773 4587 2787
rect 4633 2973 4647 2987
rect 4693 3013 4707 3027
rect 4713 3013 4727 3027
rect 4673 2973 4687 2987
rect 4673 2953 4687 2967
rect 4653 2893 4667 2907
rect 4613 2873 4627 2887
rect 4973 3753 4987 3767
rect 4993 3733 5007 3747
rect 4993 3693 5007 3707
rect 4953 3553 4967 3567
rect 4953 3533 4967 3547
rect 4953 3493 4967 3507
rect 4973 3493 4987 3507
rect 4893 3213 4907 3227
rect 4853 3193 4867 3207
rect 4833 3173 4847 3187
rect 4813 3153 4827 3167
rect 4853 3153 4867 3167
rect 4793 3133 4807 3147
rect 4793 3093 4807 3107
rect 4813 3093 4827 3107
rect 4793 3073 4807 3087
rect 4833 3053 4847 3067
rect 5133 4233 5147 4247
rect 5113 4153 5127 4167
rect 5093 4013 5107 4027
rect 5033 3933 5047 3947
rect 5033 3913 5047 3927
rect 5033 3573 5047 3587
rect 5033 3513 5047 3527
rect 4973 3473 4987 3487
rect 5013 3473 5027 3487
rect 4913 3153 4927 3167
rect 4913 3113 4927 3127
rect 4893 3073 4907 3087
rect 4773 3013 4787 3027
rect 4853 3013 4867 3027
rect 4793 2973 4807 2987
rect 4753 2953 4767 2967
rect 4713 2933 4727 2947
rect 4693 2873 4707 2887
rect 4693 2853 4707 2867
rect 4673 2833 4687 2847
rect 4653 2773 4667 2787
rect 4593 2753 4607 2767
rect 4613 2753 4627 2767
rect 4553 2733 4567 2747
rect 4673 2753 4687 2767
rect 4593 2693 4607 2707
rect 4573 2633 4587 2647
rect 4553 2573 4567 2587
rect 4533 2493 4547 2507
rect 4493 2433 4507 2447
rect 4473 2313 4487 2327
rect 4513 2293 4527 2307
rect 4493 2273 4507 2287
rect 4353 2213 4367 2227
rect 4333 2113 4347 2127
rect 4293 2093 4307 2107
rect 4313 2093 4327 2107
rect 4273 2073 4287 2087
rect 4293 2053 4307 2067
rect 4273 2033 4287 2047
rect 4233 2013 4247 2027
rect 4253 2013 4267 2027
rect 4293 2013 4307 2027
rect 4233 1973 4247 1987
rect 4273 1973 4287 1987
rect 4213 1953 4227 1967
rect 4193 1853 4207 1867
rect 4213 1833 4227 1847
rect 4173 1813 4187 1827
rect 4133 1793 4147 1807
rect 4093 1753 4107 1767
rect 4133 1753 4147 1767
rect 4173 1773 4187 1787
rect 4133 1733 4147 1747
rect 4153 1733 4167 1747
rect 4113 1713 4127 1727
rect 4113 1693 4127 1707
rect 4133 1693 4147 1707
rect 4093 1653 4107 1667
rect 4073 1633 4087 1647
rect 4013 1593 4027 1607
rect 4093 1593 4107 1607
rect 4033 1573 4047 1587
rect 4073 1573 4087 1587
rect 4013 1553 4027 1567
rect 4053 1553 4067 1567
rect 3973 1513 3987 1527
rect 3973 1473 3987 1487
rect 3953 1413 3967 1427
rect 3953 1393 3967 1407
rect 3993 1393 4007 1407
rect 3873 1373 3887 1387
rect 3933 1353 3947 1367
rect 3773 1333 3787 1347
rect 3813 1333 3827 1347
rect 3853 1333 3867 1347
rect 3893 1333 3907 1347
rect 3793 1233 3807 1247
rect 3913 1293 3927 1307
rect 3873 1273 3887 1287
rect 3833 1253 3847 1267
rect 3813 1193 3827 1207
rect 3773 1173 3787 1187
rect 3713 1073 3727 1087
rect 3673 1033 3687 1047
rect 3813 1113 3827 1127
rect 3993 1373 4007 1387
rect 3973 1333 3987 1347
rect 4073 1513 4087 1527
rect 4073 1433 4087 1447
rect 4033 1413 4047 1427
rect 4053 1353 4067 1367
rect 4013 1333 4027 1347
rect 4033 1333 4047 1347
rect 3993 1293 4007 1307
rect 3953 1253 3967 1267
rect 4033 1253 4047 1267
rect 4013 1213 4027 1227
rect 3933 1193 3947 1207
rect 3913 1173 3927 1187
rect 3933 1173 3947 1187
rect 3993 1173 4007 1187
rect 3793 1093 3807 1107
rect 3873 1093 3887 1107
rect 3913 1093 3927 1107
rect 3833 1073 3847 1087
rect 3773 993 3787 1007
rect 3753 893 3767 907
rect 3793 893 3807 907
rect 3653 873 3667 887
rect 3633 833 3647 847
rect 3493 773 3507 787
rect 3413 753 3427 767
rect 3553 813 3567 827
rect 3573 813 3587 827
rect 3653 813 3667 827
rect 3673 813 3687 827
rect 3613 753 3627 767
rect 3513 733 3527 747
rect 3273 673 3287 687
rect 3353 673 3367 687
rect 3433 673 3447 687
rect 3273 653 3287 667
rect 3293 593 3307 607
rect 3333 553 3347 567
rect 3213 533 3227 547
rect 3073 513 3087 527
rect 2933 393 2947 407
rect 2893 373 2907 387
rect 3033 373 3047 387
rect 3093 473 3107 487
rect 2713 333 2727 347
rect 2693 213 2707 227
rect 2693 173 2707 187
rect 2873 333 2887 347
rect 2833 313 2847 327
rect 2753 293 2767 307
rect 2933 353 2947 367
rect 2973 353 2987 367
rect 2913 313 2927 327
rect 2933 273 2947 287
rect 2753 253 2767 267
rect 2893 253 2907 267
rect 2753 213 2767 227
rect 2733 173 2747 187
rect 2873 173 2887 187
rect 2833 153 2847 167
rect 2993 333 3007 347
rect 2993 213 3007 227
rect 2953 193 2967 207
rect 3033 353 3047 367
rect 3013 173 3027 187
rect 2853 133 2867 147
rect 2993 153 3007 167
rect 3113 453 3127 467
rect 3213 413 3227 427
rect 3373 653 3387 667
rect 3393 633 3407 647
rect 3453 653 3467 667
rect 3513 653 3527 667
rect 3613 653 3627 667
rect 3733 853 3747 867
rect 3773 853 3787 867
rect 3813 853 3827 867
rect 3853 853 3867 867
rect 3713 833 3727 847
rect 3753 833 3767 847
rect 3673 793 3687 807
rect 3693 793 3707 807
rect 3793 813 3807 827
rect 3693 773 3707 787
rect 3773 773 3787 787
rect 3673 693 3687 707
rect 3653 673 3667 687
rect 3413 613 3427 627
rect 3433 593 3447 607
rect 3493 613 3507 627
rect 3573 633 3587 647
rect 3593 613 3607 627
rect 3513 593 3527 607
rect 3553 593 3567 607
rect 3433 513 3447 527
rect 3633 593 3647 607
rect 3633 573 3647 587
rect 3613 513 3627 527
rect 3593 433 3607 447
rect 3133 373 3147 387
rect 3173 373 3187 387
rect 3213 373 3227 387
rect 3253 373 3267 387
rect 3293 373 3307 387
rect 3313 373 3327 387
rect 3333 373 3347 387
rect 3353 373 3367 387
rect 3413 373 3427 387
rect 3113 353 3127 367
rect 3153 353 3167 367
rect 3093 333 3107 347
rect 3173 313 3187 327
rect 3153 293 3167 307
rect 3173 293 3187 307
rect 3053 273 3067 287
rect 3093 273 3107 287
rect 3133 173 3147 187
rect 3013 133 3027 147
rect 3073 133 3087 147
rect 3113 133 3127 147
rect 3373 353 3387 367
rect 3273 333 3287 347
rect 3313 333 3327 347
rect 3253 313 3267 327
rect 3353 313 3367 327
rect 3193 253 3207 267
rect 3233 253 3247 267
rect 3393 253 3407 267
rect 3433 353 3447 367
rect 3493 373 3507 387
rect 3553 373 3567 387
rect 3513 353 3527 367
rect 3553 353 3567 367
rect 3593 353 3607 367
rect 3473 333 3487 347
rect 3453 313 3467 327
rect 3433 293 3447 307
rect 3953 1153 3967 1167
rect 4013 1133 4027 1147
rect 4033 1113 4047 1127
rect 4093 1353 4107 1367
rect 4073 1333 4087 1347
rect 4253 1953 4267 1967
rect 4193 1733 4207 1747
rect 4193 1713 4207 1727
rect 4133 1653 4147 1667
rect 4173 1653 4187 1667
rect 4153 1633 4167 1647
rect 4133 1613 4147 1627
rect 4133 1573 4147 1587
rect 4133 1553 4147 1567
rect 4133 1353 4147 1367
rect 4133 1313 4147 1327
rect 4073 1273 4087 1287
rect 4113 1213 4127 1227
rect 4133 1173 4147 1187
rect 4113 1153 4127 1167
rect 4133 1133 4147 1147
rect 3993 1093 4007 1107
rect 4013 1093 4027 1107
rect 4053 1093 4067 1107
rect 4093 1093 4107 1107
rect 3953 1033 3967 1047
rect 3973 1033 3987 1047
rect 3893 953 3907 967
rect 3893 933 3907 947
rect 3933 933 3947 947
rect 3833 833 3847 847
rect 3873 833 3887 847
rect 4093 1073 4107 1087
rect 4113 1073 4127 1087
rect 3993 993 4007 1007
rect 4053 993 4067 1007
rect 3973 953 3987 967
rect 3933 893 3947 907
rect 3953 893 3967 907
rect 3933 853 3947 867
rect 4093 973 4107 987
rect 4093 933 4107 947
rect 4053 873 4067 887
rect 4013 833 4027 847
rect 3833 673 3847 687
rect 3713 653 3727 667
rect 3773 653 3787 667
rect 3813 653 3827 667
rect 3753 633 3767 647
rect 3693 613 3707 627
rect 3733 613 3747 627
rect 3653 413 3667 427
rect 3793 613 3807 627
rect 3773 593 3787 607
rect 3753 573 3767 587
rect 3813 493 3827 507
rect 3813 433 3827 447
rect 3633 353 3647 367
rect 3693 373 3707 387
rect 3733 373 3747 387
rect 3753 373 3767 387
rect 3613 333 3627 347
rect 3653 333 3667 347
rect 3713 353 3727 367
rect 3753 353 3767 367
rect 3673 313 3687 327
rect 3533 293 3547 307
rect 3533 273 3547 287
rect 3673 273 3687 287
rect 3773 333 3787 347
rect 3753 313 3767 327
rect 3733 293 3747 307
rect 3513 253 3527 267
rect 3713 253 3727 267
rect 3573 233 3587 247
rect 3253 213 3267 227
rect 3413 213 3427 227
rect 3533 213 3547 227
rect 3213 173 3227 187
rect 3393 193 3407 207
rect 3513 193 3527 207
rect 3313 173 3327 187
rect 3273 153 3287 167
rect 3353 153 3367 167
rect 3293 133 3307 147
rect 2713 113 2727 127
rect 2953 113 2967 127
rect 3113 113 3127 127
rect 3153 113 3167 127
rect 3193 113 3207 127
rect 3213 113 3227 127
rect 3453 173 3467 187
rect 3493 173 3507 187
rect 3413 153 3427 167
rect 3473 153 3487 167
rect 3653 213 3667 227
rect 3593 173 3607 187
rect 3733 173 3747 187
rect 3453 133 3467 147
rect 3553 133 3567 147
rect 3893 793 3907 807
rect 3853 653 3867 667
rect 3873 653 3887 667
rect 3913 733 3927 747
rect 3993 813 4007 827
rect 4013 813 4027 827
rect 3953 673 3967 687
rect 3993 653 4007 667
rect 3973 633 3987 647
rect 3953 613 3967 627
rect 3973 593 3987 607
rect 3993 573 4007 587
rect 3913 553 3927 567
rect 3913 433 3927 447
rect 3893 413 3907 427
rect 3913 393 3927 407
rect 3853 373 3867 387
rect 3813 333 3827 347
rect 3833 333 3847 347
rect 3873 313 3887 327
rect 3813 293 3827 307
rect 3873 293 3887 307
rect 3793 233 3807 247
rect 3873 193 3887 207
rect 3973 313 3987 327
rect 4073 853 4087 867
rect 4073 813 4087 827
rect 4053 793 4067 807
rect 4033 733 4047 747
rect 4073 693 4087 707
rect 4173 1613 4187 1627
rect 4293 1933 4307 1947
rect 4413 2233 4427 2247
rect 4473 2233 4487 2247
rect 4393 2153 4407 2167
rect 4373 2073 4387 2087
rect 4533 2273 4547 2287
rect 4533 2253 4547 2267
rect 4513 2213 4527 2227
rect 4473 2193 4487 2207
rect 4433 2093 4447 2107
rect 4453 2093 4467 2107
rect 4413 2073 4427 2087
rect 4373 2033 4387 2047
rect 4453 2073 4467 2087
rect 4513 2093 4527 2107
rect 4433 2053 4447 2067
rect 4433 1993 4447 2007
rect 4313 1913 4327 1927
rect 4353 1913 4367 1927
rect 4293 1893 4307 1907
rect 4293 1873 4307 1887
rect 4433 1893 4447 1907
rect 4373 1873 4387 1887
rect 4353 1853 4367 1867
rect 4333 1813 4347 1827
rect 4353 1813 4367 1827
rect 4493 2053 4507 2067
rect 4473 2033 4487 2047
rect 4533 2033 4547 2047
rect 4513 2013 4527 2027
rect 4473 1993 4487 2007
rect 4493 1913 4507 1927
rect 4293 1773 4307 1787
rect 4273 1733 4287 1747
rect 4373 1793 4387 1807
rect 4413 1793 4427 1807
rect 4333 1773 4347 1787
rect 4313 1753 4327 1767
rect 4293 1713 4307 1727
rect 4253 1653 4267 1667
rect 4253 1633 4267 1647
rect 4293 1633 4307 1647
rect 4193 1533 4207 1547
rect 4213 1513 4227 1527
rect 4253 1533 4267 1547
rect 4233 1493 4247 1507
rect 4253 1473 4267 1487
rect 4273 1473 4287 1487
rect 4173 1373 4187 1387
rect 4213 1373 4227 1387
rect 4193 1313 4207 1327
rect 4273 1393 4287 1407
rect 4253 1353 4267 1367
rect 4353 1693 4367 1707
rect 4413 1733 4427 1747
rect 4393 1673 4407 1687
rect 4333 1613 4347 1627
rect 4373 1613 4387 1627
rect 4373 1593 4387 1607
rect 4333 1573 4347 1587
rect 4313 1553 4327 1567
rect 4453 1833 4467 1847
rect 4473 1793 4487 1807
rect 4453 1753 4467 1767
rect 4473 1753 4487 1767
rect 4473 1713 4487 1727
rect 4473 1673 4487 1687
rect 4493 1673 4507 1687
rect 4653 2713 4667 2727
rect 4693 2713 4707 2727
rect 4673 2693 4687 2707
rect 4653 2633 4667 2647
rect 4633 2593 4647 2607
rect 4593 2573 4607 2587
rect 4613 2573 4627 2587
rect 4573 2493 4587 2507
rect 4633 2513 4647 2527
rect 4633 2493 4647 2507
rect 4613 2453 4627 2467
rect 4593 2433 4607 2447
rect 4793 2913 4807 2927
rect 4753 2893 4767 2907
rect 4773 2873 4787 2887
rect 4793 2833 4807 2847
rect 4813 2833 4827 2847
rect 4713 2693 4727 2707
rect 4773 2773 4787 2787
rect 4893 3013 4907 3027
rect 4873 2913 4887 2927
rect 4953 3233 4967 3247
rect 4893 2893 4907 2907
rect 4853 2873 4867 2887
rect 4893 2813 4907 2827
rect 4833 2793 4847 2807
rect 4853 2773 4867 2787
rect 4793 2753 4807 2767
rect 4813 2753 4827 2767
rect 4853 2753 4867 2767
rect 4733 2593 4747 2607
rect 4733 2573 4747 2587
rect 4693 2553 4707 2567
rect 4733 2533 4747 2547
rect 4673 2513 4687 2527
rect 4713 2513 4727 2527
rect 4673 2453 4687 2467
rect 4653 2313 4667 2327
rect 4593 2293 4607 2307
rect 4573 2193 4587 2207
rect 4653 2273 4667 2287
rect 4633 2253 4647 2267
rect 4613 2173 4627 2187
rect 4613 2133 4627 2147
rect 4573 2113 4587 2127
rect 4773 2633 4787 2647
rect 4773 2613 4787 2627
rect 4773 2573 4787 2587
rect 4833 2693 4847 2707
rect 4873 2733 4887 2747
rect 4873 2713 4887 2727
rect 4853 2613 4867 2627
rect 4833 2533 4847 2547
rect 4793 2453 4807 2467
rect 4793 2433 4807 2447
rect 4753 2413 4767 2427
rect 4793 2393 4807 2407
rect 4713 2333 4727 2347
rect 4733 2333 4747 2347
rect 4693 2313 4707 2327
rect 4753 2293 4767 2307
rect 4813 2333 4827 2347
rect 4753 2273 4767 2287
rect 4793 2273 4807 2287
rect 4733 2253 4747 2267
rect 4693 2153 4707 2167
rect 4693 2133 4707 2147
rect 4633 2093 4647 2107
rect 4653 2073 4667 2087
rect 4613 2053 4627 2067
rect 4653 2053 4667 2067
rect 4713 2113 4727 2127
rect 4713 2073 4727 2087
rect 4633 2033 4647 2047
rect 4673 2033 4687 2047
rect 4613 1993 4627 2007
rect 4553 1973 4567 1987
rect 4533 1953 4547 1967
rect 4593 1853 4607 1867
rect 4553 1813 4567 1827
rect 4553 1793 4567 1807
rect 4633 1853 4647 1867
rect 4613 1813 4627 1827
rect 4413 1593 4427 1607
rect 4513 1633 4527 1647
rect 4453 1613 4467 1627
rect 4473 1613 4487 1627
rect 4493 1613 4507 1627
rect 4573 1753 4587 1767
rect 4793 2153 4807 2167
rect 4773 2093 4787 2107
rect 4933 2893 4947 2907
rect 4953 2813 4967 2827
rect 5013 3453 5027 3467
rect 5073 3933 5087 3947
rect 5073 3893 5087 3907
rect 5073 3833 5087 3847
rect 5073 3513 5087 3527
rect 5133 4073 5147 4087
rect 5133 4033 5147 4047
rect 5133 3913 5147 3927
rect 5133 3893 5147 3907
rect 5113 3633 5127 3647
rect 5133 3453 5147 3467
rect 5093 3433 5107 3447
rect 5053 3413 5067 3427
rect 5133 3313 5147 3327
rect 5113 3273 5127 3287
rect 5013 3233 5027 3247
rect 4993 3213 5007 3227
rect 5053 3213 5067 3227
rect 5073 3213 5087 3227
rect 5013 3173 5027 3187
rect 5033 3173 5047 3187
rect 5053 3153 5067 3167
rect 4993 3033 5007 3047
rect 5033 3033 5047 3047
rect 5113 3193 5127 3207
rect 5093 3093 5107 3107
rect 5073 3053 5087 3067
rect 4993 2993 5007 3007
rect 5053 3013 5067 3027
rect 5013 2973 5027 2987
rect 5033 2953 5047 2967
rect 4993 2893 5007 2907
rect 5013 2873 5027 2887
rect 4993 2833 5007 2847
rect 4933 2793 4947 2807
rect 4973 2793 4987 2807
rect 4913 2693 4927 2707
rect 4893 2673 4907 2687
rect 4973 2753 4987 2767
rect 4993 2733 5007 2747
rect 4953 2673 4967 2687
rect 4933 2653 4947 2667
rect 4893 2593 4907 2607
rect 4913 2593 4927 2607
rect 4913 2573 4927 2587
rect 4973 2613 4987 2627
rect 5013 2653 5027 2667
rect 5013 2573 5027 2587
rect 4973 2553 4987 2567
rect 4913 2533 4927 2547
rect 4893 2513 4907 2527
rect 4893 2493 4907 2507
rect 4873 2313 4887 2327
rect 5013 2533 5027 2547
rect 4933 2513 4947 2527
rect 4953 2513 4967 2527
rect 4913 2473 4927 2487
rect 4993 2413 5007 2427
rect 4893 2293 4907 2307
rect 4933 2293 4947 2307
rect 4833 2273 4847 2287
rect 4873 2273 4887 2287
rect 4933 2273 4947 2287
rect 4853 2213 4867 2227
rect 4813 2113 4827 2127
rect 4833 2093 4847 2107
rect 4873 2093 4887 2107
rect 4793 2053 4807 2067
rect 4813 2053 4827 2067
rect 4953 2233 4967 2247
rect 4953 2193 4967 2207
rect 4933 2093 4947 2107
rect 4913 2073 4927 2087
rect 4853 2053 4867 2067
rect 4773 2033 4787 2047
rect 4753 1973 4767 1987
rect 4713 1953 4727 1967
rect 4733 1953 4747 1967
rect 4673 1833 4687 1847
rect 4713 1813 4727 1827
rect 4693 1793 4707 1807
rect 4673 1773 4687 1787
rect 4573 1733 4587 1747
rect 4593 1733 4607 1747
rect 4353 1513 4367 1527
rect 4313 1453 4327 1467
rect 4293 1373 4307 1387
rect 4233 1333 4247 1347
rect 4273 1333 4287 1347
rect 4313 1353 4327 1367
rect 4333 1333 4347 1347
rect 4433 1553 4447 1567
rect 4413 1513 4427 1527
rect 4433 1493 4447 1507
rect 4413 1473 4427 1487
rect 4393 1453 4407 1467
rect 4173 1273 4187 1287
rect 4193 1273 4207 1287
rect 4173 1253 4187 1267
rect 4193 1133 4207 1147
rect 4213 1133 4227 1147
rect 4193 1093 4207 1107
rect 4173 1053 4187 1067
rect 4333 1313 4347 1327
rect 4313 1293 4327 1307
rect 4253 1273 4267 1287
rect 4293 1273 4307 1287
rect 4293 1233 4307 1247
rect 4313 1233 4327 1247
rect 4373 1293 4387 1307
rect 4353 1253 4367 1267
rect 4353 1233 4367 1247
rect 4253 1193 4267 1207
rect 4333 1193 4347 1207
rect 4233 993 4247 1007
rect 4233 973 4247 987
rect 4193 953 4207 967
rect 4113 873 4127 887
rect 4153 873 4167 887
rect 4113 833 4127 847
rect 4153 833 4167 847
rect 4133 773 4147 787
rect 4173 813 4187 827
rect 4153 753 4167 767
rect 4213 853 4227 867
rect 4293 1173 4307 1187
rect 4333 1113 4347 1127
rect 4273 1093 4287 1107
rect 4333 1073 4347 1087
rect 4313 1053 4327 1067
rect 4313 913 4327 927
rect 4293 873 4307 887
rect 4213 833 4227 847
rect 4253 853 4267 867
rect 4233 773 4247 787
rect 4193 733 4207 747
rect 4253 693 4267 707
rect 4193 673 4207 687
rect 4093 633 4107 647
rect 4053 613 4067 627
rect 4033 593 4047 607
rect 4073 573 4087 587
rect 4033 433 4047 447
rect 3953 293 3967 307
rect 3993 293 4007 307
rect 4013 293 4027 307
rect 3953 253 3967 267
rect 3673 133 3687 147
rect 3713 133 3727 147
rect 3913 153 3927 167
rect 3753 133 3767 147
rect 3833 133 3847 147
rect 3773 113 3787 127
rect 3973 113 3987 127
rect 4173 653 4187 667
rect 4213 653 4227 667
rect 4273 653 4287 667
rect 4193 633 4207 647
rect 4193 613 4207 627
rect 4233 613 4247 627
rect 4253 613 4267 627
rect 4173 593 4187 607
rect 4133 573 4147 587
rect 4193 573 4207 587
rect 4273 593 4287 607
rect 4253 473 4267 487
rect 4273 393 4287 407
rect 4173 373 4187 387
rect 4053 333 4067 347
rect 4113 333 4127 347
rect 4093 313 4107 327
rect 4173 353 4187 367
rect 4133 293 4147 307
rect 4033 253 4047 267
rect 4073 253 4087 267
rect 4033 133 4047 147
rect 4113 173 4127 187
rect 4113 153 4127 167
rect 4193 333 4207 347
rect 4213 253 4227 267
rect 4213 173 4227 187
rect 4253 173 4267 187
rect 4173 153 4187 167
rect 4153 133 4167 147
rect 4373 1213 4387 1227
rect 4393 1173 4407 1187
rect 4433 1353 4447 1367
rect 4513 1593 4527 1607
rect 4553 1593 4567 1607
rect 4493 1573 4507 1587
rect 4513 1513 4527 1527
rect 4493 1433 4507 1447
rect 4473 1393 4487 1407
rect 4493 1333 4507 1347
rect 4433 1313 4447 1327
rect 4453 1313 4467 1327
rect 4473 1313 4487 1327
rect 4553 1553 4567 1567
rect 4553 1513 4567 1527
rect 4593 1653 4607 1667
rect 4613 1653 4627 1667
rect 4573 1493 4587 1507
rect 4533 1473 4547 1487
rect 4673 1733 4687 1747
rect 4653 1693 4667 1707
rect 4733 1753 4747 1767
rect 4733 1713 4747 1727
rect 4713 1673 4727 1687
rect 4733 1673 4747 1687
rect 4673 1633 4687 1647
rect 4613 1613 4627 1627
rect 4633 1613 4647 1627
rect 4633 1593 4647 1607
rect 4733 1613 4747 1627
rect 4833 1973 4847 1987
rect 4773 1833 4787 1847
rect 4933 2053 4947 2067
rect 4893 2033 4907 2047
rect 5073 2933 5087 2947
rect 5053 2913 5067 2927
rect 5073 2813 5087 2827
rect 5073 2753 5087 2767
rect 5053 2613 5067 2627
rect 5073 2533 5087 2547
rect 5073 2513 5087 2527
rect 5053 2433 5067 2447
rect 5033 2393 5047 2407
rect 5113 3033 5127 3047
rect 5113 3013 5127 3027
rect 5113 2813 5127 2827
rect 5113 2793 5127 2807
rect 5113 2713 5127 2727
rect 5113 2693 5127 2707
rect 5093 2453 5107 2467
rect 5093 2433 5107 2447
rect 5073 2333 5087 2347
rect 5073 2313 5087 2327
rect 5013 2273 5027 2287
rect 4993 2233 5007 2247
rect 5013 2233 5027 2247
rect 5053 2273 5067 2287
rect 5073 2253 5087 2267
rect 5053 2233 5067 2247
rect 5033 2213 5047 2227
rect 4973 2173 4987 2187
rect 4993 2173 5007 2187
rect 5013 2093 5027 2107
rect 5033 2073 5047 2087
rect 4973 2053 4987 2067
rect 4993 2053 5007 2067
rect 4873 2013 4887 2027
rect 4953 2013 4967 2027
rect 4973 2013 4987 2027
rect 4853 1913 4867 1927
rect 4853 1893 4867 1907
rect 4793 1793 4807 1807
rect 4773 1773 4787 1787
rect 4773 1713 4787 1727
rect 4753 1593 4767 1607
rect 4693 1553 4707 1567
rect 4653 1533 4667 1547
rect 4673 1513 4687 1527
rect 4593 1453 4607 1467
rect 4673 1433 4687 1447
rect 4653 1413 4667 1427
rect 4613 1393 4627 1407
rect 4613 1373 4627 1387
rect 4633 1373 4647 1387
rect 4553 1333 4567 1347
rect 4593 1333 4607 1347
rect 4493 1293 4507 1307
rect 4513 1293 4527 1307
rect 4433 1273 4447 1287
rect 4433 1233 4447 1247
rect 4473 1253 4487 1267
rect 4513 1253 4527 1267
rect 4453 1213 4467 1227
rect 4373 1133 4387 1147
rect 4433 1113 4447 1127
rect 4553 1313 4567 1327
rect 4533 1213 4547 1227
rect 4513 1193 4527 1207
rect 4593 1293 4607 1307
rect 4573 1273 4587 1287
rect 4633 1333 4647 1347
rect 4653 1313 4667 1327
rect 4753 1573 4767 1587
rect 4793 1693 4807 1707
rect 4833 1773 4847 1787
rect 4833 1693 4847 1707
rect 4793 1653 4807 1667
rect 4813 1653 4827 1667
rect 4793 1633 4807 1647
rect 4813 1613 4827 1627
rect 4973 1933 4987 1947
rect 4913 1873 4927 1887
rect 5013 2033 5027 2047
rect 5033 2033 5047 2047
rect 4993 1853 5007 1867
rect 4893 1833 4907 1847
rect 4913 1833 4927 1847
rect 4933 1813 4947 1827
rect 4913 1793 4927 1807
rect 4873 1733 4887 1747
rect 4873 1693 4887 1707
rect 4853 1613 4867 1627
rect 4733 1553 4747 1567
rect 4773 1553 4787 1567
rect 4813 1553 4827 1567
rect 4713 1533 4727 1547
rect 4713 1413 4727 1427
rect 4833 1533 4847 1547
rect 4753 1413 4767 1427
rect 4733 1353 4747 1367
rect 4933 1773 4947 1787
rect 5093 2213 5107 2227
rect 5073 2033 5087 2047
rect 5053 1973 5067 1987
rect 5073 1953 5087 1967
rect 5053 1933 5067 1947
rect 5013 1793 5027 1807
rect 4993 1773 5007 1787
rect 5033 1773 5047 1787
rect 4973 1753 4987 1767
rect 5013 1733 5027 1747
rect 4913 1673 4927 1687
rect 4893 1633 4907 1647
rect 4913 1613 4927 1627
rect 4973 1593 4987 1607
rect 4913 1573 4927 1587
rect 4953 1573 4967 1587
rect 4993 1573 5007 1587
rect 4953 1533 4967 1547
rect 4853 1493 4867 1507
rect 4813 1373 4827 1387
rect 4773 1333 4787 1347
rect 4573 1213 4587 1227
rect 4593 1213 4607 1227
rect 4553 1173 4567 1187
rect 4513 1153 4527 1167
rect 4553 1153 4567 1167
rect 4493 1133 4507 1147
rect 4393 1073 4407 1087
rect 4353 973 4367 987
rect 4333 853 4347 867
rect 4433 1073 4447 1087
rect 4413 1053 4427 1067
rect 4513 1093 4527 1107
rect 4493 1073 4507 1087
rect 4433 1033 4447 1047
rect 4453 1033 4467 1047
rect 4473 1013 4487 1027
rect 4493 1013 4507 1027
rect 4413 953 4427 967
rect 4333 833 4347 847
rect 4373 833 4387 847
rect 4393 833 4407 847
rect 4473 873 4487 887
rect 4313 773 4327 787
rect 4333 753 4347 767
rect 4313 733 4327 747
rect 4553 993 4567 1007
rect 4513 973 4527 987
rect 4533 933 4547 947
rect 4533 893 4547 907
rect 4513 853 4527 867
rect 4473 833 4487 847
rect 4513 813 4527 827
rect 4393 793 4407 807
rect 4453 793 4467 807
rect 4653 1233 4667 1247
rect 4653 1193 4667 1207
rect 4753 1273 4767 1287
rect 4713 1233 4727 1247
rect 4753 1233 4767 1247
rect 4613 1133 4627 1147
rect 4633 1133 4647 1147
rect 4653 1133 4667 1147
rect 4653 1113 4667 1127
rect 4593 1093 4607 1107
rect 4613 1093 4627 1107
rect 4653 1053 4667 1067
rect 4633 1033 4647 1047
rect 4613 1013 4627 1027
rect 4573 913 4587 927
rect 4693 1173 4707 1187
rect 4753 1153 4767 1167
rect 4713 1133 4727 1147
rect 4733 1113 4747 1127
rect 4713 1093 4727 1107
rect 4673 873 4687 887
rect 4713 873 4727 887
rect 4593 853 4607 867
rect 4653 853 4667 867
rect 4573 833 4587 847
rect 4693 833 4707 847
rect 4613 813 4627 827
rect 4633 813 4647 827
rect 4593 793 4607 807
rect 4693 813 4707 827
rect 4673 773 4687 787
rect 4633 733 4647 747
rect 4353 713 4367 727
rect 4533 713 4547 727
rect 4413 673 4427 687
rect 4513 673 4527 687
rect 4553 673 4567 687
rect 4453 653 4467 667
rect 4493 653 4507 667
rect 4353 613 4367 627
rect 4433 613 4447 627
rect 4473 613 4487 627
rect 4393 573 4407 587
rect 4393 453 4407 467
rect 4333 393 4347 407
rect 4693 713 4707 727
rect 4653 693 4667 707
rect 4533 613 4547 627
rect 4633 613 4647 627
rect 4593 573 4607 587
rect 4693 553 4707 567
rect 4633 473 4647 487
rect 4673 473 4687 487
rect 4613 393 4627 407
rect 4393 373 4407 387
rect 4493 373 4507 387
rect 4333 353 4347 367
rect 4433 353 4447 367
rect 4513 353 4527 367
rect 4553 353 4567 367
rect 4913 1413 4927 1427
rect 4893 1393 4907 1407
rect 4873 1353 4887 1367
rect 4793 1273 4807 1287
rect 4813 1273 4827 1287
rect 4813 1253 4827 1267
rect 4833 1173 4847 1187
rect 4873 1313 4887 1327
rect 4893 1293 4907 1307
rect 4873 1273 4887 1287
rect 4873 1253 4887 1267
rect 4873 1173 4887 1187
rect 4853 1153 4867 1167
rect 4813 1133 4827 1147
rect 4993 1533 5007 1547
rect 4973 1473 4987 1487
rect 4973 1453 4987 1467
rect 5013 1453 5027 1467
rect 4993 1433 5007 1447
rect 5133 2633 5147 2647
rect 5133 2613 5147 2627
rect 5113 1933 5127 1947
rect 5093 1833 5107 1847
rect 5093 1753 5107 1767
rect 5093 1733 5107 1747
rect 5053 1713 5067 1727
rect 5073 1713 5087 1727
rect 5073 1613 5087 1627
rect 5073 1593 5087 1607
rect 5133 1773 5147 1787
rect 5133 1713 5147 1727
rect 5113 1653 5127 1667
rect 5093 1573 5107 1587
rect 5113 1573 5127 1587
rect 5053 1553 5067 1567
rect 5073 1533 5087 1547
rect 5113 1533 5127 1547
rect 5053 1513 5067 1527
rect 5053 1493 5067 1507
rect 4993 1413 5007 1427
rect 4973 1393 4987 1407
rect 4953 1373 4967 1387
rect 4933 1353 4947 1367
rect 4973 1353 4987 1367
rect 4953 1313 4967 1327
rect 4953 1273 4967 1287
rect 4933 1153 4947 1167
rect 4813 1113 4827 1127
rect 4833 1113 4847 1127
rect 4913 1113 4927 1127
rect 4793 933 4807 947
rect 4873 1093 4887 1107
rect 4853 1053 4867 1067
rect 4893 1073 4907 1087
rect 4913 913 4927 927
rect 4873 893 4887 907
rect 4813 873 4827 887
rect 4733 853 4747 867
rect 4773 853 4787 867
rect 4813 833 4827 847
rect 4853 833 4867 847
rect 4873 833 4887 847
rect 4793 793 4807 807
rect 4833 793 4847 807
rect 4753 693 4767 707
rect 4733 613 4747 627
rect 4773 633 4787 647
rect 4813 633 4827 647
rect 4793 593 4807 607
rect 4773 573 4787 587
rect 4713 393 4727 407
rect 4653 373 4667 387
rect 4693 373 4707 387
rect 4633 353 4647 367
rect 4673 353 4687 367
rect 4713 353 4727 367
rect 4373 333 4387 347
rect 4333 313 4347 327
rect 4313 293 4327 307
rect 4293 153 4307 167
rect 4593 333 4607 347
rect 4533 313 4547 327
rect 4533 293 4547 307
rect 4493 273 4507 287
rect 4413 193 4427 207
rect 4573 193 4587 207
rect 4293 133 4307 147
rect 4333 133 4347 147
rect 4473 173 4487 187
rect 4553 153 4567 167
rect 4433 133 4447 147
rect 4493 133 4507 147
rect 4753 333 4767 347
rect 4633 313 4647 327
rect 4673 313 4687 327
rect 4993 1293 5007 1307
rect 4973 1253 4987 1267
rect 4973 1193 4987 1207
rect 5033 1373 5047 1387
rect 5093 1433 5107 1447
rect 5073 1413 5087 1427
rect 5093 1353 5107 1367
rect 5133 1493 5147 1507
rect 5133 1413 5147 1427
rect 5033 1273 5047 1287
rect 5113 1333 5127 1347
rect 5053 1253 5067 1267
rect 5073 1253 5087 1267
rect 5113 1233 5127 1247
rect 5013 1193 5027 1207
rect 5033 1173 5047 1187
rect 4993 1133 5007 1147
rect 4953 1113 4967 1127
rect 4973 1093 4987 1107
rect 4953 1073 4967 1087
rect 5033 1073 5047 1087
rect 5093 1213 5107 1227
rect 5113 1213 5127 1227
rect 5073 1193 5087 1207
rect 4993 1013 5007 1027
rect 5053 1013 5067 1027
rect 4953 873 4967 887
rect 4913 813 4927 827
rect 4933 813 4947 827
rect 4853 653 4867 667
rect 4893 653 4907 667
rect 4933 653 4947 667
rect 4853 633 4867 647
rect 4933 633 4947 647
rect 4913 613 4927 627
rect 5053 973 5067 987
rect 5033 913 5047 927
rect 4973 813 4987 827
rect 5013 793 5027 807
rect 5053 793 5067 807
rect 5013 753 5027 767
rect 4973 673 4987 687
rect 4973 613 4987 627
rect 4873 593 4887 607
rect 4953 593 4967 607
rect 4993 553 5007 567
rect 4773 273 4787 287
rect 4773 233 4787 247
rect 4733 193 4747 207
rect 4593 173 4607 187
rect 4673 153 4687 167
rect 4733 153 4747 167
rect 4833 393 4847 407
rect 4973 393 4987 407
rect 4813 373 4827 387
rect 4833 353 4847 367
rect 4793 153 4807 167
rect 4853 333 4867 347
rect 4873 293 4887 307
rect 4873 273 4887 287
rect 4853 193 4867 207
rect 4753 133 4767 147
rect 4793 133 4807 147
rect 4833 133 4847 147
rect 4953 373 4967 387
rect 4933 353 4947 367
rect 5093 1093 5107 1107
rect 5113 1053 5127 1067
rect 5133 973 5147 987
rect 5113 933 5127 947
rect 5093 893 5107 907
rect 5073 373 5087 387
rect 4913 333 4927 347
rect 4893 193 4907 207
rect 4913 153 4927 167
rect 4933 153 4947 167
rect 5013 353 5027 367
rect 5033 353 5047 367
rect 5053 333 5067 347
rect 5093 353 5107 367
rect 5013 313 5027 327
rect 5073 313 5087 327
rect 4993 293 5007 307
rect 4893 133 4907 147
rect 4953 133 4967 147
rect 4133 113 4147 127
rect 4193 113 4207 127
rect 3933 93 3947 107
rect 4093 93 4107 107
rect 4413 113 4427 127
rect 4573 113 4587 127
rect 4613 113 4627 127
rect 4693 113 4707 127
rect 4093 73 4107 87
rect 4653 73 4667 87
rect 2713 33 2727 47
rect 2673 13 2687 27
rect 2873 13 2887 27
rect 5033 13 5047 27
rect 5113 13 5127 27
<< metal3 >>
rect 1927 4816 2433 4824
rect 2987 4816 3173 4824
rect 4687 4816 4793 4824
rect 707 4756 773 4764
rect 787 4756 2473 4764
rect 1607 4736 2393 4744
rect 227 4716 733 4724
rect 747 4716 993 4724
rect 1007 4716 1453 4724
rect 1467 4716 1853 4724
rect 1867 4716 1993 4724
rect 2067 4716 2193 4724
rect 2307 4716 2713 4724
rect 3327 4716 3373 4724
rect 3387 4716 3873 4724
rect 3887 4716 4013 4724
rect 1127 4696 1253 4704
rect 1327 4696 1753 4704
rect 2036 4696 2233 4704
rect 187 4676 273 4684
rect 327 4676 353 4684
rect 367 4676 493 4684
rect 547 4676 573 4684
rect 667 4676 733 4684
rect 767 4676 953 4684
rect 107 4656 173 4664
rect 407 4656 473 4664
rect 496 4664 504 4673
rect 836 4667 844 4676
rect 1347 4676 1433 4684
rect 1476 4676 1533 4684
rect 496 4656 553 4664
rect 576 4656 633 4664
rect 47 4636 193 4644
rect 576 4644 584 4656
rect 656 4656 673 4664
rect 247 4636 584 4644
rect 656 4644 664 4656
rect 907 4656 973 4664
rect 1027 4656 1073 4664
rect 1196 4664 1204 4673
rect 1476 4667 1484 4676
rect 1667 4676 1864 4684
rect 1736 4667 1744 4676
rect 1087 4656 1233 4664
rect 1307 4656 1353 4664
rect 1367 4656 1453 4664
rect 1496 4656 1633 4664
rect 627 4636 664 4644
rect 687 4636 713 4644
rect 727 4636 1013 4644
rect 1227 4636 1273 4644
rect 1496 4644 1504 4656
rect 1787 4656 1833 4664
rect 1856 4664 1864 4676
rect 1856 4656 1873 4664
rect 2036 4647 2044 4696
rect 2287 4696 2313 4704
rect 2456 4696 2553 4704
rect 2187 4676 2253 4684
rect 2347 4676 2433 4684
rect 2096 4664 2104 4673
rect 2096 4656 2113 4664
rect 1427 4636 1504 4644
rect 1567 4636 1713 4644
rect 1767 4636 1953 4644
rect 2136 4644 2144 4673
rect 2456 4667 2464 4696
rect 2687 4696 3493 4704
rect 3507 4696 3593 4704
rect 3607 4696 3633 4704
rect 2487 4676 2513 4684
rect 2607 4676 2653 4684
rect 2707 4676 2853 4684
rect 3207 4676 3233 4684
rect 3307 4676 3433 4684
rect 3447 4676 3533 4684
rect 3827 4676 4573 4684
rect 4596 4676 4653 4684
rect 2167 4656 2193 4664
rect 2247 4656 2333 4664
rect 2507 4656 2833 4664
rect 2967 4656 3073 4664
rect 3087 4656 3193 4664
rect 3487 4656 3573 4664
rect 3727 4656 4033 4664
rect 2087 4636 2144 4644
rect 2347 4636 2373 4644
rect 2496 4644 2504 4653
rect 3876 4647 3884 4656
rect 4047 4656 4153 4664
rect 4167 4656 4173 4664
rect 4596 4664 4604 4676
rect 4467 4656 4604 4664
rect 5056 4664 5064 4713
rect 5147 4676 5184 4684
rect 5047 4656 5064 4664
rect 2387 4636 2504 4644
rect 2627 4636 2753 4644
rect 2847 4636 2873 4644
rect 3467 4636 3753 4644
rect 3927 4636 4593 4644
rect 607 4616 773 4624
rect 1127 4616 1133 4624
rect 1147 4616 1173 4624
rect 1307 4616 1493 4624
rect 1507 4616 1613 4624
rect 1987 4616 1993 4624
rect 2007 4616 2173 4624
rect 2287 4616 2533 4624
rect 2787 4616 2813 4624
rect 2827 4616 3413 4624
rect 3527 4616 5113 4624
rect 547 4596 613 4604
rect 767 4596 793 4604
rect 1047 4596 1473 4604
rect 1927 4596 2093 4604
rect 2387 4596 2493 4604
rect 2527 4596 2613 4604
rect 2627 4596 3773 4604
rect 4187 4596 4733 4604
rect 147 4576 333 4584
rect 347 4576 453 4584
rect 467 4576 2573 4584
rect 2847 4576 5133 4584
rect 947 4556 993 4564
rect 1507 4556 1813 4564
rect 1827 4556 1933 4564
rect 1947 4556 2073 4564
rect 2087 4556 2913 4564
rect 4147 4556 5184 4564
rect 147 4536 373 4544
rect 387 4536 593 4544
rect 607 4536 793 4544
rect 987 4536 1093 4544
rect 1127 4536 1253 4544
rect 1267 4536 1393 4544
rect 1407 4536 1993 4544
rect 2027 4536 2273 4544
rect 4487 4536 5053 4544
rect 5067 4536 5073 4544
rect 5176 4536 5184 4556
rect 207 4516 573 4524
rect 687 4516 733 4524
rect 747 4516 773 4524
rect 787 4516 1153 4524
rect 1187 4516 1373 4524
rect 1847 4516 2113 4524
rect 2367 4516 2713 4524
rect 3247 4516 3373 4524
rect 67 4496 113 4504
rect 527 4496 833 4504
rect 847 4496 953 4504
rect 967 4496 1233 4504
rect 1247 4496 1313 4504
rect 1347 4496 1513 4504
rect 1527 4496 1584 4504
rect 107 4476 153 4484
rect 507 4476 613 4484
rect 667 4476 713 4484
rect 727 4476 753 4484
rect 787 4476 824 4484
rect 76 4447 84 4473
rect 816 4467 824 4476
rect 987 4476 1024 4484
rect 247 4456 273 4464
rect 487 4456 533 4464
rect 647 4456 813 4464
rect 127 4436 213 4444
rect 267 4436 313 4444
rect 336 4444 344 4453
rect 336 4436 413 4444
rect 436 4427 444 4453
rect 856 4447 864 4473
rect 1016 4467 1024 4476
rect 1167 4476 1193 4484
rect 1207 4476 1273 4484
rect 1296 4476 1333 4484
rect 887 4456 913 4464
rect 1076 4464 1084 4473
rect 1076 4456 1173 4464
rect 1296 4464 1304 4476
rect 1427 4476 1553 4484
rect 1576 4484 1584 4496
rect 1607 4496 1633 4504
rect 1707 4496 1753 4504
rect 2147 4496 2313 4504
rect 2396 4496 2493 4504
rect 1576 4476 1893 4484
rect 1947 4476 2013 4484
rect 2087 4476 2213 4484
rect 2296 4476 2353 4484
rect 2296 4467 2304 4476
rect 2396 4467 2404 4496
rect 2507 4496 2553 4504
rect 2887 4496 3013 4504
rect 3236 4496 3513 4504
rect 3236 4484 3244 4496
rect 2547 4476 3244 4484
rect 3256 4476 3333 4484
rect 1187 4456 1304 4464
rect 1387 4456 1433 4464
rect 1447 4456 1564 4464
rect 587 4436 733 4444
rect 907 4436 933 4444
rect 976 4444 984 4453
rect 976 4436 1153 4444
rect 1227 4436 1253 4444
rect 1267 4436 1313 4444
rect 1367 4436 1473 4444
rect 1556 4444 1564 4456
rect 1587 4456 1713 4464
rect 1747 4456 1793 4464
rect 1807 4456 1873 4464
rect 1927 4456 1973 4464
rect 2107 4456 2124 4464
rect 1556 4436 1713 4444
rect 2007 4436 2093 4444
rect 47 4416 53 4424
rect 67 4416 93 4424
rect 767 4416 1553 4424
rect 1667 4416 1773 4424
rect 1827 4416 1913 4424
rect 2116 4424 2124 4456
rect 2187 4456 2253 4464
rect 2316 4456 2353 4464
rect 2316 4447 2324 4456
rect 2147 4436 2193 4444
rect 2227 4436 2293 4444
rect 2416 4444 2424 4473
rect 2607 4456 2633 4464
rect 2807 4456 3093 4464
rect 3256 4464 3264 4476
rect 3627 4476 3833 4484
rect 4356 4467 4364 4513
rect 4716 4496 4813 4504
rect 4616 4476 4693 4484
rect 3107 4456 3264 4464
rect 3307 4456 3353 4464
rect 3407 4456 3453 4464
rect 3647 4456 3713 4464
rect 4187 4456 4213 4464
rect 4387 4456 4593 4464
rect 2416 4436 2433 4444
rect 2687 4436 2733 4444
rect 2867 4436 3053 4444
rect 3207 4436 3253 4444
rect 3487 4436 3593 4444
rect 3607 4436 3693 4444
rect 3747 4436 3953 4444
rect 4036 4427 4044 4453
rect 4616 4447 4624 4476
rect 4716 4467 4724 4496
rect 4847 4496 4933 4504
rect 4947 4496 4973 4504
rect 5127 4496 5184 4504
rect 4927 4476 5013 4484
rect 4736 4447 4744 4473
rect 4827 4456 4893 4464
rect 4947 4456 5113 4464
rect 4747 4436 4853 4444
rect 4927 4436 4953 4444
rect 2087 4416 2453 4424
rect 2667 4416 3113 4424
rect 3127 4416 3433 4424
rect 4647 4416 4793 4424
rect 427 4396 913 4404
rect 1407 4396 1533 4404
rect 1647 4396 1673 4404
rect 1767 4396 2053 4404
rect 2176 4396 2313 4404
rect 187 4376 553 4384
rect 567 4376 1413 4384
rect 1467 4376 1833 4384
rect 1847 4376 1953 4384
rect 2176 4384 2184 4396
rect 2907 4396 3173 4404
rect 3407 4396 3493 4404
rect 4487 4396 4773 4404
rect 1967 4376 2184 4384
rect 2207 4376 2553 4384
rect 2947 4376 3953 4384
rect 4067 4376 4273 4384
rect 1147 4356 1753 4364
rect 1807 4356 2033 4364
rect 2516 4356 2833 4364
rect 887 4336 1053 4344
rect 2516 4344 2524 4356
rect 4376 4356 4813 4364
rect 1067 4336 2524 4344
rect 4376 4344 4384 4356
rect 2927 4336 4384 4344
rect 4407 4336 4873 4344
rect 2167 4316 2653 4324
rect 2727 4316 3733 4324
rect 3747 4316 4233 4324
rect 4567 4316 4913 4324
rect 1587 4296 1613 4304
rect 1987 4296 2093 4304
rect 2107 4296 2253 4304
rect 2267 4296 2513 4304
rect 2687 4296 4133 4304
rect 4527 4296 4573 4304
rect 4787 4296 4993 4304
rect 1147 4276 2413 4284
rect 2447 4276 3453 4284
rect 3727 4276 4953 4284
rect 267 4256 393 4264
rect 567 4256 933 4264
rect 947 4256 1353 4264
rect 1387 4256 1533 4264
rect 1547 4256 1793 4264
rect 1867 4256 2753 4264
rect 3067 4256 3253 4264
rect 4587 4256 4653 4264
rect 4687 4256 4833 4264
rect 287 4236 713 4244
rect 827 4236 953 4244
rect 1167 4236 1213 4244
rect 1427 4236 1493 4244
rect 1527 4236 1613 4244
rect 1627 4236 1653 4244
rect 1707 4236 1833 4244
rect 1947 4236 2173 4244
rect 2427 4236 2773 4244
rect 2787 4236 3113 4244
rect 3427 4236 3593 4244
rect 4007 4236 4613 4244
rect 4767 4236 4804 4244
rect 87 4216 113 4224
rect 127 4216 133 4224
rect 267 4216 284 4224
rect 276 4207 284 4216
rect 307 4216 373 4224
rect 387 4216 613 4224
rect 907 4216 1033 4224
rect 1156 4216 1453 4224
rect 1156 4207 1164 4216
rect 1547 4216 1584 4224
rect 36 4196 53 4204
rect 36 4187 44 4196
rect 307 4196 413 4204
rect 427 4196 444 4204
rect 47 4176 93 4184
rect 207 4176 313 4184
rect 436 4184 444 4196
rect 467 4196 504 4204
rect 436 4176 484 4184
rect 476 4167 484 4176
rect 87 4156 113 4164
rect 496 4144 504 4196
rect 547 4196 573 4204
rect 687 4196 773 4204
rect 927 4196 993 4204
rect 1207 4196 1313 4204
rect 1347 4196 1413 4204
rect 627 4176 653 4184
rect 776 4184 784 4193
rect 776 4176 833 4184
rect 876 4184 884 4193
rect 876 4176 933 4184
rect 1096 4184 1104 4193
rect 1576 4187 1584 4216
rect 1627 4216 1853 4224
rect 1907 4216 2073 4224
rect 2187 4216 2313 4224
rect 2427 4216 2473 4224
rect 2527 4216 2613 4224
rect 2627 4216 2853 4224
rect 3087 4216 3153 4224
rect 3167 4216 3353 4224
rect 3567 4216 3673 4224
rect 3687 4216 3693 4224
rect 3787 4216 4293 4224
rect 4427 4216 4453 4224
rect 4536 4216 4773 4224
rect 1607 4196 1653 4204
rect 2067 4196 2113 4204
rect 2127 4196 2204 4204
rect 1096 4176 1153 4184
rect 1176 4176 1333 4184
rect 607 4156 633 4164
rect 647 4156 753 4164
rect 887 4156 913 4164
rect 1176 4164 1184 4176
rect 1756 4184 1764 4193
rect 1627 4176 1724 4184
rect 1756 4176 1913 4184
rect 927 4156 1184 4164
rect 1227 4156 1233 4164
rect 1247 4156 1293 4164
rect 1327 4156 1473 4164
rect 1547 4156 1693 4164
rect 1716 4164 1724 4176
rect 2007 4176 2033 4184
rect 2196 4184 2204 4196
rect 2507 4196 2573 4204
rect 3047 4196 3133 4204
rect 3587 4196 3633 4204
rect 2196 4176 2273 4184
rect 2647 4176 2813 4184
rect 2907 4176 3053 4184
rect 3127 4176 3213 4184
rect 3227 4176 3413 4184
rect 3487 4176 3533 4184
rect 3736 4184 3744 4213
rect 4536 4207 4544 4216
rect 3767 4196 3813 4204
rect 3876 4196 3953 4204
rect 3856 4184 3864 4193
rect 3876 4187 3884 4196
rect 4356 4196 4393 4204
rect 3736 4176 3864 4184
rect 1716 4156 1753 4164
rect 1767 4156 2173 4164
rect 2207 4156 2293 4164
rect 2347 4156 2673 4164
rect 2867 4156 2953 4164
rect 3347 4156 3653 4164
rect 3856 4164 3864 4176
rect 3996 4184 4004 4193
rect 4356 4187 4364 4196
rect 4487 4196 4513 4204
rect 4587 4196 4664 4204
rect 3947 4176 4004 4184
rect 4027 4176 4153 4184
rect 4287 4176 4313 4184
rect 4507 4176 4553 4184
rect 4656 4167 4664 4196
rect 3856 4156 4173 4164
rect 4407 4156 4453 4164
rect 4547 4156 4573 4164
rect 247 4136 504 4144
rect 707 4136 733 4144
rect 747 4136 1073 4144
rect 1127 4136 1173 4144
rect 1287 4136 1353 4144
rect 1567 4136 1673 4144
rect 1727 4136 1773 4144
rect 1847 4136 1993 4144
rect 2147 4136 2553 4144
rect 2567 4136 2693 4144
rect 4067 4136 4093 4144
rect 4696 4144 4704 4193
rect 4796 4164 4804 4236
rect 4847 4236 5133 4244
rect 4856 4204 4864 4213
rect 4816 4196 4864 4204
rect 4816 4187 4824 4196
rect 4896 4196 4953 4204
rect 4796 4156 4813 4164
rect 4876 4164 4884 4193
rect 4896 4187 4904 4196
rect 4987 4196 5013 4204
rect 5056 4167 5064 4193
rect 4847 4156 4884 4164
rect 5087 4156 5113 4164
rect 4187 4136 4933 4144
rect 987 4116 1013 4124
rect 1167 4116 1393 4124
rect 1427 4116 1433 4124
rect 1447 4116 1593 4124
rect 1607 4116 1733 4124
rect 1747 4116 2353 4124
rect 2747 4116 3593 4124
rect 3867 4116 3913 4124
rect 4467 4116 4513 4124
rect 4567 4116 4773 4124
rect 427 4096 1613 4104
rect 1647 4096 2153 4104
rect 2187 4096 2873 4104
rect 3387 4096 3433 4104
rect 3467 4096 3753 4104
rect 3767 4096 4313 4104
rect 4387 4096 4673 4104
rect 4727 4096 4833 4104
rect 1147 4076 1313 4084
rect 1347 4076 2413 4084
rect 2507 4076 3113 4084
rect 3447 4076 3893 4084
rect 3907 4076 4153 4084
rect 4387 4076 4413 4084
rect 4647 4076 4664 4084
rect 647 4056 713 4064
rect 727 4056 773 4064
rect 1407 4056 1673 4064
rect 1707 4056 1833 4064
rect 2027 4056 2153 4064
rect 2167 4056 2213 4064
rect 2447 4056 2713 4064
rect 2727 4056 2953 4064
rect 3847 4056 3913 4064
rect 4247 4056 4473 4064
rect 4607 4056 4633 4064
rect 4656 4064 4664 4076
rect 4687 4076 5133 4084
rect 4656 4056 4733 4064
rect 107 4036 433 4044
rect 447 4036 593 4044
rect 607 4036 1733 4044
rect 1927 4036 2193 4044
rect 2667 4036 2973 4044
rect 2987 4036 3173 4044
rect 3307 4036 3673 4044
rect 3707 4036 3893 4044
rect 4147 4036 4353 4044
rect 4427 4036 4493 4044
rect 4667 4036 4733 4044
rect 4887 4036 4913 4044
rect 5047 4036 5133 4044
rect 207 4016 273 4024
rect 367 4016 453 4024
rect 687 4016 753 4024
rect 1227 4016 1253 4024
rect 1467 4016 1713 4024
rect 1727 4016 1973 4024
rect 2087 4016 2133 4024
rect 2207 4016 2293 4024
rect 2327 4016 2373 4024
rect 3107 4016 3153 4024
rect 3527 4016 3573 4024
rect 3687 4016 3693 4024
rect 3707 4016 3953 4024
rect 4276 4016 4353 4024
rect 87 3996 133 4004
rect 267 3996 333 4004
rect 347 3996 433 4004
rect 487 3996 553 4004
rect 907 3996 933 4004
rect 67 3976 153 3984
rect 216 3984 224 3993
rect 1136 3987 1144 4013
rect 1156 3996 1353 4004
rect 187 3976 224 3984
rect 387 3976 593 3984
rect 687 3976 713 3984
rect 167 3956 233 3964
rect 407 3956 453 3964
rect 587 3956 653 3964
rect 747 3956 1093 3964
rect 1156 3964 1164 3996
rect 1376 3996 1453 4004
rect 1376 3987 1384 3996
rect 1507 3996 1553 4004
rect 1656 3996 1773 4004
rect 1267 3976 1333 3984
rect 1576 3984 1584 3993
rect 1656 3987 1664 3996
rect 1847 3996 1893 4004
rect 1947 3996 2033 4004
rect 2047 3996 2493 4004
rect 2647 3996 2853 4004
rect 2907 3996 3093 4004
rect 3116 3996 3153 4004
rect 1487 3976 1644 3984
rect 1636 3967 1644 3976
rect 1907 3976 1953 3984
rect 1127 3956 1164 3964
rect 1287 3956 1313 3964
rect 1327 3956 1393 3964
rect 1547 3956 1613 3964
rect 1767 3956 1793 3964
rect 1827 3956 1873 3964
rect 707 3936 753 3944
rect 767 3936 913 3944
rect 1087 3936 1233 3944
rect 1447 3936 1753 3944
rect 1936 3944 1944 3976
rect 2127 3976 2173 3984
rect 2247 3976 2353 3984
rect 2407 3976 2453 3984
rect 2487 3976 2733 3984
rect 3027 3976 3093 3984
rect 1967 3956 2673 3964
rect 3116 3964 3124 3996
rect 3176 3996 3253 4004
rect 3176 3984 3184 3996
rect 3307 3996 3493 4004
rect 3547 3996 3733 4004
rect 3147 3976 3184 3984
rect 3467 3976 3513 3984
rect 3907 3976 3933 3984
rect 3947 3976 4093 3984
rect 4207 3976 4253 3984
rect 4276 3967 4284 4016
rect 4367 4016 4413 4024
rect 4447 4016 4593 4024
rect 4647 4016 4813 4024
rect 4867 4016 4924 4024
rect 4387 3996 4404 4004
rect 4336 3984 4344 3993
rect 4336 3976 4353 3984
rect 3116 3956 3193 3964
rect 3387 3956 3413 3964
rect 3447 3956 3553 3964
rect 4087 3956 4233 3964
rect 4396 3964 4404 3996
rect 4416 3996 4453 4004
rect 4416 3987 4424 3996
rect 4547 3996 4684 4004
rect 4447 3976 4513 3984
rect 4676 3984 4684 3996
rect 4707 3996 4773 4004
rect 4787 3996 4853 4004
rect 4867 3996 4893 4004
rect 4676 3976 4713 3984
rect 4916 3984 4924 4016
rect 4947 4016 4993 4024
rect 5027 4016 5093 4024
rect 5036 3996 5053 4004
rect 4847 3976 4924 3984
rect 4987 3976 5013 3984
rect 4396 3956 4453 3964
rect 4607 3956 4653 3964
rect 4956 3964 4964 3973
rect 5036 3964 5044 3996
rect 4947 3956 4964 3964
rect 5016 3956 5044 3964
rect 1936 3936 1973 3944
rect 2027 3936 2133 3944
rect 2227 3936 2293 3944
rect 2347 3936 2753 3944
rect 3127 3936 3213 3944
rect 3567 3936 3713 3944
rect 4287 3936 4393 3944
rect 4427 3936 4913 3944
rect 147 3916 733 3924
rect 767 3916 1124 3924
rect 547 3896 1093 3904
rect 1116 3904 1124 3916
rect 1247 3916 1513 3924
rect 1587 3916 1653 3924
rect 1676 3916 1944 3924
rect 1676 3904 1684 3916
rect 1116 3896 1684 3904
rect 1727 3896 1913 3904
rect 1936 3904 1944 3916
rect 2167 3916 2173 3924
rect 2187 3916 2413 3924
rect 2467 3916 2713 3924
rect 2787 3916 2993 3924
rect 3007 3916 3273 3924
rect 3507 3916 3713 3924
rect 4747 3916 4993 3924
rect 5016 3924 5024 3956
rect 5047 3936 5073 3944
rect 5016 3916 5033 3924
rect 5056 3916 5133 3924
rect 1936 3896 3513 3904
rect 4047 3896 4293 3904
rect 4307 3896 4393 3904
rect 5056 3904 5064 3916
rect 5007 3896 5064 3904
rect 5087 3896 5133 3904
rect 127 3876 1113 3884
rect 1147 3876 1253 3884
rect 1287 3876 1713 3884
rect 1747 3876 2373 3884
rect 2727 3876 2813 3884
rect 2827 3876 3033 3884
rect 3047 3876 3433 3884
rect 3807 3876 3873 3884
rect 3907 3876 3973 3884
rect 3987 3876 4493 3884
rect 4887 3876 4953 3884
rect 807 3856 1233 3864
rect 1527 3856 2053 3864
rect 2327 3856 3473 3864
rect 3667 3856 4873 3864
rect 607 3836 713 3844
rect 1047 3836 1273 3844
rect 1567 3836 1693 3844
rect 1767 3836 1833 3844
rect 1867 3836 1893 3844
rect 2047 3836 3033 3844
rect 3307 3836 3353 3844
rect 4527 3836 5073 3844
rect 27 3816 753 3824
rect 947 3816 1133 3824
rect 1207 3816 2073 3824
rect 2367 3816 2533 3824
rect 2547 3816 3653 3824
rect 3727 3816 4193 3824
rect 4207 3816 4253 3824
rect -24 3796 33 3804
rect 547 3796 593 3804
rect 727 3796 1293 3804
rect 1307 3796 2493 3804
rect 4667 3796 4913 3804
rect 327 3776 413 3784
rect 1027 3776 1033 3784
rect 1047 3776 1113 3784
rect 1147 3776 1313 3784
rect 1487 3776 1513 3784
rect 1627 3776 1773 3784
rect 1787 3776 1953 3784
rect 1987 3776 2313 3784
rect 2487 3776 2913 3784
rect 4056 3784 4064 3793
rect 4056 3776 4133 3784
rect 4587 3776 4613 3784
rect 4687 3776 4753 3784
rect -24 3756 53 3764
rect 407 3756 444 3764
rect 436 3744 444 3756
rect 527 3756 613 3764
rect 847 3756 1213 3764
rect 1287 3756 3393 3764
rect 3827 3756 4053 3764
rect 4167 3756 4313 3764
rect 4347 3756 4404 3764
rect 4396 3747 4404 3756
rect 4656 3756 4793 3764
rect 367 3736 424 3744
rect 436 3736 833 3744
rect -24 3716 13 3724
rect 36 3707 44 3733
rect 187 3716 233 3724
rect 416 3724 424 3736
rect 867 3736 993 3744
rect 1107 3736 1204 3744
rect 416 3716 444 3724
rect 147 3696 213 3704
rect 236 3704 244 3713
rect 236 3696 333 3704
rect 396 3704 404 3713
rect 396 3696 413 3704
rect 436 3704 444 3716
rect 487 3716 533 3724
rect 567 3716 584 3724
rect 436 3696 453 3704
rect 576 3704 584 3716
rect 607 3716 733 3724
rect 787 3716 813 3724
rect 576 3696 644 3704
rect 167 3676 273 3684
rect 327 3676 373 3684
rect 547 3676 613 3684
rect 636 3684 644 3696
rect 836 3704 844 3733
rect 1196 3727 1204 3736
rect 1447 3736 1533 3744
rect 1727 3736 1793 3744
rect 1807 3736 2033 3744
rect 2087 3736 2124 3744
rect 907 3716 933 3724
rect 1127 3716 1144 3724
rect 807 3696 844 3704
rect 887 3696 953 3704
rect 996 3704 1004 3713
rect 996 3696 1053 3704
rect 636 3676 864 3684
rect 207 3656 593 3664
rect 607 3656 833 3664
rect 856 3664 864 3676
rect 947 3676 1013 3684
rect 1076 3684 1084 3713
rect 1136 3707 1144 3716
rect 1287 3716 1304 3724
rect 1076 3676 1133 3684
rect 856 3656 933 3664
rect 947 3656 973 3664
rect 1156 3664 1164 3713
rect 1296 3707 1304 3716
rect 1467 3716 1513 3724
rect 1596 3707 1604 3733
rect 1207 3696 1273 3704
rect 1327 3696 1533 3704
rect 1636 3704 1644 3733
rect 1887 3716 1913 3724
rect 1927 3716 2044 3724
rect 1636 3696 1753 3704
rect 1836 3704 1844 3713
rect 2036 3707 2044 3716
rect 2056 3716 2093 3724
rect 1836 3696 1933 3704
rect 1247 3676 1333 3684
rect 1356 3676 1493 3684
rect 1107 3656 1173 3664
rect 1356 3664 1364 3676
rect 2056 3684 2064 3716
rect 2116 3704 2124 3736
rect 2167 3736 2353 3744
rect 2427 3736 2633 3744
rect 2747 3736 2764 3744
rect 2256 3716 2473 3724
rect 2087 3696 2124 3704
rect 2256 3704 2264 3716
rect 2527 3716 2544 3724
rect 2147 3696 2264 3704
rect 2287 3696 2333 3704
rect 2496 3704 2504 3713
rect 2536 3704 2544 3716
rect 2627 3716 2644 3724
rect 2496 3696 2524 3704
rect 2536 3696 2553 3704
rect 1567 3676 2213 3684
rect 2436 3676 2493 3684
rect 1196 3656 1364 3664
rect 807 3636 813 3644
rect 827 3636 853 3644
rect 887 3636 913 3644
rect 1007 3636 1073 3644
rect 1196 3644 1204 3656
rect 1407 3656 1613 3664
rect 1647 3656 1693 3664
rect 1787 3656 1833 3664
rect 1887 3656 2333 3664
rect 2436 3664 2444 3676
rect 2516 3684 2524 3696
rect 2576 3704 2584 3713
rect 2576 3696 2613 3704
rect 2636 3704 2644 3716
rect 2707 3716 2733 3724
rect 2636 3696 2673 3704
rect 2756 3704 2764 3736
rect 2907 3736 2973 3744
rect 3047 3736 3213 3744
rect 4227 3736 4353 3744
rect 4416 3736 4473 3744
rect 2947 3716 3013 3724
rect 3587 3716 3913 3724
rect 2756 3696 2833 3704
rect 2847 3696 2873 3704
rect 2927 3696 3133 3704
rect 3227 3696 3253 3704
rect 3547 3696 3573 3704
rect 3767 3696 3793 3704
rect 3936 3704 3944 3733
rect 4416 3727 4424 3736
rect 4656 3744 4664 3756
rect 4916 3756 4973 3764
rect 4556 3736 4664 3744
rect 3967 3716 4044 3724
rect 4036 3707 4044 3716
rect 4087 3716 4113 3724
rect 4167 3716 4293 3724
rect 4327 3716 4373 3724
rect 4436 3716 4453 3724
rect 4436 3707 4444 3716
rect 3927 3696 3944 3704
rect 4047 3696 4153 3704
rect 4187 3696 4324 3704
rect 2516 3676 2773 3684
rect 2867 3676 2933 3684
rect 3187 3676 3293 3684
rect 3467 3676 3713 3684
rect 3787 3676 3833 3684
rect 3887 3676 3973 3684
rect 4007 3676 4073 3684
rect 4087 3676 4193 3684
rect 4316 3684 4324 3696
rect 4347 3696 4433 3704
rect 4536 3684 4544 3713
rect 4316 3676 4544 3684
rect 4556 3667 4564 3736
rect 4687 3736 4753 3744
rect 4916 3744 4924 3756
rect 4807 3736 4924 3744
rect 5007 3736 5024 3744
rect 4587 3716 4733 3724
rect 4787 3716 4873 3724
rect 4607 3696 4673 3704
rect 4896 3704 4904 3713
rect 4747 3696 4904 3704
rect 4936 3704 4944 3733
rect 4936 3696 4993 3704
rect 4587 3676 4613 3684
rect 5016 3684 5024 3736
rect 4667 3676 5024 3684
rect 2347 3656 2444 3664
rect 2467 3656 2493 3664
rect 2627 3656 2913 3664
rect 2927 3656 4013 3664
rect 4067 3656 4273 3664
rect 4287 3656 4473 3664
rect 4647 3656 4753 3664
rect 4827 3656 4933 3664
rect 1127 3636 1204 3644
rect 1327 3636 2653 3644
rect 2707 3636 2793 3644
rect 2987 3636 3133 3644
rect 3147 3636 3353 3644
rect 3407 3636 3533 3644
rect 3787 3636 3933 3644
rect 4087 3636 4153 3644
rect 4367 3636 4453 3644
rect 4627 3636 5113 3644
rect 87 3616 1873 3624
rect 2127 3616 2393 3624
rect 2467 3616 2533 3624
rect 2607 3616 2633 3624
rect 2667 3616 2753 3624
rect 3527 3616 3753 3624
rect 3807 3616 3853 3624
rect 3947 3616 4133 3624
rect 4527 3616 4813 3624
rect 4827 3616 4833 3624
rect 587 3596 1413 3604
rect 1547 3596 2413 3604
rect 2487 3596 2593 3604
rect 2627 3596 2673 3604
rect 2867 3596 4093 3604
rect 4107 3596 4233 3604
rect 4247 3596 4633 3604
rect 667 3576 1013 3584
rect 1027 3576 1373 3584
rect 1387 3576 1513 3584
rect 1587 3576 1853 3584
rect 2107 3576 2233 3584
rect 2267 3576 3513 3584
rect 3847 3576 3904 3584
rect 267 3556 293 3564
rect 307 3556 393 3564
rect 407 3556 493 3564
rect 1047 3556 1064 3564
rect 167 3536 193 3544
rect 207 3536 333 3544
rect 556 3536 573 3544
rect 447 3516 533 3524
rect 307 3496 333 3504
rect 356 3484 364 3513
rect 556 3507 564 3536
rect 587 3536 664 3544
rect 587 3516 613 3524
rect 387 3496 413 3504
rect 436 3496 453 3504
rect 356 3476 373 3484
rect 436 3484 444 3496
rect 476 3496 513 3504
rect 476 3487 484 3496
rect 407 3476 444 3484
rect 616 3484 624 3493
rect 507 3476 624 3484
rect 636 3484 644 3513
rect 656 3507 664 3536
rect 687 3536 873 3544
rect 907 3536 1004 3544
rect 836 3516 953 3524
rect 767 3496 813 3504
rect 636 3476 693 3484
rect 716 3484 724 3493
rect 716 3476 753 3484
rect 836 3484 844 3516
rect 996 3507 1004 3536
rect 1016 3507 1024 3533
rect 887 3496 893 3504
rect 907 3496 973 3504
rect 807 3476 844 3484
rect 1036 3484 1044 3533
rect 1056 3504 1064 3556
rect 1367 3556 1393 3564
rect 1447 3556 1553 3564
rect 1627 3556 1673 3564
rect 1887 3556 2013 3564
rect 2087 3556 2133 3564
rect 2167 3556 2333 3564
rect 2547 3556 2713 3564
rect 2847 3556 3073 3564
rect 3207 3556 3433 3564
rect 3447 3556 3473 3564
rect 3487 3556 3673 3564
rect 3687 3556 3873 3564
rect 1087 3536 1333 3544
rect 1367 3536 1424 3544
rect 1116 3516 1153 3524
rect 1116 3507 1124 3516
rect 1176 3516 1253 3524
rect 1056 3496 1093 3504
rect 1176 3504 1184 3516
rect 1147 3496 1184 3504
rect 947 3476 1044 3484
rect 1416 3484 1424 3536
rect 1487 3536 1544 3544
rect 1436 3507 1444 3533
rect 1536 3507 1544 3536
rect 1607 3536 1973 3544
rect 2047 3536 2173 3544
rect 2207 3536 2273 3544
rect 2287 3536 2313 3544
rect 2447 3536 2513 3544
rect 2607 3536 2653 3544
rect 2687 3536 2873 3544
rect 2967 3536 2993 3544
rect 3367 3536 3493 3544
rect 3767 3536 3844 3544
rect 1556 3516 1613 3524
rect 1556 3487 1564 3516
rect 1667 3516 1713 3524
rect 1767 3516 1793 3524
rect 1927 3516 1944 3524
rect 1416 3476 1473 3484
rect 1607 3476 1793 3484
rect 1807 3476 1813 3484
rect 287 3456 473 3464
rect 787 3456 1193 3464
rect 1547 3456 1633 3464
rect 1687 3456 1693 3464
rect 1707 3456 1733 3464
rect 1856 3464 1864 3513
rect 1936 3504 1944 3516
rect 1967 3516 1984 3524
rect 1976 3504 1984 3516
rect 2067 3516 2133 3524
rect 2436 3516 2453 3524
rect 2156 3504 2164 3513
rect 1936 3496 1964 3504
rect 1976 3496 2164 3504
rect 1956 3487 1964 3496
rect 1887 3476 1933 3484
rect 2067 3476 2113 3484
rect 2296 3484 2304 3513
rect 2436 3507 2444 3516
rect 2536 3516 2573 3524
rect 2127 3476 2304 3484
rect 1856 3456 1973 3464
rect 2107 3456 2153 3464
rect 2356 3464 2364 3493
rect 2536 3484 2544 3516
rect 2667 3516 2733 3524
rect 2787 3516 2953 3524
rect 2996 3507 3004 3533
rect 3056 3516 3133 3524
rect 2816 3484 2824 3493
rect 2427 3476 2744 3484
rect 2816 3476 2853 3484
rect 2187 3456 2364 3464
rect 2467 3456 2693 3464
rect 2736 3464 2744 3476
rect 3036 3484 3044 3513
rect 3056 3507 3064 3516
rect 3427 3516 3453 3524
rect 3476 3516 3613 3524
rect 3476 3507 3484 3516
rect 3696 3524 3704 3533
rect 3836 3527 3844 3536
rect 3896 3527 3904 3576
rect 3967 3576 4113 3584
rect 4147 3576 4653 3584
rect 4947 3576 5033 3584
rect 3927 3556 4073 3564
rect 4667 3556 4953 3564
rect 4027 3536 4693 3544
rect 4707 3536 4733 3544
rect 4887 3536 4953 3544
rect 3696 3516 3753 3524
rect 3907 3516 4013 3524
rect 4147 3516 4193 3524
rect 4247 3516 4293 3524
rect 4647 3516 4773 3524
rect 4787 3516 4833 3524
rect 4956 3516 5033 3524
rect 3107 3496 3153 3504
rect 3527 3496 3573 3504
rect 3627 3496 4093 3504
rect 4107 3496 4233 3504
rect 4347 3496 4373 3504
rect 2987 3476 3044 3484
rect 3087 3476 3233 3484
rect 3247 3476 3353 3484
rect 3387 3476 3473 3484
rect 3507 3476 3533 3484
rect 3767 3476 3833 3484
rect 3927 3476 3973 3484
rect 4027 3476 4093 3484
rect 4436 3484 4444 3513
rect 4956 3507 4964 3516
rect 5056 3516 5073 3524
rect 4507 3496 4533 3504
rect 4747 3496 4913 3504
rect 5056 3504 5064 3516
rect 4987 3496 5064 3504
rect 4407 3476 4444 3484
rect 4456 3484 4464 3493
rect 4456 3476 4533 3484
rect 4547 3476 4813 3484
rect 4987 3476 5013 3484
rect 2736 3456 2893 3464
rect 2907 3456 2973 3464
rect 3007 3456 3033 3464
rect 3167 3456 3273 3464
rect 3347 3456 3813 3464
rect 3847 3456 4033 3464
rect 4047 3456 4073 3464
rect 4087 3456 4173 3464
rect 4367 3456 4413 3464
rect 4707 3456 4893 3464
rect 5027 3456 5133 3464
rect 227 3436 273 3444
rect 287 3436 413 3444
rect 447 3436 793 3444
rect 1007 3436 1313 3444
rect 1487 3436 1593 3444
rect 1647 3436 2033 3444
rect 2087 3436 2113 3444
rect 2147 3436 2373 3444
rect 2387 3436 2953 3444
rect 3027 3436 3193 3444
rect 3227 3436 3273 3444
rect 3387 3436 3653 3444
rect 3807 3436 4113 3444
rect 4187 3436 4433 3444
rect 4907 3436 5093 3444
rect 407 3416 733 3424
rect 887 3416 1473 3424
rect 2027 3416 2253 3424
rect 2407 3416 2753 3424
rect 3067 3416 3173 3424
rect 3247 3416 3333 3424
rect 3367 3416 3553 3424
rect 3587 3416 3733 3424
rect 4027 3416 4733 3424
rect 4847 3416 5053 3424
rect 1627 3396 1773 3404
rect 1807 3396 3153 3404
rect 3207 3396 3293 3404
rect 3547 3396 4053 3404
rect 4107 3396 4353 3404
rect 4367 3396 4473 3404
rect 1087 3376 1233 3384
rect 1247 3376 1493 3384
rect 1507 3376 2013 3384
rect 2227 3376 2573 3384
rect 2627 3376 2844 3384
rect 127 3356 1773 3364
rect 1847 3356 2013 3364
rect 2167 3356 2313 3364
rect 2836 3364 2844 3376
rect 2867 3376 3133 3384
rect 3487 3376 3793 3384
rect 3827 3376 4673 3384
rect 2836 3356 3573 3364
rect 3607 3356 4053 3364
rect 607 3336 953 3344
rect 967 3336 1333 3344
rect 1867 3336 2433 3344
rect 2607 3336 2913 3344
rect 3047 3336 3693 3344
rect 3707 3336 4513 3344
rect 327 3316 393 3324
rect 427 3316 513 3324
rect 1187 3316 1813 3324
rect 1827 3316 2313 3324
rect 2387 3316 2473 3324
rect 2747 3316 3533 3324
rect 3567 3316 3713 3324
rect 3767 3316 3993 3324
rect 4187 3316 5133 3324
rect 107 3296 133 3304
rect 387 3296 413 3304
rect 427 3296 693 3304
rect 1387 3296 1953 3304
rect 1987 3296 2273 3304
rect 2447 3296 2553 3304
rect 2687 3296 2773 3304
rect 2827 3296 2993 3304
rect 3087 3296 3153 3304
rect 3267 3296 4013 3304
rect 4036 3296 4413 3304
rect 127 3276 393 3284
rect 407 3276 453 3284
rect 767 3276 924 3284
rect 67 3256 113 3264
rect 167 3256 353 3264
rect 147 3236 173 3244
rect 207 3236 233 3244
rect 316 3227 324 3256
rect 376 3256 413 3264
rect 376 3244 384 3256
rect 467 3256 493 3264
rect 516 3247 524 3273
rect 547 3256 673 3264
rect 827 3256 853 3264
rect 867 3256 893 3264
rect 347 3236 384 3244
rect 567 3236 593 3244
rect 787 3236 824 3244
rect 767 3216 793 3224
rect 816 3224 824 3236
rect 916 3244 924 3276
rect 1047 3276 1113 3284
rect 1247 3276 1293 3284
rect 1847 3276 2193 3284
rect 2507 3276 2553 3284
rect 2727 3276 2913 3284
rect 2947 3276 3073 3284
rect 3096 3276 3413 3284
rect 1096 3256 1373 3264
rect 1096 3247 1104 3256
rect 1407 3256 1633 3264
rect 1707 3256 1753 3264
rect 1787 3256 2073 3264
rect 2376 3256 2613 3264
rect 867 3236 924 3244
rect 1147 3236 1184 3244
rect 816 3216 913 3224
rect 1067 3216 1093 3224
rect 1176 3207 1184 3236
rect 1327 3236 1353 3244
rect 1376 3236 1453 3244
rect 1276 3224 1284 3233
rect 1376 3224 1384 3236
rect 1467 3236 1513 3244
rect 2376 3244 2384 3256
rect 2647 3256 2713 3264
rect 3096 3264 3104 3276
rect 3496 3276 3633 3284
rect 2907 3256 3104 3264
rect 3127 3256 3473 3264
rect 2056 3236 2384 3244
rect 1276 3216 1384 3224
rect 1407 3216 1533 3224
rect 1647 3216 1864 3224
rect 267 3196 293 3204
rect 307 3196 473 3204
rect 547 3196 573 3204
rect 587 3196 773 3204
rect 887 3196 953 3204
rect 1007 3196 1113 3204
rect 1227 3196 1293 3204
rect 1447 3196 1693 3204
rect 1856 3204 1864 3216
rect 1887 3216 1933 3224
rect 1976 3207 1984 3233
rect 2056 3224 2064 3236
rect 2407 3236 2473 3244
rect 2527 3236 2673 3244
rect 2827 3236 2833 3244
rect 2967 3236 3093 3244
rect 3107 3236 3193 3244
rect 3347 3236 3393 3244
rect 3496 3244 3504 3276
rect 3676 3276 3753 3284
rect 3676 3267 3684 3276
rect 4036 3284 4044 3296
rect 3807 3276 4044 3284
rect 4127 3276 4593 3284
rect 4767 3276 5113 3284
rect 3527 3256 3613 3264
rect 3696 3256 3713 3264
rect 3696 3247 3704 3256
rect 3876 3256 3913 3264
rect 3436 3236 3504 3244
rect 2007 3216 2064 3224
rect 2547 3216 2613 3224
rect 2667 3216 2753 3224
rect 2816 3224 2824 3233
rect 2816 3216 2864 3224
rect 1856 3196 1913 3204
rect 2076 3204 2084 3213
rect 2027 3196 2084 3204
rect 2167 3196 2193 3204
rect 2447 3196 2533 3204
rect 2556 3196 2833 3204
rect 87 3176 193 3184
rect 207 3176 753 3184
rect 847 3176 933 3184
rect 947 3176 1393 3184
rect 1587 3176 1673 3184
rect 1707 3176 2053 3184
rect 2556 3184 2564 3196
rect 2856 3187 2864 3216
rect 2987 3196 3253 3204
rect 3336 3204 3344 3233
rect 3436 3227 3444 3236
rect 3527 3236 3553 3244
rect 3607 3236 3653 3244
rect 3716 3236 3733 3244
rect 3367 3216 3384 3224
rect 3336 3196 3353 3204
rect 3376 3204 3384 3216
rect 3576 3216 3673 3224
rect 3576 3207 3584 3216
rect 3716 3224 3724 3236
rect 3707 3216 3724 3224
rect 3767 3216 3813 3224
rect 3876 3224 3884 3256
rect 3947 3256 3973 3264
rect 4067 3256 4193 3264
rect 4407 3256 4553 3264
rect 3947 3236 4113 3244
rect 4247 3236 4273 3244
rect 3847 3216 3884 3224
rect 3376 3196 3533 3204
rect 3607 3196 3713 3204
rect 3896 3204 3904 3233
rect 3987 3216 4013 3224
rect 4107 3216 4253 3224
rect 4396 3224 4404 3233
rect 4267 3216 4404 3224
rect 3807 3196 3904 3204
rect 3927 3196 4093 3204
rect 4227 3196 4333 3204
rect 4347 3196 4373 3204
rect 4416 3204 4424 3256
rect 4727 3256 5104 3264
rect 4587 3236 4653 3244
rect 4707 3236 4753 3244
rect 4807 3236 4953 3244
rect 5027 3236 5084 3244
rect 4436 3224 4444 3233
rect 5076 3227 5084 3236
rect 4436 3216 4513 3224
rect 4647 3216 4773 3224
rect 4907 3216 4993 3224
rect 5007 3216 5053 3224
rect 4516 3204 4524 3213
rect 4407 3196 4424 3204
rect 4496 3196 4524 3204
rect 2067 3176 2564 3184
rect 2927 3176 3644 3184
rect 647 3156 993 3164
rect 1307 3156 1433 3164
rect 1907 3156 1933 3164
rect 2047 3156 3313 3164
rect 3636 3164 3644 3176
rect 4496 3184 4504 3196
rect 4667 3196 4733 3204
rect 4776 3196 4853 3204
rect 4776 3187 4784 3196
rect 5096 3204 5104 3256
rect 5096 3196 5113 3204
rect 3727 3176 4504 3184
rect 4567 3176 4673 3184
rect 4727 3176 4773 3184
rect 4847 3176 5013 3184
rect 5027 3176 5033 3184
rect 3636 3156 3753 3164
rect 3887 3156 3953 3164
rect 3987 3156 4113 3164
rect 4207 3156 4413 3164
rect 4467 3156 4533 3164
rect 4607 3156 4753 3164
rect 4827 3156 4853 3164
rect 4927 3156 5053 3164
rect 867 3136 913 3144
rect 927 3136 953 3144
rect 967 3136 1913 3144
rect 2467 3136 2573 3144
rect 2967 3136 3053 3144
rect 3107 3136 3453 3144
rect 3467 3136 3593 3144
rect 3627 3136 3733 3144
rect 3787 3136 3933 3144
rect 4007 3136 4293 3144
rect 4367 3136 4493 3144
rect 4607 3136 4793 3144
rect 287 3116 493 3124
rect 507 3116 553 3124
rect 567 3116 1013 3124
rect 1036 3116 1793 3124
rect 1036 3104 1044 3116
rect 1887 3116 1953 3124
rect 2027 3116 2053 3124
rect 2407 3116 2633 3124
rect 2647 3116 2733 3124
rect 2747 3116 2793 3124
rect 3007 3116 3213 3124
rect 3527 3116 3713 3124
rect 3847 3116 3913 3124
rect 3967 3116 4013 3124
rect 4147 3116 4233 3124
rect 4247 3116 4473 3124
rect 4547 3116 4733 3124
rect 4747 3116 4913 3124
rect 416 3096 1044 3104
rect 127 3076 173 3084
rect 416 3084 424 3096
rect 1087 3096 1473 3104
rect 1507 3096 1653 3104
rect 1667 3096 1773 3104
rect 1787 3096 2173 3104
rect 2527 3096 2553 3104
rect 2807 3096 2893 3104
rect 3207 3096 3493 3104
rect 3667 3096 3813 3104
rect 4027 3096 4193 3104
rect 4307 3096 4793 3104
rect 4827 3096 5093 3104
rect 387 3076 424 3084
rect 887 3076 1153 3084
rect 1247 3076 1404 3084
rect 67 3056 373 3064
rect 407 3056 613 3064
rect 687 3056 793 3064
rect 987 3056 1033 3064
rect 1047 3056 1093 3064
rect 1187 3056 1233 3064
rect 1256 3056 1293 3064
rect 107 3036 144 3044
rect 136 3027 144 3036
rect 396 3044 404 3053
rect 167 3036 404 3044
rect 727 3036 813 3044
rect 956 3036 1013 3044
rect 956 3027 964 3036
rect 1127 3036 1193 3044
rect 1256 3044 1264 3056
rect 1396 3064 1404 3076
rect 1427 3076 1493 3084
rect 1536 3076 1653 3084
rect 1396 3056 1453 3064
rect 1536 3064 1544 3076
rect 1787 3076 2033 3084
rect 2047 3076 2213 3084
rect 2267 3076 2673 3084
rect 2767 3076 3093 3084
rect 3407 3076 3453 3084
rect 3567 3076 3693 3084
rect 3747 3076 3784 3084
rect 1487 3056 1544 3064
rect 1567 3056 1613 3064
rect 1767 3056 1813 3064
rect 1847 3056 1973 3064
rect 2096 3056 2253 3064
rect 1227 3036 1264 3044
rect 1327 3036 1373 3044
rect 1396 3036 1433 3044
rect 47 3016 93 3024
rect 447 3016 573 3024
rect 776 3016 793 3024
rect 227 2996 313 3004
rect 367 2996 413 3004
rect 756 2984 764 3013
rect 776 3007 784 3016
rect 847 3016 933 3024
rect 1276 3024 1284 3033
rect 1276 3016 1293 3024
rect 1396 3024 1404 3036
rect 1687 3036 1733 3044
rect 1807 3036 1853 3044
rect 2096 3044 2104 3056
rect 2307 3056 2433 3064
rect 2547 3056 2653 3064
rect 2787 3056 2853 3064
rect 3027 3056 3133 3064
rect 3147 3056 3293 3064
rect 3387 3056 3433 3064
rect 3776 3064 3784 3076
rect 4007 3076 4093 3084
rect 4107 3076 4553 3084
rect 4587 3076 4693 3084
rect 4807 3076 4893 3084
rect 3776 3056 4053 3064
rect 1936 3036 2104 3044
rect 1376 3016 1404 3024
rect 867 2996 1113 3004
rect 1136 2987 1144 3013
rect 1376 3007 1384 3016
rect 1536 3024 1544 3033
rect 1447 3016 1544 3024
rect 1567 3016 1633 3024
rect 1656 3007 1664 3033
rect 1936 3027 1944 3036
rect 2227 3036 2353 3044
rect 2776 3036 2833 3044
rect 1967 3016 1993 3024
rect 2116 3024 2124 3033
rect 2087 3016 2124 3024
rect 2196 3007 2204 3033
rect 2776 3027 2784 3036
rect 3107 3036 3153 3044
rect 3256 3036 3413 3044
rect 2427 3016 2493 3024
rect 2827 3016 2944 3024
rect 2287 2996 2353 3004
rect 2567 2996 2913 3004
rect 2936 3004 2944 3016
rect 3007 3016 3053 3024
rect 3076 3016 3153 3024
rect 3076 3004 3084 3016
rect 3176 3016 3233 3024
rect 2936 2996 3084 3004
rect 3176 3004 3184 3016
rect 3256 3007 3264 3036
rect 3547 3036 3624 3044
rect 3616 3027 3624 3036
rect 3276 3016 3313 3024
rect 3147 2996 3184 3004
rect 756 2976 993 2984
rect 1207 2976 1433 2984
rect 1527 2976 2053 2984
rect 2187 2976 2213 2984
rect 2287 2976 2313 2984
rect 2327 2976 2453 2984
rect 2587 2976 2653 2984
rect 2747 2976 3033 2984
rect 3276 2984 3284 3016
rect 3507 3016 3593 3024
rect 3396 3004 3404 3013
rect 3307 2996 3473 3004
rect 3527 2996 3573 3004
rect 3636 3004 3644 3053
rect 3607 2996 3644 3004
rect 3756 3004 3764 3053
rect 3836 3027 3844 3056
rect 4087 3056 4153 3064
rect 4187 3056 4253 3064
rect 4447 3056 4573 3064
rect 4747 3056 4833 3064
rect 4936 3056 5073 3064
rect 3867 3036 3893 3044
rect 3987 3036 4033 3044
rect 4096 3036 4193 3044
rect 3956 3024 3964 3033
rect 4096 3027 4104 3036
rect 4247 3036 4313 3044
rect 3956 3016 3984 3024
rect 3876 3004 3884 3013
rect 3707 2996 3953 3004
rect 3227 2976 3284 2984
rect 3347 2976 3453 2984
rect 3467 2976 3633 2984
rect 3976 2984 3984 3016
rect 4027 3016 4073 3024
rect 4236 3024 4244 3033
rect 4236 3016 4304 3024
rect 4067 2996 4133 3004
rect 4187 2996 4273 3004
rect 4296 3004 4304 3016
rect 4396 3024 4404 3053
rect 4487 3036 4533 3044
rect 4636 3044 4644 3053
rect 4636 3036 4664 3044
rect 4656 3027 4664 3036
rect 4696 3036 4733 3044
rect 4696 3027 4704 3036
rect 4936 3044 4944 3056
rect 4876 3036 4944 3044
rect 4956 3036 4993 3044
rect 4347 3016 4404 3024
rect 4436 3016 4533 3024
rect 4436 3007 4444 3016
rect 4567 3016 4633 3024
rect 4727 3016 4773 3024
rect 4876 3024 4884 3036
rect 4867 3016 4884 3024
rect 4956 3024 4964 3036
rect 5047 3036 5104 3044
rect 4907 3016 4964 3024
rect 4976 3016 5053 3024
rect 4296 2996 4313 3004
rect 4507 2996 4544 3004
rect 3847 2976 3984 2984
rect 4047 2976 4113 2984
rect 4127 2976 4513 2984
rect 1007 2956 1973 2964
rect 2027 2956 2233 2964
rect 2687 2956 3093 2964
rect 3187 2956 3413 2964
rect 3587 2956 3693 2964
rect 3747 2956 4053 2964
rect 4147 2956 4313 2964
rect 4536 2964 4544 2996
rect 4976 3004 4984 3016
rect 5096 3024 5104 3036
rect 5127 3036 5144 3044
rect 5096 3016 5113 3024
rect 4627 2996 4984 3004
rect 5136 3004 5144 3036
rect 5007 2996 5144 3004
rect 4647 2976 4673 2984
rect 4807 2976 5013 2984
rect 4487 2956 4544 2964
rect 4567 2956 4673 2964
rect 4767 2956 5033 2964
rect 547 2936 633 2944
rect 647 2936 1173 2944
rect 1627 2936 1713 2944
rect 1907 2936 2164 2944
rect 1307 2916 1693 2924
rect 2156 2924 2164 2936
rect 3027 2936 3073 2944
rect 3307 2936 4413 2944
rect 4447 2936 4593 2944
rect 4727 2936 5073 2944
rect 2156 2916 2973 2924
rect 3487 2916 3913 2924
rect 4067 2916 4553 2924
rect 4607 2916 4793 2924
rect 4887 2916 5053 2924
rect 307 2896 473 2904
rect 1087 2896 1333 2904
rect 1607 2896 1693 2904
rect 1767 2896 2833 2904
rect 2947 2896 3793 2904
rect 3887 2896 4133 2904
rect 4167 2896 4293 2904
rect 4347 2896 4513 2904
rect 4587 2896 4653 2904
rect 4767 2896 4893 2904
rect 4947 2896 4993 2904
rect 187 2876 1053 2884
rect 1147 2876 1593 2884
rect 1716 2876 1873 2884
rect 267 2856 1013 2864
rect 1716 2864 1724 2876
rect 1927 2876 2133 2884
rect 2247 2876 2333 2884
rect 2367 2876 2873 2884
rect 3287 2876 3333 2884
rect 3347 2876 4213 2884
rect 4327 2876 4613 2884
rect 4707 2876 4773 2884
rect 4867 2876 5013 2884
rect 1507 2856 1724 2864
rect 1747 2856 1853 2864
rect 1867 2856 2013 2864
rect 2067 2856 2293 2864
rect 2487 2856 2513 2864
rect 2547 2856 2873 2864
rect 2987 2856 3593 2864
rect 3727 2856 3873 2864
rect 4267 2856 4693 2864
rect 367 2836 1133 2844
rect 1887 2836 2033 2844
rect 2067 2836 2393 2844
rect 2607 2836 2653 2844
rect 2667 2836 3033 2844
rect 3207 2836 3933 2844
rect 3967 2836 4533 2844
rect 4687 2836 4793 2844
rect 4827 2836 4993 2844
rect 87 2816 513 2824
rect 96 2776 293 2784
rect 96 2767 104 2776
rect 356 2767 364 2793
rect 387 2776 393 2784
rect 407 2776 413 2784
rect 436 2767 444 2793
rect 476 2767 484 2816
rect 1147 2816 1293 2824
rect 1547 2816 1793 2824
rect 2007 2816 2673 2824
rect 3067 2816 3133 2824
rect 3187 2816 3313 2824
rect 4127 2816 4253 2824
rect 4467 2816 4893 2824
rect 4967 2816 5073 2824
rect 5127 2816 5184 2824
rect 516 2796 533 2804
rect 516 2787 524 2796
rect 607 2796 653 2804
rect 687 2796 704 2804
rect 696 2787 704 2796
rect 907 2796 1113 2804
rect 1167 2796 1184 2804
rect 1176 2787 1184 2796
rect 1247 2796 1893 2804
rect 2147 2796 2253 2804
rect 2267 2796 2373 2804
rect 2387 2796 2413 2804
rect 2427 2796 2573 2804
rect 2587 2796 2733 2804
rect 2747 2796 2753 2804
rect 3107 2796 3273 2804
rect 3947 2796 4173 2804
rect 4567 2796 4684 2804
rect 667 2776 684 2784
rect 676 2767 684 2776
rect 747 2776 793 2784
rect 807 2776 913 2784
rect 1027 2776 1044 2784
rect 1036 2767 1044 2776
rect 1227 2776 1253 2784
rect 1407 2776 1433 2784
rect 1567 2776 1613 2784
rect 1967 2776 2024 2784
rect 47 2756 84 2764
rect 76 2744 84 2756
rect 147 2756 213 2764
rect 967 2756 993 2764
rect 1296 2764 1304 2773
rect 1107 2756 1304 2764
rect 1387 2756 1464 2764
rect 76 2736 153 2744
rect 167 2736 193 2744
rect 307 2736 453 2744
rect 647 2736 973 2744
rect 1047 2736 1153 2744
rect 1187 2736 1413 2744
rect 1456 2744 1464 2756
rect 1696 2764 1704 2773
rect 2016 2767 2024 2776
rect 2047 2776 2224 2784
rect 2216 2767 2224 2776
rect 2347 2776 2593 2784
rect 2607 2776 2613 2784
rect 2627 2776 2893 2784
rect 3196 2776 3373 2784
rect 1487 2756 1544 2764
rect 1456 2736 1513 2744
rect 1536 2744 1544 2756
rect 1596 2756 1704 2764
rect 1536 2736 1553 2744
rect 247 2716 313 2724
rect 327 2716 533 2724
rect 587 2716 853 2724
rect 867 2716 873 2724
rect 1027 2716 1053 2724
rect 1287 2716 1353 2724
rect 1596 2724 1604 2756
rect 1967 2756 2004 2764
rect 1627 2736 1693 2744
rect 1827 2736 1973 2744
rect 1996 2744 2004 2756
rect 1996 2736 2033 2744
rect 2156 2744 2164 2753
rect 2156 2736 2213 2744
rect 1596 2716 1633 2724
rect 1687 2716 1773 2724
rect 1867 2716 2073 2724
rect 2147 2716 2193 2724
rect 2276 2724 2284 2773
rect 2336 2756 2433 2764
rect 2336 2747 2344 2756
rect 2776 2756 2813 2764
rect 2456 2744 2464 2753
rect 2776 2747 2784 2756
rect 2456 2736 2513 2744
rect 2567 2736 2593 2744
rect 2847 2736 2893 2744
rect 2267 2716 2284 2724
rect 2327 2716 2444 2724
rect 127 2696 593 2704
rect 607 2696 713 2704
rect 827 2696 1193 2704
rect 1787 2696 1853 2704
rect 1987 2696 2113 2704
rect 2307 2696 2353 2704
rect 2436 2704 2444 2716
rect 2807 2716 2833 2724
rect 2847 2716 2853 2724
rect 2956 2724 2964 2773
rect 3096 2744 3104 2773
rect 3196 2767 3204 2776
rect 3387 2776 3413 2784
rect 3467 2776 3553 2784
rect 3707 2776 3753 2784
rect 3807 2776 3873 2784
rect 4216 2776 4273 2784
rect 3247 2756 3364 2764
rect 3356 2747 3364 2756
rect 3407 2756 3493 2764
rect 3547 2756 3593 2764
rect 3607 2756 3653 2764
rect 3787 2756 3913 2764
rect 3927 2756 3984 2764
rect 3976 2747 3984 2756
rect 4007 2756 4053 2764
rect 4127 2756 4173 2764
rect 4216 2764 4224 2776
rect 4307 2776 4353 2784
rect 4376 2776 4424 2784
rect 4196 2756 4224 2764
rect 3096 2736 3213 2744
rect 3367 2736 3384 2744
rect 3376 2727 3384 2736
rect 3527 2736 3953 2744
rect 4196 2744 4204 2756
rect 4267 2756 4304 2764
rect 4027 2736 4204 2744
rect 4296 2744 4304 2756
rect 4376 2764 4384 2776
rect 4327 2756 4384 2764
rect 4296 2736 4333 2744
rect 4356 2736 4373 2744
rect 2907 2716 2964 2724
rect 3007 2716 3324 2724
rect 2436 2696 2493 2704
rect 2667 2696 3293 2704
rect 3316 2704 3324 2716
rect 3416 2724 3424 2733
rect 3416 2716 3664 2724
rect 3316 2696 3433 2704
rect 3447 2696 3633 2704
rect 3656 2704 3664 2716
rect 3687 2716 3713 2724
rect 3787 2716 4093 2724
rect 4356 2724 4364 2736
rect 4167 2716 4364 2724
rect 4396 2724 4404 2753
rect 4416 2747 4424 2776
rect 4496 2744 4504 2793
rect 4587 2776 4653 2784
rect 4676 2784 4684 2796
rect 4847 2796 4884 2804
rect 4676 2776 4704 2784
rect 4516 2747 4524 2773
rect 4536 2756 4593 2764
rect 4487 2736 4504 2744
rect 4387 2716 4404 2724
rect 4536 2724 4544 2756
rect 4627 2756 4673 2764
rect 4696 2744 4704 2776
rect 4787 2776 4853 2784
rect 4567 2736 4704 2744
rect 4716 2756 4793 2764
rect 4536 2716 4653 2724
rect 4716 2724 4724 2756
rect 4827 2756 4844 2764
rect 4836 2744 4844 2756
rect 4876 2764 4884 2796
rect 4987 2796 5113 2804
rect 4867 2756 4884 2764
rect 4836 2736 4873 2744
rect 4936 2744 4944 2793
rect 4987 2756 5073 2764
rect 4936 2736 4993 2744
rect 4707 2716 4724 2724
rect 4887 2716 5113 2724
rect 3656 2696 3853 2704
rect 3907 2696 4133 2704
rect 4207 2696 4253 2704
rect 4267 2696 4453 2704
rect 4607 2696 4673 2704
rect 4727 2696 4833 2704
rect 4927 2696 5113 2704
rect 1007 2676 1093 2684
rect 1107 2676 1433 2684
rect 1467 2676 1993 2684
rect 2067 2676 2253 2684
rect 2547 2676 2573 2684
rect 2867 2676 2933 2684
rect 3007 2676 3113 2684
rect 3267 2676 3413 2684
rect 3447 2676 3573 2684
rect 3587 2676 3613 2684
rect 3827 2676 3893 2684
rect 4016 2676 4213 2684
rect 887 2656 1573 2664
rect 1587 2656 1833 2664
rect 1847 2656 2233 2664
rect 2267 2656 2433 2664
rect 2447 2656 2633 2664
rect 2887 2656 3073 2664
rect 4016 2664 4024 2676
rect 4407 2676 4513 2684
rect 4907 2676 4953 2684
rect 3487 2656 4024 2664
rect 4127 2656 4184 2664
rect 847 2636 1753 2644
rect 2387 2636 2933 2644
rect 2967 2636 3104 2644
rect 927 2616 1813 2624
rect 1867 2616 2073 2624
rect 2427 2616 2673 2624
rect 3096 2624 3104 2636
rect 3127 2636 3413 2644
rect 3427 2636 3813 2644
rect 3827 2636 3993 2644
rect 4016 2636 4153 2644
rect 3096 2616 3353 2624
rect 3387 2616 3513 2624
rect 3527 2616 3753 2624
rect 3887 2616 3913 2624
rect 4016 2624 4024 2636
rect 4176 2644 4184 2656
rect 4427 2656 4453 2664
rect 4467 2656 4493 2664
rect 4507 2656 4933 2664
rect 5027 2656 5164 2664
rect 4176 2636 4513 2644
rect 4587 2636 4653 2644
rect 4787 2636 5133 2644
rect 3927 2616 4024 2624
rect 4107 2616 4253 2624
rect 4456 2616 4473 2624
rect 27 2596 173 2604
rect 307 2596 633 2604
rect 987 2596 1013 2604
rect 1047 2596 1233 2604
rect 1447 2596 1533 2604
rect 1547 2596 1873 2604
rect 1887 2596 1993 2604
rect 2127 2596 2353 2604
rect 2367 2596 2633 2604
rect 2647 2596 2873 2604
rect 2887 2596 2913 2604
rect 3187 2596 3253 2604
rect 3287 2596 3373 2604
rect 3747 2596 3793 2604
rect 3847 2596 3893 2604
rect 3947 2596 4033 2604
rect 4456 2604 4464 2616
rect 4527 2616 4773 2624
rect 4867 2616 4973 2624
rect 5067 2616 5133 2624
rect 4416 2596 4464 2604
rect 247 2576 293 2584
rect 467 2576 493 2584
rect 607 2576 653 2584
rect 1196 2576 1453 2584
rect 87 2556 193 2564
rect 407 2556 513 2564
rect 327 2536 373 2544
rect 556 2544 564 2573
rect 1196 2567 1204 2576
rect 1607 2576 1653 2584
rect 1836 2576 1893 2584
rect 627 2556 673 2564
rect 787 2556 813 2564
rect 1267 2556 1304 2564
rect 1296 2547 1304 2556
rect 1567 2556 1613 2564
rect 1676 2556 1733 2564
rect 487 2536 564 2544
rect 587 2536 633 2544
rect 667 2536 684 2544
rect 47 2516 253 2524
rect 487 2516 653 2524
rect 547 2496 593 2504
rect 607 2496 613 2504
rect 676 2504 684 2536
rect 727 2536 733 2544
rect 747 2536 853 2544
rect 1227 2536 1273 2544
rect 1376 2544 1384 2553
rect 1676 2547 1684 2556
rect 1836 2547 1844 2576
rect 1927 2576 2253 2584
rect 2307 2576 2333 2584
rect 2527 2576 2564 2584
rect 1947 2556 2013 2564
rect 2027 2556 2193 2564
rect 2347 2556 2373 2564
rect 1327 2536 1384 2544
rect 1896 2544 1904 2553
rect 2396 2547 2404 2573
rect 2556 2567 2564 2576
rect 2747 2576 2913 2584
rect 3187 2576 3233 2584
rect 3307 2576 3333 2584
rect 3367 2576 3384 2584
rect 2567 2556 2593 2564
rect 2807 2556 2833 2564
rect 2856 2556 3053 2564
rect 1896 2536 1953 2544
rect 2456 2544 2464 2553
rect 2456 2536 2493 2544
rect 2856 2544 2864 2556
rect 3107 2556 3133 2564
rect 2516 2536 2864 2544
rect 707 2516 753 2524
rect 807 2516 913 2524
rect 947 2516 1033 2524
rect 647 2496 684 2504
rect 1056 2504 1064 2533
rect 1087 2516 1584 2524
rect 1056 2496 1073 2504
rect 1576 2504 1584 2516
rect 1607 2516 1913 2524
rect 2227 2516 2253 2524
rect 2516 2524 2524 2536
rect 3167 2536 3253 2544
rect 3376 2544 3384 2576
rect 3407 2576 3484 2584
rect 3407 2556 3453 2564
rect 3476 2564 3484 2576
rect 3567 2576 3653 2584
rect 3676 2576 3953 2584
rect 3476 2556 3584 2564
rect 3376 2536 3553 2544
rect 2327 2516 2524 2524
rect 2687 2516 3013 2524
rect 3347 2516 3433 2524
rect 3467 2516 3533 2524
rect 3576 2524 3584 2556
rect 3676 2564 3684 2576
rect 4127 2576 4213 2584
rect 4287 2576 4313 2584
rect 4327 2576 4353 2584
rect 3627 2556 3684 2564
rect 3747 2556 3833 2564
rect 4007 2556 4153 2564
rect 3667 2536 3693 2544
rect 3867 2536 3933 2544
rect 3987 2536 4033 2544
rect 4047 2536 4173 2544
rect 3547 2516 3584 2524
rect 3647 2516 4093 2524
rect 4147 2516 4193 2524
rect 1576 2496 2333 2504
rect 2447 2496 2533 2504
rect 527 2476 813 2484
rect 1587 2476 1713 2484
rect 1887 2476 2213 2484
rect 2227 2476 2273 2484
rect 2287 2476 2433 2484
rect 2467 2476 2613 2484
rect 2907 2476 3093 2484
rect 3107 2476 3213 2484
rect 3236 2484 3244 2513
rect 3287 2496 3373 2504
rect 3687 2496 4093 2504
rect 3236 2476 3593 2484
rect 3807 2476 4033 2484
rect 4196 2484 4204 2513
rect 4216 2504 4224 2533
rect 4216 2496 4313 2504
rect 4336 2504 4344 2553
rect 4396 2544 4404 2573
rect 4416 2564 4424 2596
rect 4487 2596 4633 2604
rect 4747 2596 4893 2604
rect 4927 2596 5044 2604
rect 4447 2576 4553 2584
rect 4627 2576 4733 2584
rect 4787 2576 4913 2584
rect 4936 2576 5013 2584
rect 4416 2556 4433 2564
rect 4396 2536 4413 2544
rect 4596 2544 4604 2573
rect 4936 2564 4944 2576
rect 4707 2556 4944 2564
rect 4956 2556 4973 2564
rect 4596 2536 4664 2544
rect 4407 2516 4633 2524
rect 4656 2524 4664 2536
rect 4847 2536 4913 2544
rect 4956 2544 4964 2556
rect 5036 2564 5044 2596
rect 4996 2556 5044 2564
rect 4996 2544 5004 2556
rect 4936 2536 4964 2544
rect 4976 2536 5004 2544
rect 4656 2516 4673 2524
rect 4736 2524 4744 2533
rect 4936 2527 4944 2536
rect 4736 2516 4893 2524
rect 4976 2524 4984 2536
rect 5027 2536 5073 2544
rect 4967 2516 4984 2524
rect 5156 2524 5164 2656
rect 5087 2516 5164 2524
rect 4336 2496 4353 2504
rect 4547 2496 4573 2504
rect 4716 2504 4724 2513
rect 4647 2496 4884 2504
rect 4196 2476 4293 2484
rect 4876 2484 4884 2496
rect 5176 2504 5184 2816
rect 4907 2496 5184 2504
rect 4876 2476 4913 2484
rect 1767 2456 3693 2464
rect 3867 2456 4213 2464
rect 4287 2456 4453 2464
rect 4627 2456 4673 2464
rect 4807 2456 5093 2464
rect 1607 2436 1633 2444
rect 1647 2436 1873 2444
rect 1927 2436 2093 2444
rect 2167 2436 2313 2444
rect 2727 2436 2993 2444
rect 3307 2436 3433 2444
rect 3507 2436 4013 2444
rect 4047 2436 4353 2444
rect 4507 2436 4593 2444
rect 4607 2436 4793 2444
rect 5067 2436 5093 2444
rect 467 2416 493 2424
rect 2947 2416 3573 2424
rect 3947 2416 4273 2424
rect 4767 2416 4993 2424
rect 3027 2396 3313 2404
rect 3467 2396 3513 2404
rect 3527 2396 4033 2404
rect 4067 2396 4133 2404
rect 4227 2396 4793 2404
rect 4807 2396 5033 2404
rect 1467 2376 1513 2384
rect 2367 2376 2413 2384
rect 3087 2376 3233 2384
rect 3247 2376 3353 2384
rect 3367 2376 3593 2384
rect 3827 2376 3973 2384
rect 4087 2376 4393 2384
rect 587 2356 1953 2364
rect 3207 2356 3713 2364
rect 3767 2356 3813 2364
rect 3967 2356 4413 2364
rect 367 2336 713 2344
rect 2187 2336 2233 2344
rect 2707 2336 2933 2344
rect 2987 2336 3253 2344
rect 3356 2336 3673 2344
rect 456 2316 753 2324
rect 456 2287 464 2316
rect 1847 2316 2413 2324
rect 2567 2316 2753 2324
rect 2787 2316 3104 2324
rect 487 2296 564 2304
rect 556 2287 564 2296
rect 747 2296 833 2304
rect 2216 2296 2373 2304
rect 67 2276 113 2284
rect 227 2276 324 2284
rect 316 2267 324 2276
rect 496 2276 533 2284
rect 107 2256 173 2264
rect 187 2256 233 2264
rect 496 2264 504 2276
rect 687 2276 713 2284
rect 827 2276 853 2284
rect 867 2276 933 2284
rect 1067 2276 1093 2284
rect 1147 2276 1284 2284
rect 387 2256 504 2264
rect 527 2256 593 2264
rect 607 2256 673 2264
rect 967 2256 993 2264
rect 1016 2264 1024 2273
rect 1016 2256 1173 2264
rect 1276 2264 1284 2276
rect 1307 2276 1373 2284
rect 2007 2276 2053 2284
rect 2107 2276 2133 2284
rect 1276 2256 1344 2264
rect 47 2236 73 2244
rect 407 2236 1053 2244
rect 1167 2236 1213 2244
rect 1336 2244 1344 2256
rect 1396 2264 1404 2273
rect 1367 2256 1404 2264
rect 1416 2264 1424 2273
rect 1416 2256 1473 2264
rect 1587 2256 1773 2264
rect 1947 2256 2033 2264
rect 2067 2256 2153 2264
rect 2216 2264 2224 2296
rect 2627 2296 2713 2304
rect 2727 2296 2793 2304
rect 2867 2296 2904 2304
rect 2236 2276 2273 2284
rect 2236 2267 2244 2276
rect 2707 2276 2733 2284
rect 2827 2276 2873 2284
rect 2207 2256 2224 2264
rect 1336 2236 1393 2244
rect 1407 2236 1433 2244
rect 1467 2236 1493 2244
rect 1536 2244 1544 2253
rect 1536 2236 1553 2244
rect 1896 2244 1904 2253
rect 2816 2247 2824 2273
rect 2896 2264 2904 2296
rect 2987 2296 3033 2304
rect 3096 2304 3104 2316
rect 3127 2316 3173 2324
rect 3216 2316 3333 2324
rect 3096 2296 3113 2304
rect 3216 2304 3224 2316
rect 3356 2307 3364 2336
rect 3727 2336 3913 2344
rect 4007 2336 4233 2344
rect 4387 2336 4713 2344
rect 4747 2336 4813 2344
rect 5087 2336 5104 2344
rect 3496 2316 3633 2324
rect 3167 2296 3224 2304
rect 3247 2296 3344 2304
rect 3336 2287 3344 2296
rect 3416 2296 3433 2304
rect 3416 2287 3424 2296
rect 2967 2276 2993 2284
rect 3047 2276 3093 2284
rect 3147 2276 3173 2284
rect 3227 2276 3324 2284
rect 2836 2256 3113 2264
rect 2836 2247 2844 2256
rect 3167 2256 3293 2264
rect 3316 2264 3324 2276
rect 3496 2284 3504 2316
rect 3687 2316 4213 2324
rect 4327 2316 4333 2324
rect 4347 2316 4473 2324
rect 4667 2316 4693 2324
rect 4756 2316 4873 2324
rect 4756 2307 4764 2316
rect 4887 2316 5073 2324
rect 3647 2296 3833 2304
rect 4087 2296 4173 2304
rect 4267 2296 4353 2304
rect 4447 2296 4513 2304
rect 4536 2296 4593 2304
rect 3536 2284 3544 2293
rect 4536 2287 4544 2296
rect 4856 2296 4893 2304
rect 3476 2276 3504 2284
rect 3516 2276 3544 2284
rect 3476 2267 3484 2276
rect 3316 2256 3333 2264
rect 1687 2236 2424 2244
rect 147 2216 613 2224
rect 1007 2216 1113 2224
rect 1147 2216 1333 2224
rect 1487 2216 1813 2224
rect 1967 2216 2053 2224
rect 2087 2216 2253 2224
rect 2416 2224 2424 2236
rect 2956 2236 3304 2244
rect 2416 2216 2553 2224
rect 2956 2224 2964 2236
rect 2587 2216 2964 2224
rect 2987 2216 3033 2224
rect 3047 2216 3093 2224
rect 3187 2216 3213 2224
rect 3296 2224 3304 2236
rect 3327 2236 3433 2244
rect 3516 2244 3524 2276
rect 3567 2276 3673 2284
rect 3796 2276 3893 2284
rect 3567 2256 3773 2264
rect 3796 2264 3804 2276
rect 3916 2276 3973 2284
rect 3787 2256 3804 2264
rect 3827 2256 3873 2264
rect 3916 2264 3924 2276
rect 4007 2276 4073 2284
rect 4127 2276 4193 2284
rect 4407 2276 4493 2284
rect 4667 2276 4753 2284
rect 4807 2276 4833 2284
rect 3896 2256 3924 2264
rect 4096 2264 4104 2273
rect 4096 2256 4213 2264
rect 3896 2247 3904 2256
rect 4276 2264 4284 2273
rect 4276 2256 4373 2264
rect 4436 2256 4533 2264
rect 3487 2236 3524 2244
rect 3627 2236 3733 2244
rect 3776 2236 3853 2244
rect 3296 2216 3353 2224
rect 3427 2216 3493 2224
rect 3776 2224 3784 2236
rect 3947 2236 3973 2244
rect 4007 2236 4073 2244
rect 4107 2236 4153 2244
rect 4436 2244 4444 2256
rect 4647 2256 4733 2264
rect 4856 2264 4864 2296
rect 4947 2296 5064 2304
rect 5056 2287 5064 2296
rect 4887 2276 4933 2284
rect 5016 2264 5024 2273
rect 4856 2256 5004 2264
rect 5016 2256 5073 2264
rect 4996 2247 5004 2256
rect 5096 2264 5104 2336
rect 5087 2256 5104 2264
rect 4427 2236 4444 2244
rect 4487 2236 4953 2244
rect 5027 2236 5053 2244
rect 3527 2216 3784 2224
rect 3807 2216 4093 2224
rect 4147 2216 4353 2224
rect 4527 2216 4853 2224
rect 5047 2216 5093 2224
rect 267 2196 413 2204
rect 667 2196 1553 2204
rect 1687 2196 1713 2204
rect 2307 2196 2533 2204
rect 2547 2196 2613 2204
rect 2747 2196 2993 2204
rect 3027 2196 3313 2204
rect 3387 2196 3613 2204
rect 3647 2196 3733 2204
rect 3767 2196 3793 2204
rect 3827 2196 4473 2204
rect 4587 2196 4953 2204
rect 807 2176 913 2184
rect 927 2176 1293 2184
rect 1787 2176 2293 2184
rect 2467 2176 2533 2184
rect 2667 2176 2853 2184
rect 2967 2176 3233 2184
rect 3367 2176 3413 2184
rect 3447 2176 4613 2184
rect 4627 2176 4973 2184
rect 4987 2176 4993 2184
rect 287 2156 393 2164
rect 407 2156 433 2164
rect 447 2156 473 2164
rect 487 2156 653 2164
rect 787 2156 873 2164
rect 887 2156 1713 2164
rect 1987 2156 2573 2164
rect 2647 2156 2773 2164
rect 2787 2156 3073 2164
rect 3107 2156 3173 2164
rect 3307 2156 3453 2164
rect 3587 2156 3713 2164
rect 3747 2156 3773 2164
rect 3787 2156 3893 2164
rect 4027 2156 4253 2164
rect 4407 2156 4644 2164
rect 667 2136 933 2144
rect 1107 2136 1213 2144
rect 1227 2136 1833 2144
rect 2027 2136 2213 2144
rect 2307 2136 2733 2144
rect 2767 2136 2953 2144
rect 3007 2136 3573 2144
rect 3627 2136 3753 2144
rect 3807 2136 3853 2144
rect 3887 2136 3953 2144
rect 4207 2136 4273 2144
rect 4307 2136 4613 2144
rect 4636 2144 4644 2156
rect 4707 2156 4793 2164
rect 4636 2136 4693 2144
rect 167 2116 433 2124
rect 447 2116 793 2124
rect 1247 2116 1513 2124
rect 1527 2116 1993 2124
rect 2067 2116 2113 2124
rect 2287 2116 2313 2124
rect 2507 2116 2713 2124
rect 2967 2116 3213 2124
rect 3336 2116 3513 2124
rect 3336 2107 3344 2116
rect 3547 2116 3633 2124
rect 3667 2116 4113 2124
rect 4167 2116 4333 2124
rect 4347 2116 4573 2124
rect 4727 2116 4813 2124
rect 147 2096 344 2104
rect 107 2076 313 2084
rect 336 2084 344 2096
rect 367 2096 413 2104
rect 427 2096 533 2104
rect 587 2096 633 2104
rect 647 2096 833 2104
rect 907 2096 953 2104
rect 1167 2096 1244 2104
rect 336 2076 453 2084
rect 487 2076 524 2084
rect 516 2067 524 2076
rect 547 2076 564 2084
rect 156 2056 193 2064
rect 156 2047 164 2056
rect 67 2036 113 2044
rect 187 2036 253 2044
rect 476 2044 484 2053
rect 556 2047 564 2076
rect 847 2076 973 2084
rect 1236 2084 1244 2096
rect 1267 2096 1284 2104
rect 987 2076 1184 2084
rect 1236 2076 1253 2084
rect 707 2056 1073 2064
rect 1176 2064 1184 2076
rect 1276 2067 1284 2096
rect 1567 2096 1593 2104
rect 1707 2096 1933 2104
rect 1987 2096 2073 2104
rect 2127 2096 2404 2104
rect 1296 2076 1473 2084
rect 1176 2056 1193 2064
rect 387 2036 484 2044
rect 727 2036 773 2044
rect 827 2036 1073 2044
rect 1127 2036 1233 2044
rect 1296 2044 1304 2076
rect 1647 2076 1693 2084
rect 1847 2076 1924 2084
rect 1327 2056 1373 2064
rect 1467 2056 1553 2064
rect 1847 2056 1873 2064
rect 1887 2056 1893 2064
rect 1247 2036 1304 2044
rect 1407 2036 1453 2044
rect 1507 2036 1613 2044
rect 1627 2036 1853 2044
rect 1916 2044 1924 2076
rect 2107 2076 2113 2084
rect 2127 2076 2333 2084
rect 2347 2076 2373 2084
rect 2027 2056 2073 2064
rect 2147 2056 2293 2064
rect 2396 2064 2404 2096
rect 2607 2096 2673 2104
rect 2736 2096 2793 2104
rect 2427 2076 2473 2084
rect 2647 2076 2693 2084
rect 2396 2056 2613 2064
rect 2736 2064 2744 2096
rect 2927 2096 2953 2104
rect 3056 2096 3193 2104
rect 2767 2076 2793 2084
rect 2816 2067 2824 2093
rect 3056 2084 3064 2096
rect 3367 2096 3444 2104
rect 2847 2076 3064 2084
rect 2736 2056 2753 2064
rect 1916 2036 1953 2044
rect 2207 2036 2313 2044
rect 2447 2036 2733 2044
rect 2856 2044 2864 2076
rect 3087 2076 3124 2084
rect 2887 2056 3013 2064
rect 3067 2056 3093 2064
rect 3116 2047 3124 2076
rect 2856 2036 2873 2044
rect 2987 2036 3033 2044
rect 296 2024 304 2033
rect 227 2016 313 2024
rect 467 2016 593 2024
rect 687 2016 853 2024
rect 1367 2016 1413 2024
rect 1427 2016 1573 2024
rect 1927 2016 2133 2024
rect 2307 2016 2353 2024
rect 2587 2016 3093 2024
rect 3156 2024 3164 2073
rect 3196 2044 3204 2093
rect 3216 2076 3233 2084
rect 3216 2067 3224 2076
rect 3316 2076 3373 2084
rect 3247 2056 3293 2064
rect 3316 2047 3324 2076
rect 3396 2076 3413 2084
rect 3396 2064 3404 2076
rect 3376 2056 3404 2064
rect 3436 2064 3444 2096
rect 3667 2096 3833 2104
rect 3847 2096 4013 2104
rect 4067 2096 4133 2104
rect 4167 2096 4184 2104
rect 3527 2076 3893 2084
rect 4027 2076 4153 2084
rect 3436 2056 3544 2064
rect 3376 2047 3384 2056
rect 3536 2047 3544 2056
rect 3776 2056 3793 2064
rect 3196 2036 3244 2044
rect 3156 2016 3193 2024
rect 287 1996 373 2004
rect 427 1996 453 2004
rect 1627 1996 2533 2004
rect 2556 1996 3193 2004
rect 247 1976 673 1984
rect 1547 1976 1713 1984
rect 2556 1984 2564 1996
rect 3236 2004 3244 2036
rect 3267 2036 3313 2044
rect 3467 2036 3493 2044
rect 3607 2036 3653 2044
rect 3687 2036 3753 2044
rect 3776 2027 3784 2056
rect 3816 2056 3853 2064
rect 3816 2044 3824 2056
rect 3867 2056 3913 2064
rect 3936 2047 3944 2073
rect 4176 2067 4184 2096
rect 4207 2096 4293 2104
rect 4327 2096 4433 2104
rect 4467 2096 4484 2104
rect 4196 2067 4204 2093
rect 4287 2076 4324 2084
rect 3967 2056 4073 2064
rect 4087 2056 4113 2064
rect 4227 2056 4293 2064
rect 3807 2036 3824 2044
rect 3967 2036 4273 2044
rect 4316 2044 4324 2076
rect 4387 2076 4413 2084
rect 4427 2076 4453 2084
rect 4447 2056 4464 2064
rect 4316 2036 4373 2044
rect 3267 2016 3353 2024
rect 3367 2016 3413 2024
rect 3427 2016 3693 2024
rect 3927 2016 4233 2024
rect 4267 2016 4293 2024
rect 4456 2024 4464 2056
rect 4476 2047 4484 2096
rect 4527 2096 4624 2104
rect 4616 2084 4624 2096
rect 4647 2096 4744 2104
rect 4616 2076 4653 2084
rect 4736 2084 4744 2096
rect 4787 2096 4833 2104
rect 4847 2096 4873 2104
rect 4896 2096 4933 2104
rect 4896 2084 4904 2096
rect 4996 2096 5013 2104
rect 4736 2076 4904 2084
rect 4507 2056 4613 2064
rect 4547 2036 4633 2044
rect 4656 2044 4664 2053
rect 4656 2036 4673 2044
rect 4456 2016 4513 2024
rect 3236 1996 3453 2004
rect 3487 1996 3513 2004
rect 3647 1996 3873 2004
rect 4127 1996 4433 2004
rect 4487 1996 4584 2004
rect 1847 1976 2564 1984
rect 2907 1976 3393 1984
rect 3407 1976 3813 1984
rect 3847 1976 3953 1984
rect 4007 1976 4033 1984
rect 4047 1976 4233 1984
rect 4287 1976 4553 1984
rect 4576 1984 4584 1996
rect 4716 2004 4724 2073
rect 4736 2044 4744 2076
rect 4827 2056 4853 2064
rect 4736 2036 4773 2044
rect 4796 2044 4804 2053
rect 4796 2036 4893 2044
rect 4916 2044 4924 2073
rect 4996 2067 5004 2096
rect 5047 2076 5104 2084
rect 4947 2056 4973 2064
rect 4916 2036 5013 2044
rect 5047 2036 5073 2044
rect 4887 2016 4953 2024
rect 5096 2024 5104 2076
rect 4987 2016 5104 2024
rect 4627 1996 4724 2004
rect 4576 1976 4753 1984
rect 4847 1976 5053 1984
rect 1747 1956 1793 1964
rect 1807 1956 2353 1964
rect 2407 1956 2493 1964
rect 2547 1956 2653 1964
rect 2667 1956 2913 1964
rect 2927 1956 3133 1964
rect 3187 1956 3413 1964
rect 3536 1956 3573 1964
rect 1167 1936 1753 1944
rect 1867 1936 2713 1944
rect 2767 1936 2973 1944
rect 3536 1944 3544 1956
rect 3727 1956 4133 1964
rect 4227 1956 4253 1964
rect 4547 1956 4713 1964
rect 4747 1956 5073 1964
rect 2987 1936 3544 1944
rect 3567 1936 3833 1944
rect 3907 1936 4073 1944
rect 4147 1936 4293 1944
rect 4307 1936 4973 1944
rect 5067 1936 5113 1944
rect 867 1916 1253 1924
rect 1267 1916 1913 1924
rect 1947 1916 1993 1924
rect 2467 1916 2593 1924
rect 2947 1916 2993 1924
rect 3027 1916 3173 1924
rect 3187 1916 3613 1924
rect 3867 1916 4313 1924
rect 4336 1916 4353 1924
rect 1107 1896 1133 1904
rect 1147 1896 1973 1904
rect 2087 1896 2173 1904
rect 2187 1896 2533 1904
rect 2547 1896 3933 1904
rect 4336 1904 4344 1916
rect 4507 1916 4853 1924
rect 4307 1896 4344 1904
rect 4447 1896 4853 1904
rect 1347 1876 1413 1884
rect 1427 1876 1553 1884
rect 1927 1876 2033 1884
rect 2387 1876 2464 1884
rect 156 1856 373 1864
rect 107 1816 144 1824
rect 56 1787 64 1813
rect 87 1796 113 1804
rect 136 1787 144 1816
rect 156 1807 164 1856
rect 487 1856 733 1864
rect 1487 1856 1633 1864
rect 1647 1856 1673 1864
rect 1707 1856 2393 1864
rect 2456 1864 2464 1876
rect 2487 1876 2513 1884
rect 3087 1876 3253 1884
rect 3287 1876 3593 1884
rect 3627 1876 4293 1884
rect 4387 1876 4913 1884
rect 2456 1856 2493 1864
rect 2707 1856 2793 1864
rect 2827 1856 3033 1864
rect 3127 1856 3333 1864
rect 3396 1856 3873 1864
rect 307 1836 333 1844
rect 447 1836 493 1844
rect 627 1836 693 1844
rect 716 1836 1013 1844
rect 176 1784 184 1833
rect 216 1816 373 1824
rect 216 1807 224 1816
rect 587 1816 653 1824
rect 716 1824 724 1836
rect 1467 1836 1593 1844
rect 2067 1836 2233 1844
rect 2327 1836 2693 1844
rect 2767 1836 2953 1844
rect 3067 1836 3113 1844
rect 3207 1836 3213 1844
rect 3227 1836 3293 1844
rect 3396 1844 3404 1856
rect 3887 1856 4013 1864
rect 4207 1856 4353 1864
rect 4607 1856 4633 1864
rect 4647 1856 4984 1864
rect 3307 1836 3404 1844
rect 3456 1836 3633 1844
rect 667 1816 724 1824
rect 807 1816 913 1824
rect 936 1816 1104 1824
rect 236 1796 253 1804
rect 167 1776 184 1784
rect 236 1784 244 1796
rect 367 1796 433 1804
rect 547 1796 593 1804
rect 727 1796 813 1804
rect 836 1796 853 1804
rect 227 1776 244 1784
rect 267 1776 393 1784
rect 747 1776 793 1784
rect 836 1784 844 1796
rect 936 1804 944 1816
rect 896 1796 944 1804
rect 896 1787 904 1796
rect 1096 1804 1104 1816
rect 1187 1816 1293 1824
rect 1307 1816 1373 1824
rect 1396 1807 1404 1833
rect 1447 1816 1473 1824
rect 1567 1816 1673 1824
rect 1807 1816 2213 1824
rect 2267 1816 2313 1824
rect 2407 1816 2873 1824
rect 2887 1816 2913 1824
rect 2967 1816 3013 1824
rect 3347 1816 3393 1824
rect 3456 1824 3464 1836
rect 3907 1836 3973 1844
rect 4027 1836 4213 1844
rect 4296 1836 4444 1844
rect 3436 1816 3464 1824
rect 1096 1796 1184 1804
rect 827 1776 844 1784
rect 47 1756 73 1764
rect 107 1756 193 1764
rect 207 1756 513 1764
rect 687 1756 833 1764
rect 47 1736 233 1744
rect 247 1736 293 1744
rect 327 1736 333 1744
rect 347 1736 413 1744
rect 567 1736 693 1744
rect 707 1736 753 1744
rect 787 1736 893 1744
rect 956 1744 964 1793
rect 1056 1764 1064 1793
rect 1076 1784 1084 1793
rect 1076 1776 1113 1784
rect 1176 1784 1184 1796
rect 1287 1796 1313 1804
rect 1587 1796 1753 1804
rect 2007 1796 2033 1804
rect 2187 1796 2233 1804
rect 2267 1796 2433 1804
rect 2487 1796 2513 1804
rect 2676 1796 2753 1804
rect 1127 1776 1164 1784
rect 1176 1776 1513 1784
rect 987 1756 1133 1764
rect 1156 1764 1164 1776
rect 1547 1776 1853 1784
rect 1636 1767 1644 1776
rect 2096 1784 2104 1793
rect 2096 1776 2153 1784
rect 2247 1776 2413 1784
rect 2436 1784 2444 1793
rect 2436 1776 2484 1784
rect 1156 1756 1213 1764
rect 1367 1756 1433 1764
rect 1787 1756 1873 1764
rect 1907 1756 1913 1764
rect 1927 1756 2113 1764
rect 2207 1756 2453 1764
rect 2476 1764 2484 1776
rect 2507 1776 2613 1784
rect 2476 1756 2573 1764
rect 2676 1764 2684 1796
rect 2996 1796 3093 1804
rect 2996 1787 3004 1796
rect 3156 1804 3164 1813
rect 3156 1796 3253 1804
rect 3436 1804 3444 1816
rect 3787 1816 3804 1824
rect 3387 1796 3444 1804
rect 2787 1776 2853 1784
rect 3027 1776 3233 1784
rect 3247 1776 3333 1784
rect 3456 1784 3464 1793
rect 3387 1776 3464 1784
rect 3476 1784 3484 1813
rect 3507 1796 3553 1804
rect 3647 1796 3704 1804
rect 3696 1787 3704 1796
rect 3747 1796 3773 1804
rect 3476 1776 3533 1784
rect 3567 1776 3613 1784
rect 3796 1767 3804 1816
rect 3947 1816 3964 1824
rect 3956 1787 3964 1816
rect 4067 1816 4173 1824
rect 4296 1804 4304 1836
rect 4147 1796 4184 1804
rect 2627 1756 2684 1764
rect 3007 1756 3033 1764
rect 3087 1756 3233 1764
rect 3247 1756 3253 1764
rect 3347 1756 3464 1764
rect 956 1736 973 1744
rect 1087 1736 1093 1744
rect 1107 1736 1153 1744
rect 1167 1736 1233 1744
rect 2367 1736 2593 1744
rect 2607 1736 2833 1744
rect 2947 1736 3173 1744
rect 3247 1736 3433 1744
rect 3456 1744 3464 1756
rect 3487 1756 3713 1764
rect 3976 1764 3984 1793
rect 4176 1787 4184 1796
rect 4256 1796 4304 1804
rect 4316 1816 4333 1824
rect 4007 1776 4124 1784
rect 3976 1756 3993 1764
rect 4027 1756 4093 1764
rect 3456 1736 3513 1744
rect 3567 1736 3593 1744
rect 3827 1736 3833 1744
rect 3847 1736 4033 1744
rect 4116 1744 4124 1776
rect 4256 1764 4264 1796
rect 4316 1784 4324 1816
rect 4436 1824 4444 1836
rect 4467 1836 4673 1844
rect 4787 1836 4893 1844
rect 4976 1844 4984 1856
rect 5007 1856 5164 1864
rect 4927 1836 4944 1844
rect 4976 1836 5093 1844
rect 4936 1827 4944 1836
rect 4436 1816 4553 1824
rect 4627 1816 4713 1824
rect 4356 1804 4364 1813
rect 4336 1796 4364 1804
rect 4336 1787 4344 1796
rect 4487 1796 4504 1804
rect 4307 1776 4324 1784
rect 4147 1756 4264 1764
rect 4376 1764 4384 1793
rect 4416 1784 4424 1793
rect 4416 1776 4484 1784
rect 4476 1767 4484 1776
rect 4327 1756 4453 1764
rect 4496 1764 4504 1796
rect 4567 1796 4693 1804
rect 4707 1796 4793 1804
rect 4927 1796 5013 1804
rect 4687 1776 4773 1784
rect 4847 1776 4933 1784
rect 4956 1776 4993 1784
rect 4496 1756 4573 1764
rect 4587 1756 4733 1764
rect 4956 1764 4964 1776
rect 5047 1776 5133 1784
rect 4747 1756 4964 1764
rect 4987 1756 5093 1764
rect 5156 1764 5164 1856
rect 5116 1756 5164 1764
rect 4116 1736 4133 1744
rect 4167 1736 4193 1744
rect 4207 1736 4273 1744
rect 4427 1736 4573 1744
rect 4607 1736 4673 1744
rect 4887 1736 5013 1744
rect 5116 1744 5124 1756
rect 5107 1736 5124 1744
rect 607 1716 973 1724
rect 1127 1716 1173 1724
rect 1196 1716 1493 1724
rect 327 1696 473 1704
rect 527 1696 673 1704
rect 687 1696 933 1704
rect 1196 1704 1204 1716
rect 1527 1716 1853 1724
rect 2287 1716 2373 1724
rect 2387 1716 2673 1724
rect 2827 1716 2913 1724
rect 3047 1716 3113 1724
rect 3267 1716 3313 1724
rect 3927 1716 4113 1724
rect 4207 1716 4293 1724
rect 4487 1716 4733 1724
rect 4787 1716 5053 1724
rect 5087 1716 5133 1724
rect 1187 1696 1204 1704
rect 1267 1696 1613 1704
rect 1807 1696 1933 1704
rect 2027 1696 2273 1704
rect 2307 1696 2733 1704
rect 2927 1696 3893 1704
rect 3947 1696 4113 1704
rect 4147 1696 4353 1704
rect 4367 1696 4653 1704
rect 4807 1696 4833 1704
rect 4847 1696 4873 1704
rect 447 1676 773 1684
rect 856 1676 1213 1684
rect 427 1656 473 1664
rect 856 1664 864 1676
rect 1227 1676 1273 1684
rect 1327 1676 1693 1684
rect 2347 1676 2493 1684
rect 2647 1676 2673 1684
rect 2707 1676 2793 1684
rect 2887 1676 3013 1684
rect 3127 1676 3153 1684
rect 3167 1676 3393 1684
rect 3547 1676 3593 1684
rect 3667 1676 3973 1684
rect 3987 1676 4053 1684
rect 4407 1676 4473 1684
rect 4507 1676 4713 1684
rect 4747 1676 4913 1684
rect 487 1656 864 1664
rect 887 1656 913 1664
rect 927 1656 1013 1664
rect 1027 1656 1193 1664
rect 1207 1656 1653 1664
rect 1667 1656 1733 1664
rect 1847 1656 1873 1664
rect 1927 1656 2073 1664
rect 2167 1656 2193 1664
rect 2207 1656 2433 1664
rect 2747 1656 2773 1664
rect 2867 1656 2964 1664
rect 287 1636 353 1644
rect 367 1636 713 1644
rect 747 1636 773 1644
rect 847 1636 1053 1644
rect 1167 1636 1433 1644
rect 1487 1636 1993 1644
rect 2007 1636 2033 1644
rect 2147 1636 2213 1644
rect 2287 1636 2373 1644
rect 2407 1636 2513 1644
rect 2627 1636 2933 1644
rect 2956 1644 2964 1656
rect 2987 1656 3213 1664
rect 3287 1656 3313 1664
rect 3747 1656 4093 1664
rect 4147 1656 4173 1664
rect 4267 1656 4593 1664
rect 4627 1656 4793 1664
rect 4827 1656 5113 1664
rect 2956 1636 3733 1644
rect 4087 1636 4153 1644
rect 4267 1636 4293 1644
rect 4476 1636 4513 1644
rect 4476 1627 4484 1636
rect 4687 1636 4784 1644
rect 127 1616 173 1624
rect 307 1616 404 1624
rect 216 1596 373 1604
rect 156 1584 164 1593
rect 216 1587 224 1596
rect 56 1576 164 1584
rect 56 1567 64 1576
rect 396 1584 404 1616
rect 547 1616 593 1624
rect 607 1616 633 1624
rect 827 1616 933 1624
rect 947 1616 953 1624
rect 1007 1616 1033 1624
rect 1047 1616 1153 1624
rect 1187 1616 1284 1624
rect 507 1596 573 1604
rect 767 1596 833 1604
rect 776 1587 784 1596
rect 856 1596 873 1604
rect 396 1576 473 1584
rect 647 1576 664 1584
rect 87 1556 153 1564
rect 167 1556 233 1564
rect 496 1564 504 1573
rect 467 1556 504 1564
rect 656 1547 664 1576
rect 856 1584 864 1596
rect 1216 1596 1233 1604
rect 796 1576 864 1584
rect 996 1584 1004 1593
rect 996 1576 1073 1584
rect 796 1564 804 1576
rect 1216 1584 1224 1596
rect 1276 1604 1284 1616
rect 1367 1616 1493 1624
rect 1507 1616 1793 1624
rect 1867 1616 2013 1624
rect 2067 1616 2093 1624
rect 2187 1616 2353 1624
rect 2507 1616 2753 1624
rect 2967 1616 3073 1624
rect 3096 1616 3164 1624
rect 1276 1596 1393 1604
rect 1547 1596 1673 1604
rect 1167 1576 1224 1584
rect 1256 1584 1264 1593
rect 1256 1576 1304 1584
rect 1296 1567 1304 1576
rect 1476 1567 1484 1593
rect 1576 1567 1584 1596
rect 1707 1596 1753 1604
rect 1787 1596 1813 1604
rect 1836 1596 1893 1604
rect 1616 1576 1793 1584
rect 1616 1567 1624 1576
rect 1836 1584 1844 1596
rect 1936 1596 2033 1604
rect 1916 1584 1924 1593
rect 1936 1587 1944 1596
rect 2087 1596 2153 1604
rect 2327 1596 2553 1604
rect 2416 1587 2424 1596
rect 2656 1596 2693 1604
rect 1807 1576 1844 1584
rect 1856 1576 1924 1584
rect 747 1556 804 1564
rect 867 1556 933 1564
rect 1067 1556 1133 1564
rect 1856 1564 1864 1576
rect 2027 1576 2413 1584
rect 2596 1576 2633 1584
rect 2596 1567 2604 1576
rect 1847 1556 2073 1564
rect 2127 1556 2433 1564
rect 2547 1556 2593 1564
rect 2656 1564 2664 1596
rect 2787 1596 2964 1604
rect 2767 1576 2844 1584
rect 2836 1567 2844 1576
rect 2876 1576 2933 1584
rect 2876 1567 2884 1576
rect 2636 1556 2664 1564
rect 2636 1547 2644 1556
rect 2747 1556 2773 1564
rect 2787 1556 2793 1564
rect 2956 1564 2964 1596
rect 3096 1604 3104 1616
rect 3007 1596 3104 1604
rect 3156 1604 3164 1616
rect 3207 1616 3273 1624
rect 3547 1616 3633 1624
rect 3667 1616 3693 1624
rect 3836 1616 3893 1624
rect 3156 1596 3293 1604
rect 3307 1596 3373 1604
rect 3387 1596 3433 1604
rect 3507 1596 3573 1604
rect 3647 1596 3693 1604
rect 2987 1576 3013 1584
rect 3136 1567 3144 1593
rect 3296 1576 3353 1584
rect 3296 1567 3304 1576
rect 3427 1576 3513 1584
rect 3756 1584 3764 1593
rect 3656 1576 3773 1584
rect 2956 1556 3093 1564
rect 3656 1564 3664 1576
rect 3836 1584 3844 1616
rect 3927 1616 3953 1624
rect 4116 1616 4133 1624
rect 3867 1596 3884 1604
rect 3836 1576 3853 1584
rect 3876 1584 3884 1596
rect 3876 1576 3933 1584
rect 4016 1584 4024 1593
rect 3956 1576 4024 1584
rect 3507 1556 3664 1564
rect 3767 1556 3793 1564
rect 3816 1564 3824 1573
rect 3956 1567 3964 1576
rect 4047 1576 4073 1584
rect 3816 1556 3873 1564
rect 3987 1556 4013 1564
rect 4096 1564 4104 1593
rect 4067 1556 4104 1564
rect 4116 1564 4124 1616
rect 4187 1616 4333 1624
rect 4387 1616 4453 1624
rect 4507 1616 4613 1624
rect 4647 1616 4733 1624
rect 4776 1624 4784 1636
rect 4807 1636 4893 1644
rect 4776 1616 4804 1624
rect 4316 1596 4373 1604
rect 4316 1584 4324 1596
rect 4427 1596 4504 1604
rect 4496 1587 4504 1596
rect 4567 1596 4633 1604
rect 4696 1596 4753 1604
rect 4147 1576 4324 1584
rect 4116 1556 4133 1564
rect 4256 1564 4264 1576
rect 4347 1576 4404 1584
rect 4256 1556 4313 1564
rect 487 1536 553 1544
rect 767 1536 813 1544
rect 827 1536 893 1544
rect 1367 1536 1373 1544
rect 1387 1536 1513 1544
rect 1527 1536 1613 1544
rect 1627 1536 1633 1544
rect 1927 1536 2013 1544
rect 2147 1536 2513 1544
rect 2707 1536 3013 1544
rect 3187 1536 3213 1544
rect 4207 1536 4253 1544
rect 4396 1544 4404 1576
rect 4516 1564 4524 1593
rect 4696 1584 4704 1596
rect 4796 1604 4804 1616
rect 4827 1616 4853 1624
rect 4927 1616 5073 1624
rect 4796 1596 4973 1604
rect 5087 1596 5144 1604
rect 4556 1576 4704 1584
rect 4716 1576 4753 1584
rect 4556 1567 4564 1576
rect 4447 1556 4524 1564
rect 4576 1556 4693 1564
rect 4576 1544 4584 1556
rect 4716 1564 4724 1576
rect 4767 1576 4913 1584
rect 5007 1576 5093 1584
rect 4707 1556 4724 1564
rect 4747 1556 4773 1564
rect 4956 1564 4964 1573
rect 4827 1556 5053 1564
rect 4836 1547 4844 1556
rect 5116 1564 5124 1573
rect 5096 1556 5124 1564
rect 4396 1536 4584 1544
rect 4667 1536 4713 1544
rect 4967 1536 4993 1544
rect 5096 1544 5104 1556
rect 5087 1536 5104 1544
rect 5136 1544 5144 1596
rect 5127 1536 5144 1544
rect 587 1516 693 1524
rect 1347 1516 1373 1524
rect 1407 1516 1493 1524
rect 1727 1516 2113 1524
rect 2136 1516 2233 1524
rect 407 1496 653 1504
rect 1047 1496 1253 1504
rect 1267 1496 1273 1504
rect 1287 1496 1733 1504
rect 1887 1496 2053 1504
rect 2136 1504 2144 1516
rect 2767 1516 3493 1524
rect 3527 1516 3673 1524
rect 3896 1516 3973 1524
rect 2067 1496 2144 1504
rect 2167 1496 2293 1504
rect 2467 1496 2713 1504
rect 2807 1496 3593 1504
rect 3896 1504 3904 1516
rect 4087 1516 4213 1524
rect 4227 1516 4353 1524
rect 4367 1516 4413 1524
rect 4527 1516 4553 1524
rect 4687 1516 5053 1524
rect 3607 1496 3904 1504
rect 3947 1496 4233 1504
rect 4247 1496 4433 1504
rect 4587 1496 4853 1504
rect 5067 1496 5133 1504
rect 907 1476 1293 1484
rect 1307 1476 1513 1484
rect 1527 1476 1693 1484
rect 2067 1476 2533 1484
rect 2587 1476 2813 1484
rect 3247 1476 3613 1484
rect 3987 1476 4253 1484
rect 4287 1476 4413 1484
rect 4547 1476 4973 1484
rect 1307 1456 1453 1464
rect 1547 1456 1833 1464
rect 1987 1456 2493 1464
rect 2587 1456 3033 1464
rect 3207 1456 3373 1464
rect 3387 1456 3473 1464
rect 3907 1456 4313 1464
rect 4407 1456 4593 1464
rect 4987 1456 5013 1464
rect 1487 1436 1593 1444
rect 2267 1436 2333 1444
rect 2467 1436 2653 1444
rect 2687 1436 2953 1444
rect 3227 1436 3393 1444
rect 3567 1436 4073 1444
rect 4507 1436 4673 1444
rect 5007 1436 5093 1444
rect 1747 1416 2033 1424
rect 2087 1416 2133 1424
rect 2347 1416 2473 1424
rect 2487 1416 2573 1424
rect 3067 1416 3693 1424
rect 3967 1416 4033 1424
rect 4047 1416 4653 1424
rect 4727 1416 4753 1424
rect 4767 1416 4913 1424
rect 5007 1416 5073 1424
rect 5087 1416 5133 1424
rect 27 1396 353 1404
rect 1427 1396 1433 1404
rect 1447 1396 1573 1404
rect 1587 1396 1824 1404
rect 1687 1376 1793 1384
rect 1816 1384 1824 1396
rect 1847 1396 2053 1404
rect 2087 1396 2313 1404
rect 2327 1396 2673 1404
rect 2707 1396 2793 1404
rect 3187 1396 3473 1404
rect 3587 1396 3653 1404
rect 3847 1396 3953 1404
rect 4007 1396 4273 1404
rect 4487 1396 4613 1404
rect 4907 1396 4973 1404
rect 1816 1376 2093 1384
rect 2107 1376 2213 1384
rect 2387 1376 2484 1384
rect 27 1356 73 1364
rect 327 1356 373 1364
rect 447 1356 633 1364
rect 996 1356 1073 1364
rect 27 1336 53 1344
rect 467 1336 553 1344
rect 927 1336 953 1344
rect 47 1316 133 1324
rect 147 1316 184 1324
rect 176 1307 184 1316
rect 27 1296 53 1304
rect 47 1276 73 1284
rect 196 1264 204 1313
rect 216 1307 224 1333
rect 247 1316 253 1324
rect 267 1316 293 1324
rect 327 1316 413 1324
rect 547 1316 613 1324
rect 727 1316 873 1324
rect 887 1316 973 1324
rect 496 1304 504 1313
rect 996 1307 1004 1356
rect 1107 1356 1313 1364
rect 1707 1356 1913 1364
rect 1967 1356 2204 1364
rect 1127 1336 1173 1344
rect 1187 1336 1253 1344
rect 1287 1336 1313 1344
rect 1467 1336 1553 1344
rect 1667 1336 1773 1344
rect 1887 1336 1904 1344
rect 1016 1307 1024 1333
rect 1087 1316 1213 1324
rect 407 1296 504 1304
rect 627 1296 693 1304
rect 747 1296 773 1304
rect 807 1296 853 1304
rect 927 1296 953 1304
rect 467 1276 513 1284
rect 647 1276 833 1284
rect 1036 1284 1044 1313
rect 1136 1307 1144 1316
rect 1227 1316 1333 1324
rect 1396 1304 1404 1333
rect 1396 1296 1553 1304
rect 1596 1304 1604 1333
rect 1667 1316 1713 1324
rect 1767 1316 1833 1324
rect 1896 1324 1904 1336
rect 1927 1336 1973 1344
rect 2027 1336 2053 1344
rect 2096 1336 2113 1344
rect 1896 1316 1924 1324
rect 1596 1296 1633 1304
rect 1736 1304 1744 1313
rect 1736 1296 1813 1304
rect 1736 1287 1744 1296
rect 1867 1296 1893 1304
rect 987 1276 1044 1284
rect 1087 1276 1173 1284
rect 1267 1276 1273 1284
rect 1287 1276 1493 1284
rect 1767 1276 1853 1284
rect 1916 1284 1924 1316
rect 2096 1307 2104 1336
rect 2196 1344 2204 1356
rect 2227 1356 2273 1364
rect 2287 1356 2453 1364
rect 2476 1364 2484 1376
rect 2507 1376 2704 1384
rect 2476 1356 2553 1364
rect 2607 1356 2673 1364
rect 2696 1364 2704 1376
rect 2727 1376 2813 1384
rect 2887 1376 2913 1384
rect 3107 1376 3133 1384
rect 3307 1376 3633 1384
rect 3676 1384 3684 1393
rect 3676 1376 3793 1384
rect 3887 1376 3993 1384
rect 4187 1376 4213 1384
rect 4307 1376 4613 1384
rect 4647 1376 4813 1384
rect 4967 1376 5033 1384
rect 2696 1356 2753 1364
rect 2787 1356 3233 1364
rect 3576 1356 3593 1364
rect 2147 1336 2184 1344
rect 2196 1336 2333 1344
rect 2176 1324 2184 1336
rect 2387 1336 2464 1344
rect 2176 1316 2344 1324
rect 2336 1307 2344 1316
rect 2396 1316 2433 1324
rect 2396 1307 2404 1316
rect 2127 1296 2133 1304
rect 2147 1296 2273 1304
rect 2456 1304 2464 1336
rect 2527 1336 2824 1344
rect 2496 1324 2504 1333
rect 2496 1316 2544 1324
rect 2456 1296 2493 1304
rect 2536 1304 2544 1316
rect 2567 1316 2593 1324
rect 2616 1316 2773 1324
rect 2616 1307 2624 1316
rect 2816 1324 2824 1336
rect 2847 1336 2893 1344
rect 2927 1336 2973 1344
rect 2996 1336 3193 1344
rect 2996 1327 3004 1336
rect 3276 1336 3313 1344
rect 3276 1327 3284 1336
rect 3347 1336 3444 1344
rect 2816 1316 2944 1324
rect 2936 1307 2944 1316
rect 3087 1316 3113 1324
rect 3167 1316 3193 1324
rect 3307 1316 3373 1324
rect 3436 1324 3444 1336
rect 3467 1336 3564 1344
rect 3556 1327 3564 1336
rect 3436 1316 3533 1324
rect 2536 1296 2573 1304
rect 2667 1296 2733 1304
rect 2847 1296 2893 1304
rect 2987 1296 3133 1304
rect 3187 1296 3213 1304
rect 3227 1296 3413 1304
rect 3576 1304 3584 1356
rect 3627 1356 3933 1364
rect 4067 1356 4093 1364
rect 4147 1356 4224 1364
rect 3727 1336 3773 1344
rect 3827 1336 3853 1344
rect 3907 1336 3973 1344
rect 3987 1336 4013 1344
rect 3607 1316 3633 1324
rect 3567 1296 3584 1304
rect 3676 1304 3684 1333
rect 4036 1324 4044 1333
rect 3707 1316 4044 1324
rect 3676 1296 3733 1304
rect 3927 1296 3993 1304
rect 4076 1304 4084 1333
rect 4147 1316 4193 1324
rect 4216 1324 4224 1356
rect 4327 1356 4344 1364
rect 4256 1344 4264 1353
rect 4336 1347 4344 1356
rect 4447 1356 4564 1364
rect 4556 1347 4564 1356
rect 4747 1356 4804 1364
rect 4247 1336 4264 1344
rect 4287 1336 4333 1344
rect 4607 1336 4633 1344
rect 4216 1316 4333 1324
rect 4076 1296 4313 1304
rect 4436 1304 4444 1313
rect 4387 1296 4444 1304
rect 1887 1276 1924 1284
rect 1936 1276 2053 1284
rect 107 1256 433 1264
rect 447 1256 473 1264
rect 507 1256 753 1264
rect 967 1256 1053 1264
rect 1156 1256 1213 1264
rect 27 1236 113 1244
rect 167 1236 273 1244
rect 296 1236 573 1244
rect 67 1216 113 1224
rect 296 1224 304 1236
rect 1156 1244 1164 1256
rect 1936 1264 1944 1276
rect 2067 1276 2133 1284
rect 2307 1276 2373 1284
rect 2527 1276 2553 1284
rect 2647 1276 2713 1284
rect 2796 1284 2804 1293
rect 2796 1276 3073 1284
rect 3127 1276 3313 1284
rect 3327 1276 3433 1284
rect 3507 1276 3533 1284
rect 3887 1276 4073 1284
rect 4187 1276 4193 1284
rect 4207 1276 4253 1284
rect 4307 1276 4433 1284
rect 1647 1256 1944 1264
rect 2047 1256 2233 1264
rect 2347 1256 2824 1264
rect 1047 1236 1164 1244
rect 1207 1236 1413 1244
rect 1436 1236 1653 1244
rect 127 1216 304 1224
rect 367 1216 533 1224
rect 587 1216 653 1224
rect 667 1216 1233 1224
rect 1287 1216 1373 1224
rect 1436 1224 1444 1236
rect 1667 1236 1753 1244
rect 1807 1236 1893 1244
rect 1907 1236 2273 1244
rect 2447 1236 2633 1244
rect 2816 1244 2824 1256
rect 2847 1256 2873 1264
rect 3036 1256 3173 1264
rect 3036 1244 3044 1256
rect 3287 1256 3833 1264
rect 3847 1256 3953 1264
rect 4047 1256 4173 1264
rect 4187 1256 4353 1264
rect 4456 1264 4464 1313
rect 4476 1284 4484 1313
rect 4496 1307 4504 1333
rect 4567 1316 4653 1324
rect 4527 1296 4593 1304
rect 4476 1276 4573 1284
rect 4776 1284 4784 1333
rect 4796 1287 4804 1356
rect 4856 1356 4873 1364
rect 4856 1304 4864 1356
rect 4987 1356 5004 1364
rect 4936 1344 4944 1353
rect 4936 1336 4984 1344
rect 4887 1316 4953 1324
rect 4856 1296 4893 1304
rect 4976 1304 4984 1336
rect 4996 1307 5004 1356
rect 5107 1356 5144 1364
rect 5076 1336 5113 1344
rect 4936 1296 4984 1304
rect 4767 1276 4784 1284
rect 4827 1276 4873 1284
rect 4456 1256 4473 1264
rect 4527 1256 4813 1264
rect 4936 1264 4944 1296
rect 4967 1276 5033 1284
rect 5076 1267 5084 1336
rect 4887 1256 4944 1264
rect 4987 1256 5053 1264
rect 2816 1236 3044 1244
rect 3807 1236 4293 1244
rect 4327 1236 4353 1244
rect 4447 1236 4653 1244
rect 4727 1236 4753 1244
rect 4767 1236 5113 1244
rect 1387 1216 1444 1224
rect 1567 1216 1813 1224
rect 1847 1216 2073 1224
rect 2167 1216 2353 1224
rect 2547 1216 2873 1224
rect 3727 1216 4013 1224
rect 4127 1216 4373 1224
rect 4467 1216 4533 1224
rect 4547 1216 4573 1224
rect 4607 1216 5093 1224
rect 5136 1224 5144 1356
rect 5127 1216 5144 1224
rect 1087 1196 1153 1204
rect 1167 1196 1253 1204
rect 1327 1196 1593 1204
rect 1627 1196 1773 1204
rect 1947 1196 2013 1204
rect 2027 1196 2053 1204
rect 2287 1196 2673 1204
rect 2687 1196 3333 1204
rect 3467 1196 3813 1204
rect 3947 1196 4253 1204
rect 4347 1196 4513 1204
rect 4667 1196 4973 1204
rect 5027 1196 5073 1204
rect 47 1176 393 1184
rect 567 1176 813 1184
rect 867 1176 1013 1184
rect 1027 1176 1133 1184
rect 1207 1176 1293 1184
rect 1427 1176 1453 1184
rect 1467 1176 1593 1184
rect 1647 1176 1953 1184
rect 2127 1176 2333 1184
rect 2467 1176 2693 1184
rect 2867 1176 3153 1184
rect 3167 1176 3193 1184
rect 3367 1176 3573 1184
rect 3787 1176 3913 1184
rect 3947 1176 3993 1184
rect 4007 1176 4133 1184
rect 4307 1176 4393 1184
rect 4567 1176 4693 1184
rect 4707 1176 4833 1184
rect 4887 1176 5033 1184
rect 347 1156 393 1164
rect 407 1156 973 1164
rect 1007 1156 1093 1164
rect 1227 1156 1873 1164
rect 1947 1156 2193 1164
rect 2327 1156 2373 1164
rect 2427 1156 2573 1164
rect 2607 1156 2613 1164
rect 2627 1156 2773 1164
rect 2787 1156 2853 1164
rect 2896 1156 3733 1164
rect 387 1136 873 1144
rect 927 1136 1093 1144
rect 1227 1136 1413 1144
rect 1467 1136 1573 1144
rect 1687 1136 1713 1144
rect 1747 1136 1773 1144
rect 2007 1136 2113 1144
rect 2167 1136 2253 1144
rect 2487 1136 2833 1144
rect 2896 1144 2904 1156
rect 3747 1156 3953 1164
rect 4127 1156 4513 1164
rect 4567 1156 4753 1164
rect 4767 1156 4853 1164
rect 4867 1156 4933 1164
rect 2867 1136 2904 1144
rect 2967 1136 3013 1144
rect 3047 1136 3173 1144
rect 3247 1136 3373 1144
rect 3667 1136 4004 1144
rect 107 1116 133 1124
rect 287 1116 433 1124
rect 567 1116 584 1124
rect 576 1107 584 1116
rect 747 1116 804 1124
rect 27 1096 73 1104
rect 187 1096 233 1104
rect 287 1096 373 1104
rect 596 1096 613 1104
rect 456 1084 464 1093
rect 596 1084 604 1096
rect 796 1104 804 1116
rect 827 1116 1133 1124
rect 1667 1116 1693 1124
rect 1876 1116 1953 1124
rect 796 1096 833 1104
rect 1027 1096 1113 1104
rect 307 1076 604 1084
rect 416 1067 424 1076
rect 776 1084 784 1093
rect 1236 1087 1244 1113
rect 1267 1096 1293 1104
rect 1347 1096 1384 1104
rect 776 1076 1053 1084
rect 1147 1076 1173 1084
rect 1376 1084 1384 1096
rect 1407 1096 1473 1104
rect 1487 1096 1553 1104
rect 1616 1104 1624 1113
rect 1596 1096 1624 1104
rect 1756 1104 1764 1113
rect 1876 1107 1884 1116
rect 2147 1116 2213 1124
rect 2247 1116 2304 1124
rect 1756 1096 1773 1104
rect 1376 1076 1573 1084
rect 756 1064 764 1073
rect 1596 1067 1604 1096
rect 1987 1096 2053 1104
rect 2107 1096 2133 1104
rect 2167 1096 2184 1104
rect 1627 1076 1713 1084
rect 2047 1076 2153 1084
rect 756 1056 893 1064
rect 1007 1056 1033 1064
rect 1207 1056 1313 1064
rect 1447 1056 1513 1064
rect 2176 1064 2184 1096
rect 2247 1096 2273 1104
rect 2296 1087 2304 1116
rect 2316 1116 2433 1124
rect 2316 1107 2324 1116
rect 2476 1116 2553 1124
rect 2347 1096 2413 1104
rect 2476 1087 2484 1116
rect 2836 1116 2873 1124
rect 2816 1104 2824 1113
rect 2836 1107 2844 1116
rect 3067 1116 3113 1124
rect 3327 1116 3444 1124
rect 3436 1107 3444 1116
rect 3527 1116 3653 1124
rect 3827 1116 3944 1124
rect 2767 1096 2824 1104
rect 2887 1096 2953 1104
rect 3056 1096 3293 1104
rect 2527 1076 2533 1084
rect 2547 1076 2653 1084
rect 2667 1076 2933 1084
rect 3056 1084 3064 1096
rect 3347 1096 3424 1104
rect 2987 1076 3064 1084
rect 3107 1076 3153 1084
rect 3267 1076 3313 1084
rect 3416 1084 3424 1096
rect 3627 1096 3693 1104
rect 3707 1096 3793 1104
rect 3807 1096 3873 1104
rect 3887 1096 3913 1104
rect 3416 1076 3484 1084
rect 2027 1056 2184 1064
rect 2267 1056 2493 1064
rect 2587 1056 2913 1064
rect 2947 1056 3213 1064
rect 3227 1056 3453 1064
rect 3476 1064 3484 1076
rect 3507 1076 3553 1084
rect 3727 1076 3833 1084
rect 3936 1084 3944 1116
rect 3996 1107 4004 1136
rect 4027 1136 4133 1144
rect 4147 1136 4193 1144
rect 4227 1136 4373 1144
rect 4047 1116 4124 1124
rect 4027 1096 4053 1104
rect 4067 1096 4093 1104
rect 4116 1087 4124 1116
rect 4207 1096 4273 1104
rect 3936 1076 4093 1084
rect 4296 1084 4304 1136
rect 4507 1136 4613 1144
rect 4667 1136 4713 1144
rect 4827 1136 4993 1144
rect 4347 1116 4433 1124
rect 4436 1104 4444 1113
rect 4416 1096 4444 1104
rect 4296 1076 4333 1084
rect 4416 1084 4424 1096
rect 4527 1096 4593 1104
rect 4636 1104 4644 1133
rect 4667 1116 4724 1124
rect 4716 1107 4724 1116
rect 4747 1116 4813 1124
rect 4847 1116 4884 1124
rect 4876 1107 4884 1116
rect 4927 1116 4953 1124
rect 4627 1096 4644 1104
rect 4987 1096 5093 1104
rect 4407 1076 4424 1084
rect 4447 1076 4493 1084
rect 4907 1076 4953 1084
rect 4967 1076 5033 1084
rect 3476 1056 3593 1064
rect 3636 1064 3644 1073
rect 3636 1056 4173 1064
rect 4327 1056 4413 1064
rect 4427 1056 4653 1064
rect 4867 1056 5113 1064
rect 547 1036 953 1044
rect 1507 1036 1893 1044
rect 2227 1036 2653 1044
rect 3647 1036 3664 1044
rect 1167 1016 2624 1024
rect 1527 996 1593 1004
rect 1867 996 2373 1004
rect 2387 996 2473 1004
rect 2616 1004 2624 1016
rect 2647 1016 3273 1024
rect 3587 1016 3633 1024
rect 3656 1024 3664 1036
rect 3687 1036 3953 1044
rect 3987 1036 4433 1044
rect 4467 1036 4633 1044
rect 3656 1016 4473 1024
rect 4507 1016 4613 1024
rect 5007 1016 5053 1024
rect 2616 996 3293 1004
rect 3347 996 3533 1004
rect 3547 996 3773 1004
rect 4007 996 4053 1004
rect 4247 996 4553 1004
rect 1387 976 2413 984
rect 2567 976 2693 984
rect 2927 976 3133 984
rect 3147 976 3253 984
rect 3287 976 4004 984
rect 307 956 333 964
rect 347 956 933 964
rect 1627 956 1653 964
rect 1827 956 1884 964
rect 947 936 1833 944
rect 1876 944 1884 956
rect 2107 956 2533 964
rect 2747 956 2773 964
rect 3356 956 3533 964
rect 1876 936 2193 944
rect 2227 936 2613 944
rect 2667 936 3033 944
rect 3356 944 3364 956
rect 3547 956 3593 964
rect 3907 956 3973 964
rect 3996 964 4004 976
rect 4107 976 4233 984
rect 4367 976 4513 984
rect 5067 976 5133 984
rect 3996 956 4124 964
rect 3187 936 3364 944
rect 3387 936 3453 944
rect 3487 936 3893 944
rect 3947 936 4093 944
rect 4116 944 4124 956
rect 4207 956 4413 964
rect 4116 936 4533 944
rect 4807 936 5113 944
rect 1007 916 1533 924
rect 1587 916 1653 924
rect 1667 916 1773 924
rect 1787 916 2233 924
rect 2247 916 2453 924
rect 2647 916 2713 924
rect 2896 916 4313 924
rect 2896 907 2904 916
rect 4516 916 4573 924
rect 607 896 793 904
rect 1547 896 1793 904
rect 2087 896 2233 904
rect 2287 896 2513 904
rect 2667 896 2753 904
rect 3367 896 3753 904
rect 3807 896 3933 904
rect 4516 904 4524 916
rect 4927 916 5033 924
rect 3967 896 4524 904
rect 4547 896 4873 904
rect 4887 896 5093 904
rect 387 876 513 884
rect 787 876 813 884
rect 1207 876 1633 884
rect 1687 876 1693 884
rect 1707 876 1753 884
rect 2067 876 2093 884
rect 2187 876 2253 884
rect 2267 876 2333 884
rect 2367 876 2824 884
rect 207 856 233 864
rect 247 856 253 864
rect 687 856 773 864
rect 836 856 853 864
rect 107 836 193 844
rect 407 836 433 844
rect 447 836 453 844
rect 836 844 844 856
rect 927 856 953 864
rect 967 856 1153 864
rect 1467 856 1533 864
rect 1676 856 1713 864
rect 767 836 844 844
rect 1187 836 1233 844
rect 256 824 264 833
rect 187 816 473 824
rect 496 824 504 833
rect 496 816 893 824
rect 1276 824 1284 833
rect 1276 816 1353 824
rect 1447 816 1593 824
rect 1676 824 1684 856
rect 1787 856 1893 864
rect 2087 856 2133 864
rect 2147 856 2153 864
rect 2327 856 2473 864
rect 2487 856 2493 864
rect 2627 856 2693 864
rect 2747 856 2793 864
rect 2816 864 2824 876
rect 3016 876 3073 884
rect 2816 856 3004 864
rect 1907 836 1953 844
rect 2027 836 2104 844
rect 2096 827 2104 836
rect 1647 816 1684 824
rect 1867 816 1993 824
rect 2007 816 2073 824
rect 2227 816 2273 824
rect 67 796 133 804
rect 247 796 273 804
rect 527 796 533 804
rect 547 796 933 804
rect 1127 796 1473 804
rect 1527 796 1593 804
rect 1687 796 1773 804
rect 1787 796 1813 804
rect 1987 796 2213 804
rect 2296 804 2304 833
rect 2316 827 2324 853
rect 2367 836 2613 844
rect 2647 836 2693 844
rect 2727 836 2753 844
rect 2816 836 2873 844
rect 2816 827 2824 836
rect 2907 836 2973 844
rect 2336 816 2573 824
rect 2336 804 2344 816
rect 2847 816 2884 824
rect 2876 807 2884 816
rect 2996 824 3004 856
rect 2967 816 3004 824
rect 3016 824 3024 876
rect 3267 876 3393 884
rect 3667 876 3824 884
rect 3816 867 3824 876
rect 4036 876 4053 884
rect 3047 856 3333 864
rect 3447 856 3664 864
rect 3067 836 3133 844
rect 3227 836 3333 844
rect 3347 836 3353 844
rect 3447 836 3633 844
rect 3656 827 3664 856
rect 3747 856 3773 864
rect 3867 856 3933 864
rect 3947 856 4024 864
rect 4016 847 4024 856
rect 3727 836 3753 844
rect 3767 836 3833 844
rect 3887 836 4004 844
rect 3996 827 4004 836
rect 3016 816 3064 824
rect 3056 807 3064 816
rect 3316 816 3473 824
rect 3316 807 3324 816
rect 3487 816 3553 824
rect 3567 816 3573 824
rect 3687 816 3793 824
rect 4036 824 4044 876
rect 4096 876 4113 884
rect 4076 827 4084 853
rect 4027 816 4044 824
rect 2296 796 2344 804
rect 2527 796 2633 804
rect 2647 796 2673 804
rect 3007 796 3033 804
rect 3147 796 3173 804
rect 3367 796 3673 804
rect 3707 796 3893 804
rect 4096 804 4104 876
rect 4167 876 4293 884
rect 4487 876 4604 884
rect 4596 867 4604 876
rect 4687 876 4713 884
rect 4827 876 4953 884
rect 4116 856 4213 864
rect 4116 847 4124 856
rect 4236 856 4253 864
rect 4167 836 4213 844
rect 4236 824 4244 856
rect 4347 856 4513 864
rect 4667 856 4733 864
rect 4787 856 4884 864
rect 4876 847 4884 856
rect 4347 836 4373 844
rect 4387 836 4393 844
rect 4487 836 4573 844
rect 4587 836 4693 844
rect 4827 836 4853 844
rect 4187 816 4244 824
rect 4527 816 4613 824
rect 4627 816 4633 824
rect 4707 816 4913 824
rect 4947 816 4973 824
rect 4067 796 4104 804
rect 4407 796 4453 804
rect 4467 796 4593 804
rect 4807 796 4833 804
rect 5027 796 5053 804
rect 227 776 333 784
rect 1267 776 1673 784
rect 1927 776 2113 784
rect 2287 776 2413 784
rect 2427 776 3153 784
rect 3207 776 3493 784
rect 3507 776 3693 784
rect 3787 776 4133 784
rect 4147 776 4233 784
rect 4327 776 4673 784
rect 127 756 313 764
rect 667 756 793 764
rect 807 756 993 764
rect 1007 756 1073 764
rect 1327 756 1573 764
rect 1747 756 1853 764
rect 1907 756 2013 764
rect 2047 756 2053 764
rect 2067 756 3413 764
rect 3627 756 4153 764
rect 4347 756 5013 764
rect 1427 736 1473 744
rect 1487 736 1613 744
rect 1647 736 1773 744
rect 1827 736 1893 744
rect 1907 736 1933 744
rect 2127 736 2533 744
rect 2567 736 2633 744
rect 2667 736 2793 744
rect 2907 736 3253 744
rect 3527 736 3913 744
rect 3927 736 4033 744
rect 4207 736 4313 744
rect 4327 736 4633 744
rect 887 716 1393 724
rect 1627 716 1753 724
rect 1867 716 2113 724
rect 2187 716 2713 724
rect 2947 716 4353 724
rect 4547 716 4693 724
rect 147 696 313 704
rect 927 696 1013 704
rect 1167 696 1273 704
rect 1307 696 1313 704
rect 1327 696 1633 704
rect 1767 696 1873 704
rect 2187 696 2293 704
rect 2327 696 2593 704
rect 2867 696 2953 704
rect 2967 696 3233 704
rect 3267 696 3673 704
rect 4087 696 4253 704
rect 4267 696 4653 704
rect 4667 696 4753 704
rect 327 676 553 684
rect 767 676 973 684
rect 1047 676 1073 684
rect 1087 676 1193 684
rect 1207 676 1693 684
rect 1847 676 1953 684
rect 1967 676 2013 684
rect 2267 676 2373 684
rect 2627 676 2753 684
rect 2947 676 3113 684
rect 3127 676 3213 684
rect 3287 676 3353 684
rect 3447 676 3644 684
rect 87 656 193 664
rect 747 656 773 664
rect 847 656 873 664
rect 987 656 1173 664
rect 1267 656 1353 664
rect 1387 656 1653 664
rect 1707 656 1833 664
rect 1867 656 1993 664
rect 2107 656 2233 664
rect 2267 656 2453 664
rect 2467 656 2493 664
rect 2507 656 2553 664
rect 2707 656 2753 664
rect 2876 656 2913 664
rect 47 636 173 644
rect 227 636 273 644
rect 387 636 433 644
rect 456 627 464 653
rect 507 636 533 644
rect 607 636 673 644
rect 987 636 1064 644
rect 76 616 93 624
rect 76 564 84 616
rect 127 616 253 624
rect 487 616 513 624
rect 627 616 653 624
rect 716 624 724 633
rect 1056 627 1064 636
rect 1167 636 1264 644
rect 716 616 853 624
rect 907 616 933 624
rect 1127 616 1213 624
rect 556 604 564 613
rect 307 596 564 604
rect 707 596 733 604
rect 767 596 773 604
rect 787 596 1153 604
rect 1256 604 1264 636
rect 1276 636 1313 644
rect 1276 627 1284 636
rect 1416 636 1493 644
rect 1416 624 1424 636
rect 1667 636 1713 644
rect 1727 636 1733 644
rect 1756 636 1913 644
rect 1756 627 1764 636
rect 2187 636 2244 644
rect 1387 616 1424 624
rect 1447 616 1513 624
rect 1547 616 1693 624
rect 1787 616 1853 624
rect 1907 616 1933 624
rect 1256 596 1273 604
rect 1316 604 1324 613
rect 1436 604 1444 613
rect 1316 596 1444 604
rect 1587 596 1913 604
rect 96 584 104 593
rect 96 576 413 584
rect 427 576 593 584
rect 1107 576 1333 584
rect 1487 576 1593 584
rect 1747 576 1993 584
rect 2036 584 2044 613
rect 2136 607 2144 633
rect 2236 627 2244 636
rect 2307 636 2333 644
rect 2467 636 2513 644
rect 2727 636 2804 644
rect 2307 616 2364 624
rect 2167 596 2313 604
rect 2356 604 2364 616
rect 2387 616 2433 624
rect 2487 616 2533 624
rect 2576 604 2584 613
rect 2356 596 2584 604
rect 2656 604 2664 633
rect 2687 616 2773 624
rect 2796 607 2804 636
rect 2876 624 2884 656
rect 2996 656 3033 664
rect 2996 644 3004 656
rect 3067 656 3073 664
rect 3087 656 3133 664
rect 3227 656 3273 664
rect 3287 656 3373 664
rect 3387 656 3453 664
rect 3527 656 3613 664
rect 2907 636 3004 644
rect 3027 636 3073 644
rect 3216 636 3393 644
rect 2876 616 2904 624
rect 2656 596 2753 604
rect 2896 604 2904 616
rect 2927 616 2953 624
rect 3096 624 3104 633
rect 3216 627 3224 636
rect 3416 636 3573 644
rect 3416 627 3424 636
rect 3636 644 3644 676
rect 3667 676 3833 684
rect 3967 676 4193 684
rect 4207 676 4413 684
rect 4427 676 4513 684
rect 4567 676 4973 684
rect 3727 656 3773 664
rect 3827 656 3853 664
rect 3887 656 3984 664
rect 3976 647 3984 656
rect 4007 656 4173 664
rect 4227 656 4264 664
rect 3636 636 3753 644
rect 3696 627 3704 636
rect 3767 636 3824 644
rect 3027 616 3104 624
rect 3127 616 3193 624
rect 3507 616 3593 624
rect 3747 616 3793 624
rect 3816 624 3824 636
rect 3987 636 4093 644
rect 4207 636 4244 644
rect 4236 627 4244 636
rect 4256 627 4264 656
rect 4287 656 4364 664
rect 4356 644 4364 656
rect 4467 656 4493 664
rect 4796 656 4853 664
rect 4356 636 4544 644
rect 4356 627 4364 636
rect 4536 627 4544 636
rect 4756 636 4773 644
rect 3816 616 3953 624
rect 4067 616 4193 624
rect 4367 616 4433 624
rect 4647 616 4733 624
rect 2896 596 2933 604
rect 2967 596 2993 604
rect 3047 596 3073 604
rect 3447 596 3513 604
rect 3567 596 3633 604
rect 3987 596 4033 604
rect 4187 596 4273 604
rect 4476 604 4484 613
rect 4756 604 4764 636
rect 4796 624 4804 656
rect 4907 656 4933 664
rect 4827 636 4853 644
rect 4896 636 4933 644
rect 4896 624 4904 636
rect 4287 596 4764 604
rect 4776 616 4804 624
rect 4856 616 4904 624
rect 2007 576 2193 584
rect 2407 576 2873 584
rect 2887 576 2973 584
rect 3296 584 3304 593
rect 3067 576 3633 584
rect 3776 584 3784 593
rect 4776 587 4784 616
rect 4856 604 4864 616
rect 4927 616 4973 624
rect 4807 596 4864 604
rect 4887 596 4953 604
rect 3767 576 3784 584
rect 4007 576 4073 584
rect 4087 576 4133 584
rect 4207 576 4393 584
rect 4407 576 4593 584
rect 67 556 84 564
rect 447 556 493 564
rect 1427 556 1713 564
rect 2667 556 2833 564
rect 2847 556 2953 564
rect 3167 556 3173 564
rect 3187 556 3333 564
rect 3347 556 3913 564
rect 4707 556 4993 564
rect 27 536 153 544
rect 167 536 353 544
rect 2247 536 2733 544
rect 2787 536 3213 544
rect 27 516 53 524
rect 227 516 693 524
rect 827 516 1073 524
rect 3087 516 3433 524
rect 3447 516 3613 524
rect 287 496 453 504
rect 2827 496 3813 504
rect 587 476 893 484
rect 927 476 1893 484
rect 2067 476 2113 484
rect 2567 476 2613 484
rect 2707 476 2793 484
rect 3107 476 4253 484
rect 4647 476 4673 484
rect 727 456 1013 464
rect 1527 456 1633 464
rect 1647 456 1673 464
rect 1707 456 1753 464
rect 2047 456 2233 464
rect 2327 456 2733 464
rect 2807 456 2853 464
rect 2867 456 3113 464
rect 3127 456 4393 464
rect 567 436 953 444
rect 1027 436 1133 444
rect 1407 436 2673 444
rect 3607 436 3813 444
rect 3927 436 4033 444
rect 107 416 293 424
rect 307 416 873 424
rect 887 416 1233 424
rect 1687 416 1793 424
rect 2087 416 2313 424
rect 2527 416 2573 424
rect 2847 416 3213 424
rect 3667 416 3893 424
rect 47 396 113 404
rect 127 396 304 404
rect 87 376 153 384
rect 176 376 273 384
rect 176 367 184 376
rect 296 384 304 396
rect 327 396 353 404
rect 367 396 393 404
rect 636 396 933 404
rect 636 384 644 396
rect 2107 396 2413 404
rect 2607 396 2833 404
rect 2947 396 3913 404
rect 4287 396 4333 404
rect 4627 396 4713 404
rect 4936 396 4973 404
rect 296 376 644 384
rect 747 376 793 384
rect 907 376 924 384
rect 27 356 53 364
rect 267 356 333 364
rect 427 356 453 364
rect 507 356 593 364
rect 916 364 924 376
rect 947 376 973 384
rect 1147 376 1193 384
rect 1207 376 1333 384
rect 1347 376 1433 384
rect 1787 376 1793 384
rect 1807 376 1873 384
rect 1967 376 2033 384
rect 2107 376 2193 384
rect 2447 376 2513 384
rect 2527 376 2564 384
rect 727 356 784 364
rect 916 356 953 364
rect 27 336 133 344
rect 216 344 224 353
rect 187 336 224 344
rect 247 336 273 344
rect 407 336 633 344
rect 676 327 684 353
rect 696 344 704 353
rect 776 347 784 356
rect 1187 356 1213 364
rect 1367 356 1933 364
rect 1987 356 2013 364
rect 2267 356 2373 364
rect 2467 356 2493 364
rect 2556 364 2564 376
rect 2587 376 2733 384
rect 2767 376 2813 384
rect 2827 376 2893 384
rect 3047 376 3133 384
rect 3187 376 3213 384
rect 3227 376 3253 384
rect 3307 376 3313 384
rect 3327 376 3333 384
rect 3367 376 3413 384
rect 3507 376 3553 384
rect 3567 376 3644 384
rect 3636 367 3644 376
rect 3707 376 3733 384
rect 3767 376 3784 384
rect 2556 356 2613 364
rect 2987 356 3033 364
rect 3127 356 3153 364
rect 3387 356 3433 364
rect 3527 356 3553 364
rect 3727 356 3753 364
rect 696 336 733 344
rect 927 336 1113 344
rect 1867 336 1993 344
rect 207 316 273 324
rect 287 316 433 324
rect 447 316 553 324
rect 707 316 753 324
rect 967 316 993 324
rect 1467 316 2033 324
rect 2056 324 2064 353
rect 2136 327 2144 353
rect 2156 327 2164 353
rect 2207 336 2333 344
rect 2347 336 2493 344
rect 2616 336 2713 344
rect 2616 327 2624 336
rect 2836 327 2844 353
rect 2936 344 2944 353
rect 2887 336 2944 344
rect 3007 336 3093 344
rect 3107 336 3273 344
rect 3327 336 3473 344
rect 2056 316 2093 324
rect 2547 316 2573 324
rect 2927 316 3173 324
rect 3267 316 3353 324
rect 3367 316 3453 324
rect 3596 324 3604 353
rect 3776 347 3784 376
rect 4187 376 4393 384
rect 4507 376 4653 384
rect 4667 376 4693 384
rect 3856 364 3864 373
rect 4716 367 4724 393
rect 4836 384 4844 393
rect 4827 376 4844 384
rect 4936 367 4944 396
rect 4967 376 5073 384
rect 3816 356 3864 364
rect 4096 356 4173 364
rect 3816 347 3824 356
rect 3627 336 3653 344
rect 3847 336 4053 344
rect 4096 344 4104 356
rect 4347 356 4433 364
rect 4567 356 4624 364
rect 4067 336 4104 344
rect 4127 336 4193 344
rect 4207 336 4373 344
rect 4516 344 4524 353
rect 4516 336 4593 344
rect 4616 344 4624 356
rect 4647 356 4673 364
rect 4847 356 4933 364
rect 5047 356 5093 364
rect 4616 336 4753 344
rect 4767 336 4853 344
rect 4867 336 4913 344
rect 5016 344 5024 353
rect 5016 336 5053 344
rect 3596 316 3673 324
rect 3767 316 3873 324
rect 3987 316 4093 324
rect 4347 316 4533 324
rect 4647 316 4673 324
rect 5027 316 5073 324
rect 347 296 473 304
rect 667 296 873 304
rect 2047 296 2273 304
rect 2287 296 2353 304
rect 2527 296 2633 304
rect 2767 296 3153 304
rect 3187 296 3433 304
rect 3547 296 3733 304
rect 3827 296 3873 304
rect 3887 296 3953 304
rect 4007 296 4013 304
rect 4027 296 4133 304
rect 4147 296 4313 304
rect 4547 296 4873 304
rect 4887 296 4993 304
rect 467 276 833 284
rect 947 276 1153 284
rect 1167 276 1233 284
rect 1567 276 1693 284
rect 1707 276 1853 284
rect 1927 276 2153 284
rect 2307 276 2473 284
rect 2947 276 3053 284
rect 3107 276 3533 284
rect 3687 276 4493 284
rect 4787 276 4873 284
rect 87 256 113 264
rect 127 256 393 264
rect 1487 256 1673 264
rect 2287 256 2513 264
rect 2627 256 2753 264
rect 2907 256 3193 264
rect 3207 256 3233 264
rect 3407 256 3513 264
rect 3527 256 3713 264
rect 3967 256 4033 264
rect 4087 256 4213 264
rect 407 236 493 244
rect 507 236 533 244
rect 1067 236 1353 244
rect 1607 236 1833 244
rect 1907 236 2073 244
rect 2187 236 2393 244
rect 2487 236 2593 244
rect 2607 236 3573 244
rect 3807 236 4773 244
rect 547 216 1013 224
rect 1027 216 1133 224
rect 1627 216 1713 224
rect 1727 216 1753 224
rect 1827 216 2373 224
rect 2427 216 2633 224
rect 2667 216 2693 224
rect 2767 216 2993 224
rect 3267 216 3413 224
rect 3427 216 3533 224
rect 3547 216 3653 224
rect 1007 196 1313 204
rect 1547 196 1913 204
rect 2007 196 2453 204
rect 2467 196 2953 204
rect 3407 196 3513 204
rect 3527 196 3873 204
rect 4427 196 4573 204
rect 4747 196 4853 204
rect 4867 196 4893 204
rect 67 176 173 184
rect 187 176 213 184
rect 347 176 653 184
rect 667 176 673 184
rect 787 176 813 184
rect 827 176 1233 184
rect 1287 176 1573 184
rect 1687 176 1773 184
rect 1967 176 2133 184
rect 2147 176 2213 184
rect 2247 176 2313 184
rect 2327 176 2404 184
rect 47 156 93 164
rect 167 156 244 164
rect 236 147 244 156
rect 267 156 373 164
rect 587 156 613 164
rect 867 156 1073 164
rect 1087 156 1493 164
rect 1596 147 1604 173
rect 1667 156 1693 164
rect 1707 156 1804 164
rect 567 136 633 144
rect 647 136 693 144
rect 767 136 853 144
rect 1047 136 1093 144
rect 1107 136 1153 144
rect 1207 136 1273 144
rect 1527 136 1553 144
rect 1656 144 1664 153
rect 1796 147 1804 156
rect 1907 156 1973 164
rect 1987 156 2193 164
rect 2396 164 2404 176
rect 2507 176 2693 184
rect 2747 176 2873 184
rect 2887 176 3013 184
rect 3036 176 3133 184
rect 2396 156 2833 164
rect 3036 164 3044 176
rect 3147 176 3213 184
rect 3327 176 3453 184
rect 3467 176 3493 184
rect 3607 176 3733 184
rect 4127 176 4213 184
rect 4227 176 4253 184
rect 4607 176 4964 184
rect 3007 156 3044 164
rect 3116 156 3273 164
rect 1647 136 1664 144
rect 1847 136 1873 144
rect 2007 136 2113 144
rect 2167 136 2193 144
rect 2376 144 2384 153
rect 3116 147 3124 156
rect 3296 156 3353 164
rect 3296 147 3304 156
rect 3427 156 3473 164
rect 3487 156 3913 164
rect 3996 156 4113 164
rect 2376 136 2413 144
rect 2627 136 2853 144
rect 3027 136 3073 144
rect 3467 136 3553 144
rect 3687 136 3713 144
rect 3767 136 3833 144
rect 3996 144 4004 156
rect 4187 156 4293 164
rect 4476 164 4484 173
rect 4307 156 4553 164
rect 4687 156 4733 164
rect 4756 156 4793 164
rect 4756 147 4764 156
rect 4807 156 4913 164
rect 4927 156 4933 164
rect 4956 147 4964 176
rect 3976 136 4004 144
rect 387 116 473 124
rect 487 116 513 124
rect 687 116 793 124
rect 807 116 833 124
rect 936 124 944 133
rect 887 116 944 124
rect 1376 124 1384 133
rect 1307 116 1384 124
rect 1687 116 1753 124
rect 1956 124 1964 133
rect 3976 127 3984 136
rect 4047 136 4124 144
rect 1807 116 1964 124
rect 2187 116 2353 124
rect 2567 116 2713 124
rect 2967 116 3113 124
rect 3127 116 3153 124
rect 3207 116 3213 124
rect 3227 116 3773 124
rect 1256 104 1264 113
rect 807 96 1264 104
rect 3947 96 4093 104
rect 4116 104 4124 136
rect 4167 136 4224 144
rect 4147 116 4193 124
rect 4216 124 4224 136
rect 4307 136 4333 144
rect 4356 136 4433 144
rect 4356 124 4364 136
rect 4447 136 4493 144
rect 4807 136 4833 144
rect 4907 136 4953 144
rect 4216 116 4364 124
rect 4427 116 4573 124
rect 4627 116 4693 124
rect 4416 104 4424 113
rect 4116 96 4424 104
rect 727 76 973 84
rect 4107 76 4653 84
rect 2087 36 2713 44
rect 2307 16 2593 24
rect 2687 16 2873 24
rect 5047 16 5113 24
use INVX1  _927_
timestamp 0
transform -1 0 4330 0 1 3610
box -6 -8 66 248
use NOR2X1  _928_
timestamp 0
transform 1 0 3990 0 1 3610
box -6 -8 86 248
use NAND2X1  _929_
timestamp 0
transform 1 0 4850 0 -1 3610
box -6 -8 86 248
use INVX1  _930_
timestamp 0
transform 1 0 4950 0 -1 3610
box -6 -8 66 248
use INVX1  _931_
timestamp 0
transform 1 0 4190 0 1 3610
box -6 -8 66 248
use INVX2  _932_
timestamp 0
transform -1 0 2830 0 1 3130
box -6 -8 66 248
use NOR2X1  _933_
timestamp 0
transform 1 0 4430 0 1 3610
box -6 -8 86 248
use NAND2X1  _934_
timestamp 0
transform 1 0 4350 0 1 3610
box -6 -8 86 248
use INVX1  _935_
timestamp 0
transform 1 0 4730 0 1 4090
box -6 -8 66 248
use NOR2X1  _936_
timestamp 0
transform -1 0 4390 0 -1 4090
box -6 -8 86 248
use AOI21X1  _937_
timestamp 0
transform 1 0 4390 0 -1 4090
box -6 -8 106 248
use NOR2X1  _938_
timestamp 0
transform -1 0 4850 0 -1 4570
box -6 -8 86 248
use OAI21X1  _939_
timestamp 0
transform -1 0 4750 0 -1 4570
box -6 -8 106 248
use INVX1  _940_
timestamp 0
transform -1 0 4650 0 -1 4090
box -6 -8 66 248
use INVX4  _941_
timestamp 0
transform -1 0 4910 0 1 3610
box -6 -8 86 248
use OAI21X1  _942_
timestamp 0
transform 1 0 4090 0 1 3610
box -6 -8 106 248
use INVX1  _943_
timestamp 0
transform 1 0 4730 0 -1 4090
box -6 -8 66 248
use NOR2X1  _944_
timestamp 0
transform 1 0 4770 0 -1 3610
box -6 -8 86 248
use INVX1  _945_
timestamp 0
transform -1 0 4770 0 -1 3610
box -6 -8 66 248
use INVX1  _946_
timestamp 0
transform 1 0 4970 0 -1 4570
box -6 -8 66 248
use OAI21X1  _947_
timestamp 0
transform 1 0 4490 0 -1 4090
box -6 -8 106 248
use OAI21X1  _948_
timestamp 0
transform 1 0 4630 0 1 3610
box -6 -8 106 248
use AOI22X1  _949_
timestamp 0
transform 1 0 4510 0 1 3610
box -6 -8 126 248
use NAND2X1  _950_
timestamp 0
transform 1 0 4570 0 -1 4570
box -6 -8 86 248
use OAI21X1  _951_
timestamp 0
transform -1 0 4610 0 1 4090
box -6 -8 106 248
use OAI21X1  _952_
timestamp 0
transform -1 0 4510 0 1 4090
box -6 -8 106 248
use NAND2X1  _953_
timestamp 0
transform 1 0 4230 0 -1 4090
box -6 -8 86 248
use NOR2X1  _954_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 86 248
use NOR2X1  _955_
timestamp 0
transform 1 0 4650 0 -1 4090
box -6 -8 86 248
use OAI22X1  _956_
timestamp 0
transform -1 0 4730 0 1 4090
box -6 -8 126 248
use OR2X2  _957_
timestamp 0
transform -1 0 4410 0 1 4090
box -6 -8 106 248
use INVX1  _958_
timestamp 0
transform 1 0 4930 0 1 4090
box -6 -8 66 248
use AOI22X1  _959_
timestamp 0
transform -1 0 4910 0 1 4090
box -6 -8 126 248
use NAND3X1  _960_
timestamp 0
transform 1 0 4730 0 1 3610
box -6 -8 106 248
use AND2X2  _961_
timestamp 0
transform 1 0 4930 0 1 3610
box -6 -8 106 248
use OAI21X1  _962_
timestamp 0
transform 1 0 4890 0 -1 4090
box -6 -8 106 248
use INVX1  _963_
timestamp 0
transform 1 0 5030 0 -1 4570
box -6 -8 66 248
use INVX1  _964_
timestamp 0
transform 1 0 3510 0 -1 4570
box -6 -8 66 248
use NAND2X1  _965_
timestamp 0
transform -1 0 3490 0 -1 4090
box -6 -8 86 248
use OAI21X1  _966_
timestamp 0
transform -1 0 3590 0 -1 4090
box -6 -8 106 248
use INVX1  _967_
timestamp 0
transform -1 0 4130 0 -1 4090
box -6 -8 66 248
use NAND2X1  _968_
timestamp 0
transform 1 0 4170 0 -1 3610
box -6 -8 86 248
use OAI21X1  _969_
timestamp 0
transform 1 0 4070 0 -1 3610
box -6 -8 106 248
use INVX1  _970_
timestamp 0
transform 1 0 2910 0 -1 4570
box -6 -8 66 248
use NAND2X1  _971_
timestamp 0
transform -1 0 3790 0 1 4090
box -6 -8 86 248
use OAI21X1  _972_
timestamp 0
transform -1 0 3890 0 1 4090
box -6 -8 106 248
use INVX1  _973_
timestamp 0
transform 1 0 2730 0 1 4570
box -6 -8 66 248
use NAND2X1  _974_
timestamp 0
transform 1 0 2470 0 1 4090
box -6 -8 86 248
use OAI21X1  _975_
timestamp 0
transform -1 0 2650 0 1 4090
box -6 -8 106 248
use INVX1  _976_
timestamp 0
transform 1 0 2450 0 -1 4090
box -6 -8 66 248
use NAND2X1  _977_
timestamp 0
transform 1 0 2670 0 1 3610
box -6 -8 86 248
use OAI21X1  _978_
timestamp 0
transform -1 0 2850 0 1 3610
box -6 -8 106 248
use INVX1  _979_
timestamp 0
transform 1 0 2770 0 -1 4570
box -6 -8 66 248
use NAND2X1  _980_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 86 248
use OAI21X1  _981_
timestamp 0
transform -1 0 3090 0 -1 4570
box -6 -8 106 248
use INVX1  _982_
timestamp 0
transform 1 0 3170 0 -1 4090
box -6 -8 66 248
use NAND2X1  _983_
timestamp 0
transform 1 0 2990 0 -1 4090
box -6 -8 86 248
use OAI21X1  _984_
timestamp 0
transform -1 0 3170 0 -1 4090
box -6 -8 106 248
use INVX4  _985_
timestamp 0
transform -1 0 2670 0 1 2650
box -6 -8 86 248
use NAND2X1  _986_
timestamp 0
transform 1 0 3550 0 -1 3610
box -6 -8 86 248
use OAI21X1  _987_
timestamp 0
transform 1 0 3450 0 -1 3610
box -6 -8 106 248
use INVX1  _988_
timestamp 0
transform 1 0 2490 0 1 3610
box -6 -8 66 248
use INVX1  _989_
timestamp 0
transform -1 0 3110 0 1 2170
box -6 -8 66 248
use INVX2  _990_
timestamp 0
transform -1 0 2430 0 -1 1690
box -6 -8 66 248
use NOR2X1  _991_
timestamp 0
transform 1 0 3190 0 1 2170
box -6 -8 86 248
use AND2X2  _992_
timestamp 0
transform 1 0 2570 0 1 2170
box -6 -8 106 248
use NAND2X1  _993_
timestamp 0
transform 1 0 3110 0 1 2170
box -6 -8 86 248
use NAND2X1  _994_
timestamp 0
transform 1 0 4430 0 -1 3610
box -6 -8 86 248
use NAND2X1  _995_
timestamp 0
transform -1 0 4330 0 -1 3130
box -6 -8 86 248
use OR2X2  _996_
timestamp 0
transform -1 0 5030 0 1 3130
box -6 -8 106 248
use NAND2X1  _997_
timestamp 0
transform 1 0 4550 0 1 3130
box -6 -8 86 248
use AND2X2  _998_
timestamp 0
transform 1 0 5030 0 1 3130
box -6 -8 106 248
use OAI21X1  _999_
timestamp 0
transform 1 0 4730 0 1 3130
box -6 -8 106 248
use NAND2X1  _1000_
timestamp 0
transform -1 0 4530 0 1 2650
box -6 -8 86 248
use INVX1  _1001_
timestamp 0
transform -1 0 4430 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1002_
timestamp 0
transform 1 0 4170 0 1 1690
box -6 -8 86 248
use OR2X2  _1003_
timestamp 0
transform 1 0 4890 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1004_
timestamp 0
transform -1 0 4250 0 -1 3130
box -6 -8 126 248
use INVX1  _1005_
timestamp 0
transform -1 0 4930 0 -1 2650
box -6 -8 66 248
use NAND3X1  _1006_
timestamp 0
transform -1 0 4750 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1007_
timestamp 0
transform 1 0 4790 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1008_
timestamp 0
transform -1 0 4530 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1009_
timestamp 0
transform 1 0 4630 0 1 2650
box -6 -8 106 248
use INVX1  _1010_
timestamp 0
transform 1 0 3570 0 1 2650
box -6 -8 66 248
use NAND2X1  _1011_
timestamp 0
transform -1 0 2770 0 1 2170
box -6 -8 86 248
use INVX2  _1012_
timestamp 0
transform -1 0 2110 0 1 1690
box -6 -8 66 248
use NAND2X1  _1013_
timestamp 0
transform 1 0 3530 0 1 1690
box -6 -8 86 248
use OAI21X1  _1014_
timestamp 0
transform 1 0 3430 0 1 1690
box -6 -8 106 248
use OAI21X1  _1015_
timestamp 0
transform -1 0 3570 0 1 2650
box -6 -8 106 248
use AOI21X1  _1016_
timestamp 0
transform -1 0 4630 0 1 2650
box -6 -8 106 248
use OAI21X1  _1017_
timestamp 0
transform 1 0 4030 0 1 2650
box -6 -8 106 248
use OAI21X1  _1018_
timestamp 0
transform 1 0 4930 0 -1 2650
box -6 -8 106 248
use AND2X2  _1019_
timestamp 0
transform 1 0 3970 0 1 1210
box -6 -8 106 248
use NAND3X1  _1020_
timestamp 0
transform 1 0 4310 0 1 1210
box -6 -8 106 248
use AOI22X1  _1021_
timestamp 0
transform 1 0 3950 0 1 1690
box -6 -8 126 248
use INVX1  _1022_
timestamp 0
transform -1 0 4670 0 1 1690
box -6 -8 66 248
use NAND2X1  _1023_
timestamp 0
transform -1 0 4350 0 1 1690
box -6 -8 86 248
use INVX1  _1024_
timestamp 0
transform 1 0 4450 0 1 1690
box -6 -8 66 248
use NAND3X1  _1025_
timestamp 0
transform 1 0 4970 0 1 1690
box -6 -8 106 248
use NAND2X1  _1026_
timestamp 0
transform -1 0 3950 0 1 1690
box -6 -8 86 248
use NOR2X1  _1027_
timestamp 0
transform -1 0 4170 0 1 1690
box -6 -8 86 248
use OAI21X1  _1028_
timestamp 0
transform 1 0 4770 0 1 1690
box -6 -8 106 248
use NAND3X1  _1029_
timestamp 0
transform 1 0 5010 0 1 2170
box -6 -8 106 248
use AOI21X1  _1030_
timestamp 0
transform -1 0 4650 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1031_
timestamp 0
transform 1 0 4670 0 1 1690
box -6 -8 106 248
use NAND3X1  _1032_
timestamp 0
transform -1 0 4970 0 1 1690
box -6 -8 106 248
use NAND3X1  _1033_
timestamp 0
transform -1 0 4850 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1034_
timestamp 0
transform -1 0 2950 0 -1 2170
box -6 -8 86 248
use INVX1  _1035_
timestamp 0
transform 1 0 2950 0 -1 2170
box -6 -8 66 248
use AND2X2  _1036_
timestamp 0
transform 1 0 3010 0 1 1690
box -6 -8 106 248
use NAND2X1  _1037_
timestamp 0
transform 1 0 3110 0 -1 2170
box -6 -8 86 248
use INVX1  _1038_
timestamp 0
transform -1 0 2850 0 1 2170
box -6 -8 66 248
use OAI21X1  _1039_
timestamp 0
transform 1 0 2850 0 1 2170
box -6 -8 106 248
use NAND3X1  _1040_
timestamp 0
transform 1 0 3010 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1041_
timestamp 0
transform -1 0 2850 0 -1 2170
box -6 -8 106 248
use INVX1  _1042_
timestamp 0
transform 1 0 3410 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1043_
timestamp 0
transform -1 0 3310 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1044_
timestamp 0
transform 1 0 3190 0 -1 2170
box -6 -8 106 248
use AND2X2  _1045_
timestamp 0
transform 1 0 3370 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1046_
timestamp 0
transform -1 0 4670 0 1 2170
box -6 -8 106 248
use AOI21X1  _1047_
timestamp 0
transform 1 0 4850 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1048_
timestamp 0
transform 1 0 4990 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1049_
timestamp 0
transform -1 0 3370 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1050_
timestamp 0
transform -1 0 4910 0 1 2170
box -6 -8 106 248
use NAND3X1  _1051_
timestamp 0
transform -1 0 4550 0 1 2170
box -6 -8 106 248
use AOI21X1  _1052_
timestamp 0
transform -1 0 4450 0 1 2170
box -6 -8 106 248
use OAI21X1  _1053_
timestamp 0
transform 1 0 4250 0 1 2170
box -6 -8 106 248
use AOI21X1  _1054_
timestamp 0
transform 1 0 4970 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1055_
timestamp 0
transform 1 0 4350 0 1 1690
box -6 -8 106 248
use AND2X2  _1056_
timestamp 0
transform 1 0 2610 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1057_
timestamp 0
transform -1 0 3650 0 -1 1210
box -6 -8 86 248
use INVX1  _1058_
timestamp 0
transform -1 0 2790 0 -1 1210
box -6 -8 66 248
use INVX2  _1059_
timestamp 0
transform 1 0 1990 0 1 1690
box -6 -8 66 248
use NAND2X1  _1060_
timestamp 0
transform -1 0 2990 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1061_
timestamp 0
transform 1 0 2810 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1062_
timestamp 0
transform 1 0 4230 0 1 1210
box -6 -8 86 248
use INVX1  _1063_
timestamp 0
transform 1 0 4170 0 1 1210
box -6 -8 66 248
use NAND3X1  _1064_
timestamp 0
transform -1 0 3970 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1065_
timestamp 0
transform -1 0 3890 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1066_
timestamp 0
transform -1 0 3970 0 -1 1690
box -6 -8 86 248
use AOI22X1  _1067_
timestamp 0
transform 1 0 3830 0 1 1210
box -6 -8 126 248
use OAI21X1  _1068_
timestamp 0
transform 1 0 4070 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1069_
timestamp 0
transform 1 0 4590 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1070_
timestamp 0
transform -1 0 4610 0 1 1690
box -6 -8 106 248
use OAI21X1  _1071_
timestamp 0
transform 1 0 4070 0 1 1210
box -6 -8 106 248
use NAND3X1  _1072_
timestamp 0
transform -1 0 3750 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1073_
timestamp 0
transform 1 0 4430 0 1 1210
box -6 -8 106 248
use NAND2X1  _1074_
timestamp 0
transform 1 0 3130 0 -1 1690
box -6 -8 86 248
use INVX1  _1075_
timestamp 0
transform 1 0 3390 0 -1 1690
box -6 -8 66 248
use AND2X2  _1076_
timestamp 0
transform 1 0 2430 0 -1 1690
box -6 -8 106 248
use AND2X2  _1077_
timestamp 0
transform 1 0 2550 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1078_
timestamp 0
transform 1 0 2830 0 -1 1690
box -6 -8 86 248
use INVX2  _1079_
timestamp 0
transform 1 0 2750 0 1 1690
box -6 -8 66 248
use NAND2X1  _1080_
timestamp 0
transform 1 0 3350 0 1 1690
box -6 -8 86 248
use OAI21X1  _1081_
timestamp 0
transform 1 0 3590 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1082_
timestamp 0
transform 1 0 3690 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1083_
timestamp 0
transform -1 0 2830 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1084_
timestamp 0
transform -1 0 3010 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1085_
timestamp 0
transform -1 0 3130 0 -1 1690
box -6 -8 106 248
use AND2X2  _1086_
timestamp 0
transform 1 0 3730 0 1 1210
box -6 -8 106 248
use OAI21X1  _1087_
timestamp 0
transform -1 0 5130 0 1 1210
box -6 -8 106 248
use NAND3X1  _1088_
timestamp 0
transform 1 0 4530 0 1 1210
box -6 -8 106 248
use NAND3X1  _1089_
timestamp 0
transform 1 0 4470 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1090_
timestamp 0
transform -1 0 3730 0 1 1210
box -6 -8 86 248
use NAND3X1  _1091_
timestamp 0
transform 1 0 4830 0 1 1210
box -6 -8 106 248
use NAND3X1  _1092_
timestamp 0
transform -1 0 5030 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1093_
timestamp 0
transform -1 0 5090 0 1 4090
box -6 -8 106 248
use NAND3X1  _1094_
timestamp 0
transform 1 0 4930 0 1 1210
box -6 -8 106 248
use OAI21X1  _1095_
timestamp 0
transform 1 0 4990 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1096_
timestamp 0
transform -1 0 5130 0 -1 1690
box -6 -8 106 248
use INVX4  _1097_
timestamp 0
transform -1 0 1990 0 1 1690
box -6 -8 86 248
use NOR2X1  _1098_
timestamp 0
transform 1 0 3710 0 1 1690
box -6 -8 86 248
use OAI21X1  _1099_
timestamp 0
transform 1 0 3610 0 1 1690
box -6 -8 106 248
use NAND2X1  _1100_
timestamp 0
transform -1 0 4070 0 -1 1690
box -6 -8 86 248
use OR2X2  _1101_
timestamp 0
transform 1 0 4070 0 -1 1690
box -6 -8 106 248
use AND2X2  _1102_
timestamp 0
transform 1 0 4370 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1103_
timestamp 0
transform 1 0 4790 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1104_
timestamp 0
transform -1 0 5050 0 1 730
box -6 -8 106 248
use AOI21X1  _1105_
timestamp 0
transform -1 0 4630 0 1 4570
box -6 -8 106 248
use NAND2X1  _1106_
timestamp 0
transform -1 0 4370 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1107_
timestamp 0
transform 1 0 4690 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1108_
timestamp 0
transform -1 0 4670 0 -1 2170
box -6 -8 106 248
use INVX1  _1109_
timestamp 0
transform -1 0 4230 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1110_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 106 248
use AOI21X1  _1111_
timestamp 0
transform 1 0 4630 0 1 1210
box -6 -8 106 248
use OAI21X1  _1112_
timestamp 0
transform -1 0 3870 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1113_
timestamp 0
transform 1 0 3290 0 -1 1210
box -6 -8 106 248
use AOI22X1  _1114_
timestamp 0
transform -1 0 3290 0 -1 1210
box -6 -8 126 248
use INVX1  _1115_
timestamp 0
transform 1 0 3310 0 1 730
box -6 -8 66 248
use NAND2X1  _1116_
timestamp 0
transform 1 0 3490 0 -1 1210
box -6 -8 86 248
use INVX1  _1117_
timestamp 0
transform 1 0 3850 0 -1 730
box -6 -8 66 248
use NAND3X1  _1118_
timestamp 0
transform 1 0 3670 0 1 730
box -6 -8 106 248
use NAND2X1  _1119_
timestamp 0
transform 1 0 3090 0 -1 1210
box -6 -8 86 248
use NOR2X1  _1120_
timestamp 0
transform 1 0 3010 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1121_
timestamp 0
transform 1 0 3570 0 1 730
box -6 -8 106 248
use AOI21X1  _1122_
timestamp 0
transform 1 0 4210 0 1 730
box -6 -8 106 248
use OAI21X1  _1123_
timestamp 0
transform -1 0 3570 0 1 730
box -6 -8 106 248
use NAND3X1  _1124_
timestamp 0
transform 1 0 3790 0 1 730
box -6 -8 106 248
use AOI22X1  _1125_
timestamp 0
transform -1 0 4010 0 1 730
box -6 -8 126 248
use NAND2X1  _1126_
timestamp 0
transform -1 0 3110 0 1 1210
box -6 -8 86 248
use INVX1  _1127_
timestamp 0
transform 1 0 3430 0 1 1210
box -6 -8 66 248
use AND2X2  _1128_
timestamp 0
transform -1 0 3010 0 1 1690
box -6 -8 106 248
use AND2X2  _1129_
timestamp 0
transform -1 0 3350 0 1 1690
box -6 -8 106 248
use NAND2X1  _1130_
timestamp 0
transform -1 0 3390 0 -1 1690
box -6 -8 86 248
use AOI22X1  _1131_
timestamp 0
transform -1 0 3250 0 1 1690
box -6 -8 126 248
use INVX1  _1132_
timestamp 0
transform 1 0 3490 0 1 1210
box -6 -8 66 248
use NAND3X1  _1133_
timestamp 0
transform 1 0 3550 0 1 1210
box -6 -8 106 248
use INVX1  _1134_
timestamp 0
transform -1 0 1890 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1135_
timestamp 0
transform 1 0 2930 0 1 1210
box -6 -8 106 248
use OAI21X1  _1136_
timestamp 0
transform 1 0 3210 0 1 1210
box -6 -8 106 248
use NAND3X1  _1137_
timestamp 0
transform 1 0 3110 0 1 1210
box -6 -8 106 248
use AND2X2  _1138_
timestamp 0
transform 1 0 4090 0 -1 730
box -6 -8 106 248
use OAI21X1  _1139_
timestamp 0
transform 1 0 4410 0 -1 730
box -6 -8 106 248
use AOI21X1  _1140_
timestamp 0
transform 1 0 3970 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1141_
timestamp 0
transform 1 0 4010 0 1 730
box -6 -8 106 248
use NAND3X1  _1142_
timestamp 0
transform 1 0 4110 0 1 730
box -6 -8 106 248
use NAND2X1  _1143_
timestamp 0
transform -1 0 4090 0 -1 730
box -6 -8 86 248
use NAND3X1  _1144_
timestamp 0
transform 1 0 4610 0 -1 730
box -6 -8 106 248
use NAND3X1  _1145_
timestamp 0
transform 1 0 4670 0 1 250
box -6 -8 106 248
use OAI21X1  _1146_
timestamp 0
transform 1 0 4690 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1147_
timestamp 0
transform 1 0 4730 0 -1 730
box -6 -8 106 248
use OAI21X1  _1148_
timestamp 0
transform 1 0 4510 0 -1 730
box -6 -8 106 248
use NAND3X1  _1149_
timestamp 0
transform 1 0 4930 0 -1 730
box -6 -8 106 248
use NAND2X1  _1150_
timestamp 0
transform -1 0 3550 0 -1 2170
box -6 -8 86 248
use INVX1  _1151_
timestamp 0
transform 1 0 4470 0 -1 250
box -6 -8 66 248
use AOI22X1  _1152_
timestamp 0
transform 1 0 3450 0 -1 1690
box -6 -8 126 248
use INVX1  _1153_
timestamp 0
transform 1 0 4310 0 1 250
box -6 -8 66 248
use OAI21X1  _1154_
timestamp 0
transform 1 0 4370 0 1 250
box -6 -8 106 248
use NOR2X1  _1155_
timestamp 0
transform -1 0 4110 0 1 250
box -6 -8 86 248
use NAND2X1  _1156_
timestamp 0
transform -1 0 4070 0 -1 250
box -6 -8 86 248
use NAND3X1  _1157_
timestamp 0
transform -1 0 4450 0 -1 250
box -6 -8 106 248
use NAND2X1  _1158_
timestamp 0
transform 1 0 4230 0 1 250
box -6 -8 86 248
use OAI21X1  _1159_
timestamp 0
transform -1 0 4210 0 1 250
box -6 -8 106 248
use NAND3X1  _1160_
timestamp 0
transform 1 0 4170 0 -1 250
box -6 -8 106 248
use NAND2X1  _1161_
timestamp 0
transform 1 0 4270 0 -1 250
box -6 -8 86 248
use NAND3X1  _1162_
timestamp 0
transform -1 0 4890 0 1 250
box -6 -8 106 248
use AOI21X1  _1163_
timestamp 0
transform -1 0 4930 0 -1 730
box -6 -8 106 248
use AOI21X1  _1164_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 106 248
use NAND3X1  _1165_
timestamp 0
transform -1 0 4170 0 -1 250
box -6 -8 106 248
use NAND3X1  _1166_
timestamp 0
transform 1 0 4550 0 -1 250
box -6 -8 106 248
use NAND2X1  _1167_
timestamp 0
transform 1 0 4650 0 -1 250
box -6 -8 86 248
use OAI21X1  _1168_
timestamp 0
transform -1 0 4930 0 -1 250
box -6 -8 106 248
use AOI21X1  _1169_
timestamp 0
transform -1 0 4830 0 1 730
box -6 -8 106 248
use AOI21X1  _1170_
timestamp 0
transform -1 0 4910 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1171_
timestamp 0
transform 1 0 4930 0 -1 250
box -6 -8 106 248
use NAND3X1  _1172_
timestamp 0
transform 1 0 4890 0 1 250
box -6 -8 106 248
use AOI21X1  _1173_
timestamp 0
transform 1 0 4990 0 1 250
box -6 -8 106 248
use OAI21X1  _1174_
timestamp 0
transform -1 0 4350 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1175_
timestamp 0
transform -1 0 4950 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1176_
timestamp 0
transform 1 0 4830 0 1 730
box -6 -8 106 248
use NAND3X1  _1177_
timestamp 0
transform -1 0 4630 0 1 730
box -6 -8 106 248
use AOI21X1  _1178_
timestamp 0
transform -1 0 4230 0 -1 2170
box -6 -8 106 248
use INVX1  _1179_
timestamp 0
transform 1 0 3830 0 -1 2170
box -6 -8 66 248
use INVX1  _1180_
timestamp 0
transform 1 0 4010 0 -1 2650
box -6 -8 66 248
use NOR2X1  _1181_
timestamp 0
transform 1 0 4830 0 1 3130
box -6 -8 86 248
use INVX1  _1182_
timestamp 0
transform -1 0 4670 0 -1 3130
box -6 -8 66 248
use INVX1  _1183_
timestamp 0
transform 1 0 4330 0 -1 3130
box -6 -8 66 248
use OAI21X1  _1184_
timestamp 0
transform 1 0 4390 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1185_
timestamp 0
transform 1 0 4670 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1186_
timestamp 0
transform 1 0 4770 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1187_
timestamp 0
transform 1 0 4930 0 1 2650
box -6 -8 106 248
use AOI21X1  _1188_
timestamp 0
transform -1 0 4830 0 1 2650
box -6 -8 106 248
use AND2X2  _1189_
timestamp 0
transform 1 0 3410 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1190_
timestamp 0
transform 1 0 4830 0 1 2650
box -6 -8 106 248
use AOI21X1  _1191_
timestamp 0
transform 1 0 4230 0 1 2650
box -6 -8 106 248
use OAI21X1  _1192_
timestamp 0
transform 1 0 4910 0 1 2170
box -6 -8 106 248
use NAND3X1  _1193_
timestamp 0
transform -1 0 4790 0 1 2170
box -6 -8 106 248
use NAND3X1  _1194_
timestamp 0
transform -1 0 4370 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1195_
timestamp 0
transform 1 0 4170 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1196_
timestamp 0
transform -1 0 4690 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1197_
timestamp 0
transform 1 0 4910 0 -1 1690
box -6 -8 106 248
use AOI22X1  _1198_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 126 248
use NAND3X1  _1199_
timestamp 0
transform 1 0 4430 0 1 730
box -6 -8 106 248
use OAI21X1  _1200_
timestamp 0
transform -1 0 4450 0 -1 1210
box -6 -8 106 248
use AOI21X1  _1201_
timestamp 0
transform -1 0 4290 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1202_
timestamp 0
transform -1 0 4230 0 1 2650
box -6 -8 106 248
use NAND3X1  _1203_
timestamp 0
transform -1 0 4590 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1204_
timestamp 0
transform 1 0 3430 0 1 3130
box -6 -8 86 248
use NAND2X1  _1205_
timestamp 0
transform 1 0 4350 0 -1 3610
box -6 -8 86 248
use AOI22X1  _1206_
timestamp 0
transform 1 0 3870 0 1 3130
box -6 -8 126 248
use OAI22X1  _1207_
timestamp 0
transform -1 0 4470 0 1 3130
box -6 -8 126 248
use OAI21X1  _1208_
timestamp 0
transform -1 0 4730 0 1 3130
box -6 -8 106 248
use NAND3X1  _1209_
timestamp 0
transform -1 0 4030 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1210_
timestamp 0
transform -1 0 4130 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1211_
timestamp 0
transform 1 0 3810 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1212_
timestamp 0
transform -1 0 4030 0 1 2650
box -6 -8 106 248
use NAND3X1  _1213_
timestamp 0
transform -1 0 3830 0 1 2650
box -6 -8 106 248
use INVX1  _1214_
timestamp 0
transform -1 0 3570 0 -1 2650
box -6 -8 66 248
use AOI22X1  _1215_
timestamp 0
transform 1 0 4330 0 1 2650
box -6 -8 126 248
use OAI21X1  _1216_
timestamp 0
transform -1 0 3890 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1217_
timestamp 0
transform -1 0 3790 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1218_
timestamp 0
transform -1 0 4550 0 -1 2170
box -6 -8 106 248
use NOR3X1  _1219_
timestamp 0
transform -1 0 3970 0 1 2170
box -6 -8 186 248
use INVX1  _1220_
timestamp 0
transform -1 0 3630 0 -1 3130
box -6 -8 66 248
use NAND3X1  _1221_
timestamp 0
transform -1 0 3550 0 -1 3130
box -6 -8 106 248
use INVX1  _1222_
timestamp 0
transform -1 0 4230 0 1 3130
box -6 -8 66 248
use NOR2X1  _1223_
timestamp 0
transform 1 0 4470 0 1 3130
box -6 -8 86 248
use NOR2X1  _1224_
timestamp 0
transform 1 0 4090 0 1 3130
box -6 -8 86 248
use NAND2X1  _1225_
timestamp 0
transform -1 0 4070 0 1 3130
box -6 -8 86 248
use NAND2X1  _1226_
timestamp 0
transform 1 0 3790 0 1 3130
box -6 -8 86 248
use NOR2X1  _1227_
timestamp 0
transform 1 0 3710 0 1 3130
box -6 -8 86 248
use OAI21X1  _1228_
timestamp 0
transform 1 0 4250 0 1 3130
box -6 -8 106 248
use NAND3X1  _1229_
timestamp 0
transform -1 0 3710 0 1 3130
box -6 -8 106 248
use INVX1  _1230_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 66 248
use INVX1  _1231_
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 66 248
use OAI21X1  _1232_
timestamp 0
transform -1 0 3750 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1233_
timestamp 0
transform 1 0 3350 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1234_
timestamp 0
transform -1 0 3930 0 1 2650
box -6 -8 106 248
use NOR3X1  _1235_
timestamp 0
transform -1 0 3450 0 1 2650
box -6 -8 186 248
use OAI21X1  _1236_
timestamp 0
transform 1 0 3910 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1237_
timestamp 0
transform -1 0 4170 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1238_
timestamp 0
transform -1 0 3670 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1239_
timestamp 0
transform 1 0 3210 0 -1 2650
box -6 -8 106 248
use INVX1  _1240_
timestamp 0
transform 1 0 3330 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1241_
timestamp 0
transform -1 0 3790 0 1 2170
box -6 -8 106 248
use AOI21X1  _1242_
timestamp 0
transform 1 0 3590 0 1 2170
box -6 -8 106 248
use OAI21X1  _1243_
timestamp 0
transform -1 0 3990 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1244_
timestamp 0
transform -1 0 4430 0 1 730
box -6 -8 106 248
use NAND2X1  _1245_
timestamp 0
transform -1 0 3990 0 -1 250
box -6 -8 86 248
use OAI21X1  _1246_
timestamp 0
transform 1 0 4730 0 -1 250
box -6 -8 106 248
use NAND2X1  _1247_
timestamp 0
transform -1 0 3310 0 1 730
box -6 -8 86 248
use INVX1  _1248_
timestamp 0
transform 1 0 3650 0 -1 250
box -6 -8 66 248
use NOR2X1  _1249_
timestamp 0
transform 1 0 3930 0 1 250
box -6 -8 86 248
use OAI21X1  _1250_
timestamp 0
transform 1 0 3310 0 1 1210
box -6 -8 106 248
use NAND2X1  _1251_
timestamp 0
transform 1 0 3850 0 1 250
box -6 -8 86 248
use OR2X2  _1252_
timestamp 0
transform -1 0 3910 0 -1 250
box -6 -8 106 248
use NAND3X1  _1253_
timestamp 0
transform 1 0 3710 0 -1 250
box -6 -8 106 248
use AND2X2  _1254_
timestamp 0
transform -1 0 3430 0 -1 250
box -6 -8 106 248
use NOR2X1  _1255_
timestamp 0
transform -1 0 3530 0 -1 250
box -6 -8 86 248
use OAI21X1  _1256_
timestamp 0
transform -1 0 3330 0 -1 250
box -6 -8 106 248
use NAND2X1  _1257_
timestamp 0
transform 1 0 3150 0 -1 250
box -6 -8 86 248
use AOI21X1  _1258_
timestamp 0
transform -1 0 4290 0 -1 730
box -6 -8 106 248
use NAND2X1  _1259_
timestamp 0
transform 1 0 1970 0 1 1210
box -6 -8 86 248
use AND2X2  _1260_
timestamp 0
transform 1 0 2190 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1261_
timestamp 0
transform -1 0 2550 0 1 1210
box -6 -8 106 248
use AND2X2  _1262_
timestamp 0
transform 1 0 2050 0 1 1210
box -6 -8 106 248
use OAI21X1  _1263_
timestamp 0
transform -1 0 2350 0 1 1210
box -6 -8 106 248
use NAND3X1  _1264_
timestamp 0
transform 1 0 2350 0 1 1210
box -6 -8 106 248
use INVX1  _1265_
timestamp 0
transform -1 0 2130 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1266_
timestamp 0
transform -1 0 2230 0 1 1210
box -6 -8 86 248
use AOI22X1  _1267_
timestamp 0
transform 1 0 1990 0 -1 1690
box -6 -8 126 248
use INVX1  _1268_
timestamp 0
transform 1 0 2010 0 -1 1210
box -6 -8 66 248
use NAND3X1  _1269_
timestamp 0
transform 1 0 2130 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1270_
timestamp 0
transform 1 0 2330 0 1 730
box -6 -8 86 248
use AOI21X1  _1271_
timestamp 0
transform -1 0 3230 0 1 730
box -6 -8 106 248
use NAND2X1  _1272_
timestamp 0
transform -1 0 2310 0 -1 1210
box -6 -8 86 248
use INVX1  _1273_
timestamp 0
transform -1 0 1570 0 1 730
box -6 -8 66 248
use AOI22X1  _1274_
timestamp 0
transform -1 0 2610 0 -1 1210
box -6 -8 126 248
use AOI21X1  _1275_
timestamp 0
transform 1 0 1790 0 1 730
box -6 -8 106 248
use NAND2X1  _1276_
timestamp 0
transform 1 0 2150 0 1 730
box -6 -8 86 248
use OAI21X1  _1277_
timestamp 0
transform -1 0 3470 0 1 730
box -6 -8 106 248
use INVX1  _1278_
timestamp 0
transform 1 0 2310 0 -1 1210
box -6 -8 66 248
use OAI21X1  _1279_
timestamp 0
transform -1 0 2490 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1280_
timestamp 0
transform 1 0 2490 0 1 730
box -6 -8 86 248
use NAND3X1  _1281_
timestamp 0
transform 1 0 2670 0 1 730
box -6 -8 106 248
use AND2X2  _1282_
timestamp 0
transform -1 0 2410 0 -1 730
box -6 -8 106 248
use NAND2X1  _1283_
timestamp 0
transform -1 0 2150 0 1 730
box -6 -8 86 248
use NAND2X1  _1284_
timestamp 0
transform -1 0 2490 0 1 730
box -6 -8 86 248
use NAND3X1  _1285_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 106 248
use NAND3X1  _1286_
timestamp 0
transform 1 0 3230 0 1 250
box -6 -8 106 248
use OAI21X1  _1287_
timestamp 0
transform -1 0 4390 0 -1 730
box -6 -8 106 248
use AOI22X1  _1288_
timestamp 0
transform 1 0 2410 0 -1 730
box -6 -8 126 248
use AOI21X1  _1289_
timestamp 0
transform -1 0 2670 0 1 730
box -6 -8 106 248
use OAI21X1  _1290_
timestamp 0
transform 1 0 2710 0 1 250
box -6 -8 106 248
use NAND3X1  _1291_
timestamp 0
transform 1 0 3430 0 1 250
box -6 -8 106 248
use AND2X2  _1292_
timestamp 0
transform -1 0 3010 0 -1 250
box -6 -8 106 248
use NAND3X1  _1293_
timestamp 0
transform -1 0 3210 0 1 250
box -6 -8 106 248
use OAI21X1  _1294_
timestamp 0
transform 1 0 2690 0 -1 250
box -6 -8 106 248
use NAND3X1  _1295_
timestamp 0
transform 1 0 3010 0 1 250
box -6 -8 106 248
use NAND3X1  _1296_
timestamp 0
transform -1 0 3550 0 -1 730
box -6 -8 106 248
use AOI21X1  _1297_
timestamp 0
transform -1 0 4570 0 1 250
box -6 -8 106 248
use AOI22X1  _1298_
timestamp 0
transform -1 0 3150 0 -1 250
box -6 -8 126 248
use AOI21X1  _1299_
timestamp 0
transform 1 0 3330 0 1 250
box -6 -8 106 248
use OAI21X1  _1300_
timestamp 0
transform 1 0 3530 0 1 250
box -6 -8 106 248
use AOI21X1  _1301_
timestamp 0
transform -1 0 3110 0 1 730
box -6 -8 106 248
use INVX1  _1302_
timestamp 0
transform 1 0 3930 0 -1 730
box -6 -8 66 248
use NAND3X1  _1303_
timestamp 0
transform 1 0 3630 0 1 250
box -6 -8 106 248
use OAI21X1  _1304_
timestamp 0
transform 1 0 3730 0 1 250
box -6 -8 106 248
use AOI21X1  _1305_
timestamp 0
transform -1 0 3750 0 -1 730
box -6 -8 106 248
use OAI21X1  _1306_
timestamp 0
transform -1 0 3010 0 1 730
box -6 -8 106 248
use OAI21X1  _1307_
timestamp 0
transform 1 0 4630 0 1 730
box -6 -8 106 248
use NAND3X1  _1308_
timestamp 0
transform 1 0 3750 0 -1 730
box -6 -8 106 248
use NAND3X1  _1309_
timestamp 0
transform -1 0 3330 0 -1 730
box -6 -8 106 248
use NAND3X1  _1310_
timestamp 0
transform -1 0 2890 0 1 730
box -6 -8 106 248
use AND2X2  _1311_
timestamp 0
transform -1 0 2750 0 1 1690
box -6 -8 106 248
use NAND2X1  _1312_
timestamp 0
transform 1 0 2490 0 1 1690
box -6 -8 86 248
use NAND3X1  _1313_
timestamp 0
transform -1 0 4350 0 -1 2170
box -6 -8 106 248
use INVX1  _1314_
timestamp 0
transform 1 0 3970 0 1 2170
box -6 -8 66 248
use NAND2X1  _1315_
timestamp 0
transform 1 0 4670 0 -1 2170
box -6 -8 86 248
use NAND3X1  _1316_
timestamp 0
transform -1 0 4450 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1317_
timestamp 0
transform 1 0 4150 0 1 2170
box -6 -8 106 248
use AOI21X1  _1318_
timestamp 0
transform -1 0 4130 0 1 2170
box -6 -8 106 248
use OAI21X1  _1319_
timestamp 0
transform 1 0 3490 0 1 2170
box -6 -8 106 248
use AOI21X1  _1320_
timestamp 0
transform -1 0 3650 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1321_
timestamp 0
transform 1 0 2310 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1322_
timestamp 0
transform 1 0 2390 0 -1 2170
box -6 -8 86 248
use AND2X2  _1323_
timestamp 0
transform 1 0 2470 0 -1 2170
box -6 -8 106 248
use NOR2X1  _1324_
timestamp 0
transform -1 0 1570 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1325_
timestamp 0
transform 1 0 2410 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1326_
timestamp 0
transform -1 0 2590 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1327_
timestamp 0
transform -1 0 3030 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1328_
timestamp 0
transform 1 0 2070 0 1 3610
box -6 -8 106 248
use OAI21X1  _1329_
timestamp 0
transform -1 0 2790 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1330_
timestamp 0
transform 1 0 2590 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1331_
timestamp 0
transform 1 0 2550 0 1 3610
box -6 -8 106 248
use INVX1  _1332_
timestamp 0
transform 1 0 2050 0 -1 3130
box -6 -8 66 248
use INVX1  _1333_
timestamp 0
transform 1 0 1630 0 1 2650
box -6 -8 66 248
use OAI21X1  _1334_
timestamp 0
transform -1 0 2290 0 1 2650
box -6 -8 106 248
use OAI21X1  _1335_
timestamp 0
transform 1 0 1770 0 1 2650
box -6 -8 106 248
use AOI21X1  _1336_
timestamp 0
transform -1 0 3650 0 -1 730
box -6 -8 106 248
use OAI21X1  _1337_
timestamp 0
transform -1 0 3450 0 -1 730
box -6 -8 106 248
use OAI21X1  _1338_
timestamp 0
transform 1 0 3530 0 -1 250
box -6 -8 106 248
use AOI21X1  _1339_
timestamp 0
transform 1 0 2810 0 1 250
box -6 -8 106 248
use OAI21X1  _1340_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 106 248
use NAND2X1  _1341_
timestamp 0
transform -1 0 1210 0 1 730
box -6 -8 86 248
use INVX1  _1342_
timestamp 0
transform 1 0 1350 0 -1 730
box -6 -8 66 248
use NOR2X1  _1343_
timestamp 0
transform -1 0 2630 0 1 1210
box -6 -8 86 248
use OAI21X1  _1344_
timestamp 0
transform -1 0 2010 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1345_
timestamp 0
transform 1 0 1410 0 -1 730
box -6 -8 86 248
use OR2X2  _1346_
timestamp 0
transform -1 0 1770 0 -1 730
box -6 -8 106 248
use NAND3X1  _1347_
timestamp 0
transform 1 0 1490 0 -1 730
box -6 -8 106 248
use AND2X2  _1348_
timestamp 0
transform -1 0 1430 0 1 730
box -6 -8 106 248
use NOR2X1  _1349_
timestamp 0
transform -1 0 1670 0 -1 730
box -6 -8 86 248
use OAI21X1  _1350_
timestamp 0
transform -1 0 1310 0 1 730
box -6 -8 106 248
use NAND2X1  _1351_
timestamp 0
transform 1 0 1510 0 1 250
box -6 -8 86 248
use NOR2X1  _1352_
timestamp 0
transform -1 0 2330 0 1 730
box -6 -8 86 248
use AOI21X1  _1353_
timestamp 0
transform -1 0 2290 0 -1 730
box -6 -8 106 248
use NAND2X1  _1354_
timestamp 0
transform 1 0 1870 0 1 1210
box -6 -8 86 248
use INVX1  _1355_
timestamp 0
transform 1 0 1370 0 -1 1210
box -6 -8 66 248
use AND2X2  _1356_
timestamp 0
transform 1 0 1470 0 -1 1690
box -6 -8 106 248
use AND2X2  _1357_
timestamp 0
transform -1 0 1970 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1358_
timestamp 0
transform 1 0 1570 0 -1 1690
box -6 -8 86 248
use AOI22X1  _1359_
timestamp 0
transform 1 0 1550 0 1 1210
box -6 -8 126 248
use INVX1  _1360_
timestamp 0
transform 1 0 1310 0 -1 1210
box -6 -8 66 248
use AOI21X1  _1361_
timestamp 0
transform 1 0 1430 0 -1 1210
box -6 -8 106 248
use INVX2  _1362_
timestamp 0
transform 1 0 1630 0 1 1690
box -6 -8 66 248
use OAI21X1  _1363_
timestamp 0
transform -1 0 1750 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1364_
timestamp 0
transform -1 0 1870 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1365_
timestamp 0
transform -1 0 1770 0 1 1210
box -6 -8 106 248
use OAI22X1  _1366_
timestamp 0
transform -1 0 1690 0 1 730
box -6 -8 126 248
use NAND3X1  _1367_
timestamp 0
transform -1 0 1870 0 1 1210
box -6 -8 106 248
use NAND3X1  _1368_
timestamp 0
transform 1 0 1550 0 -1 1210
box -6 -8 106 248
use NOR2X1  _1369_
timestamp 0
transform 1 0 1750 0 -1 1210
box -6 -8 86 248
use NAND3X1  _1370_
timestamp 0
transform -1 0 1750 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1371_
timestamp 0
transform -1 0 1770 0 1 730
box -6 -8 86 248
use NOR2X1  _1372_
timestamp 0
transform 1 0 1810 0 1 250
box -6 -8 86 248
use NOR2X1  _1373_
timestamp 0
transform 1 0 1990 0 1 730
box -6 -8 86 248
use OAI21X1  _1374_
timestamp 0
transform -1 0 1990 0 1 730
box -6 -8 106 248
use AOI21X1  _1375_
timestamp 0
transform -1 0 1990 0 -1 730
box -6 -8 106 248
use OAI21X1  _1376_
timestamp 0
transform 1 0 1850 0 -1 250
box -6 -8 106 248
use AND2X2  _1377_
timestamp 0
transform 1 0 1590 0 1 250
box -6 -8 106 248
use NAND3X1  _1378_
timestamp 0
transform -1 0 1870 0 -1 730
box -6 -8 106 248
use NAND2X1  _1379_
timestamp 0
transform -1 0 1790 0 1 250
box -6 -8 86 248
use NAND3X1  _1380_
timestamp 0
transform 1 0 1650 0 -1 250
box -6 -8 106 248
use NAND3X1  _1381_
timestamp 0
transform 1 0 1950 0 -1 250
box -6 -8 106 248
use NOR3X1  _1382_
timestamp 0
transform 1 0 2490 0 -1 250
box -6 -8 186 248
use AOI21X1  _1383_
timestamp 0
transform -1 0 2910 0 -1 250
box -6 -8 106 248
use AOI21X1  _1384_
timestamp 0
transform 1 0 1750 0 -1 250
box -6 -8 106 248
use NAND3X1  _1385_
timestamp 0
transform 1 0 1990 0 -1 730
box -6 -8 106 248
use OAI21X1  _1386_
timestamp 0
transform -1 0 2190 0 -1 730
box -6 -8 106 248
use AOI21X1  _1387_
timestamp 0
transform 1 0 2110 0 1 250
box -6 -8 106 248
use OAI21X1  _1388_
timestamp 0
transform -1 0 2390 0 -1 250
box -6 -8 106 248
use NAND3X1  _1389_
timestamp 0
transform -1 0 2310 0 1 250
box -6 -8 106 248
use INVX1  _1390_
timestamp 0
transform -1 0 2490 0 1 250
box -6 -8 66 248
use NAND3X1  _1391_
timestamp 0
transform 1 0 2190 0 -1 250
box -6 -8 106 248
use OAI21X1  _1392_
timestamp 0
transform 1 0 2390 0 -1 250
box -6 -8 106 248
use NAND3X1  _1393_
timestamp 0
transform 1 0 2490 0 1 250
box -6 -8 106 248
use AOI21X1  _1394_
timestamp 0
transform 1 0 2730 0 -1 730
box -6 -8 106 248
use NAND3X1  _1395_
timestamp 0
transform 1 0 2330 0 1 250
box -6 -8 106 248
use NAND3X1  _1396_
timestamp 0
transform 1 0 2590 0 1 250
box -6 -8 106 248
use AOI22X1  _1397_
timestamp 0
transform -1 0 2950 0 -1 730
box -6 -8 126 248
use NOR2X1  _1398_
timestamp 0
transform -1 0 2810 0 1 1210
box -6 -8 86 248
use AOI21X1  _1399_
timestamp 0
transform -1 0 2490 0 1 1690
box -6 -8 106 248
use OAI21X1  _1400_
timestamp 0
transform 1 0 2110 0 -1 2170
box -6 -8 106 248
use INVX1  _1401_
timestamp 0
transform -1 0 3230 0 -1 730
box -6 -8 66 248
use AOI21X1  _1402_
timestamp 0
transform -1 0 3170 0 -1 730
box -6 -8 106 248
use NAND3X1  _1403_
timestamp 0
transform 1 0 2970 0 -1 730
box -6 -8 106 248
use NAND3X1  _1404_
timestamp 0
transform -1 0 2730 0 -1 730
box -6 -8 106 248
use NAND2X1  _1405_
timestamp 0
transform 1 0 2650 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1406_
timestamp 0
transform -1 0 2130 0 1 2170
box -6 -8 106 248
use OAI21X1  _1407_
timestamp 0
transform -1 0 2190 0 1 2650
box -6 -8 106 248
use AND2X2  _1408_
timestamp 0
transform -1 0 2770 0 1 3130
box -6 -8 106 248
use NAND2X1  _1409_
timestamp 0
transform 1 0 2370 0 1 3130
box -6 -8 86 248
use OAI21X1  _1410_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 106 248
use OAI21X1  _1411_
timestamp 0
transform -1 0 2550 0 1 3130
box -6 -8 106 248
use AOI21X1  _1412_
timestamp 0
transform -1 0 2430 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1413_
timestamp 0
transform 1 0 2110 0 -1 3130
box -6 -8 126 248
use OAI21X1  _1414_
timestamp 0
transform -1 0 3990 0 1 3610
box -6 -8 106 248
use NAND3X1  _1415_
timestamp 0
transform -1 0 2290 0 1 1690
box -6 -8 106 248
use AOI21X1  _1416_
timestamp 0
transform -1 0 2730 0 1 1210
box -6 -8 106 248
use INVX1  _1417_
timestamp 0
transform 1 0 1870 0 -1 2170
box -6 -8 66 248
use OAI21X1  _1418_
timestamp 0
transform 1 0 1250 0 -1 730
box -6 -8 106 248
use INVX1  _1419_
timestamp 0
transform 1 0 1270 0 1 250
box -6 -8 66 248
use AOI21X1  _1420_
timestamp 0
transform -1 0 1650 0 -1 250
box -6 -8 106 248
use NAND2X1  _1421_
timestamp 0
transform -1 0 1010 0 1 730
box -6 -8 86 248
use INVX1  _1422_
timestamp 0
transform -1 0 450 0 1 250
box -6 -8 66 248
use NOR2X1  _1423_
timestamp 0
transform 1 0 530 0 1 730
box -6 -8 86 248
use OAI21X1  _1424_
timestamp 0
transform -1 0 1290 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1425_
timestamp 0
transform -1 0 370 0 1 250
box -6 -8 86 248
use OR2X2  _1426_
timestamp 0
transform -1 0 670 0 1 250
box -6 -8 106 248
use NAND3X1  _1427_
timestamp 0
transform 1 0 450 0 1 250
box -6 -8 106 248
use AND2X2  _1428_
timestamp 0
transform 1 0 90 0 -1 250
box -6 -8 106 248
use NOR2X1  _1429_
timestamp 0
transform -1 0 90 0 -1 250
box -6 -8 86 248
use OAI21X1  _1430_
timestamp 0
transform 1 0 210 0 -1 250
box -6 -8 106 248
use NAND2X1  _1431_
timestamp 0
transform -1 0 490 0 -1 250
box -6 -8 86 248
use NAND2X1  _1432_
timestamp 0
transform -1 0 1510 0 1 730
box -6 -8 86 248
use NAND2X1  _1433_
timestamp 0
transform 1 0 1470 0 1 1210
box -6 -8 86 248
use INVX1  _1434_
timestamp 0
transform -1 0 1090 0 -1 1210
box -6 -8 66 248
use NAND2X1  _1435_
timestamp 0
transform 1 0 1390 0 1 1210
box -6 -8 86 248
use NAND2X1  _1436_
timestamp 0
transform 1 0 1310 0 1 1210
box -6 -8 86 248
use NOR2X1  _1437_
timestamp 0
transform -1 0 1190 0 1 1210
box -6 -8 86 248
use INVX1  _1438_
timestamp 0
transform -1 0 870 0 -1 1210
box -6 -8 66 248
use AOI22X1  _1439_
timestamp 0
transform -1 0 1450 0 -1 1690
box -6 -8 126 248
use INVX1  _1440_
timestamp 0
transform -1 0 930 0 -1 1210
box -6 -8 66 248
use NAND3X1  _1441_
timestamp 0
transform -1 0 790 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1442_
timestamp 0
transform 1 0 1090 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1443_
timestamp 0
transform -1 0 790 0 1 730
box -6 -8 86 248
use AOI21X1  _1444_
timestamp 0
transform -1 0 1110 0 -1 730
box -6 -8 106 248
use NAND3X1  _1445_
timestamp 0
transform -1 0 1230 0 -1 730
box -6 -8 106 248
use INVX1  _1446_
timestamp 0
transform 1 0 730 0 -1 730
box -6 -8 66 248
use OAI21X1  _1447_
timestamp 0
transform 1 0 770 0 1 250
box -6 -8 106 248
use AND2X2  _1448_
timestamp 0
transform -1 0 410 0 -1 250
box -6 -8 106 248
use NAND2X1  _1449_
timestamp 0
transform -1 0 1110 0 1 730
box -6 -8 86 248
use NAND3X1  _1450_
timestamp 0
transform -1 0 710 0 1 730
box -6 -8 106 248
use NAND3X1  _1451_
timestamp 0
transform 1 0 610 0 -1 250
box -6 -8 106 248
use NAND3X1  _1452_
timestamp 0
transform 1 0 1230 0 -1 250
box -6 -8 106 248
use OAI21X1  _1453_
timestamp 0
transform -1 0 1550 0 -1 250
box -6 -8 106 248
use AOI22X1  _1454_
timestamp 0
transform 1 0 490 0 -1 250
box -6 -8 126 248
use OR2X2  _1455_
timestamp 0
transform -1 0 1010 0 -1 730
box -6 -8 106 248
use NAND2X1  _1456_
timestamp 0
transform -1 0 870 0 1 730
box -6 -8 86 248
use AOI21X1  _1457_
timestamp 0
transform -1 0 910 0 -1 730
box -6 -8 106 248
use OAI21X1  _1458_
timestamp 0
transform 1 0 1010 0 -1 250
box -6 -8 106 248
use NAND3X1  _1459_
timestamp 0
transform 1 0 1330 0 -1 250
box -6 -8 106 248
use NAND3X1  _1460_
timestamp 0
transform 1 0 810 0 -1 250
box -6 -8 106 248
use OAI21X1  _1461_
timestamp 0
transform 1 0 1130 0 -1 250
box -6 -8 106 248
use NAND3X1  _1462_
timestamp 0
transform -1 0 1270 0 1 250
box -6 -8 106 248
use NAND2X1  _1463_
timestamp 0
transform 1 0 1330 0 1 250
box -6 -8 86 248
use NAND3X1  _1464_
timestamp 0
transform -1 0 1990 0 1 250
box -6 -8 106 248
use AOI21X1  _1465_
timestamp 0
transform -1 0 2170 0 -1 250
box -6 -8 106 248
use OAI21X1  _1466_
timestamp 0
transform -1 0 2090 0 1 250
box -6 -8 106 248
use NAND3X1  _1467_
timestamp 0
transform 1 0 1410 0 1 250
box -6 -8 106 248
use NAND2X1  _1468_
timestamp 0
transform 1 0 1550 0 1 1690
box -6 -8 86 248
use AOI21X1  _1469_
timestamp 0
transform -1 0 1810 0 1 1690
box -6 -8 106 248
use NAND2X1  _1470_
timestamp 0
transform -1 0 2370 0 1 1690
box -6 -8 86 248
use OAI21X1  _1471_
timestamp 0
transform 1 0 1770 0 -1 2170
box -6 -8 106 248
use INVX1  _1472_
timestamp 0
transform -1 0 1170 0 1 2170
box -6 -8 66 248
use NOR2X1  _1473_
timestamp 0
transform 1 0 1430 0 1 2170
box -6 -8 86 248
use OAI21X1  _1474_
timestamp 0
transform 1 0 1470 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1475_
timestamp 0
transform -1 0 1790 0 -1 3130
box -6 -8 86 248
use NOR2X1  _1476_
timestamp 0
transform 1 0 1810 0 -1 3130
box -6 -8 86 248
use AOI21X1  _1477_
timestamp 0
transform -1 0 3610 0 1 3130
box -6 -8 106 248
use OAI21X1  _1478_
timestamp 0
transform -1 0 3370 0 1 3130
box -6 -8 106 248
use NOR2X1  _1479_
timestamp 0
transform -1 0 1390 0 1 3610
box -6 -8 86 248
use NOR2X1  _1480_
timestamp 0
transform -1 0 1930 0 1 3130
box -6 -8 86 248
use AOI22X1  _1481_
timestamp 0
transform -1 0 2050 0 1 3130
box -6 -8 126 248
use OAI21X1  _1482_
timestamp 0
transform 1 0 3710 0 -1 3610
box -6 -8 106 248
use INVX1  _1483_
timestamp 0
transform 1 0 2790 0 1 2650
box -6 -8 66 248
use INVX1  _1484_
timestamp 0
transform 1 0 1350 0 1 2650
box -6 -8 66 248
use OAI21X1  _1485_
timestamp 0
transform 1 0 1510 0 1 2650
box -6 -8 106 248
use INVX1  _1486_
timestamp 0
transform -1 0 1330 0 1 2170
box -6 -8 66 248
use OAI21X1  _1487_
timestamp 0
transform 1 0 190 0 1 250
box -6 -8 106 248
use INVX1  _1488_
timestamp 0
transform 1 0 450 0 -1 730
box -6 -8 66 248
use AOI21X1  _1489_
timestamp 0
transform 1 0 670 0 1 250
box -6 -8 106 248
use NAND2X1  _1490_
timestamp 0
transform -1 0 1010 0 -1 1210
box -6 -8 86 248
use INVX1  _1491_
timestamp 0
transform 1 0 330 0 -1 1210
box -6 -8 66 248
use NOR2X1  _1492_
timestamp 0
transform -1 0 850 0 1 1210
box -6 -8 86 248
use OAI22X1  _1493_
timestamp 0
transform 1 0 1190 0 1 1210
box -6 -8 126 248
use NAND2X1  _1494_
timestamp 0
transform 1 0 590 0 -1 1210
box -6 -8 86 248
use OR2X2  _1495_
timestamp 0
transform -1 0 590 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1496_
timestamp 0
transform -1 0 330 0 -1 1210
box -6 -8 106 248
use INVX2  _1497_
timestamp 0
transform -1 0 930 0 1 730
box -6 -8 66 248
use NAND2X1  _1498_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 86 248
use OAI21X1  _1499_
timestamp 0
transform -1 0 530 0 1 730
box -6 -8 106 248
use NAND2X1  _1500_
timestamp 0
transform 1 0 1470 0 1 1690
box -6 -8 86 248
use NAND2X1  _1501_
timestamp 0
transform 1 0 1250 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1502_
timestamp 0
transform -1 0 1250 0 -1 1690
box -6 -8 86 248
use INVX1  _1503_
timestamp 0
transform -1 0 1110 0 -1 1690
box -6 -8 66 248
use INVX1  _1504_
timestamp 0
transform -1 0 910 0 1 1210
box -6 -8 66 248
use OAI21X1  _1505_
timestamp 0
transform 1 0 1010 0 1 1210
box -6 -8 106 248
use AND2X2  _1506_
timestamp 0
transform -1 0 1010 0 1 1210
box -6 -8 106 248
use AOI21X1  _1507_
timestamp 0
transform 1 0 250 0 1 730
box -6 -8 106 248
use INVX1  _1508_
timestamp 0
transform -1 0 130 0 1 730
box -6 -8 66 248
use NAND3X1  _1509_
timestamp 0
transform -1 0 230 0 1 730
box -6 -8 106 248
use NAND3X1  _1510_
timestamp 0
transform 1 0 230 0 -1 730
box -6 -8 106 248
use OAI21X1  _1511_
timestamp 0
transform -1 0 730 0 -1 730
box -6 -8 106 248
use INVX1  _1512_
timestamp 0
transform -1 0 70 0 1 730
box -6 -8 66 248
use OAI21X1  _1513_
timestamp 0
transform 1 0 330 0 -1 730
box -6 -8 106 248
use NAND3X1  _1514_
timestamp 0
transform 1 0 510 0 -1 730
box -6 -8 106 248
use NAND3X1  _1515_
timestamp 0
transform -1 0 130 0 -1 730
box -6 -8 106 248
use OAI21X1  _1516_
timestamp 0
transform 1 0 130 0 -1 730
box -6 -8 106 248
use NAND3X1  _1517_
timestamp 0
transform -1 0 190 0 1 250
box -6 -8 106 248
use NAND2X1  _1518_
timestamp 0
transform -1 0 950 0 1 250
box -6 -8 86 248
use NAND3X1  _1519_
timestamp 0
transform -1 0 1170 0 1 250
box -6 -8 106 248
use AOI21X1  _1520_
timestamp 0
transform -1 0 810 0 -1 250
box -6 -8 106 248
use OAI21X1  _1521_
timestamp 0
transform -1 0 1010 0 -1 250
box -6 -8 106 248
use NAND3X1  _1522_
timestamp 0
transform 1 0 950 0 1 250
box -6 -8 106 248
use NAND2X1  _1523_
timestamp 0
transform 1 0 1290 0 1 1690
box -6 -8 86 248
use NOR3X1  _1524_
timestamp 0
transform -1 0 1290 0 -1 2650
box -6 -8 186 248
use AOI21X1  _1525_
timestamp 0
transform -1 0 1430 0 1 2170
box -6 -8 106 248
use INVX1  _1526_
timestamp 0
transform 1 0 1290 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1527_
timestamp 0
transform 1 0 1370 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1528_
timestamp 0
transform 1 0 1410 0 1 2650
box -6 -8 106 248
use NAND2X1  _1529_
timestamp 0
transform -1 0 3350 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1530_
timestamp 0
transform -1 0 3270 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1531_
timestamp 0
transform -1 0 3190 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1532_
timestamp 0
transform 1 0 2850 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1533_
timestamp 0
transform 1 0 2790 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1534_
timestamp 0
transform -1 0 2790 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1535_
timestamp 0
transform -1 0 2790 0 1 2650
box -6 -8 126 248
use INVX1  _1536_
timestamp 0
transform -1 0 2530 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1537_
timestamp 0
transform -1 0 90 0 1 250
box -6 -8 86 248
use INVX1  _1538_
timestamp 0
transform -1 0 90 0 -1 2170
box -6 -8 66 248
use OAI21X1  _1539_
timestamp 0
transform 1 0 390 0 -1 1210
box -6 -8 106 248
use INVX1  _1540_
timestamp 0
transform -1 0 170 0 1 1210
box -6 -8 66 248
use INVX1  _1541_
timestamp 0
transform -1 0 1170 0 -1 1690
box -6 -8 66 248
use NOR2X1  _1542_
timestamp 0
transform -1 0 790 0 1 1690
box -6 -8 86 248
use NOR2X1  _1543_
timestamp 0
transform 1 0 1190 0 1 1690
box -6 -8 86 248
use NOR2X1  _1544_
timestamp 0
transform 1 0 1110 0 1 1690
box -6 -8 86 248
use AOI21X1  _1545_
timestamp 0
transform -1 0 1110 0 1 1690
box -6 -8 106 248
use NAND2X1  _1546_
timestamp 0
transform 1 0 610 0 1 1690
box -6 -8 86 248
use NOR2X1  _1547_
timestamp 0
transform 1 0 950 0 -1 1690
box -6 -8 86 248
use OAI22X1  _1548_
timestamp 0
transform 1 0 890 0 1 1690
box -6 -8 126 248
use NAND2X1  _1549_
timestamp 0
transform -1 0 670 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1550_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 106 248
use INVX1  _1551_
timestamp 0
transform -1 0 490 0 -1 1690
box -6 -8 66 248
use NAND3X1  _1552_
timestamp 0
transform 1 0 490 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1553_
timestamp 0
transform 1 0 550 0 1 1210
box -6 -8 86 248
use NOR2X1  _1554_
timestamp 0
transform -1 0 110 0 -1 1210
box -6 -8 86 248
use AOI21X1  _1555_
timestamp 0
transform -1 0 550 0 1 1210
box -6 -8 106 248
use OAI21X1  _1556_
timestamp 0
transform -1 0 110 0 1 1210
box -6 -8 106 248
use OR2X2  _1557_
timestamp 0
transform 1 0 110 0 -1 1210
box -6 -8 106 248
use INVX1  _1558_
timestamp 0
transform -1 0 450 0 1 1210
box -6 -8 66 248
use NAND3X1  _1559_
timestamp 0
transform 1 0 270 0 1 1210
box -6 -8 106 248
use NAND2X1  _1560_
timestamp 0
transform 1 0 170 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1561_
timestamp 0
transform -1 0 170 0 -1 2170
box -6 -8 86 248
use NAND3X1  _1562_
timestamp 0
transform 1 0 270 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1563_
timestamp 0
transform 1 0 550 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1564_
timestamp 0
transform -1 0 2110 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1565_
timestamp 0
transform -1 0 1270 0 1 2170
box -6 -8 86 248
use NAND3X1  _1566_
timestamp 0
transform -1 0 2030 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1567_
timestamp 0
transform 1 0 1370 0 1 1690
box -6 -8 86 248
use AOI22X1  _1568_
timestamp 0
transform 1 0 1430 0 -1 2170
box -6 -8 126 248
use AOI21X1  _1569_
timestamp 0
transform -1 0 1250 0 -1 2170
box -6 -8 106 248
use INVX1  _1570_
timestamp 0
transform 1 0 830 0 1 2170
box -6 -8 66 248
use NAND2X1  _1571_
timestamp 0
transform 1 0 1350 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1572_
timestamp 0
transform 1 0 1250 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1573_
timestamp 0
transform 1 0 1570 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1574_
timestamp 0
transform -1 0 1770 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1575_
timestamp 0
transform 1 0 890 0 1 2170
box -6 -8 106 248
use OAI21X1  _1576_
timestamp 0
transform 1 0 990 0 1 2170
box -6 -8 106 248
use OR2X2  _1577_
timestamp 0
transform -1 0 1010 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1578_
timestamp 0
transform 1 0 1010 0 -1 2650
box -6 -8 106 248
use INVX1  _1579_
timestamp 0
transform -1 0 3170 0 1 2650
box -6 -8 66 248
use OAI21X1  _1580_
timestamp 0
transform -1 0 3270 0 1 2650
box -6 -8 106 248
use NAND2X1  _1581_
timestamp 0
transform -1 0 3110 0 1 2650
box -6 -8 86 248
use NAND2X1  _1582_
timestamp 0
transform 1 0 2290 0 1 2650
box -6 -8 86 248
use OAI21X1  _1583_
timestamp 0
transform -1 0 2570 0 1 2650
box -6 -8 106 248
use AOI21X1  _1584_
timestamp 0
transform -1 0 2470 0 1 2650
box -6 -8 106 248
use AOI22X1  _1585_
timestamp 0
transform -1 0 2470 0 -1 2650
box -6 -8 126 248
use INVX1  _1586_
timestamp 0
transform -1 0 2310 0 1 2170
box -6 -8 66 248
use AOI21X1  _1587_
timestamp 0
transform -1 0 590 0 1 1690
box -6 -8 106 248
use NOR2X1  _1588_
timestamp 0
transform 1 0 750 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1589_
timestamp 0
transform -1 0 830 0 -1 2170
box -6 -8 86 248
use OAI22X1  _1590_
timestamp 0
transform 1 0 830 0 -1 1690
box -6 -8 126 248
use NAND2X1  _1591_
timestamp 0
transform -1 0 750 0 -1 1690
box -6 -8 86 248
use OR2X2  _1592_
timestamp 0
transform -1 0 310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1593_
timestamp 0
transform -1 0 430 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1594_
timestamp 0
transform -1 0 210 0 -1 1690
box -6 -8 86 248
use NAND2X1  _1595_
timestamp 0
transform -1 0 190 0 1 1690
box -6 -8 86 248
use OR2X2  _1596_
timestamp 0
transform -1 0 130 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1597_
timestamp 0
transform -1 0 390 0 1 1690
box -6 -8 86 248
use NAND3X1  _1598_
timestamp 0
transform 1 0 390 0 1 1690
box -6 -8 106 248
use OAI21X1  _1599_
timestamp 0
transform 1 0 170 0 1 1210
box -6 -8 106 248
use NAND3X1  _1600_
timestamp 0
transform 1 0 210 0 1 1690
box -6 -8 106 248
use NAND2X1  _1601_
timestamp 0
transform 1 0 370 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1602_
timestamp 0
transform 1 0 930 0 -1 2170
box -6 -8 86 248
use NAND3X1  _1603_
timestamp 0
transform -1 0 930 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1604_
timestamp 0
transform -1 0 830 0 1 2170
box -6 -8 106 248
use NAND3X1  _1605_
timestamp 0
transform 1 0 410 0 1 2170
box -6 -8 106 248
use INVX1  _1606_
timestamp 0
transform -1 0 890 0 -1 2650
box -6 -8 66 248
use OR2X2  _1607_
timestamp 0
transform -1 0 290 0 1 2170
box -6 -8 106 248
use AND2X2  _1608_
timestamp 0
transform 1 0 310 0 1 2170
box -6 -8 106 248
use NAND3X1  _1609_
timestamp 0
transform 1 0 510 0 1 2170
box -6 -8 106 248
use AOI21X1  _1610_
timestamp 0
transform -1 0 3210 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1611_
timestamp 0
transform -1 0 3110 0 -1 2650
box -6 -8 106 248
use INVX1  _1612_
timestamp 0
transform 1 0 1910 0 -1 3130
box -6 -8 66 248
use AOI21X1  _1613_
timestamp 0
transform 1 0 2230 0 -1 3130
box -6 -8 106 248
use AOI21X1  _1614_
timestamp 0
transform -1 0 2330 0 -1 2650
box -6 -8 106 248
use AOI22X1  _1615_
timestamp 0
transform -1 0 2250 0 1 2170
box -6 -8 126 248
use INVX1  _1616_
timestamp 0
transform -1 0 1990 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1617_
timestamp 0
transform -1 0 550 0 -1 2170
box -6 -8 106 248
use INVX1  _1618_
timestamp 0
transform -1 0 510 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1619_
timestamp 0
transform -1 0 110 0 1 1690
box -6 -8 106 248
use INVX1  _1620_
timestamp 0
transform -1 0 90 0 1 2170
box -6 -8 66 248
use OAI21X1  _1621_
timestamp 0
transform -1 0 890 0 1 1690
box -6 -8 106 248
use OR2X2  _1622_
timestamp 0
transform -1 0 110 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1623_
timestamp 0
transform -1 0 190 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1624_
timestamp 0
transform 1 0 210 0 -1 2650
box -6 -8 86 248
use NAND3X1  _1625_
timestamp 0
transform 1 0 630 0 -1 2650
box -6 -8 106 248
use OR2X2  _1626_
timestamp 0
transform 1 0 630 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1627_
timestamp 0
transform -1 0 1130 0 -1 2170
box -6 -8 106 248
use INVX1  _1628_
timestamp 0
transform 1 0 290 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1629_
timestamp 0
transform -1 0 450 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1630_
timestamp 0
transform 1 0 730 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1631_
timestamp 0
transform -1 0 3390 0 1 2170
box -6 -8 106 248
use OAI21X1  _1632_
timestamp 0
transform -1 0 3490 0 1 2170
box -6 -8 106 248
use NAND2X1  _1633_
timestamp 0
transform -1 0 3030 0 1 2170
box -6 -8 86 248
use NAND2X1  _1634_
timestamp 0
transform 1 0 1970 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1635_
timestamp 0
transform -1 0 2090 0 1 2650
box -6 -8 106 248
use AOI21X1  _1636_
timestamp 0
transform -1 0 1970 0 1 2650
box -6 -8 106 248
use AOI22X1  _1637_
timestamp 0
transform -1 0 1910 0 -1 2650
box -6 -8 126 248
use INVX1  _1638_
timestamp 0
transform -1 0 1690 0 1 2170
box -6 -8 66 248
use AOI21X1  _1639_
timestamp 0
transform 1 0 530 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1640_
timestamp 0
transform 1 0 90 0 1 2170
box -6 -8 106 248
use OAI21X1  _1641_
timestamp 0
transform 1 0 610 0 1 2170
box -6 -8 106 248
use NAND3X1  _1642_
timestamp 0
transform -1 0 3830 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1643_
timestamp 0
transform 1 0 4010 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1644_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1645_
timestamp 0
transform 1 0 1690 0 1 2650
box -6 -8 86 248
use OAI21X1  _1646_
timestamp 0
transform -1 0 1790 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1647_
timestamp 0
transform -1 0 1690 0 -1 2650
box -6 -8 106 248
use AOI22X1  _1648_
timestamp 0
transform -1 0 1630 0 1 2170
box -6 -8 126 248
use NAND2X1  _1649_
timestamp 0
transform -1 0 3750 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1650_
timestamp 0
transform 1 0 3570 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1651_
timestamp 0
transform -1 0 3610 0 1 4090
box -6 -8 86 248
use OAI21X1  _1652_
timestamp 0
transform -1 0 3710 0 1 4090
box -6 -8 106 248
use NAND2X1  _1653_
timestamp 0
transform -1 0 4070 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1654_
timestamp 0
transform 1 0 3970 0 1 4090
box -6 -8 106 248
use NAND2X1  _1655_
timestamp 0
transform -1 0 3610 0 1 4570
box -6 -8 86 248
use OAI21X1  _1656_
timestamp 0
transform 1 0 3410 0 1 4570
box -6 -8 106 248
use NAND2X1  _1657_
timestamp 0
transform -1 0 3050 0 1 3610
box -6 -8 86 248
use OAI21X1  _1658_
timestamp 0
transform 1 0 2870 0 1 3610
box -6 -8 106 248
use NAND2X1  _1659_
timestamp 0
transform 1 0 3430 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1660_
timestamp 0
transform 1 0 3330 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1661_
timestamp 0
transform 1 0 3110 0 1 4090
box -6 -8 86 248
use OAI21X1  _1662_
timestamp 0
transform -1 0 3110 0 1 4090
box -6 -8 106 248
use NAND2X1  _1663_
timestamp 0
transform 1 0 3130 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1664_
timestamp 0
transform 1 0 3030 0 -1 3610
box -6 -8 106 248
use DFFPOSX1  _1665_
timestamp 0
transform -1 0 3830 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1666_
timestamp 0
transform -1 0 4050 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1667_
timestamp 0
transform 1 0 3830 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1668_
timestamp 0
transform 1 0 2510 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1669_
timestamp 0
transform -1 0 2670 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1670_
timestamp 0
transform 1 0 2950 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1671_
timestamp 0
transform -1 0 2990 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1672_
timestamp 0
transform -1 0 3450 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1673_
timestamp 0
transform -1 0 2490 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1674_
timestamp 0
transform -1 0 2290 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1675_
timestamp 0
transform -1 0 3790 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1676_
timestamp 0
transform -1 0 3010 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1677_
timestamp 0
transform -1 0 2770 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1678_
timestamp 0
transform 1 0 2310 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1679_
timestamp 0
transform 1 0 1990 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1680_
timestamp 0
transform 1 0 1690 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1681_
timestamp 0
transform 1 0 3750 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1682_
timestamp 0
transform -1 0 3430 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1683_
timestamp 0
transform 1 0 4070 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1684_
timestamp 0
transform -1 0 3850 0 1 4570
box -6 -8 246 248
use DFFPOSX1  _1685_
timestamp 0
transform 1 0 3050 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1686_
timestamp 0
transform -1 0 3330 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1687_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1688_
timestamp 0
transform -1 0 3070 0 1 3130
box -6 -8 246 248
use DFFSR  _1689_
timestamp 0
transform -1 0 4550 0 -1 4570
box -6 -8 486 248
use DFFSR  _1690_
timestamp 0
transform -1 0 4530 0 1 4570
box -6 -8 486 248
use DFFSR  _1691_
timestamp 0
transform -1 0 5110 0 1 4570
box -6 -8 486 248
use INVX1  _1692_
timestamp 0
transform -1 0 1830 0 1 4570
box -6 -8 66 248
use INVX4  _1693_
timestamp 0
transform -1 0 2310 0 1 4570
box -6 -8 86 248
use OAI21X1  _1694_
timestamp 0
transform 1 0 1830 0 1 4570
box -6 -8 106 248
use NOR2X1  _1695_
timestamp 0
transform 1 0 1690 0 1 4570
box -6 -8 86 248
use INVX1  _1696_
timestamp 0
transform -1 0 1570 0 1 4570
box -6 -8 66 248
use INVX2  _1697_
timestamp 0
transform -1 0 2870 0 1 4570
box -6 -8 66 248
use NAND2X1  _1698_
timestamp 0
transform 1 0 2310 0 1 4570
box -6 -8 86 248
use INVX2  _1699_
timestamp 0
transform -1 0 1990 0 1 4090
box -6 -8 66 248
use NAND2X1  _1700_
timestamp 0
transform -1 0 2210 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1701_
timestamp 0
transform 1 0 2690 0 -1 4570
box -6 -8 86 248
use AOI22X1  _1702_
timestamp 0
transform -1 0 2330 0 -1 4570
box -6 -8 126 248
use INVX2  _1703_
timestamp 0
transform -1 0 2070 0 1 3610
box -6 -8 66 248
use INVX1  _1704_
timestamp 0
transform -1 0 2150 0 1 4090
box -6 -8 66 248
use INVX1  _1705_
timestamp 0
transform -1 0 2450 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1706_
timestamp 0
transform -1 0 2090 0 1 4090
box -6 -8 106 248
use NAND2X1  _1707_
timestamp 0
transform 1 0 1950 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1708_
timestamp 0
transform -1 0 1830 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1709_
timestamp 0
transform -1 0 1950 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1710_
timestamp 0
transform 1 0 2110 0 1 4570
box -6 -8 106 248
use AOI21X1  _1711_
timestamp 0
transform -1 0 2110 0 1 4570
box -6 -8 106 248
use NOR2X1  _1712_
timestamp 0
transform 1 0 1930 0 1 4570
box -6 -8 86 248
use OAI21X1  _1713_
timestamp 0
transform -1 0 1250 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1714_
timestamp 0
transform -1 0 1350 0 -1 4570
box -6 -8 106 248
use OR2X2  _1715_
timestamp 0
transform -1 0 1510 0 1 4570
box -6 -8 106 248
use OAI21X1  _1716_
timestamp 0
transform -1 0 1690 0 1 4570
box -6 -8 106 248
use NAND2X1  _1717_
timestamp 0
transform -1 0 1410 0 1 4570
box -6 -8 86 248
use INVX1  _1718_
timestamp 0
transform -1 0 1230 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1719_
timestamp 0
transform -1 0 1130 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1720_
timestamp 0
transform -1 0 1050 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1721_
timestamp 0
transform -1 0 1630 0 1 4090
box -6 -8 86 248
use NAND3X1  _1722_
timestamp 0
transform -1 0 1950 0 -1 4090
box -6 -8 106 248
use AOI22X1  _1723_
timestamp 0
transform 1 0 1730 0 1 4090
box -6 -8 126 248
use INVX1  _1724_
timestamp 0
transform -1 0 2210 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1725_
timestamp 0
transform 1 0 2050 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1726_
timestamp 0
transform -1 0 2050 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1727_
timestamp 0
transform -1 0 1730 0 1 4090
box -6 -8 106 248
use OAI21X1  _1728_
timestamp 0
transform 1 0 1230 0 1 4570
box -6 -8 106 248
use AOI21X1  _1729_
timestamp 0
transform -1 0 1210 0 1 4570
box -6 -8 106 248
use INVX1  _1730_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 66 248
use OAI21X1  _1731_
timestamp 0
transform -1 0 1030 0 1 4570
box -6 -8 106 248
use MUX2X1  _1732_
timestamp 0
transform 1 0 810 0 1 4570
box -6 -8 126 248
use NAND2X1  _1733_
timestamp 0
transform 1 0 850 0 -1 4570
box -6 -8 86 248
use INVX1  _1734_
timestamp 0
transform -1 0 1410 0 -1 4570
box -6 -8 66 248
use OAI21X1  _1735_
timestamp 0
transform -1 0 1510 0 -1 4570
box -6 -8 106 248
use MUX2X1  _1736_
timestamp 0
transform 1 0 2250 0 1 4090
box -6 -8 126 248
use OAI21X1  _1737_
timestamp 0
transform 1 0 2210 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1738_
timestamp 0
transform -1 0 2230 0 1 4090
box -6 -8 86 248
use NAND3X1  _1739_
timestamp 0
transform -1 0 2130 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1740_
timestamp 0
transform -1 0 1750 0 -1 4570
box -6 -8 106 248
use AOI22X1  _1741_
timestamp 0
transform 1 0 1510 0 -1 4570
box -6 -8 126 248
use OAI21X1  _1742_
timestamp 0
transform -1 0 850 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1743_
timestamp 0
transform -1 0 670 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1744_
timestamp 0
transform -1 0 570 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1745_
timestamp 0
transform -1 0 470 0 -1 4570
box -6 -8 86 248
use INVX1  _1746_
timestamp 0
transform 1 0 2310 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1747_
timestamp 0
transform 1 0 670 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1748_
timestamp 0
transform -1 0 210 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1749_
timestamp 0
transform 1 0 2630 0 1 4570
box -6 -8 86 248
use INVX1  _1750_
timestamp 0
transform 1 0 2610 0 -1 4570
box -6 -8 66 248
use NOR2X1  _1751_
timestamp 0
transform 1 0 2530 0 -1 4570
box -6 -8 86 248
use NAND2X1  _1752_
timestamp 0
transform 1 0 2430 0 -1 4570
box -6 -8 86 248
use AOI22X1  _1753_
timestamp 0
transform -1 0 2510 0 1 4570
box -6 -8 126 248
use OAI21X1  _1754_
timestamp 0
transform -1 0 2430 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1755_
timestamp 0
transform 1 0 2530 0 1 4570
box -6 -8 106 248
use OAI21X1  _1756_
timestamp 0
transform -1 0 730 0 1 4570
box -6 -8 106 248
use AOI21X1  _1757_
timestamp 0
transform -1 0 630 0 1 4570
box -6 -8 106 248
use INVX1  _1758_
timestamp 0
transform -1 0 310 0 1 4570
box -6 -8 66 248
use OAI21X1  _1759_
timestamp 0
transform -1 0 250 0 1 4570
box -6 -8 106 248
use MUX2X1  _1760_
timestamp 0
transform -1 0 130 0 1 4570
box -6 -8 126 248
use NAND2X1  _1761_
timestamp 0
transform -1 0 90 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1762_
timestamp 0
transform -1 0 530 0 1 4570
box -6 -8 106 248
use OAI21X1  _1763_
timestamp 0
transform 1 0 330 0 1 4570
box -6 -8 106 248
use NAND3X1  _1764_
timestamp 0
transform -1 0 390 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1765_
timestamp 0
transform 1 0 210 0 -1 4570
box -6 -8 86 248
use INVX1  _1766_
timestamp 0
transform 1 0 770 0 -1 4090
box -6 -8 66 248
use INVX1  _1767_
timestamp 0
transform -1 0 210 0 -1 4090
box -6 -8 66 248
use AND2X2  _1768_
timestamp 0
transform 1 0 90 0 1 4090
box -6 -8 106 248
use NAND2X1  _1769_
timestamp 0
transform -1 0 1090 0 -1 4090
box -6 -8 86 248
use AND2X2  _1770_
timestamp 0
transform -1 0 1550 0 1 4090
box -6 -8 106 248
use NAND2X1  _1771_
timestamp 0
transform 1 0 1250 0 1 4090
box -6 -8 86 248
use AOI22X1  _1772_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 126 248
use OAI21X1  _1773_
timestamp 0
transform -1 0 1230 0 1 4090
box -6 -8 106 248
use OAI21X1  _1774_
timestamp 0
transform -1 0 1130 0 1 4090
box -6 -8 106 248
use OAI21X1  _1775_
timestamp 0
transform -1 0 1030 0 1 4090
box -6 -8 106 248
use AOI21X1  _1776_
timestamp 0
transform -1 0 910 0 1 4090
box -6 -8 106 248
use OAI21X1  _1777_
timestamp 0
transform -1 0 810 0 1 4090
box -6 -8 106 248
use OAI21X1  _1778_
timestamp 0
transform -1 0 710 0 1 4090
box -6 -8 106 248
use INVX1  _1779_
timestamp 0
transform 1 0 390 0 1 4090
box -6 -8 66 248
use OAI21X1  _1780_
timestamp 0
transform 1 0 210 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1781_
timestamp 0
transform 1 0 270 0 1 4090
box -6 -8 106 248
use NAND2X1  _1782_
timestamp 0
transform -1 0 410 0 -1 4090
box -6 -8 86 248
use INVX1  _1783_
timestamp 0
transform 1 0 2790 0 -1 3610
box -6 -8 66 248
use INVX1  _1784_
timestamp 0
transform -1 0 690 0 -1 4090
box -6 -8 66 248
use AOI21X1  _1785_
timestamp 0
transform -1 0 630 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1786_
timestamp 0
transform 1 0 430 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1787_
timestamp 0
transform -1 0 270 0 1 4090
box -6 -8 86 248
use INVX1  _1788_
timestamp 0
transform -1 0 610 0 1 4090
box -6 -8 66 248
use AOI21X1  _1789_
timestamp 0
transform 1 0 450 0 1 4090
box -6 -8 106 248
use NAND2X1  _1790_
timestamp 0
transform -1 0 1490 0 1 3610
box -6 -8 86 248
use AND2X2  _1791_
timestamp 0
transform -1 0 2010 0 1 3610
box -6 -8 106 248
use NAND2X1  _1792_
timestamp 0
transform 1 0 1710 0 1 3610
box -6 -8 86 248
use AOI22X1  _1793_
timestamp 0
transform 1 0 1590 0 1 3610
box -6 -8 126 248
use OAI21X1  _1794_
timestamp 0
transform 1 0 1810 0 1 3610
box -6 -8 106 248
use OAI21X1  _1795_
timestamp 0
transform -1 0 1590 0 1 3610
box -6 -8 106 248
use OAI21X1  _1796_
timestamp 0
transform 1 0 1130 0 1 3610
box -6 -8 106 248
use AOI21X1  _1797_
timestamp 0
transform -1 0 1130 0 1 3610
box -6 -8 106 248
use OAI21X1  _1798_
timestamp 0
transform 1 0 830 0 1 3610
box -6 -8 106 248
use OAI21X1  _1799_
timestamp 0
transform -1 0 1030 0 1 3610
box -6 -8 106 248
use AOI21X1  _1800_
timestamp 0
transform 1 0 510 0 1 3610
box -6 -8 106 248
use NOR2X1  _1801_
timestamp 0
transform -1 0 90 0 1 4090
box -6 -8 86 248
use OAI21X1  _1802_
timestamp 0
transform 1 0 30 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1803_
timestamp 0
transform 1 0 690 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1804_
timestamp 0
transform -1 0 710 0 1 3610
box -6 -8 106 248
use INVX1  _1805_
timestamp 0
transform 1 0 1030 0 -1 3610
box -6 -8 66 248
use NOR2X1  _1806_
timestamp 0
transform 1 0 1330 0 -1 3610
box -6 -8 86 248
use NOR2X1  _1807_
timestamp 0
transform 1 0 1410 0 -1 3610
box -6 -8 86 248
use INVX1  _1808_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 66 248
use NAND2X1  _1809_
timestamp 0
transform 1 0 1230 0 -1 4090
box -6 -8 86 248
use AND2X2  _1810_
timestamp 0
transform -1 0 1850 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1811_
timestamp 0
transform 1 0 1530 0 -1 4090
box -6 -8 86 248
use AOI22X1  _1812_
timestamp 0
transform 1 0 1410 0 -1 4090
box -6 -8 126 248
use OAI21X1  _1813_
timestamp 0
transform 1 0 1630 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1814_
timestamp 0
transform -1 0 1410 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1815_
timestamp 0
transform 1 0 410 0 1 3610
box -6 -8 106 248
use AOI21X1  _1816_
timestamp 0
transform -1 0 410 0 1 3610
box -6 -8 106 248
use OAI21X1  _1817_
timestamp 0
transform -1 0 210 0 1 3610
box -6 -8 106 248
use OAI21X1  _1818_
timestamp 0
transform 1 0 210 0 1 3610
box -6 -8 106 248
use OAI21X1  _1819_
timestamp 0
transform -1 0 690 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1820_
timestamp 0
transform -1 0 1030 0 -1 3610
box -6 -8 106 248
use INVX1  _1821_
timestamp 0
transform -1 0 310 0 -1 3610
box -6 -8 66 248
use NAND2X1  _1822_
timestamp 0
transform -1 0 490 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1823_
timestamp 0
transform 1 0 690 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1824_
timestamp 0
transform -1 0 410 0 -1 3610
box -6 -8 106 248
use INVX1  _1825_
timestamp 0
transform 1 0 1430 0 1 3130
box -6 -8 66 248
use AND2X2  _1826_
timestamp 0
transform -1 0 1870 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1827_
timestamp 0
transform 1 0 1690 0 -1 3610
box -6 -8 86 248
use AOI22X1  _1828_
timestamp 0
transform 1 0 1570 0 -1 3610
box -6 -8 126 248
use OAI21X1  _1829_
timestamp 0
transform -1 0 1730 0 1 3130
box -6 -8 106 248
use OAI22X1  _1830_
timestamp 0
transform 1 0 1490 0 1 3130
box -6 -8 126 248
use OAI21X1  _1831_
timestamp 0
transform -1 0 810 0 1 3610
box -6 -8 106 248
use AOI21X1  _1832_
timestamp 0
transform 1 0 770 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1833_
timestamp 0
transform 1 0 870 0 1 3130
box -6 -8 106 248
use OAI21X1  _1834_
timestamp 0
transform -1 0 850 0 1 3130
box -6 -8 106 248
use NAND2X1  _1835_
timestamp 0
transform -1 0 750 0 1 3130
box -6 -8 86 248
use OAI21X1  _1836_
timestamp 0
transform -1 0 590 0 -1 3610
box -6 -8 106 248
use INVX1  _1837_
timestamp 0
transform -1 0 90 0 1 3130
box -6 -8 66 248
use NAND3X1  _1838_
timestamp 0
transform 1 0 470 0 1 3130
box -6 -8 106 248
use NAND2X1  _1839_
timestamp 0
transform -1 0 790 0 -1 3130
box -6 -8 86 248
use INVX1  _1840_
timestamp 0
transform -1 0 70 0 1 2650
box -6 -8 66 248
use AOI21X1  _1841_
timestamp 0
transform -1 0 290 0 1 3130
box -6 -8 106 248
use NAND2X1  _1842_
timestamp 0
transform 1 0 1850 0 1 4090
box -6 -8 86 248
use AND2X2  _1843_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1844_
timestamp 0
transform 1 0 2110 0 -1 3610
box -6 -8 86 248
use AOI22X1  _1845_
timestamp 0
transform 1 0 1970 0 -1 3610
box -6 -8 126 248
use OAI21X1  _1846_
timestamp 0
transform 1 0 2290 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1847_
timestamp 0
transform -1 0 1970 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1848_
timestamp 0
transform 1 0 1210 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1849_
timestamp 0
transform 1 0 1090 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1850_
timestamp 0
transform -1 0 1170 0 1 3130
box -6 -8 106 248
use OAI21X1  _1851_
timestamp 0
transform -1 0 1070 0 1 3130
box -6 -8 106 248
use OAI21X1  _1852_
timestamp 0
transform 1 0 190 0 1 2650
box -6 -8 106 248
use NAND2X1  _1853_
timestamp 0
transform -1 0 470 0 1 3130
box -6 -8 86 248
use INVX1  _1854_
timestamp 0
transform -1 0 510 0 -1 3130
box -6 -8 66 248
use NAND3X1  _1855_
timestamp 0
transform -1 0 490 0 1 2650
box -6 -8 106 248
use NAND2X1  _1856_
timestamp 0
transform -1 0 390 0 1 2650
box -6 -8 86 248
use NOR2X1  _1857_
timestamp 0
transform -1 0 1170 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1858_
timestamp 0
transform -1 0 1310 0 1 3610
box -6 -8 86 248
use NOR2X1  _1859_
timestamp 0
transform 1 0 1450 0 -1 3130
box -6 -8 86 248
use INVX1  _1860_
timestamp 0
transform 1 0 910 0 -1 3130
box -6 -8 66 248
use NAND3X1  _1861_
timestamp 0
transform 1 0 790 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1862_
timestamp 0
transform 1 0 1530 0 -1 3130
box -6 -8 86 248
use AND2X2  _1863_
timestamp 0
transform 1 0 1610 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1864_
timestamp 0
transform 1 0 530 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1865_
timestamp 0
transform -1 0 170 0 1 2650
box -6 -8 106 248
use NAND2X1  _1866_
timestamp 0
transform -1 0 670 0 1 2650
box -6 -8 86 248
use OAI21X1  _1867_
timestamp 0
transform 1 0 970 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1868_
timestamp 0
transform -1 0 1830 0 1 3130
box -6 -8 86 248
use OAI21X1  _1869_
timestamp 0
transform 1 0 570 0 1 3130
box -6 -8 106 248
use INVX1  _1870_
timestamp 0
transform 1 0 390 0 -1 3130
box -6 -8 66 248
use NAND3X1  _1871_
timestamp 0
transform -1 0 390 0 1 3130
box -6 -8 106 248
use NAND3X1  _1872_
timestamp 0
transform -1 0 390 0 -1 3130
box -6 -8 106 248
use INVX1  _1873_
timestamp 0
transform -1 0 70 0 -1 3130
box -6 -8 66 248
use NAND2X1  _1874_
timestamp 0
transform -1 0 170 0 1 3130
box -6 -8 86 248
use AOI21X1  _1875_
timestamp 0
transform -1 0 230 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1876_
timestamp 0
transform -1 0 170 0 -1 3130
box -6 -8 106 248
use AND2X2  _1877_
timestamp 0
transform 1 0 170 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1878_
timestamp 0
transform 1 0 970 0 1 2650
box -6 -8 106 248
use NAND3X1  _1879_
timestamp 0
transform 1 0 1090 0 -1 3130
box -6 -8 106 248
use INVX1  _1880_
timestamp 0
transform 1 0 1170 0 1 3130
box -6 -8 66 248
use NAND2X1  _1881_
timestamp 0
transform 1 0 1330 0 1 3130
box -6 -8 86 248
use AOI21X1  _1882_
timestamp 0
transform -1 0 1330 0 1 3130
box -6 -8 106 248
use NAND2X1  _1883_
timestamp 0
transform 1 0 1370 0 -1 3130
box -6 -8 86 248
use NOR2X1  _1884_
timestamp 0
transform 1 0 1270 0 -1 3130
box -6 -8 86 248
use NOR2X1  _1885_
timestamp 0
transform -1 0 1270 0 -1 3130
box -6 -8 86 248
use NAND3X1  _1886_
timestamp 0
transform 1 0 490 0 1 2650
box -6 -8 106 248
use INVX1  _1887_
timestamp 0
transform 1 0 650 0 -1 3130
box -6 -8 66 248
use NAND3X1  _1888_
timestamp 0
transform 1 0 670 0 1 2650
box -6 -8 106 248
use NAND2X1  _1889_
timestamp 0
transform -1 0 850 0 1 2650
box -6 -8 86 248
use NAND3X1  _1890_
timestamp 0
transform 1 0 1150 0 1 2650
box -6 -8 106 248
use AND2X2  _1891_
timestamp 0
transform 1 0 870 0 1 2650
box -6 -8 106 248
use NAND2X1  _1892_
timestamp 0
transform 1 0 1070 0 1 2650
box -6 -8 86 248
use NAND2X1  _1893_
timestamp 0
transform 1 0 1250 0 1 2650
box -6 -8 86 248
use BUFX2  _1894_
timestamp 0
transform -1 0 90 0 1 3610
box -6 -8 86 248
use BUFX2  _1895_
timestamp 0
transform -1 0 110 0 -1 3610
box -6 -8 86 248
use BUFX2  _1896_
timestamp 0
transform -1 0 3550 0 1 3610
box -6 -8 86 248
use BUFX2  _1897_
timestamp 0
transform 1 0 2850 0 1 2650
box -6 -8 86 248
use BUFX2  _1898_
timestamp 0
transform 1 0 2670 0 -1 2170
box -6 -8 86 248
use BUFX2  _1899_
timestamp 0
transform 1 0 2590 0 -1 2170
box -6 -8 86 248
use BUFX2  _1900_
timestamp 0
transform 1 0 2210 0 -1 2170
box -6 -8 86 248
use BUFX2  _1901_
timestamp 0
transform 1 0 2570 0 1 1690
box -6 -8 86 248
use BUFX2  _1902_
timestamp 0
transform -1 0 5090 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 2390 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform -1 0 2190 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 2370 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 2830 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 3630 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform -1 0 3010 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform 1 0 3630 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform -1 0 2750 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform 1 0 3430 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform 1 0 3890 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 3310 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 3310 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 3470 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 4230 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 4250 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 1930 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform 1 0 2290 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 1910 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 2110 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform -1 0 2250 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert26
timestamp 0
transform 1 0 3790 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 2910 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert28
timestamp 0
transform 1 0 3790 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert29
timestamp 0
transform 1 0 2870 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert30
timestamp 0
transform 1 0 1030 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert31
timestamp 0
transform 1 0 930 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert32
timestamp 0
transform -1 0 910 0 -1 4090
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform 1 0 3850 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform -1 0 3090 0 -1 3130
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform -1 0 4710 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert15
timestamp 0
transform -1 0 3410 0 1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert16
timestamp 0
transform -1 0 3270 0 1 3130
box -6 -8 206 248
use FILL  FILL75450x150
timestamp 0
transform -1 0 5050 0 -1 250
box -6 -8 26 248
use FILL  FILL75450x7350
timestamp 0
transform -1 0 5050 0 -1 730
box -6 -8 26 248
use FILL  FILL75450x14550
timestamp 0
transform -1 0 5050 0 -1 1210
box -6 -8 26 248
use FILL  FILL75450x36150
timestamp 0
transform -1 0 5050 0 -1 2650
box -6 -8 26 248
use FILL  FILL75450x39750
timestamp 0
transform 1 0 5030 0 1 2650
box -6 -8 26 248
use FILL  FILL75450x54150
timestamp 0
transform 1 0 5030 0 1 3610
box -6 -8 26 248
use FILL  FILL75750x150
timestamp 0
transform -1 0 5070 0 -1 250
box -6 -8 26 248
use FILL  FILL75750x7350
timestamp 0
transform -1 0 5070 0 -1 730
box -6 -8 26 248
use FILL  FILL75750x10950
timestamp 0
transform 1 0 5050 0 1 730
box -6 -8 26 248
use FILL  FILL75750x14550
timestamp 0
transform -1 0 5070 0 -1 1210
box -6 -8 26 248
use FILL  FILL75750x36150
timestamp 0
transform -1 0 5070 0 -1 2650
box -6 -8 26 248
use FILL  FILL75750x39750
timestamp 0
transform 1 0 5050 0 1 2650
box -6 -8 26 248
use FILL  FILL75750x54150
timestamp 0
transform 1 0 5050 0 1 3610
box -6 -8 26 248
use FILL  FILL76050x150
timestamp 0
transform -1 0 5090 0 -1 250
box -6 -8 26 248
use FILL  FILL76050x7350
timestamp 0
transform -1 0 5090 0 -1 730
box -6 -8 26 248
use FILL  FILL76050x10950
timestamp 0
transform 1 0 5070 0 1 730
box -6 -8 26 248
use FILL  FILL76050x14550
timestamp 0
transform -1 0 5090 0 -1 1210
box -6 -8 26 248
use FILL  FILL76050x25350
timestamp 0
transform 1 0 5070 0 1 1690
box -6 -8 26 248
use FILL  FILL76050x28950
timestamp 0
transform -1 0 5090 0 -1 2170
box -6 -8 26 248
use FILL  FILL76050x36150
timestamp 0
transform -1 0 5090 0 -1 2650
box -6 -8 26 248
use FILL  FILL76050x39750
timestamp 0
transform 1 0 5070 0 1 2650
box -6 -8 26 248
use FILL  FILL76050x54150
timestamp 0
transform 1 0 5070 0 1 3610
box -6 -8 26 248
use FILL  FILL76350x150
timestamp 0
transform -1 0 5110 0 -1 250
box -6 -8 26 248
use FILL  FILL76350x3750
timestamp 0
transform 1 0 5090 0 1 250
box -6 -8 26 248
use FILL  FILL76350x7350
timestamp 0
transform -1 0 5110 0 -1 730
box -6 -8 26 248
use FILL  FILL76350x10950
timestamp 0
transform 1 0 5090 0 1 730
box -6 -8 26 248
use FILL  FILL76350x14550
timestamp 0
transform -1 0 5110 0 -1 1210
box -6 -8 26 248
use FILL  FILL76350x25350
timestamp 0
transform 1 0 5090 0 1 1690
box -6 -8 26 248
use FILL  FILL76350x28950
timestamp 0
transform -1 0 5110 0 -1 2170
box -6 -8 26 248
use FILL  FILL76350x36150
timestamp 0
transform -1 0 5110 0 -1 2650
box -6 -8 26 248
use FILL  FILL76350x39750
timestamp 0
transform 1 0 5090 0 1 2650
box -6 -8 26 248
use FILL  FILL76350x43350
timestamp 0
transform -1 0 5110 0 -1 3130
box -6 -8 26 248
use FILL  FILL76350x50550
timestamp 0
transform -1 0 5110 0 -1 3610
box -6 -8 26 248
use FILL  FILL76350x54150
timestamp 0
transform 1 0 5090 0 1 3610
box -6 -8 26 248
use FILL  FILL76350x57750
timestamp 0
transform -1 0 5110 0 -1 4090
box -6 -8 26 248
use FILL  FILL76350x61350
timestamp 0
transform 1 0 5090 0 1 4090
box -6 -8 26 248
use FILL  FILL76350x64950
timestamp 0
transform -1 0 5110 0 -1 4570
box -6 -8 26 248
use FILL  FILL76650x150
timestamp 0
transform -1 0 5130 0 -1 250
box -6 -8 26 248
use FILL  FILL76650x3750
timestamp 0
transform 1 0 5110 0 1 250
box -6 -8 26 248
use FILL  FILL76650x7350
timestamp 0
transform -1 0 5130 0 -1 730
box -6 -8 26 248
use FILL  FILL76650x10950
timestamp 0
transform 1 0 5110 0 1 730
box -6 -8 26 248
use FILL  FILL76650x14550
timestamp 0
transform -1 0 5130 0 -1 1210
box -6 -8 26 248
use FILL  FILL76650x25350
timestamp 0
transform 1 0 5110 0 1 1690
box -6 -8 26 248
use FILL  FILL76650x28950
timestamp 0
transform -1 0 5130 0 -1 2170
box -6 -8 26 248
use FILL  FILL76650x32550
timestamp 0
transform 1 0 5110 0 1 2170
box -6 -8 26 248
use FILL  FILL76650x36150
timestamp 0
transform -1 0 5130 0 -1 2650
box -6 -8 26 248
use FILL  FILL76650x39750
timestamp 0
transform 1 0 5110 0 1 2650
box -6 -8 26 248
use FILL  FILL76650x43350
timestamp 0
transform -1 0 5130 0 -1 3130
box -6 -8 26 248
use FILL  FILL76650x50550
timestamp 0
transform -1 0 5130 0 -1 3610
box -6 -8 26 248
use FILL  FILL76650x54150
timestamp 0
transform 1 0 5110 0 1 3610
box -6 -8 26 248
use FILL  FILL76650x57750
timestamp 0
transform -1 0 5130 0 -1 4090
box -6 -8 26 248
use FILL  FILL76650x61350
timestamp 0
transform 1 0 5110 0 1 4090
box -6 -8 26 248
use FILL  FILL76650x64950
timestamp 0
transform -1 0 5130 0 -1 4570
box -6 -8 26 248
use FILL  FILL76650x68550
timestamp 0
transform 1 0 5110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__927_
timestamp 0
transform -1 0 4270 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__930_
timestamp 0
transform 1 0 4930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__934_
timestamp 0
transform 1 0 4330 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__938_
timestamp 0
transform -1 0 4770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__942_
timestamp 0
transform 1 0 4070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__946_
timestamp 0
transform 1 0 4950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__950_
timestamp 0
transform 1 0 4550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__954_
timestamp 0
transform 1 0 4790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__958_
timestamp 0
transform 1 0 4910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__961_
timestamp 0
transform 1 0 4910 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__965_
timestamp 0
transform -1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__969_
timestamp 0
transform 1 0 4050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__973_
timestamp 0
transform 1 0 2710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__977_
timestamp 0
transform 1 0 2650 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__981_
timestamp 0
transform -1 0 2990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__985_
timestamp 0
transform -1 0 2590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__989_
timestamp 0
transform -1 0 3050 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__992_
timestamp 0
transform 1 0 2550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__996_
timestamp 0
transform -1 0 4930 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1003_
timestamp 0
transform 1 0 4870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1007_
timestamp 0
transform 1 0 4770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1011_
timestamp 0
transform -1 0 2690 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1015_
timestamp 0
transform -1 0 3470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1019_
timestamp 0
transform 1 0 3950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 4270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1027_
timestamp 0
transform -1 0 4090 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 4550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1034_
timestamp 0
transform -1 0 2870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1038_
timestamp 0
transform -1 0 2790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 3390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1046_
timestamp 0
transform -1 0 4570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1050_
timestamp 0
transform -1 0 4810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1054_
timestamp 0
transform 1 0 4950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 2730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1061_
timestamp 0
transform 1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1065_
timestamp 0
transform -1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 4570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 4410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 2530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 3570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 3030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 4450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1092_
timestamp 0
transform -1 0 4930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 5030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1100_
timestamp 0
transform -1 0 3990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1104_
timestamp 0
transform -1 0 4950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1108_
timestamp 0
transform -1 0 4570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1112_
timestamp 0
transform -1 0 3770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1116_
timestamp 0
transform 1 0 3470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1120_
timestamp 0
transform 1 0 2990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 3770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1127_
timestamp 0
transform 1 0 3410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1131_
timestamp 0
transform -1 0 3130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 2910 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 4390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 4010 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1147_
timestamp 0
transform 1 0 4710 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1151_
timestamp 0
transform 1 0 4450 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1155_
timestamp 0
transform -1 0 4030 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1158_
timestamp 0
transform 1 0 4210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1162_
timestamp 0
transform -1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1166_
timestamp 0
transform 1 0 4530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1170_
timestamp 0
transform -1 0 4810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1174_
timestamp 0
transform -1 0 4250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1178_
timestamp 0
transform -1 0 4130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 4610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1186_
timestamp 0
transform 1 0 4750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1189_
timestamp 0
transform 1 0 3390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 4690 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1197_
timestamp 0
transform 1 0 4890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1201_
timestamp 0
transform -1 0 4190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1205_
timestamp 0
transform 1 0 4330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 3930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1213_
timestamp 0
transform -1 0 3730 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1217_
timestamp 0
transform -1 0 3690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1220_
timestamp 0
transform -1 0 3570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 4070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1228_
timestamp 0
transform 1 0 4230 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 3650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1236_
timestamp 0
transform 1 0 3890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1240_
timestamp 0
transform 1 0 3310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1244_
timestamp 0
transform -1 0 4330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 3630 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1251_
timestamp 0
transform 1 0 3830 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1255_
timestamp 0
transform -1 0 3450 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1259_
timestamp 0
transform 1 0 1950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 2250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1267_
timestamp 0
transform 1 0 1970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1271_
timestamp 0
transform -1 0 3130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1275_
timestamp 0
transform 1 0 1770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1282_
timestamp 0
transform -1 0 2310 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1286_
timestamp 0
transform 1 0 3210 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 2690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1294_
timestamp 0
transform 1 0 2670 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1298_
timestamp 0
transform -1 0 3030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1302_
timestamp 0
transform 1 0 3910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1306_
timestamp 0
transform -1 0 2910 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1310_
timestamp 0
transform -1 0 2790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1313_
timestamp 0
transform -1 0 4250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1317_
timestamp 0
transform 1 0 4130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1321_
timestamp 0
transform 1 0 2290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 2390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 2690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1337_
timestamp 0
transform -1 0 3350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 1130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1344_
timestamp 0
transform -1 0 1910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 1330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 2250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1356_
timestamp 0
transform 1 0 1450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 1290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1364_
timestamp 0
transform -1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1368_
timestamp 0
transform 1 0 1530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1372_
timestamp 0
transform 1 0 1790 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 2810 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1387_
timestamp 0
transform 1 0 2090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 2170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1395_
timestamp 0
transform 1 0 2310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1399_
timestamp 0
transform -1 0 2390 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1403_
timestamp 0
transform 1 0 2950 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1406_
timestamp 0
transform -1 0 2030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 2570 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1414_
timestamp 0
transform -1 0 3890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1418_
timestamp 0
transform 1 0 1230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1422_
timestamp 0
transform -1 0 390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1426_
timestamp 0
transform -1 0 570 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1434_
timestamp 0
transform -1 0 1030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1441_
timestamp 0
transform -1 0 690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1445_
timestamp 0
transform -1 0 1130 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1449_
timestamp 0
transform -1 0 1030 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1453_
timestamp 0
transform -1 0 1450 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1457_
timestamp 0
transform -1 0 810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1461_
timestamp 0
transform 1 0 1110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1465_
timestamp 0
transform -1 0 2070 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__1469_
timestamp 0
transform -1 0 1710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1472_
timestamp 0
transform -1 0 1110 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1476_
timestamp 0
transform 1 0 1790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1480_
timestamp 0
transform -1 0 1850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1484_
timestamp 0
transform 1 0 1330 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1488_
timestamp 0
transform 1 0 430 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1492_
timestamp 0
transform -1 0 770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1496_
timestamp 0
transform -1 0 230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1500_
timestamp 0
transform 1 0 1450 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1503_
timestamp 0
transform -1 0 1050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1507_
timestamp 0
transform 1 0 230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__1511_
timestamp 0
transform -1 0 630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1515_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__1519_
timestamp 0
transform -1 0 1070 0 1 250
box -6 -8 26 248
use FILL  FILL_0__1523_
timestamp 0
transform 1 0 1270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 1350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1531_
timestamp 0
transform -1 0 3110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 2690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1538_
timestamp 0
transform -1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1542_
timestamp 0
transform -1 0 710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1546_
timestamp 0
transform 1 0 590 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1550_
timestamp 0
transform -1 0 650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1554_
timestamp 0
transform -1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__1558_
timestamp 0
transform -1 0 390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__1562_
timestamp 0
transform 1 0 250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1565_
timestamp 0
transform -1 0 1190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1569_
timestamp 0
transform -1 0 1150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1573_
timestamp 0
transform 1 0 1550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1577_
timestamp 0
transform -1 0 910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1581_
timestamp 0
transform -1 0 3030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1585_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1589_
timestamp 0
transform -1 0 750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1593_
timestamp 0
transform -1 0 330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1596_
timestamp 0
transform -1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__1600_
timestamp 0
transform 1 0 190 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__1604_
timestamp 0
transform -1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1608_
timestamp 0
transform 1 0 290 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1612_
timestamp 0
transform 1 0 1890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1616_
timestamp 0
transform -1 0 1930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1620_
timestamp 0
transform -1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1624_
timestamp 0
transform 1 0 190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1627_
timestamp 0
transform -1 0 1030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1631_
timestamp 0
transform -1 0 3290 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__1635_
timestamp 0
transform -1 0 1990 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1639_
timestamp 0
transform 1 0 510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1643_
timestamp 0
transform 1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__1647_
timestamp 0
transform -1 0 1590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__1651_
timestamp 0
transform -1 0 3530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1655_
timestamp 0
transform -1 0 3530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1658_
timestamp 0
transform 1 0 2850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1662_
timestamp 0
transform -1 0 3010 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1693_
timestamp 0
transform -1 0 2230 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1697_
timestamp 0
transform -1 0 2810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1701_
timestamp 0
transform 1 0 2670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1705_
timestamp 0
transform -1 0 2390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1709_
timestamp 0
transform -1 0 1850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1713_
timestamp 0
transform -1 0 1150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1716_
timestamp 0
transform -1 0 1590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1720_
timestamp 0
transform -1 0 950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1724_
timestamp 0
transform -1 0 2150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1728_
timestamp 0
transform 1 0 1210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1732_
timestamp 0
transform 1 0 790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1736_
timestamp 0
transform 1 0 2230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1740_
timestamp 0
transform -1 0 1650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1744_
timestamp 0
transform -1 0 490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1748_
timestamp 0
transform -1 0 110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1751_
timestamp 0
transform 1 0 2510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__1755_
timestamp 0
transform 1 0 2510 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1759_
timestamp 0
transform -1 0 150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1763_
timestamp 0
transform 1 0 310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__1767_
timestamp 0
transform -1 0 150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1771_
timestamp 0
transform 1 0 1230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1775_
timestamp 0
transform -1 0 930 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1779_
timestamp 0
transform 1 0 370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__1782_
timestamp 0
transform -1 0 330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1786_
timestamp 0
transform 1 0 410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1790_
timestamp 0
transform -1 0 1410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1794_
timestamp 0
transform 1 0 1790 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1798_
timestamp 0
transform 1 0 810 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1802_
timestamp 0
transform 1 0 10 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1806_
timestamp 0
transform 1 0 1310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1810_
timestamp 0
transform -1 0 1750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1813_
timestamp 0
transform 1 0 1610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__1817_
timestamp 0
transform -1 0 110 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__1821_
timestamp 0
transform -1 0 250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1825_
timestamp 0
transform 1 0 1410 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1829_
timestamp 0
transform -1 0 1630 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1833_
timestamp 0
transform 1 0 850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1837_
timestamp 0
transform -1 0 30 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1841_
timestamp 0
transform -1 0 190 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1844_
timestamp 0
transform 1 0 2090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1848_
timestamp 0
transform 1 0 1190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1852_
timestamp 0
transform 1 0 170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1856_
timestamp 0
transform -1 0 310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1860_
timestamp 0
transform 1 0 890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1864_
timestamp 0
transform 1 0 510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1868_
timestamp 0
transform -1 0 1750 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__1872_
timestamp 0
transform -1 0 290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1875_
timestamp 0
transform -1 0 130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1879_
timestamp 0
transform 1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1883_
timestamp 0
transform 1 0 1350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1887_
timestamp 0
transform 1 0 630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__1891_
timestamp 0
transform 1 0 850 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__1895_
timestamp 0
transform -1 0 30 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__1899_
timestamp 0
transform 1 0 2570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform 1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform 1 0 2810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform -1 0 2670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 3290 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 4150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 1830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 2830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform 1 0 910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert15
timestamp 0
transform -1 0 3210 0 1 4570
box -6 -8 26 248
<< labels >>
flabel metal1 s 5142 2 5202 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 3217 4857 3223 4863 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 3177 4857 3183 4863 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 2637 4857 2643 4863 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 2437 4857 2443 4863 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 2277 4857 2283 4863 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 5176 4676 5184 4684 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal3 s 5176 4536 5184 4544 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 5176 4496 5184 4504 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal2 s 2597 -23 2603 -17 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 2637 -23 2643 -17 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 2677 -23 2683 -17 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 2717 -23 2723 -17 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 2877 -23 2883 -17 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -24 3716 -16 3724 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -24 3756 -16 3764 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal3 s -24 3796 -16 3804 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 5037 -23 5043 -17 7 FreeSans 16 270 0 0 Done_o
port 18 nsew
flabel metal2 s 4757 4857 4763 4863 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 4797 4857 4803 4863 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal2 s 4957 4857 4963 4863 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal2 s 4017 4857 4023 4863 3 FreeSans 16 90 0 0 clk
port 22 nsew
flabel metal2 s 5057 4857 5063 4863 3 FreeSans 16 90 0 0 reset
port 23 nsew
<< properties >>
string FIXED_BBOX -40 -40 5180 4860
<< end >>
