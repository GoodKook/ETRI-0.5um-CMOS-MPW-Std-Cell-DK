magic
tech scmos
magscale 1 2
timestamp 1727422626
<< nwell >>
rect -12 154 92 272
<< ntransistor >>
rect 20 14 24 34
rect 42 14 46 54
<< ptransistor >>
rect 20 206 24 246
rect 42 166 46 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 28 34
rect 40 14 42 54
rect 46 14 48 54
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 28 246
rect 40 166 42 246
rect 46 166 48 246
<< ndcontact >>
rect 6 14 18 34
rect 28 14 40 54
rect 48 14 60 54
<< pdcontact >>
rect 6 206 18 246
rect 28 166 40 246
rect 48 166 60 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 20 246 24 250
rect 42 246 46 250
rect 20 129 24 206
rect 42 160 46 166
rect 44 148 46 160
rect 16 117 24 129
rect 20 34 24 117
rect 44 60 46 72
rect 42 54 46 60
rect 20 10 24 14
rect 42 10 46 14
<< polycontact >>
rect 32 148 44 160
rect 4 117 16 129
rect 32 60 44 72
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 28 246 40 252
rect 6 160 14 206
rect 6 154 32 160
rect 31 148 32 154
rect 3 103 17 117
rect 31 72 37 148
rect 50 97 58 166
rect 43 83 58 97
rect 31 66 32 72
rect 10 60 32 66
rect 10 34 18 60
rect 50 54 58 83
rect 28 8 40 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect 3 103 17 117
rect 43 83 57 97
<< labels >>
rlabel metal1 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal1 -6 252 86 268 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 43 83 57 97 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
