magic
tech scmos
magscale 1 3
timestamp 1725342160
<< nwell >>
rect 110 110 330 330
<< diffusion >>
rect 76 376 364 394
rect 46 76 64 364
rect 151 291 289 309
rect 131 151 149 289
rect 196 196 244 244
rect 291 151 309 289
rect 151 131 289 149
rect 376 76 394 364
rect 76 46 364 64
<< pdiffusion >>
rect 195 244 245 245
rect 195 196 196 244
rect 244 196 245 244
rect 195 195 245 196
<< psubstratepdiff >>
rect 45 394 395 395
rect 45 376 76 394
rect 364 376 395 394
rect 45 375 395 376
rect 45 364 65 375
rect 45 76 46 364
rect 64 76 65 364
rect 375 364 395 375
rect 45 65 65 76
rect 375 76 376 364
rect 394 76 395 364
rect 375 65 395 76
rect 45 64 395 65
rect 45 46 76 64
rect 364 46 395 64
rect 45 45 395 46
<< nsubstratendiff >>
rect 130 309 310 310
rect 130 291 151 309
rect 289 291 310 309
rect 130 290 310 291
rect 130 289 150 290
rect 130 151 131 289
rect 149 151 150 289
rect 290 289 310 290
rect 130 150 150 151
rect 290 151 291 289
rect 309 151 310 289
rect 290 150 310 151
rect 130 149 310 150
rect 130 131 151 149
rect 289 131 310 149
rect 130 130 310 131
<< metal1 >>
rect 45 375 395 395
rect 45 65 65 375
rect 130 290 310 310
rect 130 150 150 290
rect 195 195 245 245
rect 290 150 310 290
rect 130 130 310 150
rect 375 65 395 375
rect 45 45 395 65
<< end >>
