magic
tech scmos
magscale 1 30
timestamp 1739362888
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal2 >>
rect 59800 130950 60120 145940
rect 62500 132310 62820 145940
rect 76000 134050 76320 145940
rect 89500 135700 89820 145870
rect 103000 137240 103320 145940
rect 116500 138080 116820 145940
rect 116500 137760 122930 138080
rect 103000 136920 122340 137240
rect 89500 135380 121750 135700
rect 76000 133730 121130 134050
rect 62500 131990 120550 132310
rect 59800 130630 119320 130950
rect 44060 129880 53820 130200
rect 119000 128970 119320 130630
rect 120230 129410 120550 131990
rect 120330 129360 120435 129410
rect 120810 129380 121130 133730
rect 120930 129360 121035 129380
rect 121430 129290 121750 135380
rect 122020 129370 122340 136920
rect 122130 129338 122235 129370
rect 122610 129360 122930 137760
rect 130000 137640 130320 145940
rect 123220 137320 130320 137640
rect 123220 129370 123540 137320
rect 123880 134180 144710 134500
rect 122730 129318 122835 129360
rect 123330 129328 123435 129370
rect 123880 129350 124200 134180
rect 127750 132450 143620 132770
rect 123930 129318 124035 129350
rect 127750 129320 128070 132450
rect 128960 130890 141910 131210
rect 128960 129330 129280 130890
rect 127830 129308 127935 129320
rect 119130 128967 119235 128970
rect 44060 116380 52350 116700
rect 44060 102880 56050 103200
rect 141590 103320 141910 130890
rect 143300 116820 143620 132450
rect 144390 130320 144710 134180
rect 144390 130000 145940 130320
rect 143300 116500 145940 116820
rect 141590 103000 145940 103320
rect 142900 86800 145940 87120
rect 44060 75880 56050 76200
rect 140890 73300 145940 73620
rect 44060 62380 47590 62700
rect 90930 59900 91035 59901
rect 81210 56720 81530 59880
rect 59800 44060 60120 56400
rect 85440 54980 85760 59870
rect 73300 44060 73620 54670
rect 87470 49050 87790 59860
rect 86800 48730 87790 49050
rect 88160 49050 88480 59870
rect 88830 59860 88935 59865
rect 88830 51500 89150 59860
rect 90830 53550 91150 59900
rect 138700 59800 145940 60120
rect 86800 44060 87120 48730
rect 100300 44060 100620 48730
rect 113800 44060 114120 51170
rect 127300 44070 127620 53230
rect 136700 46330 141120 46650
rect 140800 44060 141120 46330
<< m3contact >>
rect 53820 129560 54140 130200
rect 52350 116060 52670 116700
rect 56050 102880 56370 103520
rect 142580 86800 142900 87500
rect 56050 75880 56370 76520
rect 140580 73300 140890 74000
rect 47590 62380 47910 63020
rect 59800 56400 60460 56720
rect 80870 56400 81530 56720
rect 73300 54670 73970 54980
rect 85090 54670 85760 54980
rect 138380 59800 138700 60460
rect 90830 53230 91470 53550
rect 127050 53230 127620 53550
rect 88830 51170 89470 51500
rect 113500 51170 114120 51500
rect 88160 48730 88800 49050
rect 99980 48730 100620 49050
rect 136380 46330 136700 46960
<< metal3 >>
rect 52350 112500 52670 116060
rect 53820 113180 54140 129560
rect 130790 119460 142900 119580
rect 132040 119250 142900 119460
rect 131945 115380 140890 115615
rect 131820 115260 140890 115380
rect 131920 115080 138700 115090
rect 131820 114960 138700 115080
rect 131920 114770 138700 114960
rect 53820 112980 58140 113180
rect 53820 112860 58260 112980
rect 52350 112380 58140 112500
rect 52350 112260 58260 112380
rect 52350 112180 58140 112260
rect 47590 111780 58160 111870
rect 47590 111660 58260 111780
rect 47590 111550 58160 111660
rect 47590 63020 47910 111550
rect 56050 104580 58110 104660
rect 56050 104460 58260 104580
rect 56050 104340 58110 104460
rect 56050 103520 56370 104340
rect 56050 100380 58140 100420
rect 56050 100260 59340 100380
rect 56050 100100 58140 100260
rect 56050 76520 56370 100100
rect 131940 79380 136700 79490
rect 131810 79260 136700 79380
rect 131940 79170 136700 79260
rect 60460 56400 80870 56720
rect 73970 54670 85090 54980
rect 91470 53230 127050 53550
rect 89470 51170 113500 51500
rect 88800 48730 99980 49050
rect 136380 46960 136700 79170
rect 138380 60460 138700 114770
rect 140580 74000 140890 115260
rect 142580 87500 142900 119250
use PIC  AUX
timestamp 1555597840
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1555597840
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1555597840
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1555597840
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1555597840
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1555597840
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_0
timestamp 1555597840
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1555597840
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1739356964
transform 1 0 59190 0 1 60120
box -1050 -360 72750 69345
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0
timestamp 1555597840
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1555597840
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1555597840
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1555597840
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1555597840
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1555597840
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1555597840
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1555597840
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PCORNER  PCORNER_0
timestamp 1555597840
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1555597840
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1555597840
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1555597840
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY
timestamp 1555597840
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PVDD  VDD
timestamp 1555597840
transform 0 1 18900 -1 0 101000
box 0 -9150 12000 25300
use POB4  VLD
timestamp 1555597840
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PVSS  VSS
timestamp 1555597840
transform 0 -1 171100 1 0 89000
box 0 -9150 12000 25300
use PIC  XIN_0
timestamp 1555597840
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1555597840
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1555597840
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1555597840
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use POB4  XOUT_0
timestamp 1555597840
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB4  XOUT_1
timestamp 1555597840
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB4  XOUT_2
timestamp 1555597840
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB4  XOUT_3
timestamp 1555597840
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1555597840
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1555597840
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1555597840
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1555597840
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use POB4  YOUT_0
timestamp 1555597840
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use POB4  YOUT_1
timestamp 1555597840
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB4  YOUT_2
timestamp 1555597840
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB4  YOUT_3
timestamp 1555597840
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
<< end >>
