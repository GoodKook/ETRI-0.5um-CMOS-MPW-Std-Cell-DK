magic
tech scmos
magscale 1 2
timestamp 1727423652
<< nwell >>
rect -12 154 132 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 166 24 246
rect 30 166 34 246
rect 60 166 64 246
rect 70 166 74 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 44 40 54
rect 24 14 26 44
rect 38 14 40 44
rect 44 14 46 54
rect 58 14 60 54
rect 64 26 66 54
rect 78 26 80 54
rect 64 14 80 26
rect 84 14 86 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 30 246
rect 34 166 36 246
rect 58 166 60 246
rect 64 166 70 246
rect 74 166 76 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 44
rect 46 14 58 54
rect 66 26 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 166 18 246
rect 36 166 58 246
rect 76 166 88 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 30 246 34 250
rect 60 246 64 250
rect 70 246 74 250
rect 20 162 24 166
rect 10 158 24 162
rect 30 162 34 166
rect 30 158 44 162
rect 10 83 16 158
rect 40 123 44 158
rect 36 111 44 123
rect 17 71 24 83
rect 20 54 24 71
rect 40 54 44 111
rect 60 123 64 166
rect 70 162 74 166
rect 70 158 88 162
rect 84 111 88 158
rect 60 54 64 111
rect 80 109 88 111
rect 80 97 83 109
rect 80 54 84 97
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 24 111 36 123
rect 5 71 17 83
rect 60 111 72 123
rect 83 97 95 109
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 6 246 18 252
rect 76 246 88 252
rect 23 123 37 137
rect 46 97 54 166
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
rect 46 72 54 83
rect 46 64 74 72
rect 6 54 58 56
rect 68 54 74 64
rect 18 50 46 54
rect 58 14 86 20
rect 26 8 38 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m1p >>
rect 23 123 37 137
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal1 -6 252 126 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal1 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal1 83 83 97 97 0 C
port 2 nsew signal input
rlabel metal1 63 123 77 137 0 D
port 3 nsew signal input
rlabel metal1 43 83 57 97 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
