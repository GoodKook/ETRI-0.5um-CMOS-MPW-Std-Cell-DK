magic
tech scmos
magscale 1 2
timestamp 1702508443
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 44
rect 38 14 42 54
rect 58 14 62 54
<< ptransistor >>
rect 18 186 22 246
rect 38 166 42 246
rect 58 166 62 246
<< ndiffusion >>
rect 24 53 38 54
rect 16 14 18 44
rect 22 14 24 44
rect 36 14 38 53
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
<< pdiffusion >>
rect 16 186 18 246
rect 22 186 24 246
rect 36 168 38 246
rect 24 166 38 168
rect 42 168 44 246
rect 56 168 58 246
rect 42 166 58 168
rect 62 166 64 246
<< ndcontact >>
rect 4 14 16 44
rect 24 14 36 53
rect 44 14 56 54
rect 64 14 76 54
<< pdcontact >>
rect 4 186 16 246
rect 24 168 36 246
rect 44 168 56 246
rect 64 166 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 44 22 186
rect 38 164 42 166
rect 58 164 62 166
rect 38 160 62 164
rect 38 152 42 160
rect 38 60 42 68
rect 38 56 62 60
rect 38 54 42 56
rect 58 54 62 56
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 6 117 18 129
rect 31 140 43 152
rect 31 68 43 80
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 24 246 36 252
rect 64 246 76 252
rect 4 162 12 186
rect 4 156 37 162
rect 31 152 37 156
rect 31 80 39 140
rect 49 117 56 168
rect 49 103 60 117
rect 31 65 37 68
rect 4 59 37 65
rect 4 44 12 59
rect 49 54 56 103
rect 24 8 36 14
rect 64 8 76 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 5 103 19 117
rect 60 103 74 117
<< metal2 >>
rect 66 117 74 134
rect 6 86 14 103
<< m1p >>
rect -6 252 86 268
rect -6 -8 86 8
<< m2p >>
rect 66 119 74 134
rect 6 86 14 101
<< labels >>
rlabel metal2 10 89 10 89 1 A
port 1 n signal input
rlabel metal2 70 131 70 131 3 Y
port 2 n signal output
rlabel metal1 -6 252 86 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
