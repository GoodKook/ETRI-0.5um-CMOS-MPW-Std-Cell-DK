magic
tech scmos
magscale 3 2
timestamp 1724157349
<< checkpaint >>
rect -36 241 240 519
rect -36 41 518 241
rect -40 -35 518 41
rect -40 -40 41 -35
<< metal1 >>
rect 99 200 100 201
rect 101 200 120 201
rect 93 199 123 200
rect 64 198 69 199
rect 88 198 125 199
rect 63 197 72 198
rect 84 197 127 198
rect 61 196 129 197
rect 61 195 130 196
rect 60 194 131 195
rect 60 193 133 194
rect 59 192 97 193
rect 104 192 134 193
rect 255 192 259 193
rect 265 192 269 193
rect 294 192 299 193
rect 306 192 308 193
rect 319 192 321 193
rect 344 192 347 193
rect 354 192 357 193
rect 362 192 368 193
rect 374 192 376 193
rect 383 192 385 193
rect 391 192 393 193
rect 60 191 68 192
rect 76 191 96 192
rect 107 191 135 192
rect 184 191 189 192
rect 196 191 201 192
rect 207 191 213 192
rect 223 191 226 192
rect 238 191 243 192
rect 255 191 260 192
rect 60 190 66 191
rect 78 190 99 191
rect 112 190 136 191
rect 183 190 190 191
rect 195 190 202 191
rect 50 189 55 190
rect 62 189 63 190
rect 80 189 102 190
rect 117 189 137 190
rect 182 189 191 190
rect 194 189 202 190
rect 206 189 214 191
rect 222 190 226 191
rect 237 190 244 191
rect 221 189 226 190
rect 48 188 57 189
rect 68 188 71 189
rect 81 188 105 189
rect 125 188 138 189
rect 181 188 185 189
rect 47 187 58 188
rect 65 187 73 188
rect 81 187 109 188
rect 129 187 139 188
rect 182 187 185 188
rect 188 187 191 189
rect 47 186 59 187
rect 63 186 75 187
rect 46 185 75 186
rect 81 186 119 187
rect 132 186 140 187
rect 187 186 191 187
rect 193 188 197 189
rect 193 186 196 188
rect 200 186 203 189
rect 205 188 209 189
rect 205 187 208 188
rect 211 187 215 189
rect 220 188 226 189
rect 236 189 245 190
rect 220 187 225 188
rect 236 187 239 189
rect 242 187 245 189
rect 211 186 214 187
rect 219 186 225 187
rect 240 186 245 187
rect 254 186 260 191
rect 264 190 269 192
rect 292 191 300 192
rect 291 190 301 191
rect 305 190 309 192
rect 318 190 322 192
rect 263 188 269 190
rect 290 189 295 190
rect 298 189 302 190
rect 271 188 273 189
rect 279 188 281 189
rect 262 186 268 188
rect 270 187 274 188
rect 278 187 281 188
rect 81 185 123 186
rect 135 185 140 186
rect 186 185 190 186
rect 192 185 196 186
rect 45 183 76 185
rect 81 184 126 185
rect 137 184 140 185
rect 185 184 189 185
rect 44 182 76 183
rect 80 183 129 184
rect 139 183 141 184
rect 184 183 188 184
rect 80 182 132 183
rect 183 182 187 183
rect 43 181 75 182
rect 80 181 135 182
rect 182 181 186 182
rect 42 180 75 181
rect 81 180 137 181
rect 181 180 185 181
rect 192 180 195 185
rect 199 184 203 186
rect 210 185 214 186
rect 218 185 221 186
rect 209 184 213 185
rect 217 184 220 185
rect 222 184 225 186
rect 239 185 244 186
rect 239 184 243 185
rect 199 182 202 184
rect 208 183 212 184
rect 216 183 219 184
rect 221 183 224 184
rect 207 182 211 183
rect 198 181 202 182
rect 206 181 210 182
rect 215 181 226 183
rect 227 181 233 184
rect 240 183 244 184
rect 234 181 237 182
rect 241 181 245 183
rect 253 181 256 186
rect 198 180 201 181
rect 205 180 209 181
rect 215 180 225 181
rect 234 180 238 181
rect 241 180 244 181
rect 41 179 74 180
rect 82 179 140 180
rect 181 179 190 180
rect 192 179 201 180
rect 39 178 73 179
rect 84 178 104 179
rect 108 178 142 179
rect 180 178 190 179
rect 193 178 200 179
rect 38 177 54 178
rect 56 177 71 178
rect 85 177 105 178
rect 110 177 143 178
rect 180 177 189 178
rect 194 177 198 178
rect 204 177 213 180
rect 221 179 224 180
rect 235 179 244 180
rect 252 180 256 181
rect 257 184 260 186
rect 261 184 264 186
rect 257 181 263 184
rect 265 183 268 186
rect 220 177 223 179
rect 235 178 243 179
rect 237 177 241 178
rect 252 177 255 180
rect 257 179 262 181
rect 257 177 261 179
rect 264 178 267 183
rect 271 182 274 187
rect 277 186 281 187
rect 289 187 293 189
rect 299 188 302 189
rect 305 188 308 190
rect 310 188 313 189
rect 319 188 320 189
rect 324 188 326 189
rect 328 188 331 189
rect 343 188 348 192
rect 353 191 358 192
rect 361 191 371 192
rect 352 189 357 191
rect 361 190 372 191
rect 361 189 364 190
rect 368 189 372 190
rect 299 187 301 188
rect 305 187 314 188
rect 318 187 321 188
rect 289 186 292 187
rect 277 185 280 186
rect 276 184 280 185
rect 276 183 279 184
rect 275 182 279 183
rect 271 181 278 182
rect 288 181 292 186
rect 304 186 314 187
rect 304 185 308 186
rect 311 185 315 186
rect 317 185 321 187
rect 323 187 333 188
rect 323 186 328 187
rect 329 186 333 187
rect 342 186 348 188
rect 351 187 357 189
rect 323 185 327 186
rect 304 182 307 185
rect 311 182 314 185
rect 317 182 320 185
rect 323 183 326 185
rect 298 181 301 182
rect 272 180 278 181
rect 289 180 293 181
rect 297 180 301 181
rect 303 181 307 182
rect 272 178 277 180
rect 289 179 300 180
rect 290 178 299 179
rect 263 177 266 178
rect 272 177 276 178
rect 291 177 298 178
rect 303 177 306 181
rect 310 180 314 182
rect 316 181 320 182
rect 310 177 313 180
rect 316 177 319 181
rect 322 180 326 183
rect 330 182 334 186
rect 342 183 345 186
rect 346 183 348 186
rect 350 186 357 187
rect 350 185 353 186
rect 354 185 357 186
rect 360 187 364 189
rect 369 187 372 189
rect 360 186 363 187
rect 368 186 372 187
rect 349 183 352 185
rect 330 181 333 182
rect 329 180 333 181
rect 322 179 327 180
rect 328 179 332 180
rect 341 179 344 183
rect 321 178 331 179
rect 340 178 344 179
rect 346 182 352 183
rect 346 180 351 182
rect 353 180 356 185
rect 360 184 371 186
rect 359 183 369 184
rect 374 183 377 192
rect 382 191 386 192
rect 381 189 386 191
rect 390 191 394 192
rect 390 190 393 191
rect 380 187 386 189
rect 389 189 393 190
rect 389 187 392 189
rect 379 185 382 187
rect 378 184 382 185
rect 378 183 381 184
rect 359 182 363 183
rect 374 182 381 183
rect 383 183 386 187
rect 388 185 391 187
rect 387 183 390 185
rect 359 180 362 182
rect 346 178 350 180
rect 321 177 325 178
rect 326 177 330 178
rect 340 177 343 178
rect 346 177 349 178
rect 352 177 355 180
rect 358 178 362 180
rect 374 180 380 182
rect 383 181 389 183
rect 374 178 379 180
rect 383 179 388 181
rect 358 177 361 178
rect 374 177 378 178
rect 383 177 387 179
rect 36 176 50 177
rect 55 176 70 177
rect 87 176 105 177
rect 112 176 144 177
rect 272 176 275 177
rect 35 175 47 176
rect 53 175 69 176
rect 88 175 105 176
rect 115 175 145 176
rect 271 175 275 176
rect 33 174 45 175
rect 51 174 69 175
rect 89 174 106 175
rect 118 174 146 175
rect 31 173 43 174
rect 50 173 68 174
rect 75 173 82 174
rect 90 173 107 174
rect 122 173 146 174
rect 269 174 274 175
rect 269 173 273 174
rect 321 173 324 177
rect 29 172 42 173
rect 49 172 69 173
rect 27 171 45 172
rect 25 170 46 171
rect 48 170 69 172
rect 75 172 84 173
rect 91 172 109 173
rect 125 172 147 173
rect 75 171 85 172
rect 92 171 110 172
rect 128 171 147 172
rect 24 169 46 170
rect 47 169 69 170
rect 76 169 86 171
rect 92 170 112 171
rect 130 170 147 171
rect 93 169 116 170
rect 132 169 148 170
rect 23 167 70 169
rect 76 168 87 169
rect 94 168 120 169
rect 133 168 148 169
rect 77 167 88 168
rect 94 167 124 168
rect 135 167 148 168
rect 22 165 70 167
rect 23 164 29 165
rect 30 164 70 165
rect 23 163 27 164
rect 29 163 70 164
rect 28 162 70 163
rect 27 161 70 162
rect 76 166 88 167
rect 95 166 126 167
rect 136 166 148 167
rect 76 163 89 166
rect 95 165 128 166
rect 137 165 148 166
rect 96 164 129 165
rect 139 164 149 165
rect 96 163 131 164
rect 140 163 149 164
rect 76 161 90 163
rect 97 162 132 163
rect 141 162 149 163
rect 98 161 133 162
rect 142 161 149 162
rect 26 160 69 161
rect 25 158 69 160
rect 76 160 91 161
rect 99 160 134 161
rect 76 159 92 160
rect 100 159 136 160
rect 143 159 149 161
rect 75 158 92 159
rect 102 158 137 159
rect 144 158 148 159
rect 26 157 68 158
rect 75 157 93 158
rect 105 157 138 158
rect 26 156 67 157
rect 75 156 95 157
rect 111 156 139 157
rect 145 156 148 158
rect 27 155 67 156
rect 74 155 96 156
rect 115 155 140 156
rect 146 155 148 156
rect 185 155 193 156
rect 27 154 44 155
rect 46 154 66 155
rect 74 154 99 155
rect 118 154 140 155
rect 28 153 43 154
rect 29 152 41 153
rect 47 152 65 154
rect 74 153 103 154
rect 120 153 141 154
rect 183 153 193 155
rect 73 152 108 153
rect 123 152 141 153
rect 31 151 36 152
rect 46 151 64 152
rect 73 151 111 152
rect 125 151 141 152
rect 182 152 192 153
rect 42 150 63 151
rect 72 150 114 151
rect 126 150 142 151
rect 36 149 63 150
rect 71 149 116 150
rect 127 149 142 150
rect 31 148 62 149
rect 71 148 118 149
rect 128 148 142 149
rect 182 148 188 152
rect 194 151 200 156
rect 301 154 305 156
rect 300 153 304 154
rect 299 151 304 153
rect 309 151 328 156
rect 298 149 303 151
rect 213 148 215 149
rect 251 148 254 149
rect 270 148 274 149
rect 31 147 61 148
rect 70 147 120 148
rect 129 147 142 148
rect 31 146 60 147
rect 69 146 121 147
rect 31 145 59 146
rect 68 145 122 146
rect 130 145 142 147
rect 32 144 58 145
rect 68 144 123 145
rect 131 144 142 145
rect 179 144 192 148
rect 32 143 57 144
rect 67 143 123 144
rect 33 142 55 143
rect 65 142 90 143
rect 97 142 124 143
rect 132 142 142 144
rect 33 141 53 142
rect 64 141 89 142
rect 99 141 124 142
rect 133 141 142 142
rect 34 140 51 141
rect 63 140 88 141
rect 100 140 125 141
rect 133 140 141 141
rect 34 139 48 140
rect 62 139 88 140
rect 101 139 125 140
rect 35 138 45 139
rect 60 138 88 139
rect 102 138 126 139
rect 35 137 42 138
rect 58 137 87 138
rect 103 137 126 138
rect 134 137 141 140
rect 36 136 39 137
rect 56 136 87 137
rect 94 136 95 137
rect 54 135 87 136
rect 93 135 96 136
rect 104 135 126 137
rect 51 134 86 135
rect 93 134 97 135
rect 49 133 86 134
rect 92 133 97 134
rect 105 134 126 135
rect 135 136 141 137
rect 135 134 140 136
rect 105 133 125 134
rect 47 132 85 133
rect 92 132 98 133
rect 45 131 85 132
rect 91 131 98 132
rect 106 131 125 133
rect 136 132 139 134
rect 136 131 138 132
rect 43 130 84 131
rect 91 130 99 131
rect 42 129 84 130
rect 90 129 99 130
rect 106 130 124 131
rect 136 130 137 131
rect 106 129 123 130
rect 41 128 83 129
rect 40 127 82 128
rect 90 127 100 129
rect 39 126 81 127
rect 89 126 100 127
rect 107 128 123 129
rect 182 128 188 144
rect 194 128 200 148
rect 205 147 210 148
rect 211 147 218 148
rect 205 146 218 147
rect 241 146 246 148
rect 248 147 256 148
rect 268 147 277 148
rect 247 146 257 147
rect 266 146 278 147
rect 297 146 302 149
rect 205 143 217 146
rect 241 145 258 146
rect 265 145 279 146
rect 296 145 302 146
rect 309 145 315 151
rect 241 144 259 145
rect 264 144 280 145
rect 241 143 248 144
rect 253 143 260 144
rect 264 143 270 144
rect 205 142 212 143
rect 205 140 211 142
rect 241 140 247 143
rect 254 141 260 143
rect 255 140 260 141
rect 263 140 269 143
rect 275 142 281 144
rect 276 140 281 142
rect 296 140 301 145
rect 205 128 210 140
rect 241 137 246 140
rect 255 137 261 140
rect 263 137 282 140
rect 295 137 301 140
rect 241 134 247 137
rect 255 135 260 137
rect 241 133 248 134
rect 254 133 260 135
rect 263 136 281 137
rect 263 133 269 136
rect 276 134 277 135
rect 241 132 249 133
rect 253 132 259 133
rect 241 131 259 132
rect 264 132 271 133
rect 275 132 281 134
rect 296 132 301 137
rect 309 140 326 145
rect 264 131 280 132
rect 296 131 302 132
rect 241 130 258 131
rect 265 130 280 131
rect 107 127 122 128
rect 107 126 121 127
rect 39 125 80 126
rect 89 125 101 126
rect 38 124 79 125
rect 88 124 101 125
rect 107 125 120 126
rect 130 125 131 126
rect 107 124 119 125
rect 129 124 131 125
rect 38 123 78 124
rect 37 122 77 123
rect 87 122 101 124
rect 37 121 76 122
rect 86 121 101 122
rect 108 123 117 124
rect 128 123 132 124
rect 108 122 116 123
rect 127 122 131 123
rect 108 121 114 122
rect 126 121 132 122
rect 216 121 239 124
rect 37 120 75 121
rect 85 120 101 121
rect 36 119 74 120
rect 84 119 101 120
rect 107 120 112 121
rect 125 120 132 121
rect 217 120 238 121
rect 241 120 246 130
rect 247 129 257 130
rect 266 129 279 130
rect 249 128 256 129
rect 268 128 277 129
rect 297 128 302 131
rect 309 128 315 140
rect 332 128 338 156
rect 343 155 360 156
rect 376 155 382 156
rect 391 155 394 156
rect 343 154 362 155
rect 373 154 384 155
rect 391 154 395 155
rect 343 153 364 154
rect 372 153 385 154
rect 391 153 396 154
rect 343 151 365 153
rect 371 151 386 153
rect 392 152 396 153
rect 392 151 397 152
rect 343 145 349 151
rect 357 150 366 151
rect 359 149 366 150
rect 360 146 366 149
rect 370 147 376 151
rect 381 150 387 151
rect 382 147 387 150
rect 393 150 397 151
rect 393 148 398 150
rect 359 145 366 146
rect 371 146 376 147
rect 381 146 387 147
rect 371 145 377 146
rect 380 145 386 146
rect 394 145 399 148
rect 343 143 365 145
rect 372 144 385 145
rect 343 142 364 143
rect 373 142 384 144
rect 394 143 400 145
rect 343 141 362 142
rect 372 141 386 142
rect 343 140 360 141
rect 371 140 377 141
rect 380 140 387 141
rect 343 139 350 140
rect 351 139 360 140
rect 370 139 376 140
rect 381 139 387 140
rect 343 128 349 139
rect 354 138 361 139
rect 355 137 362 138
rect 355 136 363 137
rect 356 135 364 136
rect 357 134 364 135
rect 370 134 375 139
rect 357 133 365 134
rect 358 132 365 133
rect 370 133 376 134
rect 382 133 388 139
rect 395 133 400 143
rect 370 132 377 133
rect 381 132 387 133
rect 359 131 366 132
rect 371 131 387 132
rect 394 132 400 133
rect 360 129 367 131
rect 372 130 386 131
rect 373 129 385 130
rect 361 128 368 129
rect 374 128 383 129
rect 394 128 399 132
rect 298 127 302 128
rect 298 125 303 127
rect 393 126 398 128
rect 393 125 397 126
rect 299 124 304 125
rect 300 122 304 124
rect 392 124 397 125
rect 392 123 396 124
rect 391 122 396 123
rect 301 121 305 122
rect 302 120 305 121
rect 391 121 395 122
rect 391 120 394 121
rect 107 119 110 120
rect 124 119 132 120
rect 36 118 72 119
rect 83 118 101 119
rect 122 118 132 119
rect 36 117 71 118
rect 82 117 101 118
rect 121 117 132 118
rect 36 116 69 117
rect 80 116 101 117
rect 119 116 132 117
rect 36 115 67 116
rect 79 115 101 116
rect 118 115 132 116
rect 36 114 65 115
rect 77 114 101 115
rect 116 114 132 115
rect 36 113 62 114
rect 76 113 101 114
rect 114 113 132 114
rect 36 112 60 113
rect 74 112 100 113
rect 112 112 131 113
rect 36 111 58 112
rect 72 111 100 112
rect 109 111 131 112
rect 36 110 56 111
rect 70 110 100 111
rect 106 110 131 111
rect 36 109 55 110
rect 68 109 100 110
rect 102 109 131 110
rect 37 108 53 109
rect 66 108 131 109
rect 37 106 52 108
rect 65 107 130 108
rect 63 106 130 107
rect 37 105 51 106
rect 62 105 130 106
rect 38 104 51 105
rect 60 104 129 105
rect 38 103 50 104
rect 59 103 129 104
rect 39 102 50 103
rect 58 102 128 103
rect 39 101 49 102
rect 40 99 49 101
rect 57 101 83 102
rect 85 101 128 102
rect 57 100 82 101
rect 85 100 127 101
rect 56 99 80 100
rect 84 99 127 100
rect 41 97 49 99
rect 55 98 78 99
rect 55 97 77 98
rect 83 97 126 99
rect 42 96 49 97
rect 54 96 75 97
rect 82 96 125 97
rect 43 95 48 96
rect 54 95 74 96
rect 81 95 124 96
rect 44 94 48 95
rect 45 93 48 94
rect 46 92 48 93
rect 53 94 73 95
rect 81 94 100 95
rect 101 94 123 95
rect 53 93 72 94
rect 80 93 98 94
rect 100 93 123 94
rect 173 94 249 105
rect 262 94 340 105
rect 351 104 425 105
rect 351 103 428 104
rect 351 102 429 103
rect 351 101 430 102
rect 351 100 431 101
rect 351 99 432 100
rect 351 94 433 99
rect 173 93 196 94
rect 53 92 71 93
rect 79 92 97 93
rect 100 92 122 93
rect 47 91 48 92
rect 52 91 70 92
rect 78 91 96 92
rect 99 91 121 92
rect 52 89 69 91
rect 78 90 95 91
rect 99 90 120 91
rect 77 89 94 90
rect 99 89 119 90
rect 52 87 68 89
rect 77 88 93 89
rect 99 88 118 89
rect 173 88 197 93
rect 76 87 93 88
rect 98 87 117 88
rect 173 87 196 88
rect 52 84 67 87
rect 76 85 92 87
rect 98 86 116 87
rect 173 86 197 87
rect 98 85 115 86
rect 53 82 66 84
rect 54 81 66 82
rect 75 83 91 85
rect 98 84 113 85
rect 98 83 112 84
rect 75 81 90 83
rect 55 79 66 81
rect 56 78 66 79
rect 57 77 66 78
rect 58 76 66 77
rect 60 75 66 76
rect 74 80 90 81
rect 98 82 111 83
rect 98 81 109 82
rect 98 80 108 81
rect 74 75 89 80
rect 98 79 107 80
rect 98 78 106 79
rect 98 77 105 78
rect 98 76 104 77
rect 173 76 249 86
rect 98 75 103 76
rect 61 74 66 75
rect 63 73 67 74
rect 64 72 67 73
rect 65 71 67 72
rect 75 71 89 75
rect 99 74 103 75
rect 173 75 198 76
rect 99 73 102 74
rect 99 71 101 73
rect 66 70 67 71
rect 76 69 89 71
rect 77 68 89 69
rect 78 67 89 68
rect 173 69 197 75
rect 173 68 196 69
rect 173 67 197 68
rect 78 66 90 67
rect 79 65 90 66
rect 80 64 90 65
rect 81 63 90 64
rect 173 63 249 67
rect 82 62 91 63
rect 83 61 91 62
rect 174 61 249 63
rect 84 60 91 61
rect 175 60 249 61
rect 86 59 92 60
rect 176 59 249 60
rect 88 58 92 59
rect 177 58 249 59
rect 90 57 93 58
rect 179 57 249 58
rect 289 57 313 94
rect 351 57 375 94
rect 409 80 433 94
rect 384 79 433 80
rect 383 78 411 79
rect 384 77 412 78
rect 385 76 413 77
rect 386 75 415 76
rect 388 74 416 75
rect 389 73 417 74
rect 390 72 418 73
rect 391 71 419 72
rect 392 70 421 71
rect 394 69 422 70
rect 395 68 423 69
rect 396 67 424 68
rect 397 66 426 67
rect 399 65 427 66
rect 400 64 428 65
rect 401 63 429 64
rect 402 62 431 63
rect 404 61 432 62
rect 405 60 433 61
rect 406 59 434 60
rect 407 58 435 59
rect 408 57 437 58
rect 450 57 474 105
rect 410 56 438 57
rect 411 55 439 56
rect 412 54 441 55
rect 413 53 441 54
rect 456 45 461 46
rect 94 44 99 45
rect 4 43 12 44
rect 14 43 22 44
rect 24 43 32 44
rect 35 43 41 44
rect 43 43 52 44
rect 55 43 63 44
rect 64 43 70 44
rect 77 43 84 44
rect 91 43 102 44
rect 112 43 121 44
rect 123 43 132 44
rect 135 43 148 44
rect 152 43 166 44
rect 178 43 187 45
rect 5 42 11 43
rect 16 42 20 43
rect 25 42 31 43
rect 6 36 10 42
rect 15 41 18 42
rect 26 41 31 42
rect 15 40 17 41
rect 27 40 31 41
rect 36 42 40 43
rect 45 42 51 43
rect 57 42 62 43
rect 66 42 71 43
rect 79 42 83 43
rect 89 42 94 43
rect 98 42 102 43
rect 113 42 119 43
rect 125 42 130 43
rect 36 41 39 42
rect 36 40 38 41
rect 14 39 16 40
rect 27 39 32 40
rect 13 38 15 39
rect 28 38 32 39
rect 35 38 37 40
rect 12 37 14 38
rect 28 37 33 38
rect 11 36 14 37
rect 29 36 33 37
rect 34 36 36 38
rect 6 34 15 36
rect 29 35 35 36
rect 6 28 10 34
rect 11 33 16 34
rect 12 31 17 33
rect 13 30 18 31
rect 14 29 19 30
rect 14 28 20 29
rect 5 27 11 28
rect 15 27 21 28
rect 30 27 35 35
rect 45 33 50 42
rect 46 30 50 33
rect 58 39 61 42
rect 67 41 72 42
rect 67 40 73 41
rect 67 39 74 40
rect 58 32 60 39
rect 67 38 75 39
rect 58 31 61 32
rect 58 30 60 31
rect 46 29 51 30
rect 57 29 60 30
rect 47 28 52 29
rect 56 28 60 29
rect 67 28 69 38
rect 70 37 75 38
rect 71 36 76 37
rect 72 35 77 36
rect 73 34 78 35
rect 74 33 79 34
rect 80 33 82 42
rect 88 41 92 42
rect 99 41 102 42
rect 87 40 91 41
rect 100 40 102 41
rect 86 39 91 40
rect 101 39 102 40
rect 114 41 119 42
rect 86 37 90 39
rect 85 33 90 37
rect 114 37 118 41
rect 126 37 130 42
rect 114 35 130 37
rect 95 34 104 35
rect 96 33 104 34
rect 114 34 119 35
rect 125 34 130 35
rect 74 32 82 33
rect 75 31 82 32
rect 76 30 82 31
rect 86 32 90 33
rect 86 30 91 32
rect 77 29 82 30
rect 87 29 92 30
rect 47 27 59 28
rect 66 27 70 28
rect 78 27 82 29
rect 88 28 92 29
rect 89 27 94 28
rect 98 27 102 33
rect 114 28 118 34
rect 126 28 130 34
rect 137 42 142 43
rect 145 42 149 43
rect 137 37 141 42
rect 147 40 149 42
rect 147 39 148 40
rect 146 37 147 38
rect 137 36 142 37
rect 145 36 147 37
rect 137 34 147 36
rect 137 28 141 34
rect 145 33 147 34
rect 146 32 147 33
rect 154 36 159 43
rect 162 42 166 43
rect 164 40 166 42
rect 175 40 191 42
rect 175 39 190 40
rect 193 39 196 45
rect 212 44 230 45
rect 211 42 231 44
rect 212 41 230 42
rect 245 41 259 44
rect 262 41 266 45
rect 296 44 299 45
rect 279 41 293 43
rect 180 38 186 39
rect 163 37 165 38
rect 177 37 188 38
rect 162 36 165 37
rect 154 34 165 36
rect 176 36 189 37
rect 193 36 199 39
rect 226 37 230 41
rect 250 39 254 41
rect 249 38 255 39
rect 248 37 255 38
rect 258 37 266 41
rect 278 40 293 41
rect 284 38 288 40
rect 209 36 233 37
rect 247 36 257 37
rect 176 35 181 36
rect 184 35 190 36
rect 175 34 180 35
rect 186 34 190 35
rect 148 29 150 31
rect 147 28 150 29
rect 154 28 159 34
rect 163 33 165 34
rect 176 33 181 34
rect 184 33 190 34
rect 163 32 164 33
rect 176 32 189 33
rect 178 31 188 32
rect 166 30 167 31
rect 165 29 167 30
rect 179 29 182 30
rect 193 29 196 36
rect 208 35 234 36
rect 246 35 258 36
rect 209 34 234 35
rect 244 34 251 35
rect 253 34 260 35
rect 209 33 233 34
rect 244 33 250 34
rect 255 33 259 34
rect 219 31 222 33
rect 245 32 248 33
rect 257 32 258 33
rect 212 30 230 31
rect 164 28 167 29
rect 114 27 119 28
rect 125 27 131 28
rect 137 27 142 28
rect 146 27 149 28
rect 154 27 160 28
rect 163 27 167 28
rect 178 27 183 29
rect 211 28 230 30
rect 212 27 230 28
rect 4 26 12 27
rect 16 26 22 27
rect 28 26 37 27
rect 48 26 58 27
rect 65 26 72 27
rect 79 26 82 27
rect 90 26 102 27
rect 112 26 121 27
rect 123 26 132 27
rect 135 26 149 27
rect 152 26 166 27
rect 178 26 196 27
rect 51 25 56 26
rect 80 25 81 26
rect 93 25 99 26
rect 178 24 197 26
rect 179 23 196 24
rect 226 23 230 27
rect 248 27 252 31
rect 262 29 266 37
rect 283 36 288 38
rect 295 37 299 44
rect 315 42 333 45
rect 315 41 319 42
rect 353 41 357 45
rect 315 39 333 41
rect 352 39 357 41
rect 315 38 319 39
rect 352 38 358 39
rect 295 36 302 37
rect 315 36 334 38
rect 351 37 359 38
rect 350 36 360 37
rect 283 34 289 36
rect 295 34 303 36
rect 315 35 333 36
rect 349 35 354 36
rect 355 35 362 36
rect 322 34 326 35
rect 347 34 353 35
rect 357 34 363 35
rect 282 33 290 34
rect 281 32 290 33
rect 295 33 302 34
rect 312 33 336 34
rect 346 33 352 34
rect 358 33 362 34
rect 280 31 285 32
rect 279 30 285 31
rect 287 31 292 32
rect 287 30 293 31
rect 278 29 284 30
rect 288 29 294 30
rect 277 28 283 29
rect 290 28 293 29
rect 278 27 282 28
rect 291 27 292 28
rect 248 26 266 27
rect 248 24 267 26
rect 295 24 299 33
rect 311 32 337 33
rect 347 32 350 33
rect 360 32 362 33
rect 312 31 336 32
rect 321 30 327 31
rect 316 29 331 30
rect 315 28 333 29
rect 314 27 320 28
rect 327 27 334 28
rect 314 26 319 27
rect 330 26 334 27
rect 314 25 320 26
rect 328 25 334 26
rect 351 27 354 31
rect 365 29 369 45
rect 387 44 390 45
rect 399 44 403 45
rect 454 44 463 45
rect 384 43 393 44
rect 399 43 404 44
rect 418 43 437 44
rect 453 43 465 44
rect 383 42 404 43
rect 417 42 437 43
rect 382 41 388 42
rect 389 41 404 42
rect 418 41 437 42
rect 382 40 386 41
rect 391 40 404 41
rect 382 38 385 40
rect 392 39 404 40
rect 392 38 396 39
rect 399 38 404 39
rect 382 37 386 38
rect 391 37 404 38
rect 382 36 387 37
rect 390 36 404 37
rect 383 35 404 36
rect 432 39 437 41
rect 452 42 457 43
rect 461 42 466 43
rect 452 41 456 42
rect 462 41 466 42
rect 452 40 457 41
rect 461 40 466 41
rect 452 39 465 40
rect 432 36 436 39
rect 453 38 464 39
rect 455 37 462 38
rect 451 36 468 37
rect 432 35 435 36
rect 384 34 394 35
rect 385 33 392 34
rect 385 27 389 31
rect 399 30 404 35
rect 415 32 440 35
rect 450 34 468 36
rect 469 34 473 45
rect 450 33 466 34
rect 468 33 473 34
rect 399 29 403 30
rect 351 26 369 27
rect 315 24 333 25
rect 351 24 370 26
rect 385 24 404 27
rect 249 23 266 24
rect 296 23 299 24
rect 317 23 332 24
rect 352 23 369 24
rect 385 23 403 24
rect 425 23 429 32
rect 456 30 459 33
rect 463 30 473 33
rect 456 29 458 30
rect 454 27 458 29
rect 469 29 473 30
rect 469 28 472 29
rect 454 24 473 27
rect 454 23 472 24
rect 321 22 328 23
rect 102 18 105 19
rect 123 18 124 19
rect 36 17 39 18
rect 36 12 38 17
rect 42 16 44 18
rect 48 16 51 18
rect 36 11 39 12
rect 42 11 43 16
rect 37 10 40 11
rect 41 10 43 11
rect 48 15 52 16
rect 54 15 56 18
rect 60 17 63 18
rect 67 17 71 18
rect 48 11 49 15
rect 50 14 53 15
rect 55 14 56 15
rect 51 13 56 14
rect 52 12 56 13
rect 53 11 56 12
rect 61 11 63 17
rect 68 16 70 17
rect 73 16 75 18
rect 79 17 82 18
rect 83 17 85 18
rect 89 17 96 18
rect 101 17 106 18
rect 109 17 113 18
rect 116 17 118 18
rect 119 17 124 18
rect 128 17 131 18
rect 68 15 71 16
rect 69 13 71 15
rect 73 14 74 16
rect 72 13 74 14
rect 80 15 82 17
rect 84 16 86 17
rect 80 13 85 15
rect 90 14 92 17
rect 94 15 96 17
rect 100 16 102 17
rect 105 16 106 17
rect 100 15 103 16
rect 93 14 96 15
rect 101 14 105 15
rect 90 13 95 14
rect 102 13 106 14
rect 38 9 42 10
rect 48 9 50 11
rect 54 9 56 11
rect 60 10 63 11
rect 70 11 73 13
rect 80 11 82 13
rect 85 11 86 12
rect 70 10 72 11
rect 60 9 61 10
rect 71 9 72 10
rect 79 10 82 11
rect 84 10 86 11
rect 90 10 92 13
rect 93 12 95 13
rect 103 12 106 13
rect 93 11 96 12
rect 100 11 101 12
rect 104 11 106 12
rect 110 11 112 17
rect 116 16 117 17
rect 119 16 121 17
rect 123 16 124 17
rect 119 12 122 16
rect 129 15 131 17
rect 133 17 135 18
rect 175 17 181 18
rect 133 16 134 17
rect 132 15 134 16
rect 175 15 178 17
rect 119 11 121 12
rect 94 10 97 11
rect 100 10 102 11
rect 104 10 105 11
rect 110 10 113 11
rect 119 10 122 11
rect 130 10 133 15
rect 175 13 181 15
rect 175 11 178 13
rect 175 10 181 11
rect 182 10 184 19
rect 198 17 200 18
rect 220 17 222 19
rect 197 16 200 17
rect 254 16 257 19
rect 260 17 267 18
rect 262 16 265 17
rect 186 15 190 16
rect 185 14 190 15
rect 192 15 206 16
rect 207 15 211 16
rect 192 14 196 15
rect 185 13 187 14
rect 188 13 193 14
rect 185 12 193 13
rect 185 11 187 12
rect 191 11 194 12
rect 197 11 200 15
rect 201 14 212 15
rect 201 11 204 14
rect 205 11 208 14
rect 210 11 212 14
rect 185 10 191 11
rect 192 10 196 11
rect 198 10 204 11
rect 206 10 212 11
rect 213 14 219 16
rect 213 10 215 14
rect 217 10 219 14
rect 220 10 222 16
rect 224 15 228 16
rect 229 15 233 16
rect 223 14 227 15
rect 228 14 233 15
rect 237 15 242 16
rect 244 15 249 16
rect 237 14 243 15
rect 223 12 225 14
rect 228 13 231 14
rect 238 13 243 14
rect 229 12 233 13
rect 223 11 226 12
rect 231 11 233 12
rect 224 10 233 11
rect 237 12 243 13
rect 237 11 239 12
rect 240 11 243 12
rect 237 10 243 11
rect 244 14 250 15
rect 251 14 257 16
rect 244 10 246 14
rect 247 11 253 14
rect 254 11 257 14
rect 247 10 250 11
rect 251 10 257 11
rect 263 10 265 16
rect 267 15 271 16
rect 266 14 272 15
rect 266 13 269 14
rect 270 13 272 14
rect 266 12 272 13
rect 266 11 269 12
rect 267 10 272 11
rect 273 10 275 19
rect 330 18 332 19
rect 330 17 333 18
rect 346 16 348 18
rect 350 17 352 19
rect 376 17 382 18
rect 277 15 281 16
rect 276 14 282 15
rect 283 14 287 16
rect 289 15 293 16
rect 295 15 304 16
rect 306 15 314 16
rect 288 14 294 15
rect 276 13 279 14
rect 280 13 285 14
rect 287 13 290 14
rect 276 12 285 13
rect 288 12 290 13
rect 276 11 278 12
rect 282 11 285 12
rect 287 11 290 12
rect 292 13 294 14
rect 295 14 315 15
rect 295 13 297 14
rect 292 12 297 13
rect 292 11 294 12
rect 276 10 282 11
rect 283 10 294 11
rect 295 10 297 12
rect 79 9 80 10
rect 81 9 83 10
rect 84 9 85 10
rect 90 9 93 10
rect 95 9 97 10
rect 101 9 104 10
rect 110 9 112 10
rect 119 9 120 10
rect 130 9 131 10
rect 176 9 177 10
rect 180 9 181 10
rect 187 9 189 10
rect 194 9 196 10
rect 202 9 203 10
rect 208 9 210 10
rect 214 9 215 10
rect 218 9 219 10
rect 226 9 227 10
rect 229 9 232 10
rect 239 9 240 10
rect 241 9 242 10
rect 244 9 245 10
rect 248 9 249 10
rect 253 9 256 10
rect 263 9 264 10
rect 268 9 271 10
rect 278 9 280 10
rect 285 9 287 10
rect 290 9 292 10
rect 296 9 297 10
rect 299 10 301 14
rect 302 11 305 14
rect 306 11 308 14
rect 302 10 308 11
rect 309 10 311 14
rect 313 10 315 14
rect 316 11 318 16
rect 320 11 322 16
rect 316 10 322 11
rect 323 14 329 16
rect 323 13 326 14
rect 323 11 325 13
rect 323 10 326 11
rect 327 10 329 14
rect 330 13 332 16
rect 334 15 338 16
rect 333 14 338 15
rect 339 14 344 16
rect 345 15 352 16
rect 354 15 359 16
rect 345 14 349 15
rect 333 13 335 14
rect 340 13 344 14
rect 330 12 335 13
rect 339 12 344 13
rect 330 11 332 12
rect 333 11 336 12
rect 338 11 341 12
rect 342 11 344 12
rect 346 11 348 14
rect 350 11 352 15
rect 330 10 333 11
rect 334 10 338 11
rect 339 10 345 11
rect 346 10 352 11
rect 353 14 359 15
rect 353 11 355 14
rect 357 13 359 14
rect 360 14 366 16
rect 368 15 372 16
rect 376 15 378 17
rect 379 16 382 17
rect 418 16 420 19
rect 380 15 382 16
rect 384 15 388 16
rect 390 15 394 16
rect 360 13 363 14
rect 357 12 360 13
rect 361 12 362 13
rect 357 11 359 12
rect 353 10 359 11
rect 360 11 362 12
rect 360 10 363 11
rect 364 10 366 14
rect 367 14 371 15
rect 376 14 382 15
rect 383 14 389 15
rect 390 14 393 15
rect 395 14 400 16
rect 402 14 407 16
rect 367 13 370 14
rect 376 13 381 14
rect 383 13 385 14
rect 387 13 392 14
rect 394 13 397 14
rect 398 13 401 14
rect 403 13 407 14
rect 368 12 372 13
rect 369 11 372 12
rect 367 10 372 11
rect 376 10 378 13
rect 379 12 389 13
rect 390 12 407 13
rect 380 11 382 12
rect 383 11 385 12
rect 392 11 397 12
rect 401 11 403 12
rect 405 11 407 12
rect 380 10 394 11
rect 395 10 400 11
rect 401 10 407 11
rect 408 15 412 16
rect 413 15 417 16
rect 408 14 416 15
rect 418 14 423 16
rect 408 10 410 14
rect 412 12 414 14
rect 412 11 415 12
rect 412 10 417 11
rect 418 10 420 14
rect 422 13 423 14
rect 421 10 423 13
rect 427 10 430 18
rect 445 17 446 18
rect 448 17 450 19
rect 444 16 446 17
rect 452 16 454 18
rect 464 17 466 18
rect 463 16 466 17
rect 431 15 437 16
rect 439 15 442 16
rect 431 14 442 15
rect 443 14 447 16
rect 431 10 433 14
rect 435 10 437 14
rect 438 13 441 14
rect 439 12 443 13
rect 440 11 443 12
rect 438 10 443 11
rect 444 11 446 14
rect 448 11 450 16
rect 451 14 455 16
rect 444 10 450 11
rect 452 11 454 14
rect 456 11 458 16
rect 460 11 462 16
rect 463 14 467 16
rect 468 14 473 16
rect 463 11 466 14
rect 467 13 470 14
rect 471 13 473 14
rect 467 12 474 13
rect 467 11 470 12
rect 452 10 462 11
rect 464 10 467 11
rect 468 10 473 11
rect 299 9 300 10
rect 303 9 304 10
rect 306 9 307 10
rect 310 9 311 10
rect 317 9 318 10
rect 320 9 321 10
rect 324 9 325 10
rect 328 9 329 10
rect 331 9 332 10
rect 336 9 337 10
rect 340 9 342 10
rect 343 9 344 10
rect 348 9 349 10
rect 356 9 357 10
rect 361 9 362 10
rect 365 9 366 10
rect 368 9 370 10
rect 376 9 377 10
rect 385 9 388 10
rect 390 9 393 10
rect 396 9 399 10
rect 402 9 404 10
rect 405 9 406 10
rect 409 9 410 10
rect 415 9 416 10
rect 418 9 419 10
rect 422 9 423 10
rect 428 9 429 10
rect 432 9 433 10
rect 436 9 437 10
rect 439 9 441 10
rect 445 9 447 10
rect 449 9 450 10
rect 453 9 455 10
rect 457 9 459 10
rect 460 9 461 10
rect 466 9 467 10
rect 470 9 472 10
<< metal2 >>
rect 101 198 102 199
rect 103 198 122 199
rect 95 197 125 198
rect 66 196 71 197
rect 90 196 127 197
rect 65 195 74 196
rect 86 195 129 196
rect 63 194 131 195
rect 63 193 132 194
rect 62 192 133 193
rect 62 191 135 192
rect 61 190 99 191
rect 106 190 136 191
rect 257 190 261 191
rect 267 190 271 191
rect 296 190 301 191
rect 308 190 310 191
rect 321 190 323 191
rect 346 190 349 191
rect 356 190 359 191
rect 364 190 370 191
rect 376 190 378 191
rect 385 190 387 191
rect 393 190 395 191
rect 62 189 70 190
rect 78 189 98 190
rect 109 189 137 190
rect 186 189 191 190
rect 198 189 203 190
rect 209 189 215 190
rect 225 189 228 190
rect 240 189 245 190
rect 257 189 262 190
rect 62 188 68 189
rect 80 188 101 189
rect 114 188 138 189
rect 185 188 192 189
rect 197 188 204 189
rect 52 187 57 188
rect 64 187 65 188
rect 82 187 104 188
rect 119 187 139 188
rect 184 187 193 188
rect 196 187 204 188
rect 208 187 216 189
rect 224 188 228 189
rect 239 188 246 189
rect 223 187 228 188
rect 50 186 59 187
rect 70 186 73 187
rect 83 186 107 187
rect 127 186 140 187
rect 183 186 187 187
rect 49 185 60 186
rect 67 185 75 186
rect 83 185 111 186
rect 131 185 141 186
rect 184 185 187 186
rect 190 185 193 187
rect 49 184 61 185
rect 65 184 77 185
rect 48 183 77 184
rect 83 184 121 185
rect 134 184 142 185
rect 189 184 193 185
rect 195 186 199 187
rect 195 184 198 186
rect 202 184 205 187
rect 207 186 211 187
rect 207 185 210 186
rect 213 185 217 187
rect 222 186 228 187
rect 238 187 247 188
rect 222 185 227 186
rect 238 185 241 187
rect 244 185 247 187
rect 213 184 216 185
rect 221 184 227 185
rect 242 184 247 185
rect 256 184 262 189
rect 266 188 271 190
rect 294 189 302 190
rect 293 188 303 189
rect 307 188 311 190
rect 320 188 324 190
rect 265 186 271 188
rect 292 187 297 188
rect 300 187 304 188
rect 273 186 275 187
rect 281 186 283 187
rect 264 184 270 186
rect 272 185 276 186
rect 280 185 283 186
rect 83 183 125 184
rect 137 183 142 184
rect 188 183 192 184
rect 194 183 198 184
rect 47 181 78 183
rect 83 182 128 183
rect 139 182 142 183
rect 187 182 191 183
rect 46 180 78 181
rect 82 181 131 182
rect 141 181 143 182
rect 186 181 190 182
rect 82 180 134 181
rect 185 180 189 181
rect 45 179 77 180
rect 82 179 137 180
rect 184 179 188 180
rect 44 178 77 179
rect 83 178 139 179
rect 183 178 187 179
rect 194 178 197 183
rect 201 182 205 184
rect 212 183 216 184
rect 220 183 223 184
rect 211 182 215 183
rect 219 182 222 183
rect 224 182 227 184
rect 241 183 246 184
rect 241 182 245 183
rect 201 180 204 182
rect 210 181 214 182
rect 218 181 221 182
rect 223 181 226 182
rect 209 180 213 181
rect 200 179 204 180
rect 208 179 212 180
rect 217 179 228 181
rect 229 179 235 182
rect 242 181 246 182
rect 236 179 239 180
rect 243 179 247 181
rect 255 179 258 184
rect 200 178 203 179
rect 207 178 211 179
rect 217 178 227 179
rect 236 178 240 179
rect 243 178 246 179
rect 43 177 76 178
rect 84 177 142 178
rect 183 177 192 178
rect 194 177 203 178
rect 41 176 75 177
rect 86 176 106 177
rect 110 176 144 177
rect 182 176 192 177
rect 195 176 202 177
rect 40 175 56 176
rect 58 175 73 176
rect 87 175 107 176
rect 112 175 145 176
rect 182 175 191 176
rect 196 175 200 176
rect 206 175 215 178
rect 223 177 226 178
rect 237 177 246 178
rect 254 178 258 179
rect 259 182 262 184
rect 263 182 266 184
rect 259 179 265 182
rect 267 181 270 184
rect 222 175 225 177
rect 237 176 245 177
rect 239 175 243 176
rect 254 175 257 178
rect 259 177 264 179
rect 259 175 263 177
rect 266 176 269 181
rect 273 180 276 185
rect 279 184 283 185
rect 291 185 295 187
rect 301 186 304 187
rect 307 186 310 188
rect 312 186 315 187
rect 321 186 322 187
rect 326 186 328 187
rect 330 186 333 187
rect 345 186 350 190
rect 355 189 360 190
rect 363 189 373 190
rect 354 187 359 189
rect 363 188 374 189
rect 363 187 366 188
rect 370 187 374 188
rect 301 185 303 186
rect 307 185 316 186
rect 320 185 323 186
rect 291 184 294 185
rect 279 183 282 184
rect 278 182 282 183
rect 278 181 281 182
rect 277 180 281 181
rect 273 179 280 180
rect 290 179 294 184
rect 306 184 316 185
rect 306 183 310 184
rect 313 183 317 184
rect 319 183 323 185
rect 325 185 335 186
rect 325 184 330 185
rect 331 184 335 185
rect 344 184 350 186
rect 353 185 359 187
rect 325 183 329 184
rect 306 180 309 183
rect 313 180 316 183
rect 319 180 322 183
rect 325 181 328 183
rect 300 179 303 180
rect 274 178 280 179
rect 291 178 295 179
rect 299 178 303 179
rect 305 179 309 180
rect 274 176 279 178
rect 291 177 302 178
rect 292 176 301 177
rect 265 175 268 176
rect 274 175 278 176
rect 293 175 300 176
rect 305 175 308 179
rect 312 178 316 180
rect 318 179 322 180
rect 312 175 315 178
rect 318 175 321 179
rect 324 178 328 181
rect 332 180 336 184
rect 344 181 347 184
rect 348 181 350 184
rect 352 184 359 185
rect 352 183 355 184
rect 356 183 359 184
rect 362 185 366 187
rect 371 185 374 187
rect 362 184 365 185
rect 370 184 374 185
rect 351 181 354 183
rect 332 179 335 180
rect 331 178 335 179
rect 324 177 329 178
rect 330 177 334 178
rect 343 177 346 181
rect 323 176 333 177
rect 342 176 346 177
rect 348 180 354 181
rect 348 178 353 180
rect 355 178 358 183
rect 362 182 373 184
rect 361 181 371 182
rect 376 181 379 190
rect 384 189 388 190
rect 383 187 388 189
rect 392 189 396 190
rect 392 188 395 189
rect 382 185 388 187
rect 391 187 395 188
rect 391 185 394 187
rect 381 183 384 185
rect 380 182 384 183
rect 380 181 383 182
rect 361 180 365 181
rect 376 180 383 181
rect 385 181 388 185
rect 390 183 393 185
rect 389 181 392 183
rect 361 178 364 180
rect 348 176 352 178
rect 323 175 327 176
rect 328 175 332 176
rect 342 175 345 176
rect 348 175 351 176
rect 354 175 357 178
rect 360 176 364 178
rect 376 178 382 180
rect 385 179 391 181
rect 376 176 381 178
rect 385 177 390 179
rect 360 175 363 176
rect 376 175 380 176
rect 385 175 389 177
rect 38 174 52 175
rect 57 174 72 175
rect 89 174 107 175
rect 114 174 146 175
rect 274 174 277 175
rect 37 173 49 174
rect 55 173 71 174
rect 90 173 107 174
rect 117 173 147 174
rect 273 173 277 174
rect 35 172 47 173
rect 53 172 71 173
rect 91 172 108 173
rect 120 172 148 173
rect 33 171 45 172
rect 52 171 70 172
rect 77 171 84 172
rect 92 171 109 172
rect 124 171 148 172
rect 271 172 276 173
rect 271 171 275 172
rect 323 171 326 175
rect 31 170 44 171
rect 51 170 71 171
rect 29 169 47 170
rect 27 168 48 169
rect 50 168 71 170
rect 77 170 86 171
rect 93 170 111 171
rect 127 170 149 171
rect 77 169 87 170
rect 94 169 112 170
rect 130 169 149 170
rect 26 167 48 168
rect 49 167 71 168
rect 78 167 88 169
rect 94 168 114 169
rect 132 168 149 169
rect 95 167 118 168
rect 134 167 150 168
rect 25 165 72 167
rect 78 166 89 167
rect 96 166 122 167
rect 135 166 150 167
rect 79 165 90 166
rect 96 165 126 166
rect 137 165 150 166
rect 24 163 72 165
rect 25 162 31 163
rect 32 162 72 163
rect 25 161 29 162
rect 31 161 72 162
rect 30 160 72 161
rect 29 159 72 160
rect 78 164 90 165
rect 97 164 128 165
rect 138 164 150 165
rect 78 161 91 164
rect 97 163 130 164
rect 139 163 150 164
rect 98 162 131 163
rect 141 162 151 163
rect 98 161 133 162
rect 142 161 151 162
rect 78 159 92 161
rect 99 160 134 161
rect 143 160 151 161
rect 100 159 135 160
rect 144 159 151 160
rect 28 158 71 159
rect 27 156 71 158
rect 78 158 93 159
rect 101 158 136 159
rect 78 157 94 158
rect 102 157 138 158
rect 145 157 151 159
rect 77 156 94 157
rect 104 156 139 157
rect 146 156 150 157
rect 28 155 70 156
rect 77 155 95 156
rect 107 155 140 156
rect 28 154 69 155
rect 77 154 97 155
rect 113 154 141 155
rect 147 154 150 156
rect 29 153 69 154
rect 76 153 98 154
rect 117 153 142 154
rect 148 153 150 154
rect 187 153 195 154
rect 29 152 46 153
rect 48 152 68 153
rect 76 152 101 153
rect 120 152 142 153
rect 30 151 45 152
rect 31 150 43 151
rect 49 150 67 152
rect 76 151 105 152
rect 122 151 143 152
rect 185 151 195 153
rect 75 150 110 151
rect 125 150 143 151
rect 33 149 38 150
rect 48 149 66 150
rect 75 149 113 150
rect 127 149 143 150
rect 184 150 194 151
rect 44 148 65 149
rect 74 148 116 149
rect 128 148 144 149
rect 38 147 65 148
rect 73 147 118 148
rect 129 147 144 148
rect 33 146 64 147
rect 73 146 120 147
rect 130 146 144 147
rect 184 146 190 150
rect 196 149 202 154
rect 303 152 307 154
rect 302 151 306 152
rect 301 149 306 151
rect 311 149 330 154
rect 300 147 305 149
rect 215 146 217 147
rect 253 146 256 147
rect 272 146 276 147
rect 33 145 63 146
rect 72 145 122 146
rect 131 145 144 146
rect 33 144 62 145
rect 71 144 123 145
rect 33 143 61 144
rect 70 143 124 144
rect 132 143 144 145
rect 34 142 60 143
rect 70 142 125 143
rect 133 142 144 143
rect 181 142 194 146
rect 34 141 59 142
rect 69 141 125 142
rect 35 140 57 141
rect 67 140 92 141
rect 99 140 126 141
rect 134 140 144 142
rect 35 139 55 140
rect 66 139 91 140
rect 101 139 126 140
rect 135 139 144 140
rect 36 138 53 139
rect 65 138 90 139
rect 102 138 127 139
rect 135 138 143 139
rect 36 137 50 138
rect 64 137 90 138
rect 103 137 127 138
rect 37 136 47 137
rect 62 136 90 137
rect 104 136 128 137
rect 37 135 44 136
rect 60 135 89 136
rect 105 135 128 136
rect 136 135 143 138
rect 38 134 41 135
rect 58 134 89 135
rect 96 134 97 135
rect 56 133 89 134
rect 95 133 98 134
rect 106 133 128 135
rect 53 132 88 133
rect 95 132 99 133
rect 51 131 88 132
rect 94 131 99 132
rect 107 132 128 133
rect 137 134 143 135
rect 137 132 142 134
rect 107 131 127 132
rect 49 130 87 131
rect 94 130 100 131
rect 47 129 87 130
rect 93 129 100 130
rect 108 129 127 131
rect 138 130 141 132
rect 138 129 140 130
rect 45 128 86 129
rect 93 128 101 129
rect 44 127 86 128
rect 92 127 101 128
rect 108 128 126 129
rect 138 128 139 129
rect 108 127 125 128
rect 43 126 85 127
rect 42 125 84 126
rect 92 125 102 127
rect 41 124 83 125
rect 91 124 102 125
rect 109 126 125 127
rect 184 126 190 142
rect 196 126 202 146
rect 207 145 212 146
rect 213 145 220 146
rect 207 144 220 145
rect 243 144 248 146
rect 250 145 258 146
rect 270 145 279 146
rect 249 144 259 145
rect 268 144 280 145
rect 299 144 304 147
rect 207 141 219 144
rect 243 143 260 144
rect 267 143 281 144
rect 298 143 304 144
rect 311 143 317 149
rect 243 142 261 143
rect 266 142 282 143
rect 243 141 250 142
rect 255 141 262 142
rect 266 141 272 142
rect 207 140 214 141
rect 207 138 213 140
rect 243 138 249 141
rect 256 139 262 141
rect 257 138 262 139
rect 265 138 271 141
rect 277 140 283 142
rect 278 138 283 140
rect 298 138 303 143
rect 207 126 212 138
rect 243 135 248 138
rect 257 135 263 138
rect 265 135 284 138
rect 297 135 303 138
rect 243 132 249 135
rect 257 133 262 135
rect 243 131 250 132
rect 256 131 262 133
rect 265 134 283 135
rect 265 131 271 134
rect 278 132 279 133
rect 243 130 251 131
rect 255 130 261 131
rect 243 129 261 130
rect 266 130 273 131
rect 277 130 283 132
rect 298 130 303 135
rect 311 138 328 143
rect 266 129 282 130
rect 298 129 304 130
rect 243 128 260 129
rect 267 128 282 129
rect 109 125 124 126
rect 109 124 123 125
rect 41 123 82 124
rect 91 123 103 124
rect 40 122 81 123
rect 90 122 103 123
rect 109 123 122 124
rect 132 123 133 124
rect 109 122 121 123
rect 131 122 133 123
rect 40 121 80 122
rect 39 120 79 121
rect 89 120 103 122
rect 39 119 78 120
rect 88 119 103 120
rect 110 121 119 122
rect 130 121 134 122
rect 110 120 118 121
rect 129 120 133 121
rect 110 119 116 120
rect 128 119 134 120
rect 218 119 241 122
rect 39 118 77 119
rect 87 118 103 119
rect 38 117 76 118
rect 86 117 103 118
rect 109 118 114 119
rect 127 118 134 119
rect 219 118 240 119
rect 243 118 248 128
rect 249 127 259 128
rect 268 127 281 128
rect 251 126 258 127
rect 270 126 279 127
rect 299 126 304 129
rect 311 126 317 138
rect 334 126 340 154
rect 345 153 362 154
rect 378 153 384 154
rect 393 153 396 154
rect 345 152 364 153
rect 375 152 386 153
rect 393 152 397 153
rect 345 151 366 152
rect 374 151 387 152
rect 393 151 398 152
rect 345 149 367 151
rect 373 149 388 151
rect 394 150 398 151
rect 394 149 399 150
rect 345 143 351 149
rect 359 148 368 149
rect 361 147 368 148
rect 362 144 368 147
rect 372 145 378 149
rect 383 148 389 149
rect 384 145 389 148
rect 395 148 399 149
rect 395 146 400 148
rect 361 143 368 144
rect 373 144 378 145
rect 383 144 389 145
rect 373 143 379 144
rect 382 143 388 144
rect 396 143 401 146
rect 345 141 367 143
rect 374 142 387 143
rect 345 140 366 141
rect 375 140 386 142
rect 396 141 402 143
rect 345 139 364 140
rect 374 139 388 140
rect 345 138 362 139
rect 373 138 379 139
rect 382 138 389 139
rect 345 137 352 138
rect 353 137 362 138
rect 372 137 378 138
rect 383 137 389 138
rect 345 126 351 137
rect 356 136 363 137
rect 357 135 364 136
rect 357 134 365 135
rect 358 133 366 134
rect 359 132 366 133
rect 372 132 377 137
rect 359 131 367 132
rect 360 130 367 131
rect 372 131 378 132
rect 384 131 390 137
rect 397 131 402 141
rect 372 130 379 131
rect 383 130 389 131
rect 361 129 368 130
rect 373 129 389 130
rect 396 130 402 131
rect 362 127 369 129
rect 374 128 388 129
rect 375 127 387 128
rect 363 126 370 127
rect 376 126 385 127
rect 396 126 401 130
rect 300 125 304 126
rect 300 123 305 125
rect 395 124 400 126
rect 395 123 399 124
rect 301 122 306 123
rect 302 120 306 122
rect 394 122 399 123
rect 394 121 398 122
rect 393 120 398 121
rect 303 119 307 120
rect 304 118 307 119
rect 393 119 397 120
rect 393 118 396 119
rect 109 117 112 118
rect 126 117 134 118
rect 38 116 74 117
rect 85 116 103 117
rect 124 116 134 117
rect 38 115 73 116
rect 84 115 103 116
rect 123 115 134 116
rect 38 114 71 115
rect 82 114 103 115
rect 121 114 134 115
rect 38 113 69 114
rect 81 113 103 114
rect 120 113 134 114
rect 38 112 67 113
rect 79 112 103 113
rect 118 112 134 113
rect 38 111 64 112
rect 78 111 103 112
rect 116 111 134 112
rect 38 110 62 111
rect 76 110 102 111
rect 114 110 133 111
rect 38 109 60 110
rect 74 109 102 110
rect 111 109 133 110
rect 38 108 58 109
rect 72 108 102 109
rect 108 108 133 109
rect 38 107 57 108
rect 70 107 102 108
rect 104 107 133 108
rect 39 106 55 107
rect 68 106 133 107
rect 39 104 54 106
rect 67 105 132 106
rect 65 104 132 105
rect 39 103 53 104
rect 64 103 132 104
rect 40 102 53 103
rect 62 102 131 103
rect 40 101 52 102
rect 61 101 131 102
rect 41 100 52 101
rect 60 100 130 101
rect 41 99 51 100
rect 42 97 51 99
rect 59 99 85 100
rect 87 99 130 100
rect 59 98 84 99
rect 87 98 129 99
rect 58 97 82 98
rect 86 97 129 98
rect 43 95 51 97
rect 57 96 80 97
rect 57 95 79 96
rect 85 95 128 97
rect 44 94 51 95
rect 56 94 77 95
rect 84 94 127 95
rect 45 93 50 94
rect 56 93 76 94
rect 83 93 126 94
rect 46 92 50 93
rect 47 91 50 92
rect 48 90 50 91
rect 55 92 75 93
rect 83 92 102 93
rect 103 92 125 93
rect 55 91 74 92
rect 82 91 100 92
rect 102 91 125 92
rect 175 92 251 103
rect 264 92 342 103
rect 353 102 427 103
rect 353 101 430 102
rect 353 100 431 101
rect 353 99 432 100
rect 353 98 433 99
rect 353 97 434 98
rect 353 92 435 97
rect 175 91 198 92
rect 55 90 73 91
rect 81 90 99 91
rect 102 90 124 91
rect 49 89 50 90
rect 54 89 72 90
rect 80 89 98 90
rect 101 89 123 90
rect 54 87 71 89
rect 80 88 97 89
rect 101 88 122 89
rect 79 87 96 88
rect 101 87 121 88
rect 54 85 70 87
rect 79 86 95 87
rect 101 86 120 87
rect 175 86 199 91
rect 78 85 95 86
rect 100 85 119 86
rect 175 85 198 86
rect 54 82 69 85
rect 78 83 94 85
rect 100 84 118 85
rect 175 84 199 85
rect 100 83 117 84
rect 55 80 68 82
rect 56 79 68 80
rect 77 81 93 83
rect 100 82 115 83
rect 100 81 114 82
rect 77 79 92 81
rect 57 77 68 79
rect 58 76 68 77
rect 59 75 68 76
rect 60 74 68 75
rect 62 73 68 74
rect 76 78 92 79
rect 100 80 113 81
rect 100 79 111 80
rect 100 78 110 79
rect 76 73 91 78
rect 100 77 109 78
rect 100 76 108 77
rect 100 75 107 76
rect 100 74 106 75
rect 175 74 251 84
rect 100 73 105 74
rect 63 72 68 73
rect 65 71 69 72
rect 66 70 69 71
rect 67 69 69 70
rect 77 69 91 73
rect 101 72 105 73
rect 175 73 200 74
rect 101 71 104 72
rect 101 69 103 71
rect 68 68 69 69
rect 78 67 91 69
rect 79 66 91 67
rect 80 65 91 66
rect 175 67 199 73
rect 175 66 198 67
rect 175 65 199 66
rect 80 64 92 65
rect 81 63 92 64
rect 82 62 92 63
rect 83 61 92 62
rect 175 61 251 65
rect 84 60 93 61
rect 85 59 93 60
rect 176 59 251 61
rect 86 58 93 59
rect 177 58 251 59
rect 88 57 94 58
rect 178 57 251 58
rect 90 56 94 57
rect 179 56 251 57
rect 92 55 95 56
rect 181 55 251 56
rect 291 55 315 92
rect 353 55 377 92
rect 411 78 435 92
rect 386 77 435 78
rect 385 76 413 77
rect 386 75 414 76
rect 387 74 415 75
rect 388 73 417 74
rect 390 72 418 73
rect 391 71 419 72
rect 392 70 420 71
rect 393 69 421 70
rect 394 68 423 69
rect 396 67 424 68
rect 397 66 425 67
rect 398 65 426 66
rect 399 64 428 65
rect 401 63 429 64
rect 402 62 430 63
rect 403 61 431 62
rect 404 60 433 61
rect 406 59 434 60
rect 407 58 435 59
rect 408 57 436 58
rect 409 56 437 57
rect 410 55 439 56
rect 452 55 476 103
rect 412 54 440 55
rect 413 53 441 54
rect 414 52 443 53
rect 415 51 443 52
rect 458 43 463 44
rect 96 42 101 43
rect 6 41 14 42
rect 16 41 24 42
rect 26 41 34 42
rect 37 41 43 42
rect 45 41 54 42
rect 57 41 65 42
rect 66 41 72 42
rect 79 41 86 42
rect 93 41 104 42
rect 114 41 123 42
rect 125 41 134 42
rect 137 41 150 42
rect 154 41 168 42
rect 180 41 189 43
rect 7 40 13 41
rect 18 40 22 41
rect 27 40 33 41
rect 8 34 12 40
rect 17 39 20 40
rect 28 39 33 40
rect 17 38 19 39
rect 29 38 33 39
rect 38 40 42 41
rect 47 40 53 41
rect 59 40 64 41
rect 68 40 73 41
rect 81 40 85 41
rect 91 40 96 41
rect 100 40 104 41
rect 115 40 121 41
rect 127 40 132 41
rect 38 39 41 40
rect 38 38 40 39
rect 16 37 18 38
rect 29 37 34 38
rect 15 36 17 37
rect 30 36 34 37
rect 37 36 39 38
rect 14 35 16 36
rect 30 35 35 36
rect 13 34 16 35
rect 31 34 35 35
rect 36 34 38 36
rect 8 32 17 34
rect 31 33 37 34
rect 8 26 12 32
rect 13 31 18 32
rect 14 29 19 31
rect 15 28 20 29
rect 16 27 21 28
rect 16 26 22 27
rect 7 25 13 26
rect 17 25 23 26
rect 32 25 37 33
rect 47 31 52 40
rect 48 28 52 31
rect 60 37 63 40
rect 69 39 74 40
rect 69 38 75 39
rect 69 37 76 38
rect 60 30 62 37
rect 69 36 77 37
rect 60 29 63 30
rect 60 28 62 29
rect 48 27 53 28
rect 59 27 62 28
rect 49 26 54 27
rect 58 26 62 27
rect 69 26 71 36
rect 72 35 77 36
rect 73 34 78 35
rect 74 33 79 34
rect 75 32 80 33
rect 76 31 81 32
rect 82 31 84 40
rect 90 39 94 40
rect 101 39 104 40
rect 89 38 93 39
rect 102 38 104 39
rect 88 37 93 38
rect 103 37 104 38
rect 116 39 121 40
rect 88 35 92 37
rect 87 31 92 35
rect 116 35 120 39
rect 128 35 132 40
rect 116 33 132 35
rect 97 32 106 33
rect 98 31 106 32
rect 116 32 121 33
rect 127 32 132 33
rect 76 30 84 31
rect 77 29 84 30
rect 78 28 84 29
rect 88 30 92 31
rect 88 28 93 30
rect 79 27 84 28
rect 89 27 94 28
rect 49 25 61 26
rect 68 25 72 26
rect 80 25 84 27
rect 90 26 94 27
rect 91 25 96 26
rect 100 25 104 31
rect 116 26 120 32
rect 128 26 132 32
rect 139 40 144 41
rect 147 40 151 41
rect 139 35 143 40
rect 149 38 151 40
rect 149 37 150 38
rect 148 35 149 36
rect 139 34 144 35
rect 147 34 149 35
rect 139 32 149 34
rect 139 26 143 32
rect 147 31 149 32
rect 148 30 149 31
rect 156 34 161 41
rect 164 40 168 41
rect 166 38 168 40
rect 177 38 193 40
rect 177 37 192 38
rect 195 37 198 43
rect 214 42 232 43
rect 213 40 233 42
rect 214 39 232 40
rect 247 39 261 42
rect 264 39 268 43
rect 298 42 301 43
rect 281 39 295 41
rect 182 36 188 37
rect 165 35 167 36
rect 179 35 190 36
rect 164 34 167 35
rect 156 32 167 34
rect 178 34 191 35
rect 195 34 201 37
rect 228 35 232 39
rect 252 37 256 39
rect 251 36 257 37
rect 250 35 257 36
rect 260 35 268 39
rect 280 38 295 39
rect 286 36 290 38
rect 211 34 235 35
rect 249 34 259 35
rect 178 33 183 34
rect 186 33 192 34
rect 177 32 182 33
rect 188 32 192 33
rect 150 27 152 29
rect 149 26 152 27
rect 156 26 161 32
rect 165 31 167 32
rect 178 31 183 32
rect 186 31 192 32
rect 165 30 166 31
rect 178 30 191 31
rect 180 29 190 30
rect 168 28 169 29
rect 167 27 169 28
rect 181 27 184 28
rect 195 27 198 34
rect 210 33 236 34
rect 248 33 260 34
rect 211 32 236 33
rect 246 32 253 33
rect 255 32 262 33
rect 211 31 235 32
rect 246 31 252 32
rect 257 31 261 32
rect 221 29 224 31
rect 247 30 250 31
rect 259 30 260 31
rect 214 28 232 29
rect 166 26 169 27
rect 116 25 121 26
rect 127 25 133 26
rect 139 25 144 26
rect 148 25 151 26
rect 156 25 162 26
rect 165 25 169 26
rect 180 25 185 27
rect 213 26 232 28
rect 214 25 232 26
rect 6 24 14 25
rect 18 24 24 25
rect 30 24 39 25
rect 50 24 60 25
rect 67 24 74 25
rect 81 24 84 25
rect 92 24 104 25
rect 114 24 123 25
rect 125 24 134 25
rect 137 24 151 25
rect 154 24 168 25
rect 180 24 198 25
rect 53 23 58 24
rect 82 23 83 24
rect 95 23 101 24
rect 180 22 199 24
rect 181 21 198 22
rect 228 21 232 25
rect 250 25 254 29
rect 264 27 268 35
rect 285 34 290 36
rect 297 35 301 42
rect 317 40 335 43
rect 317 39 321 40
rect 355 39 359 43
rect 317 37 335 39
rect 354 37 359 39
rect 317 36 321 37
rect 354 36 360 37
rect 297 34 304 35
rect 317 34 336 36
rect 353 35 361 36
rect 352 34 362 35
rect 285 32 291 34
rect 297 32 305 34
rect 317 33 335 34
rect 351 33 356 34
rect 357 33 364 34
rect 324 32 328 33
rect 349 32 355 33
rect 359 32 365 33
rect 284 31 292 32
rect 283 30 292 31
rect 297 31 304 32
rect 314 31 338 32
rect 348 31 354 32
rect 360 31 364 32
rect 282 29 287 30
rect 281 28 287 29
rect 289 29 294 30
rect 289 28 295 29
rect 280 27 286 28
rect 290 27 296 28
rect 279 26 285 27
rect 292 26 295 27
rect 280 25 284 26
rect 293 25 294 26
rect 250 24 268 25
rect 250 22 269 24
rect 297 22 301 31
rect 313 30 339 31
rect 349 30 352 31
rect 362 30 364 31
rect 314 29 338 30
rect 323 28 329 29
rect 318 27 333 28
rect 317 26 335 27
rect 316 25 322 26
rect 329 25 336 26
rect 316 24 321 25
rect 332 24 336 25
rect 316 23 322 24
rect 330 23 336 24
rect 353 25 356 29
rect 367 27 371 43
rect 389 42 392 43
rect 401 42 405 43
rect 456 42 465 43
rect 386 41 395 42
rect 401 41 406 42
rect 420 41 439 42
rect 455 41 467 42
rect 385 40 406 41
rect 419 40 439 41
rect 384 39 390 40
rect 391 39 406 40
rect 420 39 439 40
rect 384 38 388 39
rect 393 38 406 39
rect 384 36 387 38
rect 394 37 406 38
rect 394 36 398 37
rect 401 36 406 37
rect 384 35 388 36
rect 393 35 406 36
rect 384 34 389 35
rect 392 34 406 35
rect 385 33 406 34
rect 434 37 439 39
rect 454 40 459 41
rect 463 40 468 41
rect 454 39 458 40
rect 464 39 468 40
rect 454 38 459 39
rect 463 38 468 39
rect 454 37 467 38
rect 434 34 438 37
rect 455 36 466 37
rect 457 35 464 36
rect 453 34 470 35
rect 434 33 437 34
rect 386 32 396 33
rect 387 31 394 32
rect 387 25 391 29
rect 401 28 406 33
rect 417 30 442 33
rect 452 32 470 34
rect 471 32 475 43
rect 452 31 468 32
rect 470 31 475 32
rect 401 27 405 28
rect 353 24 371 25
rect 317 22 335 23
rect 353 22 372 24
rect 387 22 406 25
rect 251 21 268 22
rect 298 21 301 22
rect 319 21 334 22
rect 354 21 371 22
rect 387 21 405 22
rect 427 21 431 30
rect 458 28 461 31
rect 465 28 475 31
rect 458 27 460 28
rect 456 25 460 27
rect 471 27 475 28
rect 471 26 474 27
rect 456 22 475 25
rect 456 21 474 22
rect 323 20 330 21
rect 104 16 107 17
rect 125 16 126 17
rect 38 15 41 16
rect 38 10 40 15
rect 44 14 46 16
rect 50 14 53 16
rect 38 9 41 10
rect 44 9 45 14
rect 39 8 42 9
rect 43 8 45 9
rect 50 13 54 14
rect 56 13 58 16
rect 62 15 65 16
rect 69 15 73 16
rect 50 9 51 13
rect 52 12 55 13
rect 57 12 58 13
rect 53 11 58 12
rect 54 10 58 11
rect 55 9 58 10
rect 63 9 65 15
rect 70 14 72 15
rect 75 14 77 16
rect 81 15 84 16
rect 85 15 87 16
rect 91 15 98 16
rect 103 15 108 16
rect 111 15 115 16
rect 118 15 120 16
rect 121 15 126 16
rect 130 15 133 16
rect 70 13 73 14
rect 71 11 73 13
rect 75 12 76 14
rect 74 11 76 12
rect 82 13 84 15
rect 86 14 88 15
rect 82 11 87 13
rect 92 12 94 15
rect 96 13 98 15
rect 102 14 104 15
rect 107 14 108 15
rect 102 13 105 14
rect 95 12 98 13
rect 103 12 107 13
rect 92 11 97 12
rect 104 11 108 12
rect 40 7 44 8
rect 50 7 52 9
rect 56 7 58 9
rect 62 8 65 9
rect 72 9 75 11
rect 82 9 84 11
rect 87 9 88 10
rect 72 8 74 9
rect 62 7 63 8
rect 73 7 74 8
rect 81 8 84 9
rect 86 8 88 9
rect 92 8 94 11
rect 95 10 97 11
rect 105 10 108 11
rect 95 9 98 10
rect 102 9 103 10
rect 106 9 108 10
rect 112 9 114 15
rect 118 14 119 15
rect 121 14 123 15
rect 125 14 126 15
rect 121 10 124 14
rect 131 13 133 15
rect 135 15 137 16
rect 177 15 183 16
rect 135 14 136 15
rect 134 13 136 14
rect 177 13 180 15
rect 121 9 123 10
rect 96 8 99 9
rect 102 8 104 9
rect 106 8 107 9
rect 112 8 115 9
rect 121 8 124 9
rect 132 8 135 13
rect 177 11 183 13
rect 177 9 180 11
rect 177 8 183 9
rect 184 8 186 17
rect 200 15 202 16
rect 222 15 224 17
rect 199 14 202 15
rect 256 14 259 17
rect 262 15 269 16
rect 264 14 267 15
rect 188 13 192 14
rect 187 12 192 13
rect 194 13 208 14
rect 209 13 213 14
rect 194 12 198 13
rect 187 11 189 12
rect 190 11 195 12
rect 187 10 195 11
rect 187 9 189 10
rect 193 9 196 10
rect 199 9 202 13
rect 203 12 214 13
rect 203 9 206 12
rect 207 9 210 12
rect 212 9 214 12
rect 187 8 193 9
rect 194 8 198 9
rect 200 8 206 9
rect 208 8 214 9
rect 215 12 221 14
rect 215 8 217 12
rect 219 8 221 12
rect 222 8 224 14
rect 226 13 230 14
rect 231 13 235 14
rect 225 12 229 13
rect 230 12 235 13
rect 239 13 244 14
rect 246 13 251 14
rect 239 12 245 13
rect 225 10 227 12
rect 230 11 233 12
rect 240 11 245 12
rect 231 10 235 11
rect 225 9 228 10
rect 233 9 235 10
rect 226 8 235 9
rect 239 10 245 11
rect 239 9 241 10
rect 242 9 245 10
rect 239 8 245 9
rect 246 12 252 13
rect 253 12 259 14
rect 246 8 248 12
rect 249 9 255 12
rect 256 9 259 12
rect 249 8 252 9
rect 253 8 259 9
rect 265 8 267 14
rect 269 13 273 14
rect 268 12 274 13
rect 268 11 271 12
rect 272 11 274 12
rect 268 10 274 11
rect 268 9 271 10
rect 269 8 274 9
rect 275 8 277 17
rect 332 16 334 17
rect 332 15 335 16
rect 348 14 350 16
rect 352 15 354 17
rect 378 15 384 16
rect 279 13 283 14
rect 278 12 284 13
rect 285 12 289 14
rect 291 13 295 14
rect 297 13 306 14
rect 308 13 316 14
rect 290 12 296 13
rect 278 11 281 12
rect 282 11 287 12
rect 289 11 292 12
rect 278 10 287 11
rect 290 10 292 11
rect 278 9 280 10
rect 284 9 287 10
rect 289 9 292 10
rect 294 11 296 12
rect 297 12 317 13
rect 297 11 299 12
rect 294 10 299 11
rect 294 9 296 10
rect 278 8 284 9
rect 285 8 296 9
rect 297 8 299 10
rect 81 7 82 8
rect 83 7 85 8
rect 86 7 87 8
rect 92 7 95 8
rect 97 7 99 8
rect 103 7 106 8
rect 112 7 114 8
rect 121 7 122 8
rect 132 7 133 8
rect 178 7 179 8
rect 182 7 183 8
rect 189 7 191 8
rect 196 7 198 8
rect 204 7 205 8
rect 210 7 212 8
rect 216 7 217 8
rect 220 7 221 8
rect 228 7 229 8
rect 231 7 234 8
rect 241 7 242 8
rect 243 7 244 8
rect 246 7 247 8
rect 250 7 251 8
rect 255 7 258 8
rect 265 7 266 8
rect 270 7 273 8
rect 280 7 282 8
rect 287 7 289 8
rect 292 7 294 8
rect 298 7 299 8
rect 301 8 303 12
rect 304 9 307 12
rect 308 9 310 12
rect 304 8 310 9
rect 311 8 313 12
rect 315 8 317 12
rect 318 9 320 14
rect 322 9 324 14
rect 318 8 324 9
rect 325 12 331 14
rect 325 11 328 12
rect 325 9 327 11
rect 325 8 328 9
rect 329 8 331 12
rect 332 11 334 14
rect 336 13 340 14
rect 335 12 340 13
rect 341 12 346 14
rect 347 13 354 14
rect 356 13 361 14
rect 347 12 351 13
rect 335 11 337 12
rect 342 11 346 12
rect 332 10 337 11
rect 341 10 346 11
rect 332 9 334 10
rect 335 9 338 10
rect 340 9 343 10
rect 344 9 346 10
rect 348 9 350 12
rect 352 9 354 13
rect 332 8 335 9
rect 336 8 340 9
rect 341 8 347 9
rect 348 8 354 9
rect 355 12 361 13
rect 355 9 357 12
rect 359 11 361 12
rect 362 12 368 14
rect 370 13 374 14
rect 378 13 380 15
rect 381 14 384 15
rect 420 14 422 17
rect 382 13 384 14
rect 386 13 390 14
rect 392 13 396 14
rect 362 11 365 12
rect 359 10 362 11
rect 363 10 364 11
rect 359 9 361 10
rect 355 8 361 9
rect 362 9 364 10
rect 362 8 365 9
rect 366 8 368 12
rect 369 12 373 13
rect 378 12 384 13
rect 385 12 391 13
rect 392 12 395 13
rect 397 12 402 14
rect 404 12 409 14
rect 369 11 372 12
rect 378 11 383 12
rect 385 11 387 12
rect 389 11 394 12
rect 396 11 399 12
rect 400 11 403 12
rect 405 11 409 12
rect 370 10 374 11
rect 371 9 374 10
rect 369 8 374 9
rect 378 8 380 11
rect 381 10 391 11
rect 392 10 409 11
rect 382 9 384 10
rect 385 9 387 10
rect 394 9 399 10
rect 403 9 405 10
rect 407 9 409 10
rect 382 8 396 9
rect 397 8 402 9
rect 403 8 409 9
rect 410 13 414 14
rect 415 13 419 14
rect 410 12 418 13
rect 420 12 425 14
rect 410 8 412 12
rect 414 10 416 12
rect 414 9 417 10
rect 414 8 419 9
rect 420 8 422 12
rect 424 11 425 12
rect 423 8 425 11
rect 429 8 432 16
rect 447 15 448 16
rect 450 15 452 17
rect 446 14 448 15
rect 454 14 456 16
rect 466 15 468 16
rect 465 14 468 15
rect 433 13 439 14
rect 441 13 444 14
rect 433 12 444 13
rect 445 12 449 14
rect 433 8 435 12
rect 437 8 439 12
rect 440 11 443 12
rect 441 10 445 11
rect 442 9 445 10
rect 440 8 445 9
rect 446 9 448 12
rect 450 9 452 14
rect 453 12 457 14
rect 446 8 452 9
rect 454 9 456 12
rect 458 9 460 14
rect 462 9 464 14
rect 465 12 469 14
rect 470 12 475 14
rect 465 9 468 12
rect 469 11 472 12
rect 473 11 475 12
rect 469 10 476 11
rect 469 9 472 10
rect 454 8 464 9
rect 466 8 469 9
rect 470 8 475 9
rect 301 7 302 8
rect 305 7 306 8
rect 308 7 309 8
rect 312 7 313 8
rect 319 7 320 8
rect 322 7 323 8
rect 326 7 327 8
rect 330 7 331 8
rect 333 7 334 8
rect 338 7 339 8
rect 342 7 344 8
rect 345 7 346 8
rect 350 7 351 8
rect 358 7 359 8
rect 363 7 364 8
rect 367 7 368 8
rect 370 7 372 8
rect 378 7 379 8
rect 387 7 390 8
rect 392 7 395 8
rect 398 7 401 8
rect 404 7 406 8
rect 407 7 408 8
rect 411 7 412 8
rect 417 7 418 8
rect 420 7 421 8
rect 424 7 425 8
rect 430 7 431 8
rect 434 7 435 8
rect 438 7 439 8
rect 441 7 443 8
rect 447 7 449 8
rect 451 7 452 8
rect 455 7 457 8
rect 459 7 461 8
rect 462 7 463 8
rect 468 7 469 8
rect 472 7 474 8
<< metal3 >>
rect 103 196 104 197
rect 105 196 124 197
rect 97 195 127 196
rect 68 194 73 195
rect 92 194 129 195
rect 67 193 76 194
rect 88 193 131 194
rect 65 192 133 193
rect 65 191 134 192
rect 64 190 135 191
rect 64 189 137 190
rect 63 188 101 189
rect 108 188 138 189
rect 259 188 263 189
rect 269 188 273 189
rect 298 188 303 189
rect 310 188 312 189
rect 323 188 325 189
rect 348 188 351 189
rect 358 188 361 189
rect 366 188 372 189
rect 378 188 380 189
rect 387 188 389 189
rect 395 188 397 189
rect 64 187 72 188
rect 80 187 100 188
rect 111 187 139 188
rect 188 187 193 188
rect 200 187 205 188
rect 211 187 217 188
rect 227 187 230 188
rect 242 187 247 188
rect 259 187 264 188
rect 64 186 70 187
rect 82 186 103 187
rect 116 186 140 187
rect 187 186 194 187
rect 199 186 206 187
rect 54 185 59 186
rect 66 185 67 186
rect 84 185 106 186
rect 121 185 141 186
rect 186 185 195 186
rect 198 185 206 186
rect 210 185 218 187
rect 226 186 230 187
rect 241 186 248 187
rect 225 185 230 186
rect 52 184 61 185
rect 72 184 75 185
rect 85 184 109 185
rect 129 184 142 185
rect 185 184 189 185
rect 51 183 62 184
rect 69 183 77 184
rect 85 183 113 184
rect 133 183 143 184
rect 186 183 189 184
rect 192 183 195 185
rect 51 182 63 183
rect 67 182 79 183
rect 50 181 79 182
rect 85 182 123 183
rect 136 182 144 183
rect 191 182 195 183
rect 197 184 201 185
rect 197 182 200 184
rect 204 182 207 185
rect 209 184 213 185
rect 209 183 212 184
rect 215 183 219 185
rect 224 184 230 185
rect 240 185 249 186
rect 224 183 229 184
rect 240 183 243 185
rect 246 183 249 185
rect 215 182 218 183
rect 223 182 229 183
rect 244 182 249 183
rect 258 182 264 187
rect 268 186 273 188
rect 296 187 304 188
rect 295 186 305 187
rect 309 186 313 188
rect 322 186 326 188
rect 267 184 273 186
rect 294 185 299 186
rect 302 185 306 186
rect 275 184 277 185
rect 283 184 285 185
rect 266 182 272 184
rect 274 183 278 184
rect 282 183 285 184
rect 85 181 127 182
rect 139 181 144 182
rect 190 181 194 182
rect 196 181 200 182
rect 49 179 80 181
rect 85 180 130 181
rect 141 180 144 181
rect 189 180 193 181
rect 48 178 80 179
rect 84 179 133 180
rect 143 179 145 180
rect 188 179 192 180
rect 84 178 136 179
rect 187 178 191 179
rect 47 177 79 178
rect 84 177 139 178
rect 186 177 190 178
rect 46 176 79 177
rect 85 176 141 177
rect 185 176 189 177
rect 196 176 199 181
rect 203 180 207 182
rect 214 181 218 182
rect 222 181 225 182
rect 213 180 217 181
rect 221 180 224 181
rect 226 180 229 182
rect 243 181 248 182
rect 243 180 247 181
rect 203 178 206 180
rect 212 179 216 180
rect 220 179 223 180
rect 225 179 228 180
rect 211 178 215 179
rect 202 177 206 178
rect 210 177 214 178
rect 219 177 230 179
rect 231 177 237 180
rect 244 179 248 180
rect 238 177 241 178
rect 245 177 249 179
rect 257 177 260 182
rect 202 176 205 177
rect 209 176 213 177
rect 219 176 229 177
rect 238 176 242 177
rect 245 176 248 177
rect 45 175 78 176
rect 86 175 144 176
rect 185 175 194 176
rect 196 175 205 176
rect 43 174 77 175
rect 88 174 108 175
rect 112 174 146 175
rect 184 174 194 175
rect 197 174 204 175
rect 42 173 58 174
rect 60 173 75 174
rect 89 173 109 174
rect 114 173 147 174
rect 184 173 193 174
rect 198 173 202 174
rect 208 173 217 176
rect 225 175 228 176
rect 239 175 248 176
rect 256 176 260 177
rect 261 180 264 182
rect 265 180 268 182
rect 261 177 267 180
rect 269 179 272 182
rect 224 173 227 175
rect 239 174 247 175
rect 241 173 245 174
rect 256 173 259 176
rect 261 175 266 177
rect 261 173 265 175
rect 268 174 271 179
rect 275 178 278 183
rect 281 182 285 183
rect 293 183 297 185
rect 303 184 306 185
rect 309 184 312 186
rect 314 184 317 185
rect 323 184 324 185
rect 328 184 330 185
rect 332 184 335 185
rect 347 184 352 188
rect 357 187 362 188
rect 365 187 375 188
rect 356 185 361 187
rect 365 186 376 187
rect 365 185 368 186
rect 372 185 376 186
rect 303 183 305 184
rect 309 183 318 184
rect 322 183 325 184
rect 293 182 296 183
rect 281 181 284 182
rect 280 180 284 181
rect 280 179 283 180
rect 279 178 283 179
rect 275 177 282 178
rect 292 177 296 182
rect 308 182 318 183
rect 308 181 312 182
rect 315 181 319 182
rect 321 181 325 183
rect 327 183 337 184
rect 327 182 332 183
rect 333 182 337 183
rect 346 182 352 184
rect 355 183 361 185
rect 327 181 331 182
rect 308 178 311 181
rect 315 178 318 181
rect 321 178 324 181
rect 327 179 330 181
rect 302 177 305 178
rect 276 176 282 177
rect 293 176 297 177
rect 301 176 305 177
rect 307 177 311 178
rect 276 174 281 176
rect 293 175 304 176
rect 294 174 303 175
rect 267 173 270 174
rect 276 173 280 174
rect 295 173 302 174
rect 307 173 310 177
rect 314 176 318 178
rect 320 177 324 178
rect 314 173 317 176
rect 320 173 323 177
rect 326 176 330 179
rect 334 178 338 182
rect 346 179 349 182
rect 350 179 352 182
rect 354 182 361 183
rect 354 181 357 182
rect 358 181 361 182
rect 364 183 368 185
rect 373 183 376 185
rect 364 182 367 183
rect 372 182 376 183
rect 353 179 356 181
rect 334 177 337 178
rect 333 176 337 177
rect 326 175 331 176
rect 332 175 336 176
rect 345 175 348 179
rect 325 174 335 175
rect 344 174 348 175
rect 350 178 356 179
rect 350 176 355 178
rect 357 176 360 181
rect 364 180 375 182
rect 363 179 373 180
rect 378 179 381 188
rect 386 187 390 188
rect 385 185 390 187
rect 394 187 398 188
rect 394 186 397 187
rect 384 183 390 185
rect 393 185 397 186
rect 393 183 396 185
rect 383 181 386 183
rect 382 180 386 181
rect 382 179 385 180
rect 363 178 367 179
rect 378 178 385 179
rect 387 179 390 183
rect 392 181 395 183
rect 391 179 394 181
rect 363 176 366 178
rect 350 174 354 176
rect 325 173 329 174
rect 330 173 334 174
rect 344 173 347 174
rect 350 173 353 174
rect 356 173 359 176
rect 362 174 366 176
rect 378 176 384 178
rect 387 177 393 179
rect 378 174 383 176
rect 387 175 392 177
rect 362 173 365 174
rect 378 173 382 174
rect 387 173 391 175
rect 40 172 54 173
rect 59 172 74 173
rect 91 172 109 173
rect 116 172 148 173
rect 276 172 279 173
rect 39 171 51 172
rect 57 171 73 172
rect 92 171 109 172
rect 119 171 149 172
rect 275 171 279 172
rect 37 170 49 171
rect 55 170 73 171
rect 93 170 110 171
rect 122 170 150 171
rect 35 169 47 170
rect 54 169 72 170
rect 79 169 86 170
rect 94 169 111 170
rect 126 169 150 170
rect 273 170 278 171
rect 273 169 277 170
rect 325 169 328 173
rect 33 168 46 169
rect 53 168 73 169
rect 31 167 49 168
rect 29 166 50 167
rect 52 166 73 168
rect 79 168 88 169
rect 95 168 113 169
rect 129 168 151 169
rect 79 167 89 168
rect 96 167 114 168
rect 132 167 151 168
rect 28 165 50 166
rect 51 165 73 166
rect 80 165 90 167
rect 96 166 116 167
rect 134 166 151 167
rect 97 165 120 166
rect 136 165 152 166
rect 27 163 74 165
rect 80 164 91 165
rect 98 164 124 165
rect 137 164 152 165
rect 81 163 92 164
rect 98 163 128 164
rect 139 163 152 164
rect 26 161 74 163
rect 27 160 33 161
rect 34 160 74 161
rect 27 159 31 160
rect 33 159 74 160
rect 32 158 74 159
rect 31 157 74 158
rect 80 162 92 163
rect 99 162 130 163
rect 140 162 152 163
rect 80 159 93 162
rect 99 161 132 162
rect 141 161 152 162
rect 100 160 133 161
rect 143 160 153 161
rect 100 159 135 160
rect 144 159 153 160
rect 80 157 94 159
rect 101 158 136 159
rect 145 158 153 159
rect 102 157 137 158
rect 146 157 153 158
rect 30 156 73 157
rect 29 154 73 156
rect 80 156 95 157
rect 103 156 138 157
rect 80 155 96 156
rect 104 155 140 156
rect 147 155 153 157
rect 79 154 96 155
rect 106 154 141 155
rect 148 154 152 155
rect 30 153 72 154
rect 79 153 97 154
rect 109 153 142 154
rect 30 152 71 153
rect 79 152 99 153
rect 115 152 143 153
rect 149 152 152 154
rect 31 151 71 152
rect 78 151 100 152
rect 119 151 144 152
rect 150 151 152 152
rect 189 151 197 152
rect 31 150 48 151
rect 50 150 70 151
rect 78 150 103 151
rect 122 150 144 151
rect 32 149 47 150
rect 33 148 45 149
rect 51 148 69 150
rect 78 149 107 150
rect 124 149 145 150
rect 187 149 197 151
rect 77 148 112 149
rect 127 148 145 149
rect 35 147 40 148
rect 50 147 68 148
rect 77 147 115 148
rect 129 147 145 148
rect 186 148 196 149
rect 46 146 67 147
rect 76 146 118 147
rect 130 146 146 147
rect 40 145 67 146
rect 75 145 120 146
rect 131 145 146 146
rect 35 144 66 145
rect 75 144 122 145
rect 132 144 146 145
rect 186 144 192 148
rect 198 147 204 152
rect 305 150 309 152
rect 304 149 308 150
rect 303 147 308 149
rect 313 147 332 152
rect 302 145 307 147
rect 217 144 219 145
rect 255 144 258 145
rect 274 144 278 145
rect 35 143 65 144
rect 74 143 124 144
rect 133 143 146 144
rect 35 142 64 143
rect 73 142 125 143
rect 35 141 63 142
rect 72 141 126 142
rect 134 141 146 143
rect 36 140 62 141
rect 72 140 127 141
rect 135 140 146 141
rect 183 140 196 144
rect 36 139 61 140
rect 71 139 127 140
rect 37 138 59 139
rect 69 138 94 139
rect 101 138 128 139
rect 136 138 146 140
rect 37 137 57 138
rect 68 137 93 138
rect 103 137 128 138
rect 137 137 146 138
rect 38 136 55 137
rect 67 136 92 137
rect 104 136 129 137
rect 137 136 145 137
rect 38 135 52 136
rect 66 135 92 136
rect 105 135 129 136
rect 39 134 49 135
rect 64 134 92 135
rect 106 134 130 135
rect 39 133 46 134
rect 62 133 91 134
rect 107 133 130 134
rect 138 133 145 136
rect 40 132 43 133
rect 60 132 91 133
rect 98 132 99 133
rect 58 131 91 132
rect 97 131 100 132
rect 108 131 130 133
rect 55 130 90 131
rect 97 130 101 131
rect 53 129 90 130
rect 96 129 101 130
rect 109 130 130 131
rect 139 132 145 133
rect 139 130 144 132
rect 109 129 129 130
rect 51 128 89 129
rect 96 128 102 129
rect 49 127 89 128
rect 95 127 102 128
rect 110 127 129 129
rect 140 128 143 130
rect 140 127 142 128
rect 47 126 88 127
rect 95 126 103 127
rect 46 125 88 126
rect 94 125 103 126
rect 110 126 128 127
rect 140 126 141 127
rect 110 125 127 126
rect 45 124 87 125
rect 44 123 86 124
rect 94 123 104 125
rect 43 122 85 123
rect 93 122 104 123
rect 111 124 127 125
rect 186 124 192 140
rect 198 124 204 144
rect 209 143 214 144
rect 215 143 222 144
rect 209 142 222 143
rect 245 142 250 144
rect 252 143 260 144
rect 272 143 281 144
rect 251 142 261 143
rect 270 142 282 143
rect 301 142 306 145
rect 209 139 221 142
rect 245 141 262 142
rect 269 141 283 142
rect 300 141 306 142
rect 313 141 319 147
rect 245 140 263 141
rect 268 140 284 141
rect 245 139 252 140
rect 257 139 264 140
rect 268 139 274 140
rect 209 138 216 139
rect 209 136 215 138
rect 245 136 251 139
rect 258 137 264 139
rect 259 136 264 137
rect 267 136 273 139
rect 279 138 285 140
rect 280 136 285 138
rect 300 136 305 141
rect 209 124 214 136
rect 245 133 250 136
rect 259 133 265 136
rect 267 133 286 136
rect 299 133 305 136
rect 245 130 251 133
rect 259 131 264 133
rect 245 129 252 130
rect 258 129 264 131
rect 267 132 285 133
rect 267 129 273 132
rect 280 130 281 131
rect 245 128 253 129
rect 257 128 263 129
rect 245 127 263 128
rect 268 128 275 129
rect 279 128 285 130
rect 300 128 305 133
rect 313 136 330 141
rect 268 127 284 128
rect 300 127 306 128
rect 245 126 262 127
rect 269 126 284 127
rect 111 123 126 124
rect 111 122 125 123
rect 43 121 84 122
rect 93 121 105 122
rect 42 120 83 121
rect 92 120 105 121
rect 111 121 124 122
rect 134 121 135 122
rect 111 120 123 121
rect 133 120 135 121
rect 42 119 82 120
rect 41 118 81 119
rect 91 118 105 120
rect 41 117 80 118
rect 90 117 105 118
rect 112 119 121 120
rect 132 119 136 120
rect 112 118 120 119
rect 131 118 135 119
rect 112 117 118 118
rect 130 117 136 118
rect 220 117 243 120
rect 41 116 79 117
rect 89 116 105 117
rect 40 115 78 116
rect 88 115 105 116
rect 111 116 116 117
rect 129 116 136 117
rect 221 116 242 117
rect 245 116 250 126
rect 251 125 261 126
rect 270 125 283 126
rect 253 124 260 125
rect 272 124 281 125
rect 301 124 306 127
rect 313 124 319 136
rect 336 124 342 152
rect 347 151 364 152
rect 380 151 386 152
rect 395 151 398 152
rect 347 150 366 151
rect 377 150 388 151
rect 395 150 399 151
rect 347 149 368 150
rect 376 149 389 150
rect 395 149 400 150
rect 347 147 369 149
rect 375 147 390 149
rect 396 148 400 149
rect 396 147 401 148
rect 347 141 353 147
rect 361 146 370 147
rect 363 145 370 146
rect 364 142 370 145
rect 374 143 380 147
rect 385 146 391 147
rect 386 143 391 146
rect 397 146 401 147
rect 397 144 402 146
rect 363 141 370 142
rect 375 142 380 143
rect 385 142 391 143
rect 375 141 381 142
rect 384 141 390 142
rect 398 141 403 144
rect 347 139 369 141
rect 376 140 389 141
rect 347 138 368 139
rect 377 138 388 140
rect 398 139 404 141
rect 347 137 366 138
rect 376 137 390 138
rect 347 136 364 137
rect 375 136 381 137
rect 384 136 391 137
rect 347 135 354 136
rect 355 135 364 136
rect 374 135 380 136
rect 385 135 391 136
rect 347 124 353 135
rect 358 134 365 135
rect 359 133 366 134
rect 359 132 367 133
rect 360 131 368 132
rect 361 130 368 131
rect 374 130 379 135
rect 361 129 369 130
rect 362 128 369 129
rect 374 129 380 130
rect 386 129 392 135
rect 399 129 404 139
rect 374 128 381 129
rect 385 128 391 129
rect 363 127 370 128
rect 375 127 391 128
rect 398 128 404 129
rect 364 125 371 127
rect 376 126 390 127
rect 377 125 389 126
rect 365 124 372 125
rect 378 124 387 125
rect 398 124 403 128
rect 302 123 306 124
rect 302 121 307 123
rect 397 122 402 124
rect 397 121 401 122
rect 303 120 308 121
rect 304 118 308 120
rect 396 120 401 121
rect 396 119 400 120
rect 395 118 400 119
rect 305 117 309 118
rect 306 116 309 117
rect 395 117 399 118
rect 395 116 398 117
rect 111 115 114 116
rect 128 115 136 116
rect 40 114 76 115
rect 87 114 105 115
rect 126 114 136 115
rect 40 113 75 114
rect 86 113 105 114
rect 125 113 136 114
rect 40 112 73 113
rect 84 112 105 113
rect 123 112 136 113
rect 40 111 71 112
rect 83 111 105 112
rect 122 111 136 112
rect 40 110 69 111
rect 81 110 105 111
rect 120 110 136 111
rect 40 109 66 110
rect 80 109 105 110
rect 118 109 136 110
rect 40 108 64 109
rect 78 108 104 109
rect 116 108 135 109
rect 40 107 62 108
rect 76 107 104 108
rect 113 107 135 108
rect 40 106 60 107
rect 74 106 104 107
rect 110 106 135 107
rect 40 105 59 106
rect 72 105 104 106
rect 106 105 135 106
rect 41 104 57 105
rect 70 104 135 105
rect 41 102 56 104
rect 69 103 134 104
rect 67 102 134 103
rect 41 101 55 102
rect 66 101 134 102
rect 42 100 55 101
rect 64 100 133 101
rect 42 99 54 100
rect 63 99 133 100
rect 43 98 54 99
rect 62 98 132 99
rect 43 97 53 98
rect 44 95 53 97
rect 61 97 87 98
rect 89 97 132 98
rect 61 96 86 97
rect 89 96 131 97
rect 60 95 84 96
rect 88 95 131 96
rect 45 93 53 95
rect 59 94 82 95
rect 59 93 81 94
rect 87 93 130 95
rect 46 92 53 93
rect 58 92 79 93
rect 86 92 129 93
rect 47 91 52 92
rect 58 91 78 92
rect 85 91 128 92
rect 48 90 52 91
rect 49 89 52 90
rect 50 88 52 89
rect 57 90 77 91
rect 85 90 104 91
rect 105 90 127 91
rect 57 89 76 90
rect 84 89 102 90
rect 104 89 127 90
rect 177 90 253 101
rect 266 90 344 101
rect 355 100 429 101
rect 355 99 432 100
rect 355 98 433 99
rect 355 97 434 98
rect 355 96 435 97
rect 355 95 436 96
rect 355 90 437 95
rect 177 89 200 90
rect 57 88 75 89
rect 83 88 101 89
rect 104 88 126 89
rect 51 87 52 88
rect 56 87 74 88
rect 82 87 100 88
rect 103 87 125 88
rect 56 85 73 87
rect 82 86 99 87
rect 103 86 124 87
rect 81 85 98 86
rect 103 85 123 86
rect 56 83 72 85
rect 81 84 97 85
rect 103 84 122 85
rect 177 84 201 89
rect 80 83 97 84
rect 102 83 121 84
rect 177 83 200 84
rect 56 80 71 83
rect 80 81 96 83
rect 102 82 120 83
rect 177 82 201 83
rect 102 81 119 82
rect 57 78 70 80
rect 58 77 70 78
rect 79 79 95 81
rect 102 80 117 81
rect 102 79 116 80
rect 79 77 94 79
rect 59 75 70 77
rect 60 74 70 75
rect 61 73 70 74
rect 62 72 70 73
rect 64 71 70 72
rect 78 76 94 77
rect 102 78 115 79
rect 102 77 113 78
rect 102 76 112 77
rect 78 71 93 76
rect 102 75 111 76
rect 102 74 110 75
rect 102 73 109 74
rect 102 72 108 73
rect 177 72 253 82
rect 102 71 107 72
rect 65 70 70 71
rect 67 69 71 70
rect 68 68 71 69
rect 69 67 71 68
rect 79 67 93 71
rect 103 70 107 71
rect 177 71 202 72
rect 103 69 106 70
rect 103 67 105 69
rect 70 66 71 67
rect 80 65 93 67
rect 81 64 93 65
rect 82 63 93 64
rect 177 65 201 71
rect 177 64 200 65
rect 177 63 201 64
rect 82 62 94 63
rect 83 61 94 62
rect 84 60 94 61
rect 85 59 94 60
rect 177 59 253 63
rect 86 58 95 59
rect 87 57 95 58
rect 178 57 253 59
rect 88 56 95 57
rect 179 56 253 57
rect 90 55 96 56
rect 180 55 253 56
rect 92 54 96 55
rect 181 54 253 55
rect 94 53 97 54
rect 183 53 253 54
rect 293 53 317 90
rect 355 53 379 90
rect 413 76 437 90
rect 388 75 437 76
rect 387 74 415 75
rect 388 73 416 74
rect 389 72 417 73
rect 390 71 419 72
rect 392 70 420 71
rect 393 69 421 70
rect 394 68 422 69
rect 395 67 423 68
rect 396 66 425 67
rect 398 65 426 66
rect 399 64 427 65
rect 400 63 428 64
rect 401 62 430 63
rect 403 61 431 62
rect 404 60 432 61
rect 405 59 433 60
rect 406 58 435 59
rect 408 57 436 58
rect 409 56 437 57
rect 410 55 438 56
rect 411 54 439 55
rect 412 53 441 54
rect 454 53 478 101
rect 414 52 442 53
rect 415 51 443 52
rect 416 50 445 51
rect 417 49 445 50
rect 460 41 465 42
rect 98 40 103 41
rect 8 39 16 40
rect 18 39 26 40
rect 28 39 36 40
rect 39 39 45 40
rect 47 39 56 40
rect 59 39 67 40
rect 68 39 74 40
rect 81 39 88 40
rect 95 39 106 40
rect 116 39 125 40
rect 127 39 136 40
rect 139 39 152 40
rect 156 39 170 40
rect 182 39 191 41
rect 9 38 15 39
rect 20 38 24 39
rect 29 38 35 39
rect 10 32 14 38
rect 19 37 22 38
rect 30 37 35 38
rect 19 36 21 37
rect 31 36 35 37
rect 40 38 44 39
rect 49 38 55 39
rect 61 38 66 39
rect 70 38 75 39
rect 83 38 87 39
rect 93 38 98 39
rect 102 38 106 39
rect 117 38 123 39
rect 129 38 134 39
rect 40 37 43 38
rect 40 36 42 37
rect 18 35 20 36
rect 31 35 36 36
rect 17 34 19 35
rect 32 34 36 35
rect 39 34 41 36
rect 16 33 18 34
rect 32 33 37 34
rect 15 32 18 33
rect 33 32 37 33
rect 38 32 40 34
rect 10 30 19 32
rect 33 31 39 32
rect 10 24 14 30
rect 15 29 20 30
rect 16 27 21 29
rect 17 26 22 27
rect 18 25 23 26
rect 18 24 24 25
rect 9 23 15 24
rect 19 23 25 24
rect 34 23 39 31
rect 49 29 54 38
rect 50 26 54 29
rect 62 35 65 38
rect 71 37 76 38
rect 71 36 77 37
rect 71 35 78 36
rect 62 28 64 35
rect 71 34 79 35
rect 62 27 65 28
rect 62 26 64 27
rect 50 25 55 26
rect 61 25 64 26
rect 51 24 56 25
rect 60 24 64 25
rect 71 24 73 34
rect 74 33 79 34
rect 75 32 80 33
rect 76 31 81 32
rect 77 30 82 31
rect 78 29 83 30
rect 84 29 86 38
rect 92 37 96 38
rect 103 37 106 38
rect 91 36 95 37
rect 104 36 106 37
rect 90 35 95 36
rect 105 35 106 36
rect 118 37 123 38
rect 90 33 94 35
rect 89 29 94 33
rect 118 33 122 37
rect 130 33 134 38
rect 118 31 134 33
rect 99 30 108 31
rect 100 29 108 30
rect 118 30 123 31
rect 129 30 134 31
rect 78 28 86 29
rect 79 27 86 28
rect 80 26 86 27
rect 90 28 94 29
rect 90 26 95 28
rect 81 25 86 26
rect 91 25 96 26
rect 51 23 63 24
rect 70 23 74 24
rect 82 23 86 25
rect 92 24 96 25
rect 93 23 98 24
rect 102 23 106 29
rect 118 24 122 30
rect 130 24 134 30
rect 141 38 146 39
rect 149 38 153 39
rect 141 33 145 38
rect 151 36 153 38
rect 151 35 152 36
rect 150 33 151 34
rect 141 32 146 33
rect 149 32 151 33
rect 141 30 151 32
rect 141 24 145 30
rect 149 29 151 30
rect 150 28 151 29
rect 158 32 163 39
rect 166 38 170 39
rect 168 36 170 38
rect 179 36 195 38
rect 179 35 194 36
rect 197 35 200 41
rect 216 40 234 41
rect 215 38 235 40
rect 216 37 234 38
rect 249 37 263 40
rect 266 37 270 41
rect 300 40 303 41
rect 283 37 297 39
rect 184 34 190 35
rect 167 33 169 34
rect 181 33 192 34
rect 166 32 169 33
rect 158 30 169 32
rect 180 32 193 33
rect 197 32 203 35
rect 230 33 234 37
rect 254 35 258 37
rect 253 34 259 35
rect 252 33 259 34
rect 262 33 270 37
rect 282 36 297 37
rect 288 34 292 36
rect 213 32 237 33
rect 251 32 261 33
rect 180 31 185 32
rect 188 31 194 32
rect 179 30 184 31
rect 190 30 194 31
rect 152 25 154 27
rect 151 24 154 25
rect 158 24 163 30
rect 167 29 169 30
rect 180 29 185 30
rect 188 29 194 30
rect 167 28 168 29
rect 180 28 193 29
rect 182 27 192 28
rect 170 26 171 27
rect 169 25 171 26
rect 183 25 186 26
rect 197 25 200 32
rect 212 31 238 32
rect 250 31 262 32
rect 213 30 238 31
rect 248 30 255 31
rect 257 30 264 31
rect 213 29 237 30
rect 248 29 254 30
rect 259 29 263 30
rect 223 27 226 29
rect 249 28 252 29
rect 261 28 262 29
rect 216 26 234 27
rect 168 24 171 25
rect 118 23 123 24
rect 129 23 135 24
rect 141 23 146 24
rect 150 23 153 24
rect 158 23 164 24
rect 167 23 171 24
rect 182 23 187 25
rect 215 24 234 26
rect 216 23 234 24
rect 8 22 16 23
rect 20 22 26 23
rect 32 22 41 23
rect 52 22 62 23
rect 69 22 76 23
rect 83 22 86 23
rect 94 22 106 23
rect 116 22 125 23
rect 127 22 136 23
rect 139 22 153 23
rect 156 22 170 23
rect 182 22 200 23
rect 55 21 60 22
rect 84 21 85 22
rect 97 21 103 22
rect 182 20 201 22
rect 183 19 200 20
rect 230 19 234 23
rect 252 23 256 27
rect 266 25 270 33
rect 287 32 292 34
rect 299 33 303 40
rect 319 38 337 41
rect 319 37 323 38
rect 357 37 361 41
rect 319 35 337 37
rect 356 35 361 37
rect 319 34 323 35
rect 356 34 362 35
rect 299 32 306 33
rect 319 32 338 34
rect 355 33 363 34
rect 354 32 364 33
rect 287 30 293 32
rect 299 30 307 32
rect 319 31 337 32
rect 353 31 358 32
rect 359 31 366 32
rect 326 30 330 31
rect 351 30 357 31
rect 361 30 367 31
rect 286 29 294 30
rect 285 28 294 29
rect 299 29 306 30
rect 316 29 340 30
rect 350 29 356 30
rect 362 29 366 30
rect 284 27 289 28
rect 283 26 289 27
rect 291 27 296 28
rect 291 26 297 27
rect 282 25 288 26
rect 292 25 298 26
rect 281 24 287 25
rect 294 24 297 25
rect 282 23 286 24
rect 295 23 296 24
rect 252 22 270 23
rect 252 20 271 22
rect 299 20 303 29
rect 315 28 341 29
rect 351 28 354 29
rect 364 28 366 29
rect 316 27 340 28
rect 325 26 331 27
rect 320 25 335 26
rect 319 24 337 25
rect 318 23 324 24
rect 331 23 338 24
rect 318 22 323 23
rect 334 22 338 23
rect 318 21 324 22
rect 332 21 338 22
rect 355 23 358 27
rect 369 25 373 41
rect 391 40 394 41
rect 403 40 407 41
rect 458 40 467 41
rect 388 39 397 40
rect 403 39 408 40
rect 422 39 441 40
rect 457 39 469 40
rect 387 38 408 39
rect 421 38 441 39
rect 386 37 392 38
rect 393 37 408 38
rect 422 37 441 38
rect 386 36 390 37
rect 395 36 408 37
rect 386 34 389 36
rect 396 35 408 36
rect 396 34 400 35
rect 403 34 408 35
rect 386 33 390 34
rect 395 33 408 34
rect 386 32 391 33
rect 394 32 408 33
rect 387 31 408 32
rect 436 35 441 37
rect 456 38 461 39
rect 465 38 470 39
rect 456 37 460 38
rect 466 37 470 38
rect 456 36 461 37
rect 465 36 470 37
rect 456 35 469 36
rect 436 32 440 35
rect 457 34 468 35
rect 459 33 466 34
rect 455 32 472 33
rect 436 31 439 32
rect 388 30 398 31
rect 389 29 396 30
rect 389 23 393 27
rect 403 26 408 31
rect 419 28 444 31
rect 454 30 472 32
rect 473 30 477 41
rect 454 29 470 30
rect 472 29 477 30
rect 403 25 407 26
rect 355 22 373 23
rect 319 20 337 21
rect 355 20 374 22
rect 389 20 408 23
rect 253 19 270 20
rect 300 19 303 20
rect 321 19 336 20
rect 356 19 373 20
rect 389 19 407 20
rect 429 19 433 28
rect 460 26 463 29
rect 467 26 477 29
rect 460 25 462 26
rect 458 23 462 25
rect 473 25 477 26
rect 473 24 476 25
rect 458 20 477 23
rect 458 19 476 20
rect 325 18 332 19
rect 106 14 109 15
rect 127 14 128 15
rect 40 13 43 14
rect 40 8 42 13
rect 46 12 48 14
rect 52 12 55 14
rect 40 7 43 8
rect 46 7 47 12
rect 41 6 44 7
rect 45 6 47 7
rect 52 11 56 12
rect 58 11 60 14
rect 64 13 67 14
rect 71 13 75 14
rect 52 7 53 11
rect 54 10 57 11
rect 59 10 60 11
rect 55 9 60 10
rect 56 8 60 9
rect 57 7 60 8
rect 65 7 67 13
rect 72 12 74 13
rect 77 12 79 14
rect 83 13 86 14
rect 87 13 89 14
rect 93 13 100 14
rect 105 13 110 14
rect 113 13 117 14
rect 120 13 122 14
rect 123 13 128 14
rect 132 13 135 14
rect 72 11 75 12
rect 73 9 75 11
rect 77 10 78 12
rect 76 9 78 10
rect 84 11 86 13
rect 88 12 90 13
rect 84 9 89 11
rect 94 10 96 13
rect 98 11 100 13
rect 104 12 106 13
rect 109 12 110 13
rect 104 11 107 12
rect 97 10 100 11
rect 105 10 109 11
rect 94 9 99 10
rect 106 9 110 10
rect 42 5 46 6
rect 52 5 54 7
rect 58 5 60 7
rect 64 6 67 7
rect 74 7 77 9
rect 84 7 86 9
rect 89 7 90 8
rect 74 6 76 7
rect 64 5 65 6
rect 75 5 76 6
rect 83 6 86 7
rect 88 6 90 7
rect 94 6 96 9
rect 97 8 99 9
rect 107 8 110 9
rect 97 7 100 8
rect 104 7 105 8
rect 108 7 110 8
rect 114 7 116 13
rect 120 12 121 13
rect 123 12 125 13
rect 127 12 128 13
rect 123 8 126 12
rect 133 11 135 13
rect 137 13 139 14
rect 179 13 185 14
rect 137 12 138 13
rect 136 11 138 12
rect 179 11 182 13
rect 123 7 125 8
rect 98 6 101 7
rect 104 6 106 7
rect 108 6 109 7
rect 114 6 117 7
rect 123 6 126 7
rect 134 6 137 11
rect 179 9 185 11
rect 179 7 182 9
rect 179 6 185 7
rect 186 6 188 15
rect 202 13 204 14
rect 224 13 226 15
rect 201 12 204 13
rect 258 12 261 15
rect 264 13 271 14
rect 266 12 269 13
rect 190 11 194 12
rect 189 10 194 11
rect 196 11 210 12
rect 211 11 215 12
rect 196 10 200 11
rect 189 9 191 10
rect 192 9 197 10
rect 189 8 197 9
rect 189 7 191 8
rect 195 7 198 8
rect 201 7 204 11
rect 205 10 216 11
rect 205 7 208 10
rect 209 7 212 10
rect 214 7 216 10
rect 189 6 195 7
rect 196 6 200 7
rect 202 6 208 7
rect 210 6 216 7
rect 217 10 223 12
rect 217 6 219 10
rect 221 6 223 10
rect 224 6 226 12
rect 228 11 232 12
rect 233 11 237 12
rect 227 10 231 11
rect 232 10 237 11
rect 241 11 246 12
rect 248 11 253 12
rect 241 10 247 11
rect 227 8 229 10
rect 232 9 235 10
rect 242 9 247 10
rect 233 8 237 9
rect 227 7 230 8
rect 235 7 237 8
rect 228 6 237 7
rect 241 8 247 9
rect 241 7 243 8
rect 244 7 247 8
rect 241 6 247 7
rect 248 10 254 11
rect 255 10 261 12
rect 248 6 250 10
rect 251 7 257 10
rect 258 7 261 10
rect 251 6 254 7
rect 255 6 261 7
rect 267 6 269 12
rect 271 11 275 12
rect 270 10 276 11
rect 270 9 273 10
rect 274 9 276 10
rect 270 8 276 9
rect 270 7 273 8
rect 271 6 276 7
rect 277 6 279 15
rect 334 14 336 15
rect 334 13 337 14
rect 350 12 352 14
rect 354 13 356 15
rect 380 13 386 14
rect 281 11 285 12
rect 280 10 286 11
rect 287 10 291 12
rect 293 11 297 12
rect 299 11 308 12
rect 310 11 318 12
rect 292 10 298 11
rect 280 9 283 10
rect 284 9 289 10
rect 291 9 294 10
rect 280 8 289 9
rect 292 8 294 9
rect 280 7 282 8
rect 286 7 289 8
rect 291 7 294 8
rect 296 9 298 10
rect 299 10 319 11
rect 299 9 301 10
rect 296 8 301 9
rect 296 7 298 8
rect 280 6 286 7
rect 287 6 298 7
rect 299 6 301 8
rect 83 5 84 6
rect 85 5 87 6
rect 88 5 89 6
rect 94 5 97 6
rect 99 5 101 6
rect 105 5 108 6
rect 114 5 116 6
rect 123 5 124 6
rect 134 5 135 6
rect 180 5 181 6
rect 184 5 185 6
rect 191 5 193 6
rect 198 5 200 6
rect 206 5 207 6
rect 212 5 214 6
rect 218 5 219 6
rect 222 5 223 6
rect 230 5 231 6
rect 233 5 236 6
rect 243 5 244 6
rect 245 5 246 6
rect 248 5 249 6
rect 252 5 253 6
rect 257 5 260 6
rect 267 5 268 6
rect 272 5 275 6
rect 282 5 284 6
rect 289 5 291 6
rect 294 5 296 6
rect 300 5 301 6
rect 303 6 305 10
rect 306 7 309 10
rect 310 7 312 10
rect 306 6 312 7
rect 313 6 315 10
rect 317 6 319 10
rect 320 7 322 12
rect 324 7 326 12
rect 320 6 326 7
rect 327 10 333 12
rect 327 9 330 10
rect 327 7 329 9
rect 327 6 330 7
rect 331 6 333 10
rect 334 9 336 12
rect 338 11 342 12
rect 337 10 342 11
rect 343 10 348 12
rect 349 11 356 12
rect 358 11 363 12
rect 349 10 353 11
rect 337 9 339 10
rect 344 9 348 10
rect 334 8 339 9
rect 343 8 348 9
rect 334 7 336 8
rect 337 7 340 8
rect 342 7 345 8
rect 346 7 348 8
rect 350 7 352 10
rect 354 7 356 11
rect 334 6 337 7
rect 338 6 342 7
rect 343 6 349 7
rect 350 6 356 7
rect 357 10 363 11
rect 357 7 359 10
rect 361 9 363 10
rect 364 10 370 12
rect 372 11 376 12
rect 380 11 382 13
rect 383 12 386 13
rect 422 12 424 15
rect 384 11 386 12
rect 388 11 392 12
rect 394 11 398 12
rect 364 9 367 10
rect 361 8 364 9
rect 365 8 366 9
rect 361 7 363 8
rect 357 6 363 7
rect 364 7 366 8
rect 364 6 367 7
rect 368 6 370 10
rect 371 10 375 11
rect 380 10 386 11
rect 387 10 393 11
rect 394 10 397 11
rect 399 10 404 12
rect 406 10 411 12
rect 371 9 374 10
rect 380 9 385 10
rect 387 9 389 10
rect 391 9 396 10
rect 398 9 401 10
rect 402 9 405 10
rect 407 9 411 10
rect 372 8 376 9
rect 373 7 376 8
rect 371 6 376 7
rect 380 6 382 9
rect 383 8 393 9
rect 394 8 411 9
rect 384 7 386 8
rect 387 7 389 8
rect 396 7 401 8
rect 405 7 407 8
rect 409 7 411 8
rect 384 6 398 7
rect 399 6 404 7
rect 405 6 411 7
rect 412 11 416 12
rect 417 11 421 12
rect 412 10 420 11
rect 422 10 427 12
rect 412 6 414 10
rect 416 8 418 10
rect 416 7 419 8
rect 416 6 421 7
rect 422 6 424 10
rect 426 9 427 10
rect 425 6 427 9
rect 431 6 434 14
rect 449 13 450 14
rect 452 13 454 15
rect 448 12 450 13
rect 456 12 458 14
rect 468 13 470 14
rect 467 12 470 13
rect 435 11 441 12
rect 443 11 446 12
rect 435 10 446 11
rect 447 10 451 12
rect 435 6 437 10
rect 439 6 441 10
rect 442 9 445 10
rect 443 8 447 9
rect 444 7 447 8
rect 442 6 447 7
rect 448 7 450 10
rect 452 7 454 12
rect 455 10 459 12
rect 448 6 454 7
rect 456 7 458 10
rect 460 7 462 12
rect 464 7 466 12
rect 467 10 471 12
rect 472 10 477 12
rect 467 7 470 10
rect 471 9 474 10
rect 475 9 477 10
rect 471 8 478 9
rect 471 7 474 8
rect 456 6 466 7
rect 468 6 471 7
rect 472 6 477 7
rect 303 5 304 6
rect 307 5 308 6
rect 310 5 311 6
rect 314 5 315 6
rect 321 5 322 6
rect 324 5 325 6
rect 328 5 329 6
rect 332 5 333 6
rect 335 5 336 6
rect 340 5 341 6
rect 344 5 346 6
rect 347 5 348 6
rect 352 5 353 6
rect 360 5 361 6
rect 365 5 366 6
rect 369 5 370 6
rect 372 5 374 6
rect 380 5 381 6
rect 389 5 392 6
rect 394 5 397 6
rect 400 5 403 6
rect 406 5 408 6
rect 409 5 410 6
rect 413 5 414 6
rect 419 5 420 6
rect 422 5 423 6
rect 426 5 427 6
rect 432 5 433 6
rect 436 5 437 6
rect 440 5 441 6
rect 443 5 445 6
rect 449 5 451 6
rect 453 5 454 6
rect 457 5 459 6
rect 461 5 463 6
rect 464 5 465 6
rect 470 5 471 6
rect 474 5 476 6
<< end >>
