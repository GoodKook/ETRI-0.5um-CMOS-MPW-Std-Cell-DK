magic
tech scmos
magscale 1 2
timestamp 1727268894
<< nwell >>
rect -12 152 92 272
<< ntransistor >>
rect 20 14 24 34
rect 40 14 44 34
<< ptransistor >>
rect 20 166 24 246
rect 34 166 38 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 46 34
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 34 246
rect 38 166 40 246
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
rect 46 14 58 34
<< pdcontact >>
rect 6 166 18 246
rect 40 166 52 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 20 246 24 250
rect 34 246 38 250
rect 20 109 24 166
rect 34 161 38 166
rect 34 156 44 161
rect 16 97 24 109
rect 20 34 24 97
rect 40 34 44 156
rect 20 10 24 14
rect 40 10 44 14
<< polycontact >>
rect 4 97 16 109
rect 44 97 56 109
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 6 246 18 252
rect 28 166 40 174
rect 28 117 34 166
rect 28 34 34 103
rect 6 8 18 14
rect 46 8 58 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 23 103 37 117
rect 3 83 17 97
rect 43 83 57 97
<< metal2 >>
rect 26 117 34 134
rect 6 66 14 83
rect 46 66 54 83
<< m1p >>
rect -6 252 86 268
rect -6 -8 86 8
<< m2p >>
rect 26 117 34 134
rect 6 66 14 83
rect 46 66 54 83
<< labels >>
rlabel metal1 -6 252 66 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 66 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 30 130 30 130 1 Y
port 3 n signal output
rlabel metal2 10 70 10 70 1 A
port 1 n signal input
rlabel metal2 50 68 50 68 5 B
port 2 n signal input
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
