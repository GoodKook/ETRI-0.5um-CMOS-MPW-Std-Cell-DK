magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 114 114
<< diffusion >>
rect 5 5 53 53
<< metal1 >>
rect 4 4 54 54
<< end >>
