#--------------------------------------------------
# LEF file for Route & Via Rile
#  Ported from osu050 by GoodKook@gmail.com
#

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.15 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.6 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH	    0.9 ;   # ETRI050 Rule: WIDTH=0.8
  SPACING	1.05 ;  # ETRI050 Rule: SPACING=0.8(1.0)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 3.2e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  SPACING	0.9 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.05 ;  # ETRI050 Rule: WIDTH=1.0
  SPACING	1.2 ;   # ETRI050 Rule: SPACING=1.0(1.2)
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 1.6e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.9 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.2 ;   # ETRI050 Rule: WIDTH=1.2
  SPACING	1.2 ;   # ETRI050 Rule: SPACING=1.0(1.2)
  RESISTANCE	RPERSQ 0.05 ;
  CAPACITANCE	CPERSQDIST 1e-05 ;
END metal3

SPACING
  SAMENET cc   via1	0.900 ;
  SAMENET via1 via2	0.900 ;
END SPACING

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via1 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal3 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M3_M2


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via1 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen32

VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	300.000 BY 300.000 ;
END  corner

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	3.000 BY 30.000 ;
END  core

# =====================================================================
#  Core MACROS
# =====================================================================
MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 21.450 8.550 23.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 0.900 30.900 2.700 37.800 ;
        RECT 6.900 30.900 8.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 5.100 1.200 6.900 8.100 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 9.900 30.900 11.700 36.900 ;
        RECT 0.600 16.650 2.400 17.400 ;
        RECT 4.050 10.800 5.100 30.900 ;
        RECT 6.600 24.600 8.400 25.350 ;
        RECT 9.900 18.600 11.100 30.900 ;
        RECT 0.900 9.600 8.400 10.800 ;
        RECT 0.900 2.100 2.700 9.600 ;
        RECT 6.600 9.000 8.400 9.600 ;
        RECT 9.450 5.850 10.500 14.400 ;
        RECT 8.400 5.100 10.500 5.850 ;
        RECT 8.400 2.100 10.200 5.100 ;
  END
END AND2X1
MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 0.900 30.900 2.700 37.800 ;
        RECT 7.500 24.900 9.300 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 5.400 1.200 7.200 8.100 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 0.600 18.600 2.400 19.350 ;
        RECT 3.900 10.800 4.950 30.900 ;
        RECT 10.500 24.900 12.300 36.900 ;
        RECT 6.600 16.650 8.400 17.400 ;
        RECT 10.500 15.600 11.550 24.900 ;
        RECT 0.900 9.900 8.400 10.800 ;
        RECT 0.900 2.100 2.700 9.900 ;
        RECT 6.600 9.000 8.400 9.900 ;
        RECT 9.450 8.100 10.350 11.400 ;
        RECT 8.400 6.300 10.350 8.100 ;
        RECT 8.400 2.100 10.200 6.300 ;
  END
END AND2X2
MACRO AOI21X1
  CLASS CORE ;
  FOREIGN AOI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 3.900 26.700 5.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.500 1.200 3.300 8.100 ;
        RECT 9.000 1.200 10.800 5.100 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.900 ;
        RECT 6.900 25.800 8.700 36.900 ;
        RECT 0.900 24.900 8.700 25.800 ;
        RECT 9.900 24.900 11.700 36.900 ;
        RECT 0.600 16.650 2.400 17.400 ;
        RECT 6.600 16.650 8.400 17.400 ;
        RECT 3.600 15.600 5.400 16.350 ;
        RECT 10.200 15.600 11.100 24.900 ;
        RECT 10.200 8.100 11.100 11.400 ;
        RECT 5.700 6.450 11.100 8.100 ;
        RECT 5.700 2.100 7.500 6.450 ;
  END
END AOI21X1
MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 18.900 40.200 ;
        RECT 3.900 27.000 5.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.500 1.200 3.300 8.100 ;
        RECT 9.900 1.200 11.700 8.100 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 26.100 2.700 36.900 ;
        RECT 6.900 36.000 14.700 36.900 ;
        RECT 6.900 26.100 8.700 36.000 ;
        RECT 0.900 25.200 8.700 26.100 ;
        RECT 9.900 24.000 11.700 35.100 ;
        RECT 12.900 24.900 14.700 36.000 ;
        RECT 7.650 23.100 11.700 24.000 ;
        RECT 7.650 21.600 8.550 23.100 ;
        RECT 7.650 17.400 8.400 21.600 ;
        RECT 3.750 16.650 5.550 17.400 ;
        RECT 0.750 15.600 2.550 16.350 ;
        RECT 7.650 15.600 8.550 17.400 ;
        RECT 9.450 16.650 11.250 17.400 ;
        RECT 12.600 15.600 14.400 16.350 ;
        RECT 6.450 8.100 7.500 11.400 ;
        RECT 5.700 2.100 7.500 8.100 ;
  END
END AOI22X1
MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
        RECT 4.200 24.900 6.000 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 4.200 1.200 6.000 8.100 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 30.900 2.700 36.900 ;
        RECT 0.900 24.000 2.100 30.900 ;
        RECT 7.200 24.900 9.000 36.900 ;
        RECT 0.900 23.100 6.600 24.000 ;
        RECT 4.650 22.200 6.600 23.100 ;
        RECT 0.600 18.600 2.400 19.350 ;
        RECT 4.650 15.600 5.550 22.200 ;
        RECT 7.500 15.600 8.700 24.900 ;
        RECT 4.650 11.400 5.400 15.600 ;
        RECT 4.650 10.800 5.550 11.400 ;
        RECT 4.650 9.900 6.600 10.800 ;
        RECT 1.500 9.000 6.600 9.900 ;
        RECT 1.500 5.100 2.700 9.000 ;
        RECT 7.500 8.100 8.700 11.400 ;
        RECT 0.900 2.100 2.700 5.100 ;
        RECT 7.200 2.100 9.000 8.100 ;
  END
END BUFX2
MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 16.050 40.200 ;
        RECT 4.200 24.900 6.000 37.800 ;
        RECT 10.200 24.900 12.000 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 4.200 1.200 6.000 8.100 ;
        RECT 10.200 1.200 12.000 8.100 ;
        RECT -0.900 -1.200 16.200 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 24.000 2.700 36.900 ;
        RECT 7.200 24.900 9.000 36.900 ;
        RECT 0.900 23.100 6.750 24.000 ;
        RECT 4.950 22.200 6.750 23.100 ;
        RECT 0.600 18.600 2.400 19.350 ;
        RECT 4.950 10.800 6.150 22.200 ;
        RECT 7.650 15.600 8.700 24.900 ;
        RECT 7.650 11.400 8.400 15.600 ;
        RECT 4.950 9.900 6.750 10.800 ;
        RECT 0.900 9.000 6.750 9.900 ;
        RECT 0.900 6.600 2.100 9.000 ;
        RECT 7.650 8.100 8.700 11.400 ;
        RECT 0.900 2.100 2.700 6.600 ;
        RECT 7.200 2.100 9.000 8.100 ;
  END
END BUFX4
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.450 15.450 26.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 30.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 6.900 24.900 8.700 37.800 ;
        RECT 12.900 24.900 14.700 37.800 ;
        RECT 18.900 24.900 20.700 37.800 ;
        RECT 24.900 24.900 26.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT 6.900 1.200 8.700 8.100 ;
        RECT 12.900 1.200 14.700 8.100 ;
        RECT 18.900 1.200 20.700 8.100 ;
        RECT 24.900 1.200 26.700 8.100 ;
        RECT -0.900 -1.200 30.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.000 5.700 36.900 ;
        RECT 9.900 24.000 11.700 36.900 ;
        RECT 15.900 24.000 17.700 36.900 ;
        RECT 21.900 24.000 23.700 36.900 ;
        RECT 3.900 22.800 7.800 24.000 ;
        RECT 9.900 22.800 13.800 24.000 ;
        RECT 15.900 22.800 19.800 24.000 ;
        RECT 21.900 22.800 24.600 24.000 ;
        RECT 3.600 13.650 5.400 14.400 ;
        RECT 6.600 12.300 7.800 22.800 ;
        RECT 9.000 12.300 10.800 12.900 ;
        RECT 6.600 11.100 10.800 12.300 ;
        RECT 12.600 12.300 13.800 22.800 ;
        RECT 15.000 12.300 16.800 12.900 ;
        RECT 12.600 11.100 16.800 12.300 ;
        RECT 18.600 12.300 19.800 22.800 ;
        RECT 23.700 18.600 24.600 22.800 ;
        RECT 21.000 12.300 22.800 12.900 ;
        RECT 18.600 11.100 22.800 12.300 ;
        RECT 6.600 10.200 7.800 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 23.700 10.200 24.600 14.400 ;
        RECT 3.900 9.000 7.800 10.200 ;
        RECT 9.900 9.000 13.800 10.200 ;
        RECT 15.900 9.000 19.800 10.200 ;
        RECT 21.900 9.000 24.600 10.200 ;
        RECT 3.900 2.100 5.700 9.000 ;
        RECT 9.900 2.100 11.700 9.000 ;
        RECT 15.900 2.100 17.700 9.000 ;
        RECT 21.900 2.100 23.700 9.000 ;
  END
END CLKBUF1
MACRO CLKBUF2
  CLASS CORE ;
  FOREIGN CLKBUF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.450 15.450 38.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 42.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 6.900 24.900 8.700 37.800 ;
        RECT 12.900 24.900 14.700 37.800 ;
        RECT 18.900 24.900 20.700 37.800 ;
        RECT 24.900 24.900 26.700 37.800 ;
        RECT 30.900 24.900 32.700 37.800 ;
        RECT 36.900 24.900 38.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT 6.900 1.200 8.700 8.100 ;
        RECT 12.900 1.200 14.700 8.100 ;
        RECT 18.900 1.200 20.700 8.100 ;
        RECT 24.900 1.200 26.700 8.100 ;
        RECT 30.900 1.200 32.700 8.100 ;
        RECT 36.900 1.200 38.700 8.100 ;
        RECT -0.900 -1.200 42.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.000 5.700 36.900 ;
        RECT 9.900 24.000 11.700 36.900 ;
        RECT 15.900 24.000 17.700 36.900 ;
        RECT 21.900 24.000 23.700 36.900 ;
        RECT 27.900 24.000 29.700 36.900 ;
        RECT 33.900 24.000 35.700 36.900 ;
        RECT 3.900 22.800 7.950 24.000 ;
        RECT 9.900 22.800 13.800 24.000 ;
        RECT 15.900 22.800 19.800 24.000 ;
        RECT 21.900 22.800 26.100 24.000 ;
        RECT 27.900 22.800 31.200 24.000 ;
        RECT 33.900 22.800 37.200 24.000 ;
        RECT 3.600 13.650 5.400 14.400 ;
        RECT 6.750 12.300 7.950 22.800 ;
        RECT 9.000 12.300 10.800 12.900 ;
        RECT 6.750 11.100 10.800 12.300 ;
        RECT 12.600 12.300 13.800 22.800 ;
        RECT 15.000 12.300 16.800 12.900 ;
        RECT 12.600 11.100 16.800 12.300 ;
        RECT 18.600 12.300 19.800 22.800 ;
        RECT 21.000 12.300 22.800 12.900 ;
        RECT 18.600 11.100 22.800 12.300 ;
        RECT 24.900 12.300 26.100 22.800 ;
        RECT 27.000 12.300 28.800 12.900 ;
        RECT 24.900 11.100 28.800 12.300 ;
        RECT 30.000 12.300 31.200 22.800 ;
        RECT 36.000 18.600 37.200 22.800 ;
        RECT 33.000 12.300 34.800 12.900 ;
        RECT 30.000 11.100 34.800 12.300 ;
        RECT 6.750 10.200 7.950 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 24.900 10.200 26.100 11.100 ;
        RECT 30.000 10.200 31.200 11.100 ;
        RECT 36.000 10.200 37.200 14.400 ;
        RECT 3.900 9.000 7.950 10.200 ;
        RECT 9.900 9.000 13.800 10.200 ;
        RECT 15.900 9.000 19.800 10.200 ;
        RECT 21.900 9.000 26.100 10.200 ;
        RECT 27.900 9.000 31.200 10.200 ;
        RECT 33.900 9.000 37.200 10.200 ;
        RECT 3.900 2.100 5.700 9.000 ;
        RECT 9.900 2.100 11.700 9.000 ;
        RECT 15.900 2.100 17.700 9.000 ;
        RECT 21.900 2.100 23.700 9.000 ;
        RECT 27.900 2.100 29.700 9.000 ;
        RECT 33.900 2.100 35.700 9.000 ;
  END
END CLKBUF2
MACRO CLKBUF3
  CLASS CORE ;
  FOREIGN CLKBUF3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.450 15.450 50.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 54.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 6.900 24.900 8.700 37.800 ;
        RECT 12.900 24.900 14.700 37.800 ;
        RECT 18.900 24.900 20.700 37.800 ;
        RECT 24.900 24.900 26.700 37.800 ;
        RECT 30.900 24.900 32.700 37.800 ;
        RECT 36.900 24.900 38.700 37.800 ;
        RECT 42.900 24.900 44.700 37.800 ;
        RECT 48.900 24.900 50.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT 6.900 1.200 8.700 8.100 ;
        RECT 12.900 1.200 14.700 8.100 ;
        RECT 18.900 1.200 20.700 8.100 ;
        RECT 24.900 1.200 26.700 8.100 ;
        RECT 30.900 1.200 32.700 8.100 ;
        RECT 36.900 1.200 38.700 8.100 ;
        RECT 42.900 1.200 44.700 8.100 ;
        RECT 48.900 1.200 50.700 8.100 ;
        RECT -0.900 -1.200 55.200 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.000 5.700 36.900 ;
        RECT 9.900 24.000 11.700 36.900 ;
        RECT 15.900 24.000 17.700 36.900 ;
        RECT 21.900 24.000 23.700 36.900 ;
        RECT 27.900 24.000 29.700 36.900 ;
        RECT 33.900 24.000 35.700 36.900 ;
        RECT 39.900 24.000 41.700 36.900 ;
        RECT 45.900 24.000 47.700 36.900 ;
        RECT 3.900 22.800 7.800 24.000 ;
        RECT 9.900 22.800 13.800 24.000 ;
        RECT 15.900 22.800 19.800 24.000 ;
        RECT 21.900 22.800 26.100 24.000 ;
        RECT 27.900 22.800 31.200 24.000 ;
        RECT 33.900 22.800 37.800 24.000 ;
        RECT 39.900 22.800 42.900 24.000 ;
        RECT 45.900 22.800 49.050 24.000 ;
        RECT 3.600 13.650 5.400 14.400 ;
        RECT 6.750 12.900 7.800 22.800 ;
        RECT 12.600 12.900 13.800 22.800 ;
        RECT 18.600 12.900 19.800 22.800 ;
        RECT 24.900 12.900 26.100 22.800 ;
        RECT 30.000 12.900 31.200 22.800 ;
        RECT 36.600 12.900 37.800 22.800 ;
        RECT 41.700 12.900 42.900 22.800 ;
        RECT 47.850 18.600 49.050 22.800 ;
        RECT 6.750 11.100 10.800 12.900 ;
        RECT 12.600 11.100 16.800 12.900 ;
        RECT 18.600 11.100 22.800 12.900 ;
        RECT 24.900 11.100 28.800 12.900 ;
        RECT 30.000 11.100 34.800 12.900 ;
        RECT 36.600 11.100 40.800 12.900 ;
        RECT 41.700 11.100 46.800 12.900 ;
        RECT 6.750 10.200 7.800 11.100 ;
        RECT 12.600 10.200 13.800 11.100 ;
        RECT 18.600 10.200 19.800 11.100 ;
        RECT 24.900 10.200 26.100 11.100 ;
        RECT 30.000 10.200 31.200 11.100 ;
        RECT 36.600 10.200 37.800 11.100 ;
        RECT 41.700 10.200 42.900 11.100 ;
        RECT 47.850 10.200 49.050 14.400 ;
        RECT 3.900 9.000 7.800 10.200 ;
        RECT 9.900 9.000 13.800 10.200 ;
        RECT 15.900 9.000 19.800 10.200 ;
        RECT 21.900 9.000 26.100 10.200 ;
        RECT 27.900 9.000 31.200 10.200 ;
        RECT 33.900 9.000 37.800 10.200 ;
        RECT 39.900 9.000 42.900 10.200 ;
        RECT 45.900 9.000 49.050 10.200 ;
        RECT 3.900 2.100 5.700 9.000 ;
        RECT 9.900 2.100 11.700 9.000 ;
        RECT 15.900 2.100 17.700 9.000 ;
        RECT 21.900 2.100 23.700 9.000 ;
        RECT 27.900 2.100 29.700 9.000 ;
        RECT 33.900 2.100 35.700 9.000 ;
        RECT 39.900 2.100 41.700 9.000 ;
        RECT 45.900 2.100 47.700 9.000 ;
  END
END CLKBUF3
MACRO DFFNEGX1
  CLASS CORE ;
  FOREIGN DFFNEGX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 15.450 12.450 17.550 14.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 15.450 32.550 17.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 36.900 40.200 ;
        RECT 3.900 30.900 5.700 37.800 ;
        RECT 13.500 30.900 15.300 37.800 ;
        RECT 20.100 30.900 21.900 37.800 ;
        RECT 29.100 33.900 30.900 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 5.100 ;
        RECT 13.200 1.200 15.000 5.100 ;
        RECT 20.100 1.200 21.900 5.100 ;
        RECT 29.100 1.200 30.900 5.100 ;
        RECT -0.900 -1.200 36.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 24.300 2.700 36.900 ;
        RECT 8.700 32.100 10.500 36.900 ;
        RECT 6.900 30.900 10.500 32.100 ;
        RECT 6.900 30.300 8.550 30.900 ;
        RECT 6.450 28.200 8.550 30.300 ;
        RECT 16.500 30.000 18.300 36.900 ;
        RECT 24.600 30.900 26.400 36.900 ;
        RECT 9.600 27.300 11.400 30.000 ;
        RECT 12.600 28.800 19.200 30.000 ;
        RECT 24.300 28.800 26.400 30.900 ;
        RECT 12.600 28.200 14.400 28.800 ;
        RECT 17.400 28.200 19.200 28.800 ;
        RECT 9.450 25.200 11.550 27.300 ;
        RECT 25.200 27.000 27.000 27.600 ;
        RECT 20.100 25.800 27.000 27.000 ;
        RECT 20.100 25.200 21.900 25.800 ;
        RECT 20.100 24.300 21.000 25.200 ;
        RECT 0.900 23.100 21.000 24.300 ;
        RECT 32.100 24.900 33.900 36.900 ;
        RECT 0.900 8.100 1.800 23.100 ;
        RECT 7.800 22.500 9.600 23.100 ;
        RECT 14.400 21.600 16.200 22.200 ;
        RECT 6.450 20.400 16.200 21.600 ;
        RECT 24.300 21.000 26.400 21.600 ;
        RECT 29.400 21.000 31.200 21.600 ;
        RECT 6.450 19.500 8.550 20.400 ;
        RECT 24.300 19.800 31.200 21.000 ;
        RECT 24.300 19.500 26.400 19.800 ;
        RECT 3.600 18.600 5.400 19.350 ;
        RECT 32.100 18.600 33.300 24.900 ;
        RECT 27.000 15.450 29.400 17.250 ;
        RECT 9.450 11.400 11.550 13.200 ;
        RECT 2.850 10.200 23.700 11.400 ;
        RECT 2.850 9.600 4.650 10.200 ;
        RECT 7.800 9.000 9.600 10.200 ;
        RECT 21.900 9.600 23.700 10.200 ;
        RECT 32.100 8.100 33.300 14.400 ;
        RECT 0.900 2.100 2.700 8.100 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 12.600 7.200 14.400 7.800 ;
        RECT 12.600 6.000 17.700 7.200 ;
        RECT 6.900 5.100 8.550 6.000 ;
        RECT 16.500 5.100 17.700 6.000 ;
        RECT 6.900 4.050 10.500 5.100 ;
        RECT 8.700 2.100 10.500 4.050 ;
        RECT 16.500 2.100 18.300 5.100 ;
        RECT 24.300 4.200 26.400 7.200 ;
        RECT 24.600 2.100 26.400 4.200 ;
        RECT 32.100 2.100 33.900 8.100 ;
      LAYER metal2 ;
        RECT 6.450 28.200 8.550 30.300 ;
        RECT 24.300 28.800 26.400 30.900 ;
        RECT 7.050 21.600 8.100 28.200 ;
        RECT 9.450 25.200 11.550 27.300 ;
        RECT 6.450 19.500 8.550 21.600 ;
        RECT 7.050 8.100 8.100 19.500 ;
        RECT 10.050 13.200 11.400 25.200 ;
        RECT 24.300 21.600 25.500 28.800 ;
        RECT 24.300 19.500 26.400 21.600 ;
        RECT 9.450 11.100 11.550 13.200 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 24.300 7.200 25.500 19.500 ;
        RECT 24.300 5.100 26.400 7.200 ;
  END
END DFFNEGX1
MACRO DFFPOSX1
  CLASS CORE ;
  FOREIGN DFFPOSX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 18.450 15.450 20.550 17.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 12.450 32.550 14.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 36.900 40.200 ;
        RECT 4.650 30.900 6.450 37.800 ;
        RECT 14.850 30.900 16.650 37.800 ;
        RECT 21.450 30.900 23.250 37.800 ;
        RECT 30.150 33.900 31.950 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 4.650 1.200 6.450 5.100 ;
        RECT 13.950 1.200 15.750 5.100 ;
        RECT 20.850 1.200 22.650 5.100 ;
        RECT 29.850 1.200 31.650 5.100 ;
        RECT -0.900 -1.200 36.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.650 24.900 3.450 36.900 ;
        RECT 10.050 30.900 11.850 36.900 ;
        RECT 10.050 30.000 11.250 30.900 ;
        RECT 17.850 30.000 19.650 36.900 ;
        RECT 25.650 30.900 27.450 36.900 ;
        RECT 6.450 27.900 11.250 30.000 ;
        RECT 13.950 28.950 20.550 30.000 ;
        RECT 13.950 28.200 15.750 28.950 ;
        RECT 18.750 28.200 20.550 28.950 ;
        RECT 25.650 28.800 29.550 30.900 ;
        RECT 10.050 27.000 11.250 27.900 ;
        RECT 22.950 27.300 24.750 27.900 ;
        RECT 10.050 25.800 17.550 27.000 ;
        RECT 15.750 25.200 17.550 25.800 ;
        RECT 18.450 26.400 24.750 27.300 ;
        RECT 1.650 24.000 2.550 24.900 ;
        RECT 18.450 24.300 19.350 26.400 ;
        RECT 22.950 26.100 24.750 26.400 ;
        RECT 25.650 26.100 28.350 27.900 ;
        RECT 25.650 25.200 26.550 26.100 ;
        RECT 10.950 24.000 19.350 24.300 ;
        RECT 1.650 23.400 19.350 24.000 ;
        RECT 20.550 24.300 26.550 25.200 ;
        RECT 27.450 24.300 29.550 25.200 ;
        RECT 33.150 24.900 34.950 36.900 ;
        RECT 1.650 22.800 12.750 23.400 ;
        RECT 1.650 8.100 2.550 22.800 ;
        RECT 10.950 22.500 12.750 22.800 ;
        RECT 6.600 17.700 11.400 18.900 ;
        RECT 20.550 18.600 21.450 24.300 ;
        RECT 27.450 23.100 31.650 24.300 ;
        RECT 30.750 21.300 32.550 23.100 ;
        RECT 6.600 17.100 8.400 17.700 ;
        RECT 3.600 13.650 5.400 15.450 ;
        RECT 33.750 14.550 34.950 24.900 ;
        RECT 4.500 12.900 5.400 13.650 ;
        RECT 20.550 13.500 21.450 14.400 ;
        RECT 9.600 12.900 11.400 13.500 ;
        RECT 20.550 12.900 22.350 13.500 ;
        RECT 4.500 11.700 22.350 12.900 ;
        RECT 28.650 12.450 29.400 14.250 ;
        RECT 33.600 12.450 34.950 14.550 ;
        RECT 10.350 8.700 11.400 11.700 ;
        RECT 1.650 2.100 3.450 8.100 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 10.050 6.900 11.850 8.700 ;
        RECT 13.350 7.950 15.150 8.700 ;
        RECT 33.750 8.100 34.950 12.450 ;
        RECT 13.350 6.900 18.300 7.950 ;
        RECT 27.450 7.200 29.550 8.100 ;
        RECT 7.500 5.100 8.550 6.000 ;
        RECT 17.250 5.100 18.300 6.900 ;
        RECT 25.800 6.000 29.550 7.200 ;
        RECT 25.800 5.100 26.850 6.000 ;
        RECT 7.500 4.200 11.250 5.100 ;
        RECT 9.450 2.100 11.250 4.200 ;
        RECT 17.250 2.100 19.050 5.100 ;
        RECT 25.050 2.100 26.850 5.100 ;
        RECT 33.150 2.100 34.950 8.100 ;
      LAYER metal2 ;
        RECT 6.450 27.900 8.550 30.000 ;
        RECT 27.450 28.800 29.550 30.900 ;
        RECT 7.200 8.100 8.400 27.900 ;
        RECT 27.450 25.200 28.650 28.800 ;
        RECT 27.450 23.100 29.550 25.200 ;
        RECT 27.450 8.100 28.650 23.100 ;
        RECT 6.450 6.000 8.550 8.100 ;
        RECT 27.450 6.000 29.550 8.100 ;
  END
END DFFPOSX1
MACRO DFFSR
  CLASS CORE ;
  FOREIGN DFFSR ;
  ORIGIN 0.000 0.000 ;
  SIZE 72.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 21.450 5.550 23.550 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END S
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.450 12.450 29.550 14.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 57.450 18.450 59.550 20.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 66.450 15.450 68.550 17.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 72.900 40.200 ;
        RECT 1.200 30.900 3.000 37.800 ;
        RECT 7.200 30.900 9.000 37.800 ;
        RECT 13.200 32.100 15.000 37.800 ;
        RECT 25.800 30.900 27.600 37.800 ;
        RECT 32.700 30.900 34.500 37.800 ;
        RECT 48.900 30.900 50.700 37.800 ;
        RECT 54.900 30.900 56.700 37.800 ;
        RECT 60.900 30.900 62.700 37.800 ;
        RECT 67.500 30.900 69.300 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 6.600 1.200 8.400 8.100 ;
        RECT 25.200 1.200 27.000 5.100 ;
        RECT 32.700 1.200 34.500 5.100 ;
        RECT 55.200 1.200 57.000 8.100 ;
        RECT 67.500 1.200 69.300 5.100 ;
        RECT -0.900 -1.200 72.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 4.200 30.900 6.000 36.900 ;
        RECT 4.200 30.000 5.250 30.900 ;
        RECT 1.200 29.100 5.250 30.000 ;
        RECT 1.200 12.900 2.400 29.100 ;
        RECT 5.700 27.900 7.500 28.200 ;
        RECT 10.200 27.900 12.000 36.900 ;
        RECT 16.350 33.900 18.600 36.900 ;
        RECT 19.500 33.900 21.600 36.900 ;
        RECT 22.650 33.900 24.600 36.900 ;
        RECT 16.350 31.200 17.250 33.900 ;
        RECT 19.500 31.200 20.550 33.900 ;
        RECT 22.650 31.200 23.850 33.900 ;
        RECT 15.150 29.100 17.250 31.200 ;
        RECT 18.450 29.100 20.550 31.200 ;
        RECT 21.750 29.100 23.850 31.200 ;
        RECT 29.700 29.400 31.500 36.900 ;
        RECT 35.700 30.900 37.500 36.900 ;
        RECT 39.300 33.900 41.100 36.900 ;
        RECT 39.000 31.800 41.100 33.900 ;
        RECT 42.300 33.900 44.100 36.900 ;
        RECT 45.300 33.900 47.100 36.900 ;
        RECT 42.300 31.800 44.400 33.900 ;
        RECT 45.750 31.800 47.850 33.900 ;
        RECT 5.700 26.700 24.900 27.900 ;
        RECT 29.700 27.300 32.550 29.400 ;
        RECT 35.400 28.650 37.500 30.900 ;
        RECT 43.350 30.000 44.400 31.800 ;
        RECT 51.900 30.000 53.700 36.900 ;
        RECT 57.900 30.900 59.700 36.900 ;
        RECT 43.350 28.800 51.000 30.000 ;
        RECT 51.900 28.800 57.600 30.000 ;
        RECT 35.400 26.850 38.400 28.650 ;
        RECT 49.200 28.200 51.000 28.800 ;
        RECT 55.800 28.200 57.600 28.800 ;
        RECT 5.700 26.400 7.500 26.700 ;
        RECT 23.700 25.950 24.900 26.700 ;
        RECT 39.450 25.950 41.550 27.000 ;
        RECT 9.000 25.200 10.800 25.800 ;
        RECT 18.450 25.200 20.550 25.800 ;
        RECT 9.000 24.000 20.550 25.200 ;
        RECT 23.700 24.900 41.550 25.950 ;
        RECT 45.450 25.800 47.550 27.000 ;
        RECT 58.500 25.800 59.700 30.900 ;
        RECT 64.500 30.900 66.300 36.900 ;
        RECT 45.450 24.900 62.400 25.800 ;
        RECT 18.450 23.700 20.550 24.000 ;
        RECT 23.700 22.800 60.600 24.000 ;
        RECT 23.700 22.200 24.900 22.800 ;
        RECT 58.800 22.200 60.600 22.800 ;
        RECT 11.550 21.600 24.900 22.200 ;
        RECT 12.600 21.300 24.900 21.600 ;
        RECT 3.600 18.750 5.400 20.400 ;
        RECT 12.600 18.750 13.350 21.300 ;
        RECT 30.450 19.800 32.550 21.900 ;
        RECT 36.450 21.600 38.550 21.900 ;
        RECT 34.650 19.800 38.550 21.600 ;
        RECT 43.200 19.800 45.000 21.600 ;
        RECT 4.200 18.600 5.400 18.750 ;
        RECT 4.200 16.950 5.550 18.600 ;
        RECT 14.250 18.300 21.000 19.350 ;
        RECT 14.250 16.950 15.450 18.300 ;
        RECT 4.200 15.750 15.450 16.950 ;
        RECT 17.250 15.600 19.050 17.400 ;
        RECT 19.950 16.800 21.000 18.300 ;
        RECT 21.900 18.600 32.550 19.800 ;
        RECT 44.100 18.600 45.000 19.800 ;
        RECT 21.900 18.000 23.700 18.600 ;
        RECT 30.450 17.700 45.000 18.600 ;
        RECT 48.300 18.300 53.400 20.100 ;
        RECT 48.300 16.800 49.200 18.300 ;
        RECT 19.950 15.600 49.200 16.800 ;
        RECT 56.100 17.400 56.400 20.550 ;
        RECT 56.100 15.600 57.300 17.400 ;
        RECT 1.200 11.700 16.500 12.900 ;
        RECT 1.200 8.100 2.400 11.700 ;
        RECT 5.400 10.200 7.200 10.800 ;
        RECT 5.400 9.000 13.800 10.200 ;
        RECT 12.300 8.100 13.800 9.000 ;
        RECT 15.450 8.100 16.500 11.700 ;
        RECT 18.000 10.500 19.050 15.600 ;
        RECT 50.400 14.400 57.300 15.600 ;
        RECT 24.300 12.450 26.400 14.250 ;
        RECT 50.400 14.100 51.900 14.400 ;
        RECT 33.600 12.600 51.900 14.100 ;
        RECT 54.000 13.200 55.800 13.500 ;
        RECT 58.800 13.200 60.600 13.500 ;
        RECT 21.300 10.500 23.100 12.300 ;
        RECT 18.000 9.300 27.900 10.500 ;
        RECT 33.600 10.200 35.400 12.600 ;
        RECT 52.800 11.700 60.600 13.200 ;
        RECT 41.400 9.900 48.000 11.700 ;
        RECT 27.000 8.100 27.900 9.300 ;
        RECT 52.800 8.100 54.300 11.700 ;
        RECT 61.500 8.100 62.400 24.900 ;
        RECT 1.200 2.100 3.000 8.100 ;
        RECT 12.000 2.100 13.800 8.100 ;
        RECT 15.150 6.000 17.550 8.100 ;
        RECT 18.450 6.000 20.550 8.100 ;
        RECT 21.750 6.000 23.850 8.100 ;
        RECT 27.000 6.300 28.800 8.100 ;
        RECT 16.200 5.100 17.550 6.000 ;
        RECT 19.200 5.100 20.550 6.000 ;
        RECT 22.200 5.100 23.850 6.000 ;
        RECT 30.450 6.000 32.550 8.100 ;
        RECT 35.850 6.000 37.950 8.100 ;
        RECT 39.150 6.000 41.250 8.100 ;
        RECT 42.450 6.000 44.550 8.100 ;
        RECT 45.750 6.000 47.850 8.100 ;
        RECT 50.100 6.900 54.300 8.100 ;
        RECT 30.450 5.100 31.500 6.000 ;
        RECT 35.850 5.100 37.500 6.000 ;
        RECT 16.200 2.100 18.000 5.100 ;
        RECT 19.200 2.100 21.000 5.100 ;
        RECT 22.200 2.100 24.000 5.100 ;
        RECT 29.700 2.100 31.500 5.100 ;
        RECT 35.700 2.100 37.500 5.100 ;
        RECT 39.300 2.100 41.100 6.000 ;
        RECT 42.450 5.100 44.100 6.000 ;
        RECT 45.750 5.100 47.100 6.000 ;
        RECT 42.300 2.100 44.100 5.100 ;
        RECT 45.300 2.100 47.100 5.100 ;
        RECT 50.100 2.100 51.900 6.900 ;
        RECT 60.600 2.100 62.400 8.100 ;
        RECT 64.500 18.600 66.000 30.900 ;
        RECT 64.500 14.400 65.400 18.600 ;
        RECT 64.500 5.100 66.000 14.400 ;
        RECT 64.500 2.100 66.300 5.100 ;
      LAYER metal2 ;
        RECT 39.000 31.800 41.100 33.900 ;
        RECT 42.300 31.800 44.400 33.900 ;
        RECT 15.150 29.100 17.250 31.200 ;
        RECT 18.450 29.100 20.550 31.200 ;
        RECT 21.750 29.100 23.850 31.200 ;
        RECT 15.900 8.100 17.100 29.100 ;
        RECT 18.900 25.800 20.100 29.100 ;
        RECT 18.450 23.700 20.550 25.800 ;
        RECT 19.350 8.100 20.550 23.700 ;
        RECT 22.350 8.100 23.550 29.100 ;
        RECT 30.450 27.300 32.550 29.400 ;
        RECT 35.400 28.800 37.650 30.900 ;
        RECT 30.450 21.900 31.650 27.300 ;
        RECT 36.450 21.900 37.650 28.800 ;
        RECT 39.900 27.000 41.100 31.800 ;
        RECT 43.350 28.800 44.400 31.800 ;
        RECT 45.750 31.800 47.850 33.900 ;
        RECT 39.450 24.900 41.550 27.000 ;
        RECT 30.450 19.800 32.550 21.900 ;
        RECT 36.450 19.800 38.550 21.900 ;
        RECT 31.050 8.100 32.250 19.800 ;
        RECT 36.450 8.100 37.650 19.800 ;
        RECT 39.750 8.100 41.250 24.900 ;
        RECT 43.350 8.100 44.550 28.800 ;
        RECT 45.750 27.000 46.950 31.800 ;
        RECT 45.450 24.900 47.550 27.000 ;
        RECT 15.150 6.000 17.250 8.100 ;
        RECT 18.450 6.000 20.550 8.100 ;
        RECT 21.750 6.000 23.850 8.100 ;
        RECT 30.450 6.000 32.550 8.100 ;
        RECT 35.850 6.000 37.950 8.100 ;
        RECT 39.150 6.000 41.250 8.100 ;
        RECT 42.450 6.000 44.550 8.100 ;
        RECT 45.750 8.100 46.950 24.900 ;
        RECT 45.750 6.000 47.850 8.100 ;
  END
END DFFSR
MACRO FAX1
  CLASS CORE ;
  FOREIGN FAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
        RECT 3.600 11.700 5.100 15.450 ;
        RECT 3.600 10.800 14.400 11.700 ;
      LAYER metal2 ;
        RECT 3.450 15.450 5.550 17.550 ;
        RECT 3.900 12.900 5.100 15.450 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 16.500 32.550 17.550 ;
        RECT 28.800 15.600 32.550 16.500 ;
        RECT 17.400 14.550 32.550 15.600 ;
      LAYER metal2 ;
        RECT 30.450 15.450 32.550 17.550 ;
        RECT 30.900 12.900 32.100 15.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
      LAYER metal2 ;
        RECT 6.900 17.550 8.100 20.100 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END C
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 35.700 32.250 37.500 36.900 ;
        RECT 35.400 30.900 37.500 32.250 ;
        RECT 35.400 23.400 36.300 30.900 ;
        RECT 35.400 22.500 38.250 23.400 ;
        RECT 37.350 17.550 38.250 22.500 ;
        RECT 36.450 15.450 38.550 17.550 ;
        RECT 37.350 7.200 38.250 15.450 ;
        RECT 36.000 6.000 38.250 7.200 ;
        RECT 36.000 5.100 36.900 6.000 ;
        RECT 35.700 2.100 37.500 5.100 ;
      LAYER metal2 ;
        RECT 36.450 15.450 38.550 17.550 ;
        RECT 36.900 12.900 38.100 15.450 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 42.300 30.900 44.100 36.900 ;
        RECT 42.300 23.400 43.500 30.900 ;
        RECT 39.450 22.200 43.500 23.400 ;
        RECT 39.450 17.550 40.650 22.200 ;
        RECT 39.450 15.450 41.550 17.550 ;
        RECT 39.450 5.100 40.500 15.450 ;
        RECT 39.300 2.100 41.100 5.100 ;
      LAYER metal2 ;
        RECT 39.900 17.550 41.100 20.100 ;
        RECT 39.450 15.450 41.550 17.550 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 45.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 45.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.750 ;
        RECT 3.900 27.000 5.700 36.750 ;
        RECT 6.900 27.000 8.700 36.750 ;
        RECT 6.900 25.800 8.250 27.000 ;
        RECT 9.900 26.100 11.700 36.750 ;
        RECT 0.900 24.900 8.250 25.800 ;
        RECT 9.450 24.000 11.550 26.100 ;
        RECT 14.400 24.900 16.200 36.750 ;
        RECT 17.400 27.000 19.200 36.750 ;
        RECT 20.400 27.900 22.200 36.750 ;
        RECT 23.400 27.000 25.200 36.750 ;
        RECT 17.400 26.100 25.200 27.000 ;
        RECT 26.400 24.000 28.350 36.750 ;
        RECT 32.700 30.900 34.500 36.750 ;
        RECT 39.300 30.900 41.100 36.750 ;
        RECT 37.500 26.400 39.600 26.550 ;
        RECT 37.500 24.600 41.400 26.400 ;
        RECT 37.500 24.450 39.600 24.600 ;
        RECT 21.450 21.900 23.550 24.000 ;
        RECT 24.450 21.900 28.350 24.000 ;
        RECT 21.900 21.300 23.550 21.900 ;
        RECT 21.900 19.500 23.700 21.300 ;
        RECT 27.450 21.150 28.350 21.900 ;
        RECT 27.450 20.250 36.300 21.150 ;
        RECT 34.500 19.350 36.300 20.250 ;
        RECT 0.900 7.200 8.100 8.100 ;
        RECT 9.450 7.800 11.550 9.900 ;
        RECT 24.450 8.700 27.450 10.800 ;
        RECT 0.900 2.250 2.700 7.200 ;
        RECT 3.900 2.250 5.700 6.300 ;
        RECT 6.900 2.250 8.700 7.200 ;
        RECT 9.900 6.900 11.550 7.800 ;
        RECT 9.900 2.250 11.700 6.900 ;
        RECT 14.400 2.250 16.200 7.500 ;
        RECT 17.400 6.900 25.200 7.800 ;
        RECT 17.400 2.250 19.200 6.900 ;
        RECT 20.400 2.250 22.200 6.000 ;
        RECT 23.400 2.250 25.200 6.900 ;
        RECT 26.400 6.600 27.450 8.700 ;
        RECT 26.400 2.250 28.350 6.600 ;
        RECT 32.700 2.250 34.500 5.100 ;
        RECT 42.300 2.250 44.100 5.100 ;
      LAYER metal2 ;
        RECT 37.500 26.100 39.600 26.550 ;
        RECT 9.450 25.200 39.600 26.100 ;
        RECT 9.450 24.000 11.550 25.200 ;
        RECT 10.050 9.900 10.950 24.000 ;
        RECT 21.450 21.900 23.550 25.200 ;
        RECT 37.500 24.450 39.600 25.200 ;
        RECT 24.450 21.900 26.550 24.000 ;
        RECT 25.050 10.800 26.250 21.900 ;
        RECT 9.450 7.800 11.550 9.900 ;
        RECT 24.450 8.700 26.550 10.800 ;
  END
END FAX1
MACRO FILL
  CLASS CORE ;
  FOREIGN FILL ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 3.900 1.200 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 3.900 40.200 ;
    END
  END vdd
END FILL
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 15.450 2.550 17.550 ;
      LAYER metal2 ;
        RECT 0.450 15.450 2.550 17.550 ;
        RECT 0.900 12.900 2.100 15.450 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.450 17.550 17.550 ;
      LAYER metal2 ;
        RECT 15.900 17.550 17.100 20.100 ;
        RECT 15.450 15.450 17.550 17.550 ;
    END
  END B
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 23.700 30.900 25.500 36.900 ;
        RECT 23.700 17.550 24.600 30.900 ;
        RECT 21.450 15.450 24.600 17.550 ;
        RECT 23.700 12.450 24.600 15.450 ;
        RECT 23.700 11.550 28.200 12.450 ;
        RECT 27.300 5.100 28.200 11.550 ;
        RECT 27.300 2.100 29.100 5.100 ;
      LAYER metal2 ;
        RECT 21.450 15.450 23.550 17.550 ;
        RECT 21.900 12.900 23.100 15.450 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.500 30.900 12.300 36.900 ;
        RECT 10.500 17.550 11.550 30.900 ;
        RECT 9.450 15.450 11.550 17.550 ;
        RECT 8.700 4.950 10.800 7.200 ;
        RECT 8.700 2.100 10.500 4.950 ;
      LAYER metal2 ;
        RECT 9.900 17.550 11.100 20.100 ;
        RECT 9.450 15.450 11.550 17.550 ;
        RECT 10.200 7.200 11.400 15.450 ;
        RECT 8.700 5.100 11.400 7.200 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 30.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 30.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 30.900 2.700 36.750 ;
        RECT 3.900 31.500 5.700 36.750 ;
        RECT 1.200 30.600 2.700 30.900 ;
        RECT 6.900 30.900 8.700 36.750 ;
        RECT 13.500 30.900 15.300 36.750 ;
        RECT 6.900 30.600 8.100 30.900 ;
        RECT 1.200 29.700 8.100 30.600 ;
        RECT 7.050 17.850 8.100 29.700 ;
        RECT 16.500 24.900 18.300 36.750 ;
        RECT 20.700 30.900 22.500 36.750 ;
        RECT 16.650 22.950 17.550 24.900 ;
        RECT 16.650 22.050 19.950 22.950 ;
        RECT 6.450 15.750 8.550 17.850 ;
        RECT 18.600 14.250 19.950 22.050 ;
        RECT 18.600 13.350 22.200 14.250 ;
        RECT 21.300 10.650 22.200 13.350 ;
        RECT 5.100 9.900 8.550 10.200 ;
        RECT 5.100 8.100 11.550 9.900 ;
        RECT 21.300 9.750 23.400 10.650 ;
        RECT 17.850 8.850 23.400 9.750 ;
        RECT 17.850 8.100 19.650 8.850 ;
        RECT 0.900 2.250 2.700 8.100 ;
        RECT 5.100 2.250 6.900 8.100 ;
        RECT 11.700 2.250 13.500 5.100 ;
        RECT 14.700 3.000 16.500 8.100 ;
        RECT 17.700 3.900 19.500 8.100 ;
        RECT 20.700 3.000 22.500 7.500 ;
        RECT 14.700 2.250 22.500 3.000 ;
        RECT 24.300 2.250 26.100 5.100 ;
      LAYER metal2 ;
        RECT 6.450 15.750 8.550 17.850 ;
        RECT 6.900 10.200 7.950 15.750 ;
        RECT 6.450 8.100 8.550 10.200 ;
  END
END HAX1
MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 9.900 40.200 ;
        RECT 0.900 30.900 2.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 5.100 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 3.900 21.600 5.100 30.900 ;
        RECT 0.600 15.600 2.400 16.350 ;
        RECT 3.900 5.100 5.100 17.400 ;
        RECT 3.900 2.100 5.700 5.100 ;
  END
END INVX1
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 9.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.900 5.700 36.900 ;
        RECT 0.600 16.650 2.400 17.400 ;
        RECT 3.900 15.600 5.100 24.900 ;
        RECT 3.900 8.100 5.100 11.400 ;
        RECT 3.900 2.100 5.700 8.100 ;
  END
END INVX2
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 15.450 2.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 6.900 24.900 8.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT 6.900 1.200 8.700 8.100 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.900 5.700 36.900 ;
        RECT 4.200 21.600 5.550 24.900 ;
        RECT 4.200 17.400 5.400 21.600 ;
        RECT 0.600 13.650 2.400 14.400 ;
        RECT 4.200 8.100 5.550 17.400 ;
        RECT 3.900 2.100 5.700 8.100 ;
  END
END INVX4
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 12.450 11.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 18.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 6.900 24.900 8.700 37.800 ;
        RECT 12.900 24.900 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 8.100 ;
        RECT 6.900 1.200 8.700 8.100 ;
        RECT 12.900 1.200 14.700 8.100 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 24.000 5.700 36.900 ;
        RECT 9.900 24.900 11.700 36.900 ;
        RECT 9.900 24.000 11.100 24.900 ;
        RECT 3.900 23.100 11.100 24.000 ;
        RECT 3.600 18.600 5.400 19.350 ;
        RECT 9.900 15.600 11.100 23.100 ;
        RECT 9.900 10.200 11.100 11.400 ;
        RECT 3.900 9.000 11.100 10.200 ;
        RECT 3.900 8.100 5.100 9.000 ;
        RECT 9.900 8.100 11.100 9.000 ;
        RECT 3.900 2.100 5.700 8.100 ;
        RECT 9.900 2.100 11.700 8.100 ;
  END
END INVX8
MACRO LATCH
  CLASS CORE ;
  FOREIGN LATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.700 18.450 14.550 20.550 ;
        RECT 6.900 17.550 12.750 18.450 ;
      LAYER metal2 ;
        RECT 12.900 20.550 14.100 23.100 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 13.050 9.900 14.550 ;
        RECT 3.450 12.450 5.550 13.050 ;
        RECT 8.550 9.900 9.600 13.050 ;
      LAYER metal2 ;
        RECT 3.900 14.550 5.100 17.100 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.000 24.900 19.800 36.900 ;
        RECT 18.600 17.550 19.800 24.900 ;
        RECT 15.450 15.450 19.800 17.550 ;
        RECT 18.600 8.100 19.800 15.450 ;
        RECT 18.000 2.100 19.800 8.100 ;
      LAYER metal2 ;
        RECT 15.450 15.450 17.550 17.550 ;
        RECT 15.900 12.900 17.100 15.450 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 24.900 3.000 36.750 ;
        RECT 4.200 24.900 6.000 36.750 ;
        RECT 9.300 30.900 11.250 36.750 ;
        RECT 9.450 28.800 11.550 30.900 ;
        RECT 15.000 24.900 16.800 36.750 ;
        RECT 1.200 21.300 2.400 24.900 ;
        RECT 9.450 24.000 11.550 24.900 ;
        RECT 9.450 22.800 17.400 24.000 ;
        RECT 15.600 22.200 17.400 22.800 ;
        RECT 1.200 20.400 9.900 21.300 ;
        RECT 1.200 8.100 2.400 20.400 ;
        RECT 8.100 19.500 9.900 20.400 ;
        RECT 1.200 2.250 3.000 8.100 ;
        RECT 9.450 5.100 11.550 7.200 ;
        RECT 4.200 2.250 6.000 5.100 ;
        RECT 9.300 2.250 11.400 5.100 ;
        RECT 15.000 2.250 16.800 8.100 ;
      LAYER metal2 ;
        RECT 9.450 28.800 11.550 30.900 ;
        RECT 9.600 24.900 10.800 28.800 ;
        RECT 9.450 22.800 11.550 24.900 ;
        RECT 9.600 7.200 10.800 22.800 ;
        RECT 9.450 5.100 11.550 7.200 ;
  END
END LATCH
MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 18.750 40.200 ;
        RECT 3.900 29.700 5.700 37.800 ;
        RECT 12.900 24.900 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 6.300 ;
        RECT 12.900 1.200 14.700 9.300 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 29.700 2.700 35.700 ;
        RECT 1.800 24.600 2.700 29.700 ;
        RECT 8.400 26.400 10.200 35.700 ;
        RECT 8.400 25.500 10.500 26.400 ;
        RECT 1.800 23.700 7.950 24.600 ;
        RECT 6.750 19.350 7.950 23.700 ;
        RECT 9.600 21.600 10.500 25.500 ;
        RECT 6.750 17.550 8.400 19.350 ;
        RECT 0.600 16.650 2.400 17.400 ;
        RECT 3.600 15.600 5.400 16.350 ;
        RECT 6.750 10.500 7.950 17.550 ;
        RECT 1.650 9.600 7.950 10.500 ;
        RECT 1.650 6.300 2.700 9.600 ;
        RECT 9.600 8.700 10.500 17.400 ;
        RECT 12.600 15.600 14.400 16.350 ;
        RECT 0.900 3.300 2.700 6.300 ;
        RECT 8.400 7.800 10.500 8.700 ;
        RECT 8.400 3.300 10.200 7.800 ;
  END
END MUX2X1
MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 21.450 2.550 23.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 21.450 8.550 23.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
        RECT 0.900 30.900 2.700 37.800 ;
        RECT 6.900 30.900 8.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.200 1.200 3.000 8.100 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 0.600 19.650 2.400 20.400 ;
        RECT 3.900 18.600 5.100 30.900 ;
        RECT 6.600 19.650 8.400 20.400 ;
        RECT 3.900 10.200 5.100 14.400 ;
        RECT 3.900 9.300 7.500 10.200 ;
        RECT 5.700 2.100 7.500 9.300 ;
  END
END NAND2X1
MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 24.450 2.550 26.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 21.450 11.550 23.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 0.900 30.900 2.700 37.800 ;
        RECT 6.900 31.500 8.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.200 1.200 3.000 11.100 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 3.900 30.900 5.700 36.900 ;
        RECT 4.200 30.600 5.700 30.900 ;
        RECT 9.900 30.900 11.700 36.900 ;
        RECT 9.900 30.600 10.800 30.900 ;
        RECT 4.200 29.700 10.800 30.600 ;
        RECT 9.900 24.600 10.800 29.700 ;
        RECT 0.600 22.650 2.400 23.400 ;
        RECT 3.600 21.600 5.400 22.350 ;
        RECT 6.600 13.650 8.400 14.400 ;
        RECT 9.900 12.150 10.800 20.400 ;
        RECT 6.600 10.500 10.800 12.150 ;
        RECT 6.600 2.100 8.400 10.500 ;
  END
END NAND3X1
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 9.450 5.550 11.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 5.100 ;
        RECT 6.900 1.200 8.700 5.100 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 5.100 24.900 6.900 36.900 ;
        RECT 4.200 23.850 6.900 24.900 ;
        RECT 0.600 21.600 2.400 22.350 ;
        RECT 4.200 18.600 5.550 23.850 ;
        RECT 6.600 18.600 8.400 19.350 ;
        RECT 4.200 14.400 5.400 18.600 ;
        RECT 4.200 12.600 5.550 14.400 ;
        RECT 3.900 5.100 5.100 8.400 ;
        RECT 3.900 2.100 5.700 5.100 ;
  END
END NOR2X1
MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 12.300 5.550 14.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.300 11.550 20.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 12.300 14.550 14.400 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.450 15.300 20.550 17.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 27.900 40.200 ;
        RECT 3.900 27.900 5.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 1.200 5.700 5.100 ;
        RECT 9.900 1.200 11.700 5.100 ;
        RECT -0.900 -1.200 27.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 27.000 2.700 36.900 ;
        RECT 6.900 36.000 14.700 36.900 ;
        RECT 6.900 27.000 8.700 36.000 ;
        RECT 0.900 26.100 8.700 27.000 ;
        RECT 9.900 27.300 11.700 35.100 ;
        RECT 12.900 28.200 14.700 36.000 ;
        RECT 16.500 36.000 24.300 36.900 ;
        RECT 16.500 27.300 18.300 36.000 ;
        RECT 9.900 26.400 18.300 27.300 ;
        RECT 19.500 27.300 21.300 35.100 ;
        RECT 19.500 24.900 20.700 27.300 ;
        RECT 22.500 26.700 24.300 36.000 ;
        RECT 17.250 23.700 20.700 24.900 ;
        RECT 17.250 18.450 18.450 23.700 ;
        RECT 9.600 16.500 11.400 17.250 ;
        RECT 3.600 15.450 5.400 16.200 ;
        RECT 12.600 15.450 14.400 16.200 ;
        RECT 17.250 14.250 17.400 18.450 ;
        RECT 17.250 6.900 18.450 14.250 ;
        RECT 7.650 6.000 18.450 6.900 ;
        RECT 7.650 5.100 8.700 6.000 ;
        RECT 13.650 5.100 14.700 6.000 ;
        RECT 6.900 2.100 8.700 5.100 ;
        RECT 12.900 2.100 14.700 5.100 ;
  END
END NOR3X1
MACRO OAI21X1
  CLASS CORE ;
  FOREIGN OAI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 1.800 24.900 3.600 37.800 ;
        RECT 9.300 30.900 11.100 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 6.300 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 6.000 24.900 7.800 36.900 ;
        RECT 6.450 21.600 7.650 24.900 ;
        RECT 6.600 17.400 7.650 21.600 ;
        RECT 3.600 16.650 5.400 17.400 ;
        RECT 0.600 15.600 2.400 16.350 ;
        RECT 6.450 15.600 7.650 17.400 ;
        RECT 9.600 16.650 11.400 17.400 ;
        RECT 7.350 11.250 8.550 11.400 ;
        RECT 7.350 10.200 11.100 11.250 ;
        RECT 0.900 7.200 8.700 8.550 ;
        RECT 0.900 2.100 2.700 7.200 ;
        RECT 6.900 2.100 8.700 7.200 ;
        RECT 9.900 8.100 11.100 10.200 ;
        RECT 9.900 2.100 11.700 8.100 ;
  END
END OAI21X1
MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 12.450 2.550 14.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 12.450 14.550 14.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 12.450 8.550 14.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 18.900 40.200 ;
        RECT 0.900 24.900 2.700 37.800 ;
        RECT 11.400 24.900 13.200 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 6.600 ;
        RECT -0.900 -1.200 18.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 5.400 24.900 8.700 36.900 ;
        RECT 3.600 16.650 5.400 17.400 ;
        RECT 6.900 15.600 8.100 24.900 ;
        RECT 9.000 16.650 10.800 17.400 ;
        RECT 12.450 15.600 14.250 16.350 ;
        RECT 0.750 10.650 2.550 11.400 ;
        RECT 6.900 10.800 8.100 11.400 ;
        RECT 6.900 9.600 11.100 10.800 ;
        RECT 0.900 7.500 8.700 8.400 ;
        RECT 10.200 8.100 11.100 9.600 ;
        RECT 0.900 2.100 2.700 7.500 ;
        RECT 6.900 3.000 8.700 7.500 ;
        RECT 9.900 3.900 11.700 8.100 ;
        RECT 12.900 3.000 14.700 8.100 ;
        RECT 6.900 2.100 14.700 3.000 ;
  END
END OAI22X1
MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 9.450 2.550 11.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 15.900 40.200 ;
        RECT 5.400 24.900 7.200 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 1.200 2.700 5.100 ;
        RECT 6.900 1.200 8.700 5.100 ;
        RECT -1.050 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 24.000 2.700 36.900 ;
        RECT 8.700 30.900 10.500 36.900 ;
        RECT 8.700 30.000 11.400 30.900 ;
        RECT 0.900 23.100 9.600 24.000 ;
        RECT 7.650 22.200 9.600 23.100 ;
        RECT 7.650 18.600 8.550 22.200 ;
        RECT 10.500 18.600 11.400 30.000 ;
        RECT 7.650 14.400 8.400 18.600 ;
        RECT 3.600 13.650 5.400 14.400 ;
        RECT 0.600 12.600 2.400 13.350 ;
        RECT 7.650 8.400 8.550 14.400 ;
        RECT 7.650 7.500 9.600 8.400 ;
        RECT 4.200 6.600 9.600 7.500 ;
        RECT 4.200 5.100 5.100 6.600 ;
        RECT 10.500 5.100 11.400 14.400 ;
        RECT 3.900 2.100 5.700 5.100 ;
        RECT 9.900 2.100 11.700 5.100 ;
  END
END OR2X1
MACRO OR2X2
  CLASS CORE ;
  FOREIGN OR2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 12.450 5.550 14.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
        RECT 5.400 24.900 7.200 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.900 2.100 2.700 5.100 ;
        RECT 0.900 1.200 2.100 2.100 ;
        RECT 6.900 1.200 8.700 5.100 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 24.900 2.700 36.900 ;
        RECT 8.400 26.400 10.200 36.900 ;
        RECT 8.400 24.900 10.800 26.400 ;
        RECT 0.900 23.700 2.100 24.900 ;
        RECT 0.900 22.500 8.100 23.700 ;
        RECT 6.300 21.900 8.100 22.500 ;
        RECT 0.600 16.650 2.400 17.400 ;
        RECT 3.600 15.600 5.400 16.350 ;
        RECT 7.200 11.100 8.100 21.900 ;
        RECT 9.450 18.600 10.800 24.900 ;
        RECT 6.450 10.200 8.250 11.100 ;
        RECT 4.800 9.300 8.250 10.200 ;
        RECT 4.800 5.100 5.700 9.300 ;
        RECT 10.500 8.100 11.550 14.400 ;
        RECT 3.900 2.100 5.700 5.100 ;
        RECT 9.900 2.100 11.700 8.100 ;
  END
END OR2X2
MACRO TBUFX1
  CLASS CORE ;
  FOREIGN TBUFX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.500 15.450 12.600 17.550 ;
      LAYER metal2 ;
        RECT 11.400 17.550 12.600 20.100 ;
        RECT 10.500 15.450 12.600 17.550 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.450 3.000 17.550 ;
      LAYER metal2 ;
        RECT 0.900 17.550 2.100 20.100 ;
        RECT 0.900 15.450 3.000 17.550 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.500 24.900 9.300 36.900 ;
        RECT 7.950 17.550 9.000 24.900 ;
        RECT 6.900 15.450 9.000 17.550 ;
        RECT 7.950 8.100 9.000 15.450 ;
        RECT 7.500 2.100 9.300 8.100 ;
      LAYER metal2 ;
        RECT 6.900 17.550 8.100 20.100 ;
        RECT 6.900 15.450 9.000 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 16.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 16.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 30.900 3.000 36.750 ;
        RECT 4.200 30.900 6.000 36.750 ;
        RECT 5.100 23.550 6.000 30.900 ;
        RECT 12.000 24.900 13.800 36.750 ;
        RECT 5.100 21.750 6.900 23.550 ;
        RECT 5.100 5.100 6.000 21.750 ;
        RECT 1.200 2.250 3.000 5.100 ;
        RECT 4.200 2.250 6.000 5.100 ;
        RECT 12.000 2.250 13.800 8.100 ;
  END
END TBUFX1
MACRO TBUFX2
  CLASS CORE ;
  FOREIGN TBUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.600 15.450 17.700 17.550 ;
      LAYER metal2 ;
        RECT 15.900 17.550 17.100 20.100 ;
        RECT 15.600 15.450 17.700 17.550 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.450 3.000 17.550 ;
      LAYER metal2 ;
        RECT 0.900 17.550 2.100 20.100 ;
        RECT 0.900 15.450 3.000 17.550 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.600 24.900 11.400 35.100 ;
        RECT 9.600 17.550 10.500 24.900 ;
        RECT 9.600 15.450 11.700 17.550 ;
        RECT 9.600 8.100 10.500 15.450 ;
        RECT 9.600 3.900 11.400 8.100 ;
      LAYER metal2 ;
        RECT 9.900 17.550 11.100 20.100 ;
        RECT 9.600 15.450 11.700 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 22.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 22.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 36.750 ;
        RECT 3.600 24.900 5.400 36.750 ;
        RECT 6.600 36.000 14.400 36.750 ;
        RECT 6.600 24.900 8.400 36.000 ;
        RECT 12.600 26.100 14.400 36.000 ;
        RECT 15.600 27.000 17.400 36.750 ;
        RECT 18.600 26.100 20.400 36.750 ;
        RECT 12.600 24.900 20.400 26.100 ;
        RECT 4.500 22.950 5.400 24.900 ;
        RECT 4.500 21.150 6.300 22.950 ;
        RECT 4.500 8.100 5.400 21.150 ;
        RECT 12.600 8.100 19.800 9.000 ;
        RECT 0.600 2.250 2.400 8.100 ;
        RECT 3.600 2.250 5.400 8.100 ;
        RECT 6.600 3.000 8.400 8.100 ;
        RECT 12.600 3.000 14.400 8.100 ;
        RECT 6.600 2.250 14.400 3.000 ;
        RECT 15.600 2.250 17.400 7.200 ;
        RECT 18.600 2.250 20.400 8.100 ;
  END
END TBUFX2
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.300 3.000 17.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.300 17.550 17.400 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.900 18.300 12.000 20.400 ;
    END
    PORT
      LAYER metal1 ;
        RECT 9.900 9.600 12.000 11.700 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.900 40.200 ;
        RECT 3.900 27.000 5.700 37.800 ;
        RECT 12.600 27.000 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 7.200 ;
        RECT 12.600 1.200 14.400 7.200 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.900 ;
        RECT 8.400 25.800 10.200 36.900 ;
        RECT 15.900 26.100 17.700 36.900 ;
        RECT 0.900 24.600 5.700 25.800 ;
        RECT 8.400 24.900 11.700 25.800 ;
        RECT 3.600 23.700 5.700 24.600 ;
        RECT 3.600 22.800 9.000 23.700 ;
        RECT 7.200 21.450 9.000 22.800 ;
        RECT 10.500 21.450 11.700 24.900 ;
        RECT 12.600 24.900 17.700 26.100 ;
        RECT 12.600 24.000 14.700 24.900 ;
        RECT 7.200 20.700 8.850 21.450 ;
        RECT 5.700 17.700 7.500 19.500 ;
        RECT 15.600 18.450 17.400 19.200 ;
        RECT 5.700 15.600 7.800 17.700 ;
        RECT 4.050 14.250 7.800 14.700 ;
        RECT 1.200 13.500 7.800 14.250 ;
        RECT 5.700 12.600 7.800 13.500 ;
        RECT 8.850 12.750 9.750 17.250 ;
        RECT 10.800 15.600 12.600 17.250 ;
        RECT 10.650 13.500 12.750 15.600 ;
        RECT 3.150 10.500 5.250 11.100 ;
        RECT 6.150 10.800 7.950 12.600 ;
        RECT 0.900 9.000 5.250 10.500 ;
        RECT 13.200 9.300 15.300 11.400 ;
        RECT 0.900 8.100 2.400 9.000 ;
        RECT 0.900 2.100 2.700 8.100 ;
        RECT 8.850 7.500 9.900 8.550 ;
        RECT 13.200 8.100 17.700 9.300 ;
        RECT 8.100 2.100 9.900 7.500 ;
        RECT 15.900 2.100 17.700 8.100 ;
      LAYER metal2 ;
        RECT 3.600 23.700 5.700 25.800 ;
        RECT 12.600 24.000 14.700 26.100 ;
        RECT 3.900 11.100 4.800 23.700 ;
        RECT 5.700 17.400 7.800 17.700 ;
        RECT 13.650 17.400 14.550 24.000 ;
        RECT 5.700 16.500 14.550 17.400 ;
        RECT 5.700 15.600 7.800 16.500 ;
        RECT 10.650 14.700 12.750 15.600 ;
        RECT 5.700 13.500 12.750 14.700 ;
        RECT 5.700 12.600 7.800 13.500 ;
        RECT 13.650 11.400 14.550 16.500 ;
        RECT 3.150 9.000 5.250 11.100 ;
        RECT 13.200 9.300 15.300 11.400 ;
  END
END XNOR2X1
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.900 15.450 3.000 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.450 17.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.600 18.300 11.700 20.400 ;
    END
    PORT
      LAYER metal1 ;
        RECT 9.600 9.600 11.700 11.700 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.750 40.200 ;
        RECT 3.900 27.000 5.700 37.800 ;
        RECT 12.900 27.000 14.700 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.900 1.200 5.700 7.200 ;
        RECT 12.900 1.200 14.700 7.200 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.900 25.800 2.700 36.900 ;
        RECT 0.900 24.900 5.400 25.800 ;
        RECT 8.400 24.900 10.200 36.900 ;
        RECT 15.900 26.100 17.700 36.900 ;
        RECT 3.300 22.800 5.400 24.900 ;
        RECT 9.000 23.400 10.200 24.900 ;
        RECT 12.900 24.900 17.700 26.100 ;
        RECT 12.900 24.000 15.000 24.900 ;
        RECT 9.000 22.500 10.500 23.400 ;
        RECT 9.600 21.450 10.500 22.500 ;
        RECT 6.600 21.000 8.550 21.300 ;
        RECT 4.800 19.200 8.550 21.000 ;
        RECT 15.600 18.600 17.400 19.350 ;
        RECT 6.000 17.400 7.800 18.000 ;
        RECT 4.050 16.200 7.800 17.400 ;
        RECT 0.900 13.650 2.700 14.400 ;
        RECT 6.000 12.900 7.800 14.700 ;
        RECT 5.700 10.800 7.800 12.900 ;
        RECT 8.700 12.750 9.750 17.250 ;
        RECT 11.100 14.700 12.900 16.500 ;
        RECT 10.650 12.750 12.750 14.700 ;
        RECT 1.500 9.900 7.800 10.800 ;
        RECT 1.500 8.100 2.700 9.900 ;
        RECT 12.900 9.000 15.000 10.200 ;
        RECT 8.700 8.100 9.900 8.550 ;
        RECT 12.900 8.100 17.700 9.000 ;
        RECT 0.900 2.100 2.700 8.100 ;
        RECT 8.400 2.100 10.200 8.100 ;
        RECT 15.900 2.100 17.700 8.100 ;
      LAYER metal2 ;
        RECT 3.300 22.800 5.400 24.900 ;
        RECT 12.900 24.000 15.000 26.100 ;
        RECT 4.200 13.800 5.100 22.800 ;
        RECT 6.600 19.200 8.700 21.300 ;
        RECT 7.800 16.800 8.700 19.200 ;
        RECT 13.500 16.800 14.550 24.000 ;
        RECT 7.800 15.600 14.550 16.800 ;
        RECT 10.650 13.800 12.750 14.700 ;
        RECT 4.200 12.600 12.750 13.800 ;
        RECT 5.700 10.800 7.800 12.600 ;
        RECT 13.650 10.200 14.550 15.600 ;
        RECT 12.900 8.100 15.000 10.200 ;
  END
END XOR2X1
END LIBRARY
