magic
tech scmos
magscale 1 3
timestamp 1555589239
<< checkpaint >>
rect -64 -64 64 64
<< gv1 >>
rect -4 -4 4 4
<< end >>
