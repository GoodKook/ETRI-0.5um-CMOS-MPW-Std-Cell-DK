magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 82 164
<< psubstratepdiff >>
rect 5 85 21 103
rect 5 79 10 85
rect 16 79 21 85
rect 5 57 21 79
rect 5 51 10 57
rect 16 51 21 57
rect 5 29 21 51
rect 5 23 10 29
rect 16 23 21 29
rect 5 5 21 23
<< psubstratepcontact >>
rect 10 79 16 85
rect 10 51 16 57
rect 10 23 16 29
<< genericcontact >>
rect 10 79 16 85
rect 10 51 16 57
rect 10 23 16 29
<< metal1 >>
rect 4 85 22 104
rect 4 79 10 85
rect 16 79 22 85
rect 4 57 22 79
rect 4 51 10 57
rect 16 51 22 57
rect 4 29 22 51
rect 4 23 10 29
rect 16 23 22 29
rect 4 4 22 23
<< end >>
