magic
tech scmos
magscale 1 2
timestamp 1702307383
<< nwell >>
rect -12 154 92 272
<< ntransistor >>
rect 24 14 28 54
rect 34 14 38 54
rect 54 14 58 34
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 34 54
rect 38 14 40 54
rect 52 14 54 34
rect 58 14 60 34
<< pdiffusion >>
rect 16 175 18 246
rect 4 166 18 175
rect 22 178 24 246
rect 36 178 38 246
rect 22 166 38 178
rect 42 166 44 246
rect 56 166 58 246
rect 62 166 64 246
<< ndcontact >>
rect 10 14 22 54
rect 40 14 52 54
rect 60 14 72 34
<< pdcontact >>
rect 4 175 16 246
rect 24 178 36 246
rect 44 166 56 246
rect 64 166 76 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 18 162 22 166
rect 38 162 42 166
rect 12 158 22 162
rect 30 158 42 162
rect 12 117 17 158
rect 12 60 17 105
rect 30 97 35 158
rect 58 117 62 166
rect 56 105 62 117
rect 30 75 37 85
rect 30 65 38 75
rect 12 56 28 60
rect 24 54 28 56
rect 34 54 38 65
rect 54 34 58 105
rect 24 10 28 14
rect 34 10 38 14
rect 54 10 58 14
<< polycontact >>
rect 5 105 17 117
rect 44 105 56 117
rect 25 85 37 97
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 24 246 36 252
rect 4 172 16 175
rect 4 166 44 172
rect 3 123 17 137
rect 43 123 57 137
rect 5 117 17 123
rect 44 117 56 123
rect 65 117 73 166
rect 23 103 37 117
rect 63 103 77 117
rect 25 97 37 103
rect 65 54 73 103
rect 52 47 73 54
rect 10 8 22 14
rect 60 8 72 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
<< labels >>
rlabel metal1 39 260 39 260 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 39 -1 39 -1 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 9 126 9 126 0 A
port 1 nsew signal input
rlabel metal1 29 105 29 105 0 B
port 2 nsew signal input
rlabel metal1 71 106 71 106 0 Y
port 4 nsew signal output
rlabel metal1 50 128 50 128 0 C
port 3 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
