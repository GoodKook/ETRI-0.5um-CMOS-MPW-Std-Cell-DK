//
// wozmon.v
//

module wozmon(clk, address, dout);
input           clk;
input  [7:0]    address;
output [7:0]    dout;

    reg [7:0]   dout;
    reg [7:0]   Memory[256];

// 1.4.2. Inferring ROM Functions from HDL Code
// Because small ROMs typically achieve the best performance when they are implemented
// using the registers in regular logic, each ROM function must meet a minimum size requirement
// for inference and placement in memory.
// https://www.intel.com/content/www/us/en/docs/programmable/683082/21-3/inferring-rom-functions-from-hdl-code.html

    always @(posedge clk)
    begin
		case (address)
            8'h00: dout <= 8'hD8;
            8'h01: dout <= 8'h58;
            8'h02: dout <= 8'hA0;
            8'h03: dout <= 8'h7F;
            8'h04: dout <= 8'h8C;
            8'h05: dout <= 8'h12;
            8'h06: dout <= 8'hD0;
            8'h07: dout <= 8'hA9;
            8'h08: dout <= 8'hA7;
            8'h09: dout <= 8'h8D;
            8'h0A: dout <= 8'h11;
            8'h0B: dout <= 8'hD0;
            8'h0C: dout <= 8'h8D;
            8'h0D: dout <= 8'h13;
            8'h0E: dout <= 8'hD0;
            8'h0F: dout <= 8'hC9;
            8'h10: dout <= 8'hDF;
            8'h11: dout <= 8'hF0;
            8'h12: dout <= 8'h13;
            8'h13: dout <= 8'hC9;
            8'h14: dout <= 8'h9B;
            8'h15: dout <= 8'hF0;
            8'h16: dout <= 8'h03;
            8'h17: dout <= 8'hC8;
            8'h18: dout <= 8'h10;
            8'h19: dout <= 8'h0F;
            8'h1A: dout <= 8'hA9;
            8'h1B: dout <= 8'hDC;
            8'h1C: dout <= 8'h20;
            8'h1D: dout <= 8'hEF;
            8'h1E: dout <= 8'hFF;
            8'h1F: dout <= 8'hA9;
            8'h20: dout <= 8'h8D;
            8'h21: dout <= 8'h20;
            8'h22: dout <= 8'hEF;
            8'h23: dout <= 8'hFF;
            8'h24: dout <= 8'hA0;
            8'h25: dout <= 8'h01;
            8'h26: dout <= 8'h88;
            8'h27: dout <= 8'h30;
            8'h28: dout <= 8'hF6;
            8'h29: dout <= 8'hAD;
            8'h2A: dout <= 8'h11;
            8'h2B: dout <= 8'hD0;
            8'h2C: dout <= 8'h10;
            8'h2D: dout <= 8'hFB;
            8'h2E: dout <= 8'hAD;
            8'h2F: dout <= 8'h10;
            8'h30: dout <= 8'hD0;
            8'h31: dout <= 8'h99;
            8'h32: dout <= 8'h00;
            8'h33: dout <= 8'h02;
            8'h34: dout <= 8'h20;
            8'h35: dout <= 8'hEF;
            8'h36: dout <= 8'hFF;
            8'h37: dout <= 8'hC9;
            8'h38: dout <= 8'h8D;
            8'h39: dout <= 8'hD0;
            8'h3A: dout <= 8'hD4;
            8'h3B: dout <= 8'hA0;
            8'h3C: dout <= 8'hFF;
            8'h3D: dout <= 8'hA9;
            8'h3E: dout <= 8'h00;
            8'h3F: dout <= 8'hAA;
            8'h40: dout <= 8'h0A;
            8'h41: dout <= 8'h85;
            8'h42: dout <= 8'h2B;
            8'h43: dout <= 8'hC8;
            8'h44: dout <= 8'hB9;
            8'h45: dout <= 8'h00;
            8'h46: dout <= 8'h02;
            8'h47: dout <= 8'hC9;
            8'h48: dout <= 8'h8D;
            8'h49: dout <= 8'hF0;
            8'h4A: dout <= 8'hD4;
            8'h4B: dout <= 8'hC9;
            8'h4C: dout <= 8'hAE;
            8'h4D: dout <= 8'h90;
            8'h4E: dout <= 8'hF4;
            8'h4F: dout <= 8'hF0;
            8'h50: dout <= 8'hF0;
            8'h51: dout <= 8'hC9;
            8'h52: dout <= 8'hBA;
            8'h53: dout <= 8'hF0;
            8'h54: dout <= 8'hEB;
            8'h55: dout <= 8'hC9;
            8'h56: dout <= 8'hD2;
            8'h57: dout <= 8'hF0;
            8'h58: dout <= 8'h3B;
            8'h59: dout <= 8'h86;
            8'h5A: dout <= 8'h28;
            8'h5B: dout <= 8'h86;
            8'h5C: dout <= 8'h29;
            8'h5D: dout <= 8'h84;
            8'h5E: dout <= 8'h2A;
            8'h5F: dout <= 8'hB9;
            8'h60: dout <= 8'h00;
            8'h61: dout <= 8'h02;
            8'h62: dout <= 8'h49;
            8'h63: dout <= 8'hB0;
            8'h64: dout <= 8'hC9;
            8'h65: dout <= 8'h0A;
            8'h66: dout <= 8'h90;
            8'h67: dout <= 8'h06;
            8'h68: dout <= 8'h69;
            8'h69: dout <= 8'h88;
            8'h6A: dout <= 8'hC9;
            8'h6B: dout <= 8'hFA;
            8'h6C: dout <= 8'h90;
            8'h6D: dout <= 8'h11;
            8'h6E: dout <= 8'h0A;
            8'h6F: dout <= 8'h0A;
            8'h70: dout <= 8'h0A;
            8'h71: dout <= 8'h0A;
            8'h72: dout <= 8'hA2;
            8'h73: dout <= 8'h04;
            8'h74: dout <= 8'h0A;
            8'h75: dout <= 8'h26;
            8'h76: dout <= 8'h28;
            8'h77: dout <= 8'h26;
            8'h78: dout <= 8'h29;
            8'h79: dout <= 8'hCA;
            8'h7A: dout <= 8'hD0;
            8'h7B: dout <= 8'hF8;
            8'h7C: dout <= 8'hC8;
            8'h7D: dout <= 8'hD0;
            8'h7E: dout <= 8'hE0;
            8'h7F: dout <= 8'hC4;
            8'h80: dout <= 8'h2A;
            8'h81: dout <= 8'hF0;
            8'h82: dout <= 8'h97;
            8'h83: dout <= 8'h24;
            8'h84: dout <= 8'h2B;
            8'h85: dout <= 8'h50;
            8'h86: dout <= 8'h10;
            8'h87: dout <= 8'hA5;
            8'h88: dout <= 8'h28;
            8'h89: dout <= 8'h81;
            8'h8A: dout <= 8'h26;
            8'h8B: dout <= 8'hE6;
            8'h8C: dout <= 8'h26;
            8'h8D: dout <= 8'hD0;
            8'h8E: dout <= 8'hB5;
            8'h8F: dout <= 8'hE6;
            8'h90: dout <= 8'h27;
            8'h91: dout <= 8'h4C;
            8'h92: dout <= 8'h44;
            8'h93: dout <= 8'hFF;
            8'h94: dout <= 8'h6C;
            8'h95: dout <= 8'h24;
            8'h96: dout <= 8'h00;
            8'h97: dout <= 8'h30;
            8'h98: dout <= 8'h2B;
            8'h99: dout <= 8'hA2;
            8'h9A: dout <= 8'h02;
            8'h9B: dout <= 8'hB5;
            8'h9C: dout <= 8'h27;
            8'h9D: dout <= 8'h95;
            8'h9E: dout <= 8'h25;
            8'h9F: dout <= 8'h95;
            8'hA0: dout <= 8'h23;
            8'hA1: dout <= 8'hCA;
            8'hA2: dout <= 8'hD0;
            8'hA3: dout <= 8'hF7;
            8'hA4: dout <= 8'hD0;
            8'hA5: dout <= 8'h14;
            8'hA6: dout <= 8'hA9;
            8'hA7: dout <= 8'h8D;
            8'hA8: dout <= 8'h20;
            8'hA9: dout <= 8'hEF;
            8'hAA: dout <= 8'hFF;
            8'hAB: dout <= 8'hA5;
            8'hAC: dout <= 8'h25;
            8'hAD: dout <= 8'h20;
            8'hAE: dout <= 8'hDC;
            8'hAF: dout <= 8'hFF;
            8'hB0: dout <= 8'hA5;
            8'hB1: dout <= 8'h24;
            8'hB2: dout <= 8'h20;
            8'hB3: dout <= 8'hDC;
            8'hB4: dout <= 8'hFF;
            8'hB5: dout <= 8'hA9;
            8'hB6: dout <= 8'hBA;
            8'hB7: dout <= 8'h20;
            8'hB8: dout <= 8'hEF;
            8'hB9: dout <= 8'hFF;
            8'hBA: dout <= 8'hA9;
            8'hBB: dout <= 8'hA0;
            8'hBC: dout <= 8'h20;
            8'hBD: dout <= 8'hEF;
            8'hBE: dout <= 8'hFF;
            8'hBF: dout <= 8'hA1;
            8'hC0: dout <= 8'h24;
            8'hC1: dout <= 8'h20;
            8'hC2: dout <= 8'hDC;
            8'hC3: dout <= 8'hFF;
            8'hC4: dout <= 8'h86;
            8'hC5: dout <= 8'h2B;
            8'hC6: dout <= 8'hA5;
            8'hC7: dout <= 8'h24;
            8'hC8: dout <= 8'hC5;
            8'hC9: dout <= 8'h28;
            8'hCA: dout <= 8'hA5;
            8'hCB: dout <= 8'h25;
            8'hCC: dout <= 8'hE5;
            8'hCD: dout <= 8'h29;
            8'hCE: dout <= 8'hB0;
            8'hCF: dout <= 8'hC1;
            8'hD0: dout <= 8'hE6;
            8'hD1: dout <= 8'h24;
            8'hD2: dout <= 8'hD0;
            8'hD3: dout <= 8'h02;
            8'hD4: dout <= 8'hE6;
            8'hD5: dout <= 8'h25;
            8'hD6: dout <= 8'hA5;
            8'hD7: dout <= 8'h24;
            8'hD8: dout <= 8'h29;
            8'hD9: dout <= 8'h07;
            8'hDA: dout <= 8'h10;
            8'hDB: dout <= 8'hC8;
            8'hDC: dout <= 8'h48;
            8'hDD: dout <= 8'h4A;
            8'hDE: dout <= 8'h4A;
            8'hDF: dout <= 8'h4A;
            8'hE0: dout <= 8'h4A;
            8'hE1: dout <= 8'h20;
            8'hE2: dout <= 8'hE5;
            8'hE3: dout <= 8'hFF;
            8'hE4: dout <= 8'h68;
            8'hE5: dout <= 8'h29;
            8'hE6: dout <= 8'h0F;
            8'hE7: dout <= 8'h09;
            8'hE8: dout <= 8'hB0;
            8'hE9: dout <= 8'hC9;
            8'hEA: dout <= 8'hBA;
            8'hEB: dout <= 8'h90;
            8'hEC: dout <= 8'h02;
            8'hED: dout <= 8'h69;
            8'hEE: dout <= 8'h06;
            8'hEF: dout <= 8'h2C;
            8'hF0: dout <= 8'h12;
            8'hF1: dout <= 8'hD0;
            8'hF2: dout <= 8'h30;
            8'hF3: dout <= 8'hFB;
            8'hF4: dout <= 8'h8D;
            8'hF5: dout <= 8'h12;
            8'hF6: dout <= 8'hD0;
            8'hF7: dout <= 8'h60;
            8'hF8: dout <= 8'h00;
            8'hF9: dout <= 8'h00;
            8'hFA: dout <= 8'h00;
            8'hFB: dout <= 8'h0F;
            8'hFC: dout <= 8'h00;
            8'hFD: dout <= 8'hFF;
            8'hFE: dout <= 8'h00;
            8'hFF: dout <= 8'h00;
        endcase
    end

 endmodule
