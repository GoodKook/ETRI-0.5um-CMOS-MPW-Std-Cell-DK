magic
tech scmos
magscale 1 6
timestamp 1727178812
<< checkpaint >>
rect 8700 8700 29300 29300
<< metal1 >>
rect 10220 29147 11560 29180
rect 10220 29129 10233 29147
rect 10251 29129 10269 29147
rect 10287 29129 10305 29147
rect 10323 29129 10341 29147
rect 10359 29129 10377 29147
rect 10395 29129 10413 29147
rect 10431 29129 10449 29147
rect 10467 29129 10485 29147
rect 10503 29129 10521 29147
rect 10539 29129 10557 29147
rect 10575 29129 10593 29147
rect 10611 29129 10629 29147
rect 10647 29129 10665 29147
rect 10683 29129 10701 29147
rect 10719 29129 10737 29147
rect 10755 29129 10773 29147
rect 10791 29129 10809 29147
rect 10827 29129 10845 29147
rect 10863 29129 10881 29147
rect 10899 29129 10917 29147
rect 10935 29129 10953 29147
rect 10971 29129 10989 29147
rect 11007 29129 11025 29147
rect 11043 29129 11061 29147
rect 11079 29129 11097 29147
rect 11115 29129 11133 29147
rect 11151 29129 11169 29147
rect 11187 29129 11205 29147
rect 11223 29129 11241 29147
rect 11259 29129 11277 29147
rect 11295 29129 11313 29147
rect 11331 29129 11349 29147
rect 11367 29129 11385 29147
rect 11403 29129 11421 29147
rect 11439 29129 11457 29147
rect 11475 29129 11493 29147
rect 11511 29129 11529 29147
rect 11547 29129 11560 29147
rect 10220 29111 11560 29129
rect 10220 29093 10233 29111
rect 10251 29093 10269 29111
rect 10287 29093 10305 29111
rect 10323 29093 10341 29111
rect 10359 29093 10377 29111
rect 10395 29093 10413 29111
rect 10431 29093 10449 29111
rect 10467 29093 10485 29111
rect 10503 29093 10521 29111
rect 10539 29093 10557 29111
rect 10575 29093 10593 29111
rect 10611 29093 10629 29111
rect 10647 29093 10665 29111
rect 10683 29093 10701 29111
rect 10719 29093 10737 29111
rect 10755 29093 10773 29111
rect 10791 29093 10809 29111
rect 10827 29093 10845 29111
rect 10863 29093 10881 29111
rect 10899 29093 10917 29111
rect 10935 29093 10953 29111
rect 10971 29093 10989 29111
rect 11007 29093 11025 29111
rect 11043 29093 11061 29111
rect 11079 29093 11097 29111
rect 11115 29093 11133 29111
rect 11151 29093 11169 29111
rect 11187 29093 11205 29111
rect 11223 29093 11241 29111
rect 11259 29093 11277 29111
rect 11295 29093 11313 29111
rect 11331 29093 11349 29111
rect 11367 29093 11385 29111
rect 11403 29093 11421 29111
rect 11439 29093 11457 29111
rect 11475 29093 11493 29111
rect 11511 29093 11529 29111
rect 11547 29093 11560 29111
rect 10220 29075 11560 29093
rect 10220 29057 10233 29075
rect 10251 29057 10269 29075
rect 10287 29057 10305 29075
rect 10323 29057 10341 29075
rect 10359 29057 10377 29075
rect 10395 29057 10413 29075
rect 10431 29057 10449 29075
rect 10467 29057 10485 29075
rect 10503 29057 10521 29075
rect 10539 29057 10557 29075
rect 10575 29057 10593 29075
rect 10611 29057 10629 29075
rect 10647 29057 10665 29075
rect 10683 29057 10701 29075
rect 10719 29057 10737 29075
rect 10755 29057 10773 29075
rect 10791 29057 10809 29075
rect 10827 29057 10845 29075
rect 10863 29057 10881 29075
rect 10899 29057 10917 29075
rect 10935 29057 10953 29075
rect 10971 29057 10989 29075
rect 11007 29057 11025 29075
rect 11043 29057 11061 29075
rect 11079 29057 11097 29075
rect 11115 29057 11133 29075
rect 11151 29057 11169 29075
rect 11187 29057 11205 29075
rect 11223 29057 11241 29075
rect 11259 29057 11277 29075
rect 11295 29057 11313 29075
rect 11331 29057 11349 29075
rect 11367 29057 11385 29075
rect 11403 29057 11421 29075
rect 11439 29057 11457 29075
rect 11475 29057 11493 29075
rect 11511 29057 11529 29075
rect 11547 29057 11560 29075
rect 10220 29039 11560 29057
rect 10220 29021 10233 29039
rect 10251 29021 10269 29039
rect 10287 29021 10305 29039
rect 10323 29021 10341 29039
rect 10359 29021 10377 29039
rect 10395 29021 10413 29039
rect 10431 29021 10449 29039
rect 10467 29021 10485 29039
rect 10503 29021 10521 29039
rect 10539 29021 10557 29039
rect 10575 29021 10593 29039
rect 10611 29021 10629 29039
rect 10647 29021 10665 29039
rect 10683 29021 10701 29039
rect 10719 29021 10737 29039
rect 10755 29021 10773 29039
rect 10791 29021 10809 29039
rect 10827 29021 10845 29039
rect 10863 29021 10881 29039
rect 10899 29021 10917 29039
rect 10935 29021 10953 29039
rect 10971 29021 10989 29039
rect 11007 29021 11025 29039
rect 11043 29021 11061 29039
rect 11079 29021 11097 29039
rect 11115 29021 11133 29039
rect 11151 29021 11169 29039
rect 11187 29021 11205 29039
rect 11223 29021 11241 29039
rect 11259 29021 11277 29039
rect 11295 29021 11313 29039
rect 11331 29021 11349 29039
rect 11367 29021 11385 29039
rect 11403 29021 11421 29039
rect 11439 29021 11457 29039
rect 11475 29021 11493 29039
rect 11511 29021 11529 29039
rect 11547 29021 11560 29039
rect 10220 29003 11560 29021
rect 10220 28985 10233 29003
rect 10251 28985 10269 29003
rect 10287 28985 10305 29003
rect 10323 28985 10341 29003
rect 10359 28985 10377 29003
rect 10395 28985 10413 29003
rect 10431 28985 10449 29003
rect 10467 28985 10485 29003
rect 10503 28985 10521 29003
rect 10539 28985 10557 29003
rect 10575 28985 10593 29003
rect 10611 28985 10629 29003
rect 10647 28985 10665 29003
rect 10683 28985 10701 29003
rect 10719 28985 10737 29003
rect 10755 28985 10773 29003
rect 10791 28985 10809 29003
rect 10827 28985 10845 29003
rect 10863 28985 10881 29003
rect 10899 28985 10917 29003
rect 10935 28985 10953 29003
rect 10971 28985 10989 29003
rect 11007 28985 11025 29003
rect 11043 28985 11061 29003
rect 11079 28985 11097 29003
rect 11115 28985 11133 29003
rect 11151 28985 11169 29003
rect 11187 28985 11205 29003
rect 11223 28985 11241 29003
rect 11259 28985 11277 29003
rect 11295 28985 11313 29003
rect 11331 28985 11349 29003
rect 11367 28985 11385 29003
rect 11403 28985 11421 29003
rect 11439 28985 11457 29003
rect 11475 28985 11493 29003
rect 11511 28985 11529 29003
rect 11547 28985 11560 29003
rect 10220 28967 11560 28985
rect 10220 28949 10233 28967
rect 10251 28949 10269 28967
rect 10287 28949 10305 28967
rect 10323 28949 10341 28967
rect 10359 28949 10377 28967
rect 10395 28949 10413 28967
rect 10431 28949 10449 28967
rect 10467 28949 10485 28967
rect 10503 28949 10521 28967
rect 10539 28949 10557 28967
rect 10575 28949 10593 28967
rect 10611 28949 10629 28967
rect 10647 28949 10665 28967
rect 10683 28949 10701 28967
rect 10719 28949 10737 28967
rect 10755 28949 10773 28967
rect 10791 28949 10809 28967
rect 10827 28949 10845 28967
rect 10863 28949 10881 28967
rect 10899 28949 10917 28967
rect 10935 28949 10953 28967
rect 10971 28949 10989 28967
rect 11007 28949 11025 28967
rect 11043 28949 11061 28967
rect 11079 28949 11097 28967
rect 11115 28949 11133 28967
rect 11151 28949 11169 28967
rect 11187 28949 11205 28967
rect 11223 28949 11241 28967
rect 11259 28949 11277 28967
rect 11295 28949 11313 28967
rect 11331 28949 11349 28967
rect 11367 28949 11385 28967
rect 11403 28949 11421 28967
rect 11439 28949 11457 28967
rect 11475 28949 11493 28967
rect 11511 28949 11529 28967
rect 11547 28949 11560 28967
rect 10220 28931 11560 28949
rect 10220 28913 10233 28931
rect 10251 28913 10269 28931
rect 10287 28913 10305 28931
rect 10323 28913 10341 28931
rect 10359 28913 10377 28931
rect 10395 28913 10413 28931
rect 10431 28913 10449 28931
rect 10467 28913 10485 28931
rect 10503 28913 10521 28931
rect 10539 28913 10557 28931
rect 10575 28913 10593 28931
rect 10611 28913 10629 28931
rect 10647 28913 10665 28931
rect 10683 28913 10701 28931
rect 10719 28913 10737 28931
rect 10755 28913 10773 28931
rect 10791 28913 10809 28931
rect 10827 28913 10845 28931
rect 10863 28913 10881 28931
rect 10899 28913 10917 28931
rect 10935 28913 10953 28931
rect 10971 28913 10989 28931
rect 11007 28913 11025 28931
rect 11043 28913 11061 28931
rect 11079 28913 11097 28931
rect 11115 28913 11133 28931
rect 11151 28913 11169 28931
rect 11187 28913 11205 28931
rect 11223 28913 11241 28931
rect 11259 28913 11277 28931
rect 11295 28913 11313 28931
rect 11331 28913 11349 28931
rect 11367 28913 11385 28931
rect 11403 28913 11421 28931
rect 11439 28913 11457 28931
rect 11475 28913 11493 28931
rect 11511 28913 11529 28931
rect 11547 28913 11560 28931
rect 10220 28900 11560 28913
rect 9700 28400 11560 28900
rect 28480 28011 29160 28040
rect 28480 27993 28941 28011
rect 28959 27993 28977 28011
rect 28995 27993 29013 28011
rect 29031 27993 29049 28011
rect 29067 27993 29085 28011
rect 29103 27993 29121 28011
rect 29139 27993 29160 28011
rect 28480 27975 29160 27993
rect 28480 27957 28941 27975
rect 28959 27957 28977 27975
rect 28995 27957 29013 27975
rect 29031 27957 29049 27975
rect 29067 27957 29085 27975
rect 29103 27957 29121 27975
rect 29139 27957 29160 27975
rect 28480 27939 29160 27957
rect 28480 27921 28941 27939
rect 28959 27921 28977 27939
rect 28995 27921 29013 27939
rect 29031 27921 29049 27939
rect 29067 27921 29085 27939
rect 29103 27921 29121 27939
rect 29139 27921 29160 27939
rect 28480 27903 29160 27921
rect 28480 27885 28941 27903
rect 28959 27885 28977 27903
rect 28995 27885 29013 27903
rect 29031 27885 29049 27903
rect 29067 27885 29085 27903
rect 29103 27885 29121 27903
rect 29139 27885 29160 27903
rect 28480 27867 29160 27885
rect 28480 27849 28941 27867
rect 28959 27849 28977 27867
rect 28995 27849 29013 27867
rect 29031 27849 29049 27867
rect 29067 27849 29085 27867
rect 29103 27849 29121 27867
rect 29139 27849 29160 27867
rect 28480 27831 29160 27849
rect 28480 27813 28941 27831
rect 28959 27813 28977 27831
rect 28995 27813 29013 27831
rect 29031 27813 29049 27831
rect 29067 27813 29085 27831
rect 29103 27813 29121 27831
rect 29139 27813 29160 27831
rect 28480 27795 29160 27813
rect 28480 27777 28941 27795
rect 28959 27777 28977 27795
rect 28995 27777 29013 27795
rect 29031 27777 29049 27795
rect 29067 27777 29085 27795
rect 29103 27777 29121 27795
rect 29139 27777 29160 27795
rect 28480 27759 29160 27777
rect 28480 27741 28941 27759
rect 28959 27741 28977 27759
rect 28995 27741 29013 27759
rect 29031 27741 29049 27759
rect 29067 27741 29085 27759
rect 29103 27741 29121 27759
rect 29139 27741 29160 27759
rect 28480 27723 29160 27741
rect 28480 27705 28941 27723
rect 28959 27705 28977 27723
rect 28995 27705 29013 27723
rect 29031 27705 29049 27723
rect 29067 27705 29085 27723
rect 29103 27705 29121 27723
rect 29139 27705 29160 27723
rect 28480 27687 29160 27705
rect 28480 27669 28941 27687
rect 28959 27669 28977 27687
rect 28995 27669 29013 27687
rect 29031 27669 29049 27687
rect 29067 27669 29085 27687
rect 29103 27669 29121 27687
rect 29139 27669 29160 27687
rect 28480 27651 29160 27669
rect 28480 27633 28941 27651
rect 28959 27633 28977 27651
rect 28995 27633 29013 27651
rect 29031 27633 29049 27651
rect 29067 27633 29085 27651
rect 29103 27633 29121 27651
rect 29139 27633 29160 27651
rect 28480 27615 29160 27633
rect 28480 27597 28941 27615
rect 28959 27597 28977 27615
rect 28995 27597 29013 27615
rect 29031 27597 29049 27615
rect 29067 27597 29085 27615
rect 29103 27597 29121 27615
rect 29139 27597 29160 27615
rect 28480 27579 29160 27597
rect 28480 27561 28941 27579
rect 28959 27561 28977 27579
rect 28995 27561 29013 27579
rect 29031 27561 29049 27579
rect 29067 27561 29085 27579
rect 29103 27561 29121 27579
rect 29139 27561 29160 27579
rect 28480 27543 29160 27561
rect 28480 27525 28941 27543
rect 28959 27525 28977 27543
rect 28995 27525 29013 27543
rect 29031 27525 29049 27543
rect 29067 27525 29085 27543
rect 29103 27525 29121 27543
rect 29139 27525 29160 27543
rect 28480 27507 29160 27525
rect 28480 27489 28941 27507
rect 28959 27489 28977 27507
rect 28995 27489 29013 27507
rect 29031 27489 29049 27507
rect 29067 27489 29085 27507
rect 29103 27489 29121 27507
rect 29139 27489 29160 27507
rect 28480 27471 29160 27489
rect 28480 27453 28941 27471
rect 28959 27453 28977 27471
rect 28995 27453 29013 27471
rect 29031 27453 29049 27471
rect 29067 27453 29085 27471
rect 29103 27453 29121 27471
rect 29139 27453 29160 27471
rect 28480 27435 29160 27453
rect 28480 27417 28941 27435
rect 28959 27417 28977 27435
rect 28995 27417 29013 27435
rect 29031 27417 29049 27435
rect 29067 27417 29085 27435
rect 29103 27417 29121 27435
rect 29139 27417 29160 27435
rect 28480 27399 29160 27417
rect 28480 27381 28941 27399
rect 28959 27381 28977 27399
rect 28995 27381 29013 27399
rect 29031 27381 29049 27399
rect 29067 27381 29085 27399
rect 29103 27381 29121 27399
rect 29139 27381 29160 27399
rect 28480 27363 29160 27381
rect 28480 27345 28941 27363
rect 28959 27345 28977 27363
rect 28995 27345 29013 27363
rect 29031 27345 29049 27363
rect 29067 27345 29085 27363
rect 29103 27345 29121 27363
rect 29139 27345 29160 27363
rect 28480 27327 29160 27345
rect 28480 27309 28941 27327
rect 28959 27309 28977 27327
rect 28995 27309 29013 27327
rect 29031 27309 29049 27327
rect 29067 27309 29085 27327
rect 29103 27309 29121 27327
rect 29139 27309 29160 27327
rect 28480 27291 29160 27309
rect 28480 27273 28941 27291
rect 28959 27273 28977 27291
rect 28995 27273 29013 27291
rect 29031 27273 29049 27291
rect 29067 27273 29085 27291
rect 29103 27273 29121 27291
rect 29139 27273 29160 27291
rect 28480 27255 29160 27273
rect 28480 27237 28941 27255
rect 28959 27237 28977 27255
rect 28995 27237 29013 27255
rect 29031 27237 29049 27255
rect 29067 27237 29085 27255
rect 29103 27237 29121 27255
rect 29139 27237 29160 27255
rect 28480 27219 29160 27237
rect 28480 27201 28941 27219
rect 28959 27201 28977 27219
rect 28995 27201 29013 27219
rect 29031 27201 29049 27219
rect 29067 27201 29085 27219
rect 29103 27201 29121 27219
rect 29139 27201 29160 27219
rect 28480 27183 29160 27201
rect 28480 27165 28941 27183
rect 28959 27165 28977 27183
rect 28995 27165 29013 27183
rect 29031 27165 29049 27183
rect 29067 27165 29085 27183
rect 29103 27165 29121 27183
rect 29139 27165 29160 27183
rect 28480 27147 29160 27165
rect 28480 27129 28941 27147
rect 28959 27129 28977 27147
rect 28995 27129 29013 27147
rect 29031 27129 29049 27147
rect 29067 27129 29085 27147
rect 29103 27129 29121 27147
rect 29139 27129 29160 27147
rect 28480 27111 29160 27129
rect 28480 27093 28941 27111
rect 28959 27093 28977 27111
rect 28995 27093 29013 27111
rect 29031 27093 29049 27111
rect 29067 27093 29085 27111
rect 29103 27093 29121 27111
rect 29139 27093 29160 27111
rect 28480 27075 29160 27093
rect 28480 27057 28941 27075
rect 28959 27057 28977 27075
rect 28995 27057 29013 27075
rect 29031 27057 29049 27075
rect 29067 27057 29085 27075
rect 29103 27057 29121 27075
rect 29139 27057 29160 27075
rect 28480 27039 29160 27057
rect 28480 27021 28941 27039
rect 28959 27021 28977 27039
rect 28995 27021 29013 27039
rect 29031 27021 29049 27039
rect 29067 27021 29085 27039
rect 29103 27021 29121 27039
rect 29139 27021 29160 27039
rect 28480 27003 29160 27021
rect 28480 26985 28941 27003
rect 28959 26985 28977 27003
rect 28995 26985 29013 27003
rect 29031 26985 29049 27003
rect 29067 26985 29085 27003
rect 29103 26985 29121 27003
rect 29139 26985 29160 27003
rect 28480 26967 29160 26985
rect 28480 26949 28941 26967
rect 28959 26949 28977 26967
rect 28995 26949 29013 26967
rect 29031 26949 29049 26967
rect 29067 26949 29085 26967
rect 29103 26949 29121 26967
rect 29139 26949 29160 26967
rect 28480 26931 29160 26949
rect 28480 26913 28941 26931
rect 28959 26913 28977 26931
rect 28995 26913 29013 26931
rect 29031 26913 29049 26931
rect 29067 26913 29085 26931
rect 29103 26913 29121 26931
rect 29139 26913 29160 26931
rect 28480 26895 29160 26913
rect 28480 26877 28941 26895
rect 28959 26877 28977 26895
rect 28995 26877 29013 26895
rect 29031 26877 29049 26895
rect 29067 26877 29085 26895
rect 29103 26877 29121 26895
rect 29139 26877 29160 26895
rect 28480 26859 29160 26877
rect 28480 26841 28941 26859
rect 28959 26841 28977 26859
rect 28995 26841 29013 26859
rect 29031 26841 29049 26859
rect 29067 26841 29085 26859
rect 29103 26841 29121 26859
rect 29139 26841 29160 26859
rect 28480 26823 29160 26841
rect 28480 26805 28941 26823
rect 28959 26805 28977 26823
rect 28995 26805 29013 26823
rect 29031 26805 29049 26823
rect 29067 26805 29085 26823
rect 29103 26805 29121 26823
rect 29139 26805 29160 26823
rect 28480 26787 29160 26805
rect 28480 26769 28941 26787
rect 28959 26769 28977 26787
rect 28995 26769 29013 26787
rect 29031 26769 29049 26787
rect 29067 26769 29085 26787
rect 29103 26769 29121 26787
rect 29139 26769 29160 26787
rect 28480 26751 29160 26769
rect 28480 26733 28941 26751
rect 28959 26733 28977 26751
rect 28995 26733 29013 26751
rect 29031 26733 29049 26751
rect 29067 26733 29085 26751
rect 29103 26733 29121 26751
rect 29139 26733 29160 26751
rect 28480 26715 29160 26733
rect 28480 26697 28941 26715
rect 28959 26697 28977 26715
rect 28995 26697 29013 26715
rect 29031 26697 29049 26715
rect 29067 26697 29085 26715
rect 29103 26697 29121 26715
rect 29139 26697 29160 26715
rect 28480 26679 29160 26697
rect 28480 26661 28941 26679
rect 28959 26661 28977 26679
rect 28995 26661 29013 26679
rect 29031 26661 29049 26679
rect 29067 26661 29085 26679
rect 29103 26661 29121 26679
rect 29139 26661 29160 26679
rect 28480 26643 29160 26661
rect 28480 26625 28941 26643
rect 28959 26625 28977 26643
rect 28995 26625 29013 26643
rect 29031 26625 29049 26643
rect 29067 26625 29085 26643
rect 29103 26625 29121 26643
rect 29139 26625 29160 26643
rect 28480 26607 29160 26625
rect 28480 26589 28941 26607
rect 28959 26589 28977 26607
rect 28995 26589 29013 26607
rect 29031 26589 29049 26607
rect 29067 26589 29085 26607
rect 29103 26589 29121 26607
rect 29139 26589 29160 26607
rect 28480 26571 29160 26589
rect 28480 26553 28941 26571
rect 28959 26553 28977 26571
rect 28995 26553 29013 26571
rect 29031 26553 29049 26571
rect 29067 26553 29085 26571
rect 29103 26553 29121 26571
rect 29139 26553 29160 26571
rect 28480 26535 29160 26553
rect 28480 26517 28941 26535
rect 28959 26517 28977 26535
rect 28995 26517 29013 26535
rect 29031 26517 29049 26535
rect 29067 26517 29085 26535
rect 29103 26517 29121 26535
rect 29139 26517 29160 26535
rect 28480 26499 29160 26517
rect 28480 26481 28941 26499
rect 28959 26481 28977 26499
rect 28995 26481 29013 26499
rect 29031 26481 29049 26499
rect 29067 26481 29085 26499
rect 29103 26481 29121 26499
rect 29139 26481 29160 26499
rect 28480 26463 29160 26481
rect 28480 26445 28941 26463
rect 28959 26445 28977 26463
rect 28995 26445 29013 26463
rect 29031 26445 29049 26463
rect 29067 26445 29085 26463
rect 29103 26445 29121 26463
rect 29139 26445 29160 26463
rect 28480 26427 29160 26445
rect 28480 26409 28941 26427
rect 28959 26409 28977 26427
rect 28995 26409 29013 26427
rect 29031 26409 29049 26427
rect 29067 26409 29085 26427
rect 29103 26409 29121 26427
rect 29139 26409 29160 26427
rect 28480 26380 29160 26409
rect 8960 25999 9500 26020
rect 8960 25981 8987 25999
rect 9005 25981 9023 25999
rect 9041 25981 9059 25999
rect 9077 25981 9095 25999
rect 9113 25981 9131 25999
rect 9149 25981 9167 25999
rect 9185 25981 9203 25999
rect 9221 25981 9239 25999
rect 9257 25981 9275 25999
rect 9293 25981 9311 25999
rect 9329 25981 9347 25999
rect 9365 25981 9383 25999
rect 9401 25981 9419 25999
rect 9437 25981 9455 25999
rect 9473 25981 9500 25999
rect 8960 25920 9500 25981
rect 9060 25763 9140 25780
rect 9060 25745 9081 25763
rect 9099 25745 9140 25763
rect 9060 25727 9140 25745
rect 9060 25709 9081 25727
rect 9099 25709 9140 25727
rect 9060 25691 9140 25709
rect 9060 25673 9081 25691
rect 9099 25673 9140 25691
rect 9060 25655 9140 25673
rect 9060 25637 9081 25655
rect 9099 25637 9140 25655
rect 9060 25619 9140 25637
rect 9060 25601 9081 25619
rect 9099 25601 9140 25619
rect 9060 25583 9140 25601
rect 9060 25565 9081 25583
rect 9099 25565 9140 25583
rect 9060 25547 9140 25565
rect 9060 25529 9081 25547
rect 9099 25529 9140 25547
rect 9060 25511 9140 25529
rect 9060 25493 9081 25511
rect 9099 25493 9140 25511
rect 9280 25643 9340 25660
rect 9280 25625 9301 25643
rect 9319 25625 9340 25643
rect 9280 25607 9340 25625
rect 9280 25589 9301 25607
rect 9319 25589 9340 25607
rect 9280 25571 9340 25589
rect 9280 25553 9301 25571
rect 9319 25553 9340 25571
rect 9280 25535 9340 25553
rect 9280 25517 9301 25535
rect 9319 25517 9340 25535
rect 9280 25500 9340 25517
rect 9060 25475 9140 25493
rect 9060 25457 9081 25475
rect 9099 25457 9140 25475
rect 9060 25440 9140 25457
rect 8820 11539 9740 11560
rect 8820 11521 8861 11539
rect 8879 11521 8897 11539
rect 8915 11521 8933 11539
rect 8951 11521 8969 11539
rect 8987 11521 9005 11539
rect 9023 11521 9041 11539
rect 9059 11521 9740 11539
rect 8820 11503 9740 11521
rect 8820 11485 8861 11503
rect 8879 11485 8897 11503
rect 8915 11485 8933 11503
rect 8951 11485 8969 11503
rect 8987 11485 9005 11503
rect 9023 11485 9041 11503
rect 9059 11485 9740 11503
rect 8820 11467 9740 11485
rect 8820 11449 8861 11467
rect 8879 11449 8897 11467
rect 8915 11449 8933 11467
rect 8951 11449 8969 11467
rect 8987 11449 9005 11467
rect 9023 11449 9041 11467
rect 9059 11449 9740 11467
rect 8820 11431 9740 11449
rect 8820 11413 8861 11431
rect 8879 11413 8897 11431
rect 8915 11413 8933 11431
rect 8951 11413 8969 11431
rect 8987 11413 9005 11431
rect 9023 11413 9041 11431
rect 9059 11413 9740 11431
rect 8820 11395 9740 11413
rect 8820 11377 8861 11395
rect 8879 11377 8897 11395
rect 8915 11377 8933 11395
rect 8951 11377 8969 11395
rect 8987 11377 9005 11395
rect 9023 11377 9041 11395
rect 9059 11377 9740 11395
rect 8820 11359 9740 11377
rect 8820 11341 8861 11359
rect 8879 11341 8897 11359
rect 8915 11341 8933 11359
rect 8951 11341 8969 11359
rect 8987 11341 9005 11359
rect 9023 11341 9041 11359
rect 9059 11341 9740 11359
rect 8820 11323 9740 11341
rect 8820 11305 8861 11323
rect 8879 11305 8897 11323
rect 8915 11305 8933 11323
rect 8951 11305 8969 11323
rect 8987 11305 9005 11323
rect 9023 11305 9041 11323
rect 9059 11305 9740 11323
rect 8820 11287 9740 11305
rect 8820 11269 8861 11287
rect 8879 11269 8897 11287
rect 8915 11269 8933 11287
rect 8951 11269 8969 11287
rect 8987 11269 9005 11287
rect 9023 11269 9041 11287
rect 9059 11269 9740 11287
rect 8820 11251 9740 11269
rect 8820 11233 8861 11251
rect 8879 11233 8897 11251
rect 8915 11233 8933 11251
rect 8951 11233 8969 11251
rect 8987 11233 9005 11251
rect 9023 11233 9041 11251
rect 9059 11233 9740 11251
rect 8820 11215 9740 11233
rect 8820 11197 8861 11215
rect 8879 11197 8897 11215
rect 8915 11197 8933 11215
rect 8951 11197 8969 11215
rect 8987 11197 9005 11215
rect 9023 11197 9041 11215
rect 9059 11197 9740 11215
rect 8820 11179 9740 11197
rect 8820 11161 8861 11179
rect 8879 11161 8897 11179
rect 8915 11161 8933 11179
rect 8951 11161 8969 11179
rect 8987 11161 9005 11179
rect 9023 11161 9041 11179
rect 9059 11161 9740 11179
rect 8820 11143 9740 11161
rect 8820 11125 8861 11143
rect 8879 11125 8897 11143
rect 8915 11125 8933 11143
rect 8951 11125 8969 11143
rect 8987 11125 9005 11143
rect 9023 11125 9041 11143
rect 9059 11125 9740 11143
rect 8820 11107 9740 11125
rect 8820 11089 8861 11107
rect 8879 11089 8897 11107
rect 8915 11089 8933 11107
rect 8951 11089 8969 11107
rect 8987 11089 9005 11107
rect 9023 11089 9041 11107
rect 9059 11089 9740 11107
rect 8820 11071 9740 11089
rect 8820 11053 8861 11071
rect 8879 11053 8897 11071
rect 8915 11053 8933 11071
rect 8951 11053 8969 11071
rect 8987 11053 9005 11071
rect 9023 11053 9041 11071
rect 9059 11053 9740 11071
rect 8820 11035 9740 11053
rect 8820 11017 8861 11035
rect 8879 11017 8897 11035
rect 8915 11017 8933 11035
rect 8951 11017 8969 11035
rect 8987 11017 9005 11035
rect 9023 11017 9041 11035
rect 9059 11017 9740 11035
rect 8820 10999 9740 11017
rect 8820 10981 8861 10999
rect 8879 10981 8897 10999
rect 8915 10981 8933 10999
rect 8951 10981 8969 10999
rect 8987 10981 9005 10999
rect 9023 10981 9041 10999
rect 9059 10981 9740 10999
rect 8820 10963 9740 10981
rect 8820 10945 8861 10963
rect 8879 10945 8897 10963
rect 8915 10945 8933 10963
rect 8951 10945 8969 10963
rect 8987 10945 9005 10963
rect 9023 10945 9041 10963
rect 9059 10945 9740 10963
rect 8820 10927 9740 10945
rect 8820 10909 8861 10927
rect 8879 10909 8897 10927
rect 8915 10909 8933 10927
rect 8951 10909 8969 10927
rect 8987 10909 9005 10927
rect 9023 10909 9041 10927
rect 9059 10909 9740 10927
rect 8820 10891 9740 10909
rect 8820 10873 8861 10891
rect 8879 10873 8897 10891
rect 8915 10873 8933 10891
rect 8951 10873 8969 10891
rect 8987 10873 9005 10891
rect 9023 10873 9041 10891
rect 9059 10873 9740 10891
rect 8820 10855 9740 10873
rect 8820 10837 8861 10855
rect 8879 10837 8897 10855
rect 8915 10837 8933 10855
rect 8951 10837 8969 10855
rect 8987 10837 9005 10855
rect 9023 10837 9041 10855
rect 9059 10837 9740 10855
rect 8820 10819 9740 10837
rect 8820 10801 8861 10819
rect 8879 10801 8897 10819
rect 8915 10801 8933 10819
rect 8951 10801 8969 10819
rect 8987 10801 9005 10819
rect 9023 10801 9041 10819
rect 9059 10801 9740 10819
rect 8820 10783 9740 10801
rect 8820 10765 8861 10783
rect 8879 10765 8897 10783
rect 8915 10765 8933 10783
rect 8951 10765 8969 10783
rect 8987 10765 9005 10783
rect 9023 10765 9041 10783
rect 9059 10765 9740 10783
rect 8820 10747 9740 10765
rect 8820 10729 8861 10747
rect 8879 10729 8897 10747
rect 8915 10729 8933 10747
rect 8951 10729 8969 10747
rect 8987 10729 9005 10747
rect 9023 10729 9041 10747
rect 9059 10729 9740 10747
rect 8820 10711 9740 10729
rect 8820 10693 8861 10711
rect 8879 10693 8897 10711
rect 8915 10693 8933 10711
rect 8951 10693 8969 10711
rect 8987 10693 9005 10711
rect 9023 10693 9041 10711
rect 9059 10693 9740 10711
rect 8820 10675 9740 10693
rect 8820 10657 8861 10675
rect 8879 10657 8897 10675
rect 8915 10657 8933 10675
rect 8951 10657 8969 10675
rect 8987 10657 9005 10675
rect 9023 10657 9041 10675
rect 9059 10657 9740 10675
rect 8820 10639 9740 10657
rect 8820 10621 8861 10639
rect 8879 10621 8897 10639
rect 8915 10621 8933 10639
rect 8951 10621 8969 10639
rect 8987 10621 9005 10639
rect 9023 10621 9041 10639
rect 9059 10621 9740 10639
rect 8820 10603 9740 10621
rect 8820 10585 8861 10603
rect 8879 10585 8897 10603
rect 8915 10585 8933 10603
rect 8951 10585 8969 10603
rect 8987 10585 9005 10603
rect 9023 10585 9041 10603
rect 9059 10585 9740 10603
rect 8820 10567 9740 10585
rect 8820 10549 8861 10567
rect 8879 10549 8897 10567
rect 8915 10549 8933 10567
rect 8951 10549 8969 10567
rect 8987 10549 9005 10567
rect 9023 10549 9041 10567
rect 9059 10549 9740 10567
rect 8820 10531 9740 10549
rect 8820 10513 8861 10531
rect 8879 10513 8897 10531
rect 8915 10513 8933 10531
rect 8951 10513 8969 10531
rect 8987 10513 9005 10531
rect 9023 10513 9041 10531
rect 9059 10513 9740 10531
rect 8820 10495 9740 10513
rect 8820 10477 8861 10495
rect 8879 10477 8897 10495
rect 8915 10477 8933 10495
rect 8951 10477 8969 10495
rect 8987 10477 9005 10495
rect 9023 10477 9041 10495
rect 9059 10477 9740 10495
rect 8820 10459 9740 10477
rect 8820 10441 8861 10459
rect 8879 10441 8897 10459
rect 8915 10441 8933 10459
rect 8951 10441 8969 10459
rect 8987 10441 9005 10459
rect 9023 10441 9041 10459
rect 9059 10441 9740 10459
rect 8820 10423 9740 10441
rect 8820 10405 8861 10423
rect 8879 10405 8897 10423
rect 8915 10405 8933 10423
rect 8951 10405 8969 10423
rect 8987 10405 9005 10423
rect 9023 10405 9041 10423
rect 9059 10405 9740 10423
rect 8820 10387 9740 10405
rect 8820 10369 8861 10387
rect 8879 10369 8897 10387
rect 8915 10369 8933 10387
rect 8951 10369 8969 10387
rect 8987 10369 9005 10387
rect 9023 10369 9041 10387
rect 9059 10369 9740 10387
rect 8820 10351 9740 10369
rect 8820 10333 8861 10351
rect 8879 10333 8897 10351
rect 8915 10333 8933 10351
rect 8951 10333 8969 10351
rect 8987 10333 9005 10351
rect 9023 10333 9041 10351
rect 9059 10333 9740 10351
rect 8820 10315 9740 10333
rect 8820 10297 8861 10315
rect 8879 10297 8897 10315
rect 8915 10297 8933 10315
rect 8951 10297 8969 10315
rect 8987 10297 9005 10315
rect 9023 10297 9041 10315
rect 9059 10297 9740 10315
rect 8820 10279 9740 10297
rect 8820 10261 8861 10279
rect 8879 10261 8897 10279
rect 8915 10261 8933 10279
rect 8951 10261 8969 10279
rect 8987 10261 9005 10279
rect 9023 10261 9041 10279
rect 9059 10261 9740 10279
rect 8820 10240 9740 10261
<< m2contact >>
rect 10233 29129 10251 29147
rect 10269 29129 10287 29147
rect 10305 29129 10323 29147
rect 10341 29129 10359 29147
rect 10377 29129 10395 29147
rect 10413 29129 10431 29147
rect 10449 29129 10467 29147
rect 10485 29129 10503 29147
rect 10521 29129 10539 29147
rect 10557 29129 10575 29147
rect 10593 29129 10611 29147
rect 10629 29129 10647 29147
rect 10665 29129 10683 29147
rect 10701 29129 10719 29147
rect 10737 29129 10755 29147
rect 10773 29129 10791 29147
rect 10809 29129 10827 29147
rect 10845 29129 10863 29147
rect 10881 29129 10899 29147
rect 10917 29129 10935 29147
rect 10953 29129 10971 29147
rect 10989 29129 11007 29147
rect 11025 29129 11043 29147
rect 11061 29129 11079 29147
rect 11097 29129 11115 29147
rect 11133 29129 11151 29147
rect 11169 29129 11187 29147
rect 11205 29129 11223 29147
rect 11241 29129 11259 29147
rect 11277 29129 11295 29147
rect 11313 29129 11331 29147
rect 11349 29129 11367 29147
rect 11385 29129 11403 29147
rect 11421 29129 11439 29147
rect 11457 29129 11475 29147
rect 11493 29129 11511 29147
rect 11529 29129 11547 29147
rect 10233 29093 10251 29111
rect 10269 29093 10287 29111
rect 10305 29093 10323 29111
rect 10341 29093 10359 29111
rect 10377 29093 10395 29111
rect 10413 29093 10431 29111
rect 10449 29093 10467 29111
rect 10485 29093 10503 29111
rect 10521 29093 10539 29111
rect 10557 29093 10575 29111
rect 10593 29093 10611 29111
rect 10629 29093 10647 29111
rect 10665 29093 10683 29111
rect 10701 29093 10719 29111
rect 10737 29093 10755 29111
rect 10773 29093 10791 29111
rect 10809 29093 10827 29111
rect 10845 29093 10863 29111
rect 10881 29093 10899 29111
rect 10917 29093 10935 29111
rect 10953 29093 10971 29111
rect 10989 29093 11007 29111
rect 11025 29093 11043 29111
rect 11061 29093 11079 29111
rect 11097 29093 11115 29111
rect 11133 29093 11151 29111
rect 11169 29093 11187 29111
rect 11205 29093 11223 29111
rect 11241 29093 11259 29111
rect 11277 29093 11295 29111
rect 11313 29093 11331 29111
rect 11349 29093 11367 29111
rect 11385 29093 11403 29111
rect 11421 29093 11439 29111
rect 11457 29093 11475 29111
rect 11493 29093 11511 29111
rect 11529 29093 11547 29111
rect 10233 29057 10251 29075
rect 10269 29057 10287 29075
rect 10305 29057 10323 29075
rect 10341 29057 10359 29075
rect 10377 29057 10395 29075
rect 10413 29057 10431 29075
rect 10449 29057 10467 29075
rect 10485 29057 10503 29075
rect 10521 29057 10539 29075
rect 10557 29057 10575 29075
rect 10593 29057 10611 29075
rect 10629 29057 10647 29075
rect 10665 29057 10683 29075
rect 10701 29057 10719 29075
rect 10737 29057 10755 29075
rect 10773 29057 10791 29075
rect 10809 29057 10827 29075
rect 10845 29057 10863 29075
rect 10881 29057 10899 29075
rect 10917 29057 10935 29075
rect 10953 29057 10971 29075
rect 10989 29057 11007 29075
rect 11025 29057 11043 29075
rect 11061 29057 11079 29075
rect 11097 29057 11115 29075
rect 11133 29057 11151 29075
rect 11169 29057 11187 29075
rect 11205 29057 11223 29075
rect 11241 29057 11259 29075
rect 11277 29057 11295 29075
rect 11313 29057 11331 29075
rect 11349 29057 11367 29075
rect 11385 29057 11403 29075
rect 11421 29057 11439 29075
rect 11457 29057 11475 29075
rect 11493 29057 11511 29075
rect 11529 29057 11547 29075
rect 10233 29021 10251 29039
rect 10269 29021 10287 29039
rect 10305 29021 10323 29039
rect 10341 29021 10359 29039
rect 10377 29021 10395 29039
rect 10413 29021 10431 29039
rect 10449 29021 10467 29039
rect 10485 29021 10503 29039
rect 10521 29021 10539 29039
rect 10557 29021 10575 29039
rect 10593 29021 10611 29039
rect 10629 29021 10647 29039
rect 10665 29021 10683 29039
rect 10701 29021 10719 29039
rect 10737 29021 10755 29039
rect 10773 29021 10791 29039
rect 10809 29021 10827 29039
rect 10845 29021 10863 29039
rect 10881 29021 10899 29039
rect 10917 29021 10935 29039
rect 10953 29021 10971 29039
rect 10989 29021 11007 29039
rect 11025 29021 11043 29039
rect 11061 29021 11079 29039
rect 11097 29021 11115 29039
rect 11133 29021 11151 29039
rect 11169 29021 11187 29039
rect 11205 29021 11223 29039
rect 11241 29021 11259 29039
rect 11277 29021 11295 29039
rect 11313 29021 11331 29039
rect 11349 29021 11367 29039
rect 11385 29021 11403 29039
rect 11421 29021 11439 29039
rect 11457 29021 11475 29039
rect 11493 29021 11511 29039
rect 11529 29021 11547 29039
rect 10233 28985 10251 29003
rect 10269 28985 10287 29003
rect 10305 28985 10323 29003
rect 10341 28985 10359 29003
rect 10377 28985 10395 29003
rect 10413 28985 10431 29003
rect 10449 28985 10467 29003
rect 10485 28985 10503 29003
rect 10521 28985 10539 29003
rect 10557 28985 10575 29003
rect 10593 28985 10611 29003
rect 10629 28985 10647 29003
rect 10665 28985 10683 29003
rect 10701 28985 10719 29003
rect 10737 28985 10755 29003
rect 10773 28985 10791 29003
rect 10809 28985 10827 29003
rect 10845 28985 10863 29003
rect 10881 28985 10899 29003
rect 10917 28985 10935 29003
rect 10953 28985 10971 29003
rect 10989 28985 11007 29003
rect 11025 28985 11043 29003
rect 11061 28985 11079 29003
rect 11097 28985 11115 29003
rect 11133 28985 11151 29003
rect 11169 28985 11187 29003
rect 11205 28985 11223 29003
rect 11241 28985 11259 29003
rect 11277 28985 11295 29003
rect 11313 28985 11331 29003
rect 11349 28985 11367 29003
rect 11385 28985 11403 29003
rect 11421 28985 11439 29003
rect 11457 28985 11475 29003
rect 11493 28985 11511 29003
rect 11529 28985 11547 29003
rect 10233 28949 10251 28967
rect 10269 28949 10287 28967
rect 10305 28949 10323 28967
rect 10341 28949 10359 28967
rect 10377 28949 10395 28967
rect 10413 28949 10431 28967
rect 10449 28949 10467 28967
rect 10485 28949 10503 28967
rect 10521 28949 10539 28967
rect 10557 28949 10575 28967
rect 10593 28949 10611 28967
rect 10629 28949 10647 28967
rect 10665 28949 10683 28967
rect 10701 28949 10719 28967
rect 10737 28949 10755 28967
rect 10773 28949 10791 28967
rect 10809 28949 10827 28967
rect 10845 28949 10863 28967
rect 10881 28949 10899 28967
rect 10917 28949 10935 28967
rect 10953 28949 10971 28967
rect 10989 28949 11007 28967
rect 11025 28949 11043 28967
rect 11061 28949 11079 28967
rect 11097 28949 11115 28967
rect 11133 28949 11151 28967
rect 11169 28949 11187 28967
rect 11205 28949 11223 28967
rect 11241 28949 11259 28967
rect 11277 28949 11295 28967
rect 11313 28949 11331 28967
rect 11349 28949 11367 28967
rect 11385 28949 11403 28967
rect 11421 28949 11439 28967
rect 11457 28949 11475 28967
rect 11493 28949 11511 28967
rect 11529 28949 11547 28967
rect 10233 28913 10251 28931
rect 10269 28913 10287 28931
rect 10305 28913 10323 28931
rect 10341 28913 10359 28931
rect 10377 28913 10395 28931
rect 10413 28913 10431 28931
rect 10449 28913 10467 28931
rect 10485 28913 10503 28931
rect 10521 28913 10539 28931
rect 10557 28913 10575 28931
rect 10593 28913 10611 28931
rect 10629 28913 10647 28931
rect 10665 28913 10683 28931
rect 10701 28913 10719 28931
rect 10737 28913 10755 28931
rect 10773 28913 10791 28931
rect 10809 28913 10827 28931
rect 10845 28913 10863 28931
rect 10881 28913 10899 28931
rect 10917 28913 10935 28931
rect 10953 28913 10971 28931
rect 10989 28913 11007 28931
rect 11025 28913 11043 28931
rect 11061 28913 11079 28931
rect 11097 28913 11115 28931
rect 11133 28913 11151 28931
rect 11169 28913 11187 28931
rect 11205 28913 11223 28931
rect 11241 28913 11259 28931
rect 11277 28913 11295 28931
rect 11313 28913 11331 28931
rect 11349 28913 11367 28931
rect 11385 28913 11403 28931
rect 11421 28913 11439 28931
rect 11457 28913 11475 28931
rect 11493 28913 11511 28931
rect 11529 28913 11547 28931
rect 28941 27993 28959 28011
rect 28977 27993 28995 28011
rect 29013 27993 29031 28011
rect 29049 27993 29067 28011
rect 29085 27993 29103 28011
rect 29121 27993 29139 28011
rect 28941 27957 28959 27975
rect 28977 27957 28995 27975
rect 29013 27957 29031 27975
rect 29049 27957 29067 27975
rect 29085 27957 29103 27975
rect 29121 27957 29139 27975
rect 28941 27921 28959 27939
rect 28977 27921 28995 27939
rect 29013 27921 29031 27939
rect 29049 27921 29067 27939
rect 29085 27921 29103 27939
rect 29121 27921 29139 27939
rect 28941 27885 28959 27903
rect 28977 27885 28995 27903
rect 29013 27885 29031 27903
rect 29049 27885 29067 27903
rect 29085 27885 29103 27903
rect 29121 27885 29139 27903
rect 28941 27849 28959 27867
rect 28977 27849 28995 27867
rect 29013 27849 29031 27867
rect 29049 27849 29067 27867
rect 29085 27849 29103 27867
rect 29121 27849 29139 27867
rect 28941 27813 28959 27831
rect 28977 27813 28995 27831
rect 29013 27813 29031 27831
rect 29049 27813 29067 27831
rect 29085 27813 29103 27831
rect 29121 27813 29139 27831
rect 28941 27777 28959 27795
rect 28977 27777 28995 27795
rect 29013 27777 29031 27795
rect 29049 27777 29067 27795
rect 29085 27777 29103 27795
rect 29121 27777 29139 27795
rect 28941 27741 28959 27759
rect 28977 27741 28995 27759
rect 29013 27741 29031 27759
rect 29049 27741 29067 27759
rect 29085 27741 29103 27759
rect 29121 27741 29139 27759
rect 28941 27705 28959 27723
rect 28977 27705 28995 27723
rect 29013 27705 29031 27723
rect 29049 27705 29067 27723
rect 29085 27705 29103 27723
rect 29121 27705 29139 27723
rect 28941 27669 28959 27687
rect 28977 27669 28995 27687
rect 29013 27669 29031 27687
rect 29049 27669 29067 27687
rect 29085 27669 29103 27687
rect 29121 27669 29139 27687
rect 28941 27633 28959 27651
rect 28977 27633 28995 27651
rect 29013 27633 29031 27651
rect 29049 27633 29067 27651
rect 29085 27633 29103 27651
rect 29121 27633 29139 27651
rect 28941 27597 28959 27615
rect 28977 27597 28995 27615
rect 29013 27597 29031 27615
rect 29049 27597 29067 27615
rect 29085 27597 29103 27615
rect 29121 27597 29139 27615
rect 28941 27561 28959 27579
rect 28977 27561 28995 27579
rect 29013 27561 29031 27579
rect 29049 27561 29067 27579
rect 29085 27561 29103 27579
rect 29121 27561 29139 27579
rect 28941 27525 28959 27543
rect 28977 27525 28995 27543
rect 29013 27525 29031 27543
rect 29049 27525 29067 27543
rect 29085 27525 29103 27543
rect 29121 27525 29139 27543
rect 28941 27489 28959 27507
rect 28977 27489 28995 27507
rect 29013 27489 29031 27507
rect 29049 27489 29067 27507
rect 29085 27489 29103 27507
rect 29121 27489 29139 27507
rect 28941 27453 28959 27471
rect 28977 27453 28995 27471
rect 29013 27453 29031 27471
rect 29049 27453 29067 27471
rect 29085 27453 29103 27471
rect 29121 27453 29139 27471
rect 28941 27417 28959 27435
rect 28977 27417 28995 27435
rect 29013 27417 29031 27435
rect 29049 27417 29067 27435
rect 29085 27417 29103 27435
rect 29121 27417 29139 27435
rect 28941 27381 28959 27399
rect 28977 27381 28995 27399
rect 29013 27381 29031 27399
rect 29049 27381 29067 27399
rect 29085 27381 29103 27399
rect 29121 27381 29139 27399
rect 28941 27345 28959 27363
rect 28977 27345 28995 27363
rect 29013 27345 29031 27363
rect 29049 27345 29067 27363
rect 29085 27345 29103 27363
rect 29121 27345 29139 27363
rect 28941 27309 28959 27327
rect 28977 27309 28995 27327
rect 29013 27309 29031 27327
rect 29049 27309 29067 27327
rect 29085 27309 29103 27327
rect 29121 27309 29139 27327
rect 28941 27273 28959 27291
rect 28977 27273 28995 27291
rect 29013 27273 29031 27291
rect 29049 27273 29067 27291
rect 29085 27273 29103 27291
rect 29121 27273 29139 27291
rect 28941 27237 28959 27255
rect 28977 27237 28995 27255
rect 29013 27237 29031 27255
rect 29049 27237 29067 27255
rect 29085 27237 29103 27255
rect 29121 27237 29139 27255
rect 28941 27201 28959 27219
rect 28977 27201 28995 27219
rect 29013 27201 29031 27219
rect 29049 27201 29067 27219
rect 29085 27201 29103 27219
rect 29121 27201 29139 27219
rect 28941 27165 28959 27183
rect 28977 27165 28995 27183
rect 29013 27165 29031 27183
rect 29049 27165 29067 27183
rect 29085 27165 29103 27183
rect 29121 27165 29139 27183
rect 28941 27129 28959 27147
rect 28977 27129 28995 27147
rect 29013 27129 29031 27147
rect 29049 27129 29067 27147
rect 29085 27129 29103 27147
rect 29121 27129 29139 27147
rect 28941 27093 28959 27111
rect 28977 27093 28995 27111
rect 29013 27093 29031 27111
rect 29049 27093 29067 27111
rect 29085 27093 29103 27111
rect 29121 27093 29139 27111
rect 28941 27057 28959 27075
rect 28977 27057 28995 27075
rect 29013 27057 29031 27075
rect 29049 27057 29067 27075
rect 29085 27057 29103 27075
rect 29121 27057 29139 27075
rect 28941 27021 28959 27039
rect 28977 27021 28995 27039
rect 29013 27021 29031 27039
rect 29049 27021 29067 27039
rect 29085 27021 29103 27039
rect 29121 27021 29139 27039
rect 28941 26985 28959 27003
rect 28977 26985 28995 27003
rect 29013 26985 29031 27003
rect 29049 26985 29067 27003
rect 29085 26985 29103 27003
rect 29121 26985 29139 27003
rect 28941 26949 28959 26967
rect 28977 26949 28995 26967
rect 29013 26949 29031 26967
rect 29049 26949 29067 26967
rect 29085 26949 29103 26967
rect 29121 26949 29139 26967
rect 28941 26913 28959 26931
rect 28977 26913 28995 26931
rect 29013 26913 29031 26931
rect 29049 26913 29067 26931
rect 29085 26913 29103 26931
rect 29121 26913 29139 26931
rect 28941 26877 28959 26895
rect 28977 26877 28995 26895
rect 29013 26877 29031 26895
rect 29049 26877 29067 26895
rect 29085 26877 29103 26895
rect 29121 26877 29139 26895
rect 28941 26841 28959 26859
rect 28977 26841 28995 26859
rect 29013 26841 29031 26859
rect 29049 26841 29067 26859
rect 29085 26841 29103 26859
rect 29121 26841 29139 26859
rect 28941 26805 28959 26823
rect 28977 26805 28995 26823
rect 29013 26805 29031 26823
rect 29049 26805 29067 26823
rect 29085 26805 29103 26823
rect 29121 26805 29139 26823
rect 28941 26769 28959 26787
rect 28977 26769 28995 26787
rect 29013 26769 29031 26787
rect 29049 26769 29067 26787
rect 29085 26769 29103 26787
rect 29121 26769 29139 26787
rect 28941 26733 28959 26751
rect 28977 26733 28995 26751
rect 29013 26733 29031 26751
rect 29049 26733 29067 26751
rect 29085 26733 29103 26751
rect 29121 26733 29139 26751
rect 28941 26697 28959 26715
rect 28977 26697 28995 26715
rect 29013 26697 29031 26715
rect 29049 26697 29067 26715
rect 29085 26697 29103 26715
rect 29121 26697 29139 26715
rect 28941 26661 28959 26679
rect 28977 26661 28995 26679
rect 29013 26661 29031 26679
rect 29049 26661 29067 26679
rect 29085 26661 29103 26679
rect 29121 26661 29139 26679
rect 28941 26625 28959 26643
rect 28977 26625 28995 26643
rect 29013 26625 29031 26643
rect 29049 26625 29067 26643
rect 29085 26625 29103 26643
rect 29121 26625 29139 26643
rect 28941 26589 28959 26607
rect 28977 26589 28995 26607
rect 29013 26589 29031 26607
rect 29049 26589 29067 26607
rect 29085 26589 29103 26607
rect 29121 26589 29139 26607
rect 28941 26553 28959 26571
rect 28977 26553 28995 26571
rect 29013 26553 29031 26571
rect 29049 26553 29067 26571
rect 29085 26553 29103 26571
rect 29121 26553 29139 26571
rect 28941 26517 28959 26535
rect 28977 26517 28995 26535
rect 29013 26517 29031 26535
rect 29049 26517 29067 26535
rect 29085 26517 29103 26535
rect 29121 26517 29139 26535
rect 28941 26481 28959 26499
rect 28977 26481 28995 26499
rect 29013 26481 29031 26499
rect 29049 26481 29067 26499
rect 29085 26481 29103 26499
rect 29121 26481 29139 26499
rect 28941 26445 28959 26463
rect 28977 26445 28995 26463
rect 29013 26445 29031 26463
rect 29049 26445 29067 26463
rect 29085 26445 29103 26463
rect 29121 26445 29139 26463
rect 28941 26409 28959 26427
rect 28977 26409 28995 26427
rect 29013 26409 29031 26427
rect 29049 26409 29067 26427
rect 29085 26409 29103 26427
rect 29121 26409 29139 26427
rect 8987 25981 9005 25999
rect 9023 25981 9041 25999
rect 9059 25981 9077 25999
rect 9095 25981 9113 25999
rect 9131 25981 9149 25999
rect 9167 25981 9185 25999
rect 9203 25981 9221 25999
rect 9239 25981 9257 25999
rect 9275 25981 9293 25999
rect 9311 25981 9329 25999
rect 9347 25981 9365 25999
rect 9383 25981 9401 25999
rect 9419 25981 9437 25999
rect 9455 25981 9473 25999
rect 9081 25745 9099 25763
rect 9081 25709 9099 25727
rect 9081 25673 9099 25691
rect 9081 25637 9099 25655
rect 9081 25601 9099 25619
rect 9081 25565 9099 25583
rect 9081 25529 9099 25547
rect 9081 25493 9099 25511
rect 9301 25625 9319 25643
rect 9301 25589 9319 25607
rect 9301 25553 9319 25571
rect 9301 25517 9319 25535
rect 9081 25457 9099 25475
rect 8861 11521 8879 11539
rect 8897 11521 8915 11539
rect 8933 11521 8951 11539
rect 8969 11521 8987 11539
rect 9005 11521 9023 11539
rect 9041 11521 9059 11539
rect 8861 11485 8879 11503
rect 8897 11485 8915 11503
rect 8933 11485 8951 11503
rect 8969 11485 8987 11503
rect 9005 11485 9023 11503
rect 9041 11485 9059 11503
rect 8861 11449 8879 11467
rect 8897 11449 8915 11467
rect 8933 11449 8951 11467
rect 8969 11449 8987 11467
rect 9005 11449 9023 11467
rect 9041 11449 9059 11467
rect 8861 11413 8879 11431
rect 8897 11413 8915 11431
rect 8933 11413 8951 11431
rect 8969 11413 8987 11431
rect 9005 11413 9023 11431
rect 9041 11413 9059 11431
rect 8861 11377 8879 11395
rect 8897 11377 8915 11395
rect 8933 11377 8951 11395
rect 8969 11377 8987 11395
rect 9005 11377 9023 11395
rect 9041 11377 9059 11395
rect 8861 11341 8879 11359
rect 8897 11341 8915 11359
rect 8933 11341 8951 11359
rect 8969 11341 8987 11359
rect 9005 11341 9023 11359
rect 9041 11341 9059 11359
rect 8861 11305 8879 11323
rect 8897 11305 8915 11323
rect 8933 11305 8951 11323
rect 8969 11305 8987 11323
rect 9005 11305 9023 11323
rect 9041 11305 9059 11323
rect 8861 11269 8879 11287
rect 8897 11269 8915 11287
rect 8933 11269 8951 11287
rect 8969 11269 8987 11287
rect 9005 11269 9023 11287
rect 9041 11269 9059 11287
rect 8861 11233 8879 11251
rect 8897 11233 8915 11251
rect 8933 11233 8951 11251
rect 8969 11233 8987 11251
rect 9005 11233 9023 11251
rect 9041 11233 9059 11251
rect 8861 11197 8879 11215
rect 8897 11197 8915 11215
rect 8933 11197 8951 11215
rect 8969 11197 8987 11215
rect 9005 11197 9023 11215
rect 9041 11197 9059 11215
rect 8861 11161 8879 11179
rect 8897 11161 8915 11179
rect 8933 11161 8951 11179
rect 8969 11161 8987 11179
rect 9005 11161 9023 11179
rect 9041 11161 9059 11179
rect 8861 11125 8879 11143
rect 8897 11125 8915 11143
rect 8933 11125 8951 11143
rect 8969 11125 8987 11143
rect 9005 11125 9023 11143
rect 9041 11125 9059 11143
rect 8861 11089 8879 11107
rect 8897 11089 8915 11107
rect 8933 11089 8951 11107
rect 8969 11089 8987 11107
rect 9005 11089 9023 11107
rect 9041 11089 9059 11107
rect 8861 11053 8879 11071
rect 8897 11053 8915 11071
rect 8933 11053 8951 11071
rect 8969 11053 8987 11071
rect 9005 11053 9023 11071
rect 9041 11053 9059 11071
rect 8861 11017 8879 11035
rect 8897 11017 8915 11035
rect 8933 11017 8951 11035
rect 8969 11017 8987 11035
rect 9005 11017 9023 11035
rect 9041 11017 9059 11035
rect 8861 10981 8879 10999
rect 8897 10981 8915 10999
rect 8933 10981 8951 10999
rect 8969 10981 8987 10999
rect 9005 10981 9023 10999
rect 9041 10981 9059 10999
rect 8861 10945 8879 10963
rect 8897 10945 8915 10963
rect 8933 10945 8951 10963
rect 8969 10945 8987 10963
rect 9005 10945 9023 10963
rect 9041 10945 9059 10963
rect 8861 10909 8879 10927
rect 8897 10909 8915 10927
rect 8933 10909 8951 10927
rect 8969 10909 8987 10927
rect 9005 10909 9023 10927
rect 9041 10909 9059 10927
rect 8861 10873 8879 10891
rect 8897 10873 8915 10891
rect 8933 10873 8951 10891
rect 8969 10873 8987 10891
rect 9005 10873 9023 10891
rect 9041 10873 9059 10891
rect 8861 10837 8879 10855
rect 8897 10837 8915 10855
rect 8933 10837 8951 10855
rect 8969 10837 8987 10855
rect 9005 10837 9023 10855
rect 9041 10837 9059 10855
rect 8861 10801 8879 10819
rect 8897 10801 8915 10819
rect 8933 10801 8951 10819
rect 8969 10801 8987 10819
rect 9005 10801 9023 10819
rect 9041 10801 9059 10819
rect 8861 10765 8879 10783
rect 8897 10765 8915 10783
rect 8933 10765 8951 10783
rect 8969 10765 8987 10783
rect 9005 10765 9023 10783
rect 9041 10765 9059 10783
rect 8861 10729 8879 10747
rect 8897 10729 8915 10747
rect 8933 10729 8951 10747
rect 8969 10729 8987 10747
rect 9005 10729 9023 10747
rect 9041 10729 9059 10747
rect 8861 10693 8879 10711
rect 8897 10693 8915 10711
rect 8933 10693 8951 10711
rect 8969 10693 8987 10711
rect 9005 10693 9023 10711
rect 9041 10693 9059 10711
rect 8861 10657 8879 10675
rect 8897 10657 8915 10675
rect 8933 10657 8951 10675
rect 8969 10657 8987 10675
rect 9005 10657 9023 10675
rect 9041 10657 9059 10675
rect 8861 10621 8879 10639
rect 8897 10621 8915 10639
rect 8933 10621 8951 10639
rect 8969 10621 8987 10639
rect 9005 10621 9023 10639
rect 9041 10621 9059 10639
rect 8861 10585 8879 10603
rect 8897 10585 8915 10603
rect 8933 10585 8951 10603
rect 8969 10585 8987 10603
rect 9005 10585 9023 10603
rect 9041 10585 9059 10603
rect 8861 10549 8879 10567
rect 8897 10549 8915 10567
rect 8933 10549 8951 10567
rect 8969 10549 8987 10567
rect 9005 10549 9023 10567
rect 9041 10549 9059 10567
rect 8861 10513 8879 10531
rect 8897 10513 8915 10531
rect 8933 10513 8951 10531
rect 8969 10513 8987 10531
rect 9005 10513 9023 10531
rect 9041 10513 9059 10531
rect 8861 10477 8879 10495
rect 8897 10477 8915 10495
rect 8933 10477 8951 10495
rect 8969 10477 8987 10495
rect 9005 10477 9023 10495
rect 9041 10477 9059 10495
rect 8861 10441 8879 10459
rect 8897 10441 8915 10459
rect 8933 10441 8951 10459
rect 8969 10441 8987 10459
rect 9005 10441 9023 10459
rect 9041 10441 9059 10459
rect 8861 10405 8879 10423
rect 8897 10405 8915 10423
rect 8933 10405 8951 10423
rect 8969 10405 8987 10423
rect 9005 10405 9023 10423
rect 9041 10405 9059 10423
rect 8861 10369 8879 10387
rect 8897 10369 8915 10387
rect 8933 10369 8951 10387
rect 8969 10369 8987 10387
rect 9005 10369 9023 10387
rect 9041 10369 9059 10387
rect 8861 10333 8879 10351
rect 8897 10333 8915 10351
rect 8933 10333 8951 10351
rect 8969 10333 8987 10351
rect 9005 10333 9023 10351
rect 9041 10333 9059 10351
rect 8861 10297 8879 10315
rect 8897 10297 8915 10315
rect 8933 10297 8951 10315
rect 8969 10297 8987 10315
rect 9005 10297 9023 10315
rect 9041 10297 9059 10315
rect 8861 10261 8879 10279
rect 8897 10261 8915 10279
rect 8933 10261 8951 10279
rect 8969 10261 8987 10279
rect 9005 10261 9023 10279
rect 9041 10261 9059 10279
<< metal2 >>
rect 10220 29147 11560 29180
rect 10220 29129 10233 29147
rect 10251 29129 10269 29147
rect 10287 29129 10305 29147
rect 10323 29129 10341 29147
rect 10359 29129 10377 29147
rect 10395 29129 10413 29147
rect 10431 29129 10449 29147
rect 10467 29129 10485 29147
rect 10503 29129 10521 29147
rect 10539 29129 10557 29147
rect 10575 29129 10593 29147
rect 10611 29129 10629 29147
rect 10647 29129 10665 29147
rect 10683 29129 10701 29147
rect 10719 29129 10737 29147
rect 10755 29129 10773 29147
rect 10791 29129 10809 29147
rect 10827 29129 10845 29147
rect 10863 29129 10881 29147
rect 10899 29129 10917 29147
rect 10935 29129 10953 29147
rect 10971 29129 10989 29147
rect 11007 29129 11025 29147
rect 11043 29129 11061 29147
rect 11079 29129 11097 29147
rect 11115 29129 11133 29147
rect 11151 29129 11169 29147
rect 11187 29129 11205 29147
rect 11223 29129 11241 29147
rect 11259 29129 11277 29147
rect 11295 29129 11313 29147
rect 11331 29129 11349 29147
rect 11367 29129 11385 29147
rect 11403 29129 11421 29147
rect 11439 29129 11457 29147
rect 11475 29129 11493 29147
rect 11511 29129 11529 29147
rect 11547 29129 11560 29147
rect 10220 29111 11560 29129
rect 10220 29093 10233 29111
rect 10251 29093 10269 29111
rect 10287 29093 10305 29111
rect 10323 29093 10341 29111
rect 10359 29093 10377 29111
rect 10395 29093 10413 29111
rect 10431 29093 10449 29111
rect 10467 29093 10485 29111
rect 10503 29093 10521 29111
rect 10539 29093 10557 29111
rect 10575 29093 10593 29111
rect 10611 29093 10629 29111
rect 10647 29093 10665 29111
rect 10683 29093 10701 29111
rect 10719 29093 10737 29111
rect 10755 29093 10773 29111
rect 10791 29093 10809 29111
rect 10827 29093 10845 29111
rect 10863 29093 10881 29111
rect 10899 29093 10917 29111
rect 10935 29093 10953 29111
rect 10971 29093 10989 29111
rect 11007 29093 11025 29111
rect 11043 29093 11061 29111
rect 11079 29093 11097 29111
rect 11115 29093 11133 29111
rect 11151 29093 11169 29111
rect 11187 29093 11205 29111
rect 11223 29093 11241 29111
rect 11259 29093 11277 29111
rect 11295 29093 11313 29111
rect 11331 29093 11349 29111
rect 11367 29093 11385 29111
rect 11403 29093 11421 29111
rect 11439 29093 11457 29111
rect 11475 29093 11493 29111
rect 11511 29093 11529 29111
rect 11547 29093 11560 29111
rect 10220 29075 11560 29093
rect 10220 29057 10233 29075
rect 10251 29057 10269 29075
rect 10287 29057 10305 29075
rect 10323 29057 10341 29075
rect 10359 29057 10377 29075
rect 10395 29057 10413 29075
rect 10431 29057 10449 29075
rect 10467 29057 10485 29075
rect 10503 29057 10521 29075
rect 10539 29057 10557 29075
rect 10575 29057 10593 29075
rect 10611 29057 10629 29075
rect 10647 29057 10665 29075
rect 10683 29057 10701 29075
rect 10719 29057 10737 29075
rect 10755 29057 10773 29075
rect 10791 29057 10809 29075
rect 10827 29057 10845 29075
rect 10863 29057 10881 29075
rect 10899 29057 10917 29075
rect 10935 29057 10953 29075
rect 10971 29057 10989 29075
rect 11007 29057 11025 29075
rect 11043 29057 11061 29075
rect 11079 29057 11097 29075
rect 11115 29057 11133 29075
rect 11151 29057 11169 29075
rect 11187 29057 11205 29075
rect 11223 29057 11241 29075
rect 11259 29057 11277 29075
rect 11295 29057 11313 29075
rect 11331 29057 11349 29075
rect 11367 29057 11385 29075
rect 11403 29057 11421 29075
rect 11439 29057 11457 29075
rect 11475 29057 11493 29075
rect 11511 29057 11529 29075
rect 11547 29057 11560 29075
rect 10220 29039 11560 29057
rect 10220 29021 10233 29039
rect 10251 29021 10269 29039
rect 10287 29021 10305 29039
rect 10323 29021 10341 29039
rect 10359 29021 10377 29039
rect 10395 29021 10413 29039
rect 10431 29021 10449 29039
rect 10467 29021 10485 29039
rect 10503 29021 10521 29039
rect 10539 29021 10557 29039
rect 10575 29021 10593 29039
rect 10611 29021 10629 29039
rect 10647 29021 10665 29039
rect 10683 29021 10701 29039
rect 10719 29021 10737 29039
rect 10755 29021 10773 29039
rect 10791 29021 10809 29039
rect 10827 29021 10845 29039
rect 10863 29021 10881 29039
rect 10899 29021 10917 29039
rect 10935 29021 10953 29039
rect 10971 29021 10989 29039
rect 11007 29021 11025 29039
rect 11043 29021 11061 29039
rect 11079 29021 11097 29039
rect 11115 29021 11133 29039
rect 11151 29021 11169 29039
rect 11187 29021 11205 29039
rect 11223 29021 11241 29039
rect 11259 29021 11277 29039
rect 11295 29021 11313 29039
rect 11331 29021 11349 29039
rect 11367 29021 11385 29039
rect 11403 29021 11421 29039
rect 11439 29021 11457 29039
rect 11475 29021 11493 29039
rect 11511 29021 11529 29039
rect 11547 29021 11560 29039
rect 10220 29003 11560 29021
rect 10220 28985 10233 29003
rect 10251 28985 10269 29003
rect 10287 28985 10305 29003
rect 10323 28985 10341 29003
rect 10359 28985 10377 29003
rect 10395 28985 10413 29003
rect 10431 28985 10449 29003
rect 10467 28985 10485 29003
rect 10503 28985 10521 29003
rect 10539 28985 10557 29003
rect 10575 28985 10593 29003
rect 10611 28985 10629 29003
rect 10647 28985 10665 29003
rect 10683 28985 10701 29003
rect 10719 28985 10737 29003
rect 10755 28985 10773 29003
rect 10791 28985 10809 29003
rect 10827 28985 10845 29003
rect 10863 28985 10881 29003
rect 10899 28985 10917 29003
rect 10935 28985 10953 29003
rect 10971 28985 10989 29003
rect 11007 28985 11025 29003
rect 11043 28985 11061 29003
rect 11079 28985 11097 29003
rect 11115 28985 11133 29003
rect 11151 28985 11169 29003
rect 11187 28985 11205 29003
rect 11223 28985 11241 29003
rect 11259 28985 11277 29003
rect 11295 28985 11313 29003
rect 11331 28985 11349 29003
rect 11367 28985 11385 29003
rect 11403 28985 11421 29003
rect 11439 28985 11457 29003
rect 11475 28985 11493 29003
rect 11511 28985 11529 29003
rect 11547 28985 11560 29003
rect 10220 28967 11560 28985
rect 10220 28949 10233 28967
rect 10251 28949 10269 28967
rect 10287 28949 10305 28967
rect 10323 28949 10341 28967
rect 10359 28949 10377 28967
rect 10395 28949 10413 28967
rect 10431 28949 10449 28967
rect 10467 28949 10485 28967
rect 10503 28949 10521 28967
rect 10539 28949 10557 28967
rect 10575 28949 10593 28967
rect 10611 28949 10629 28967
rect 10647 28949 10665 28967
rect 10683 28949 10701 28967
rect 10719 28949 10737 28967
rect 10755 28949 10773 28967
rect 10791 28949 10809 28967
rect 10827 28949 10845 28967
rect 10863 28949 10881 28967
rect 10899 28949 10917 28967
rect 10935 28949 10953 28967
rect 10971 28949 10989 28967
rect 11007 28949 11025 28967
rect 11043 28949 11061 28967
rect 11079 28949 11097 28967
rect 11115 28949 11133 28967
rect 11151 28949 11169 28967
rect 11187 28949 11205 28967
rect 11223 28949 11241 28967
rect 11259 28949 11277 28967
rect 11295 28949 11313 28967
rect 11331 28949 11349 28967
rect 11367 28949 11385 28967
rect 11403 28949 11421 28967
rect 11439 28949 11457 28967
rect 11475 28949 11493 28967
rect 11511 28949 11529 28967
rect 11547 28949 11560 28967
rect 10220 28931 11560 28949
rect 10220 28913 10233 28931
rect 10251 28913 10269 28931
rect 10287 28913 10305 28931
rect 10323 28913 10341 28931
rect 10359 28913 10377 28931
rect 10395 28913 10413 28931
rect 10431 28913 10449 28931
rect 10467 28913 10485 28931
rect 10503 28913 10521 28931
rect 10539 28913 10557 28931
rect 10575 28913 10593 28931
rect 10611 28913 10629 28931
rect 10647 28913 10665 28931
rect 10683 28913 10701 28931
rect 10719 28913 10737 28931
rect 10755 28913 10773 28931
rect 10791 28913 10809 28931
rect 10827 28913 10845 28931
rect 10863 28913 10881 28931
rect 10899 28913 10917 28931
rect 10935 28913 10953 28931
rect 10971 28913 10989 28931
rect 11007 28913 11025 28931
rect 11043 28913 11061 28931
rect 11079 28913 11097 28931
rect 11115 28913 11133 28931
rect 11151 28913 11169 28931
rect 11187 28913 11205 28931
rect 11223 28913 11241 28931
rect 11259 28913 11277 28931
rect 11295 28913 11313 28931
rect 11331 28913 11349 28931
rect 11367 28913 11385 28931
rect 11403 28913 11421 28931
rect 11439 28913 11457 28931
rect 11475 28913 11493 28931
rect 11511 28913 11529 28931
rect 11547 28913 11560 28931
rect 10220 28900 11560 28913
rect 14660 28600 14740 29180
rect 17360 28720 17440 29180
rect 20060 28840 20140 29180
rect 22760 28960 22840 29180
rect 25460 29080 25540 29180
rect 28160 29080 28240 29180
rect 25460 29059 25620 29080
rect 25460 29041 25477 29059
rect 25495 29041 25513 29059
rect 25531 29041 25549 29059
rect 25567 29041 25585 29059
rect 25603 29041 25620 29059
rect 25460 29020 25620 29041
rect 27240 29059 27400 29080
rect 27240 29041 27257 29059
rect 27275 29041 27293 29059
rect 27311 29041 27329 29059
rect 27347 29041 27365 29059
rect 27383 29041 27400 29059
rect 27240 29020 27400 29041
rect 22760 28939 22940 28960
rect 22760 28921 22787 28939
rect 22805 28921 22823 28939
rect 22841 28921 22859 28939
rect 22877 28921 22895 28939
rect 22913 28921 22940 28939
rect 22760 28900 22940 28921
rect 25140 28939 25300 28960
rect 25140 28921 25157 28939
rect 25175 28921 25193 28939
rect 25211 28921 25229 28939
rect 25247 28921 25265 28939
rect 25283 28921 25300 28939
rect 25140 28900 25300 28921
rect 20060 28819 21680 28840
rect 20060 28801 21527 28819
rect 21545 28801 21563 28819
rect 21581 28801 21599 28819
rect 21617 28801 21635 28819
rect 21653 28801 21680 28819
rect 20060 28780 21680 28801
rect 23440 28819 24820 28840
rect 23440 28801 23467 28819
rect 23485 28801 23503 28819
rect 23521 28801 23539 28819
rect 23557 28801 23575 28819
rect 23593 28801 24820 28819
rect 23440 28780 24820 28801
rect 17360 28699 17540 28720
rect 17360 28681 17387 28699
rect 17405 28681 17423 28699
rect 17441 28681 17459 28699
rect 17477 28681 17495 28699
rect 17513 28681 17540 28699
rect 17360 28660 17540 28681
rect 19120 28699 21200 28720
rect 19120 28681 19147 28699
rect 19165 28681 19183 28699
rect 19201 28681 19219 28699
rect 19237 28681 19255 28699
rect 19273 28681 21047 28699
rect 21065 28681 21083 28699
rect 21101 28681 21119 28699
rect 21137 28681 21155 28699
rect 21173 28681 21200 28699
rect 19120 28660 21200 28681
rect 23180 28699 24520 28720
rect 23180 28681 23207 28699
rect 23225 28681 23243 28699
rect 23261 28681 23279 28699
rect 23297 28681 23315 28699
rect 23333 28681 24520 28699
rect 23180 28660 24520 28681
rect 14660 28579 16400 28600
rect 14660 28561 14687 28579
rect 14705 28561 14723 28579
rect 14741 28561 14759 28579
rect 14777 28561 14795 28579
rect 14813 28561 16247 28579
rect 16265 28561 16283 28579
rect 16301 28561 16319 28579
rect 16337 28561 16355 28579
rect 16373 28561 16400 28579
rect 14660 28540 16400 28561
rect 18380 28579 19940 28600
rect 18380 28561 18407 28579
rect 18425 28561 18443 28579
rect 18461 28561 18479 28579
rect 18497 28561 18515 28579
rect 18533 28561 19940 28579
rect 18380 28540 19940 28561
rect 24440 28540 24520 28660
rect 24740 28540 24820 28780
rect 25220 28540 25300 28900
rect 27320 28540 27400 29020
rect 27440 29020 28240 29080
rect 27440 28540 27520 29020
rect 27620 28813 28840 28840
rect 27620 28795 28801 28813
rect 28819 28795 28840 28813
rect 27620 28777 28840 28795
rect 27620 28760 28801 28777
rect 27620 28540 27700 28760
rect 28780 28759 28801 28760
rect 28819 28759 28840 28777
rect 28780 28741 28840 28759
rect 28780 28723 28801 28741
rect 28819 28723 28840 28741
rect 28780 28705 28840 28723
rect 27880 28673 28720 28700
rect 27880 28655 28681 28673
rect 28699 28655 28720 28673
rect 28780 28687 28801 28705
rect 28819 28687 28840 28705
rect 28780 28660 28840 28687
rect 27880 28637 28720 28655
rect 27880 28620 28681 28637
rect 27880 28540 27960 28620
rect 28660 28619 28681 28620
rect 28699 28619 28720 28637
rect 28660 28601 28720 28619
rect 28660 28583 28681 28601
rect 28699 28583 28720 28601
rect 28660 28565 28720 28583
rect 28660 28547 28681 28565
rect 28699 28547 28720 28565
rect 28660 28520 28720 28547
rect 28920 28011 29180 28040
rect 28920 27993 28941 28011
rect 28959 27993 28977 28011
rect 28995 27993 29013 28011
rect 29031 27993 29049 28011
rect 29067 27993 29085 28011
rect 29103 27993 29121 28011
rect 29139 27993 29180 28011
rect 28920 27975 29180 27993
rect 28920 27957 28941 27975
rect 28959 27957 28977 27975
rect 28995 27957 29013 27975
rect 29031 27957 29049 27975
rect 29067 27957 29085 27975
rect 29103 27957 29121 27975
rect 29139 27957 29180 27975
rect 28920 27939 29180 27957
rect 28920 27921 28941 27939
rect 28959 27921 28977 27939
rect 28995 27921 29013 27939
rect 29031 27921 29049 27939
rect 29067 27921 29085 27939
rect 29103 27921 29121 27939
rect 29139 27921 29180 27939
rect 28920 27903 29180 27921
rect 28920 27885 28941 27903
rect 28959 27885 28977 27903
rect 28995 27885 29013 27903
rect 29031 27885 29049 27903
rect 29067 27885 29085 27903
rect 29103 27885 29121 27903
rect 29139 27885 29180 27903
rect 28920 27867 29180 27885
rect 28920 27849 28941 27867
rect 28959 27849 28977 27867
rect 28995 27849 29013 27867
rect 29031 27849 29049 27867
rect 29067 27849 29085 27867
rect 29103 27849 29121 27867
rect 29139 27849 29180 27867
rect 28920 27831 29180 27849
rect 28920 27813 28941 27831
rect 28959 27813 28977 27831
rect 28995 27813 29013 27831
rect 29031 27813 29049 27831
rect 29067 27813 29085 27831
rect 29103 27813 29121 27831
rect 29139 27813 29180 27831
rect 28920 27795 29180 27813
rect 28920 27777 28941 27795
rect 28959 27777 28977 27795
rect 28995 27777 29013 27795
rect 29031 27777 29049 27795
rect 29067 27777 29085 27795
rect 29103 27777 29121 27795
rect 29139 27777 29180 27795
rect 28920 27759 29180 27777
rect 28920 27741 28941 27759
rect 28959 27741 28977 27759
rect 28995 27741 29013 27759
rect 29031 27741 29049 27759
rect 29067 27741 29085 27759
rect 29103 27741 29121 27759
rect 29139 27741 29180 27759
rect 28920 27723 29180 27741
rect 28920 27705 28941 27723
rect 28959 27705 28977 27723
rect 28995 27705 29013 27723
rect 29031 27705 29049 27723
rect 29067 27705 29085 27723
rect 29103 27705 29121 27723
rect 29139 27705 29180 27723
rect 28920 27687 29180 27705
rect 28920 27669 28941 27687
rect 28959 27669 28977 27687
rect 28995 27669 29013 27687
rect 29031 27669 29049 27687
rect 29067 27669 29085 27687
rect 29103 27669 29121 27687
rect 29139 27669 29180 27687
rect 28920 27651 29180 27669
rect 28920 27633 28941 27651
rect 28959 27633 28977 27651
rect 28995 27633 29013 27651
rect 29031 27633 29049 27651
rect 29067 27633 29085 27651
rect 29103 27633 29121 27651
rect 29139 27633 29180 27651
rect 28920 27615 29180 27633
rect 28920 27597 28941 27615
rect 28959 27597 28977 27615
rect 28995 27597 29013 27615
rect 29031 27597 29049 27615
rect 29067 27597 29085 27615
rect 29103 27597 29121 27615
rect 29139 27597 29180 27615
rect 28920 27579 29180 27597
rect 28920 27561 28941 27579
rect 28959 27561 28977 27579
rect 28995 27561 29013 27579
rect 29031 27561 29049 27579
rect 29067 27561 29085 27579
rect 29103 27561 29121 27579
rect 29139 27561 29180 27579
rect 28920 27543 29180 27561
rect 28920 27525 28941 27543
rect 28959 27525 28977 27543
rect 28995 27525 29013 27543
rect 29031 27525 29049 27543
rect 29067 27525 29085 27543
rect 29103 27525 29121 27543
rect 29139 27525 29180 27543
rect 28920 27507 29180 27525
rect 28920 27489 28941 27507
rect 28959 27489 28977 27507
rect 28995 27489 29013 27507
rect 29031 27489 29049 27507
rect 29067 27489 29085 27507
rect 29103 27489 29121 27507
rect 29139 27489 29180 27507
rect 28920 27471 29180 27489
rect 28920 27453 28941 27471
rect 28959 27453 28977 27471
rect 28995 27453 29013 27471
rect 29031 27453 29049 27471
rect 29067 27453 29085 27471
rect 29103 27453 29121 27471
rect 29139 27453 29180 27471
rect 28920 27435 29180 27453
rect 28920 27417 28941 27435
rect 28959 27417 28977 27435
rect 28995 27417 29013 27435
rect 29031 27417 29049 27435
rect 29067 27417 29085 27435
rect 29103 27417 29121 27435
rect 29139 27417 29180 27435
rect 28920 27399 29180 27417
rect 28920 27381 28941 27399
rect 28959 27381 28977 27399
rect 28995 27381 29013 27399
rect 29031 27381 29049 27399
rect 29067 27381 29085 27399
rect 29103 27381 29121 27399
rect 29139 27381 29180 27399
rect 28920 27363 29180 27381
rect 28920 27345 28941 27363
rect 28959 27345 28977 27363
rect 28995 27345 29013 27363
rect 29031 27345 29049 27363
rect 29067 27345 29085 27363
rect 29103 27345 29121 27363
rect 29139 27345 29180 27363
rect 28920 27327 29180 27345
rect 28920 27309 28941 27327
rect 28959 27309 28977 27327
rect 28995 27309 29013 27327
rect 29031 27309 29049 27327
rect 29067 27309 29085 27327
rect 29103 27309 29121 27327
rect 29139 27309 29180 27327
rect 28920 27291 29180 27309
rect 28920 27273 28941 27291
rect 28959 27273 28977 27291
rect 28995 27273 29013 27291
rect 29031 27273 29049 27291
rect 29067 27273 29085 27291
rect 29103 27273 29121 27291
rect 29139 27273 29180 27291
rect 28920 27255 29180 27273
rect 28920 27237 28941 27255
rect 28959 27237 28977 27255
rect 28995 27237 29013 27255
rect 29031 27237 29049 27255
rect 29067 27237 29085 27255
rect 29103 27237 29121 27255
rect 29139 27237 29180 27255
rect 8840 26280 9060 27220
rect 28920 27219 29180 27237
rect 28920 27201 28941 27219
rect 28959 27201 28977 27219
rect 28995 27201 29013 27219
rect 29031 27201 29049 27219
rect 29067 27201 29085 27219
rect 29103 27201 29121 27219
rect 29139 27201 29180 27219
rect 28920 27183 29180 27201
rect 28920 27165 28941 27183
rect 28959 27165 28977 27183
rect 28995 27165 29013 27183
rect 29031 27165 29049 27183
rect 29067 27165 29085 27183
rect 29103 27165 29121 27183
rect 29139 27165 29180 27183
rect 28920 27147 29180 27165
rect 28920 27129 28941 27147
rect 28959 27129 28977 27147
rect 28995 27129 29013 27147
rect 29031 27129 29049 27147
rect 29067 27129 29085 27147
rect 29103 27129 29121 27147
rect 29139 27129 29180 27147
rect 28920 27111 29180 27129
rect 28920 27093 28941 27111
rect 28959 27093 28977 27111
rect 28995 27093 29013 27111
rect 29031 27093 29049 27111
rect 29067 27093 29085 27111
rect 29103 27093 29121 27111
rect 29139 27093 29180 27111
rect 28920 27075 29180 27093
rect 28920 27057 28941 27075
rect 28959 27057 28977 27075
rect 28995 27057 29013 27075
rect 29031 27057 29049 27075
rect 29067 27057 29085 27075
rect 29103 27057 29121 27075
rect 29139 27057 29180 27075
rect 28920 27039 29180 27057
rect 28920 27021 28941 27039
rect 28959 27021 28977 27039
rect 28995 27021 29013 27039
rect 29031 27021 29049 27039
rect 29067 27021 29085 27039
rect 29103 27021 29121 27039
rect 29139 27021 29180 27039
rect 28920 27003 29180 27021
rect 28920 26985 28941 27003
rect 28959 26985 28977 27003
rect 28995 26985 29013 27003
rect 29031 26985 29049 27003
rect 29067 26985 29085 27003
rect 29103 26985 29121 27003
rect 29139 26985 29180 27003
rect 28920 26967 29180 26985
rect 28920 26949 28941 26967
rect 28959 26949 28977 26967
rect 28995 26949 29013 26967
rect 29031 26949 29049 26967
rect 29067 26949 29085 26967
rect 29103 26949 29121 26967
rect 29139 26949 29180 26967
rect 28920 26931 29180 26949
rect 28920 26913 28941 26931
rect 28959 26913 28977 26931
rect 28995 26913 29013 26931
rect 29031 26913 29049 26931
rect 29067 26913 29085 26931
rect 29103 26913 29121 26931
rect 29139 26913 29180 26931
rect 28920 26895 29180 26913
rect 28920 26877 28941 26895
rect 28959 26877 28977 26895
rect 28995 26877 29013 26895
rect 29031 26877 29049 26895
rect 29067 26877 29085 26895
rect 29103 26877 29121 26895
rect 29139 26877 29180 26895
rect 28920 26859 29180 26877
rect 28920 26841 28941 26859
rect 28959 26841 28977 26859
rect 28995 26841 29013 26859
rect 29031 26841 29049 26859
rect 29067 26841 29085 26859
rect 29103 26841 29121 26859
rect 29139 26841 29180 26859
rect 28920 26823 29180 26841
rect 28920 26805 28941 26823
rect 28959 26805 28977 26823
rect 28995 26805 29013 26823
rect 29031 26805 29049 26823
rect 29067 26805 29085 26823
rect 29103 26805 29121 26823
rect 29139 26805 29180 26823
rect 28920 26787 29180 26805
rect 28920 26769 28941 26787
rect 28959 26769 28977 26787
rect 28995 26769 29013 26787
rect 29031 26769 29049 26787
rect 29067 26769 29085 26787
rect 29103 26769 29121 26787
rect 29139 26769 29180 26787
rect 28920 26751 29180 26769
rect 28920 26733 28941 26751
rect 28959 26733 28977 26751
rect 28995 26733 29013 26751
rect 29031 26733 29049 26751
rect 29067 26733 29085 26751
rect 29103 26733 29121 26751
rect 29139 26733 29180 26751
rect 28920 26715 29180 26733
rect 28920 26697 28941 26715
rect 28959 26697 28977 26715
rect 28995 26697 29013 26715
rect 29031 26697 29049 26715
rect 29067 26697 29085 26715
rect 29103 26697 29121 26715
rect 29139 26697 29180 26715
rect 28920 26679 29180 26697
rect 28920 26661 28941 26679
rect 28959 26661 28977 26679
rect 28995 26661 29013 26679
rect 29031 26661 29049 26679
rect 29067 26661 29085 26679
rect 29103 26661 29121 26679
rect 29139 26661 29180 26679
rect 28920 26643 29180 26661
rect 28920 26625 28941 26643
rect 28959 26625 28977 26643
rect 28995 26625 29013 26643
rect 29031 26625 29049 26643
rect 29067 26625 29085 26643
rect 29103 26625 29121 26643
rect 29139 26625 29180 26643
rect 28920 26607 29180 26625
rect 28920 26589 28941 26607
rect 28959 26589 28977 26607
rect 28995 26589 29013 26607
rect 29031 26589 29049 26607
rect 29067 26589 29085 26607
rect 29103 26589 29121 26607
rect 29139 26589 29180 26607
rect 28920 26571 29180 26589
rect 28920 26553 28941 26571
rect 28959 26553 28977 26571
rect 28995 26553 29013 26571
rect 29031 26553 29049 26571
rect 29067 26553 29085 26571
rect 29103 26553 29121 26571
rect 29139 26553 29180 26571
rect 28920 26535 29180 26553
rect 28920 26517 28941 26535
rect 28959 26517 28977 26535
rect 28995 26517 29013 26535
rect 29031 26517 29049 26535
rect 29067 26517 29085 26535
rect 29103 26517 29121 26535
rect 29139 26517 29180 26535
rect 28920 26499 29180 26517
rect 28920 26481 28941 26499
rect 28959 26481 28977 26499
rect 28995 26481 29013 26499
rect 29031 26481 29049 26499
rect 29067 26481 29085 26499
rect 29103 26481 29121 26499
rect 29139 26481 29180 26499
rect 28920 26463 29180 26481
rect 28920 26445 28941 26463
rect 28959 26445 28977 26463
rect 28995 26445 29013 26463
rect 29031 26445 29049 26463
rect 29067 26445 29085 26463
rect 29103 26445 29121 26463
rect 29139 26445 29180 26463
rect 28920 26427 29180 26445
rect 28920 26409 28941 26427
rect 28959 26409 28977 26427
rect 28995 26409 29013 26427
rect 29031 26409 29049 26427
rect 29067 26409 29085 26427
rect 29103 26409 29121 26427
rect 29139 26409 29180 26427
rect 28920 26380 29180 26409
rect 8960 26020 9060 26280
rect 28780 26279 29020 26300
rect 28780 26261 28801 26279
rect 28819 26261 28837 26279
rect 28855 26261 28873 26279
rect 28891 26261 28909 26279
rect 28927 26261 28945 26279
rect 28963 26261 28981 26279
rect 28999 26261 29020 26279
rect 28780 26240 29020 26261
rect 28660 26159 28900 26180
rect 28660 26141 28681 26159
rect 28699 26141 28717 26159
rect 28735 26141 28753 26159
rect 28771 26141 28789 26159
rect 28807 26141 28825 26159
rect 28843 26141 28861 26159
rect 28879 26141 28900 26159
rect 28660 26120 28900 26141
rect 8960 25999 9500 26020
rect 8960 25981 8987 25999
rect 9005 25981 9023 25999
rect 9041 25981 9059 25999
rect 9077 25981 9095 25999
rect 9113 25981 9131 25999
rect 9149 25981 9167 25999
rect 9185 25981 9203 25999
rect 9221 25981 9239 25999
rect 9257 25981 9275 25999
rect 9293 25981 9311 25999
rect 9329 25981 9347 25999
rect 9365 25981 9383 25999
rect 9401 25981 9419 25999
rect 9437 25981 9455 25999
rect 9473 25981 9500 25999
rect 8960 25960 9500 25981
rect 9060 25763 9120 25780
rect 9060 25745 9081 25763
rect 9099 25745 9120 25763
rect 9060 25727 9120 25745
rect 9060 25709 9081 25727
rect 9099 25709 9120 25727
rect 9060 25691 9120 25709
rect 9060 25673 9081 25691
rect 9099 25673 9120 25691
rect 9060 25655 9120 25673
rect 9060 25637 9081 25655
rect 9099 25637 9120 25655
rect 9060 25619 9120 25637
rect 9060 25601 9081 25619
rect 9099 25601 9120 25619
rect 9060 25583 9120 25601
rect 9060 25565 9081 25583
rect 9099 25565 9120 25583
rect 9060 25547 9120 25565
rect 9060 25529 9081 25547
rect 9099 25529 9120 25547
rect 9060 25511 9120 25529
rect 9060 25493 9081 25511
rect 9099 25493 9120 25511
rect 9060 25475 9120 25493
rect 9060 25457 9081 25475
rect 9099 25457 9120 25475
rect 9060 24520 9120 25457
rect 8820 23580 9120 24520
rect 9280 25643 9340 25660
rect 9280 25625 9301 25643
rect 9319 25625 9340 25643
rect 9280 25607 9340 25625
rect 9280 25589 9301 25607
rect 9319 25589 9340 25607
rect 9280 25571 9340 25589
rect 9280 25553 9301 25571
rect 9319 25553 9340 25571
rect 9280 25535 9340 25553
rect 9280 25517 9301 25535
rect 9319 25517 9340 25535
rect 9280 21820 9340 25517
rect 28840 25260 28900 26120
rect 28960 25540 29020 26240
rect 28960 25460 29180 25540
rect 28840 25200 29020 25260
rect 28760 24393 28820 24420
rect 28760 24375 28781 24393
rect 28799 24375 28820 24393
rect 28760 24357 28820 24375
rect 28760 24339 28781 24357
rect 28799 24339 28820 24357
rect 28760 24321 28820 24339
rect 28760 24303 28781 24321
rect 28799 24303 28820 24321
rect 28760 24285 28820 24303
rect 28760 24267 28781 24285
rect 28799 24267 28820 24285
rect 28640 24093 28700 24120
rect 28640 24075 28661 24093
rect 28679 24075 28700 24093
rect 28640 24057 28700 24075
rect 28640 24039 28661 24057
rect 28679 24039 28700 24057
rect 28640 24021 28700 24039
rect 28640 24003 28661 24021
rect 28679 24003 28700 24021
rect 28640 23985 28700 24003
rect 28640 23967 28661 23985
rect 28679 23967 28700 23985
rect 8820 20880 9340 21820
rect 28520 22793 28580 22820
rect 28520 22775 28541 22793
rect 28559 22775 28580 22793
rect 28520 22757 28580 22775
rect 28520 22739 28541 22757
rect 28559 22739 28580 22757
rect 28520 22721 28580 22739
rect 28520 22703 28541 22721
rect 28559 22703 28580 22721
rect 28520 22685 28580 22703
rect 28520 22667 28541 22685
rect 28559 22667 28580 22685
rect 8820 20020 9480 20100
rect 9420 18041 9480 20020
rect 28520 19833 28580 22667
rect 28640 21833 28700 23967
rect 28760 22153 28820 24267
rect 28960 22840 29020 25200
rect 28960 22760 29180 22840
rect 28760 22135 28781 22153
rect 28799 22135 28820 22153
rect 28760 22117 28820 22135
rect 28760 22099 28781 22117
rect 28799 22099 28820 22117
rect 28760 22081 28820 22099
rect 28760 22063 28781 22081
rect 28799 22063 28820 22081
rect 28760 22045 28820 22063
rect 28760 22027 28781 22045
rect 28799 22027 28820 22045
rect 28760 22000 28820 22027
rect 28640 21815 28661 21833
rect 28679 21815 28700 21833
rect 28640 21797 28700 21815
rect 28640 21779 28661 21797
rect 28679 21779 28700 21797
rect 28640 21761 28700 21779
rect 28640 21743 28661 21761
rect 28679 21743 28700 21761
rect 28640 21725 28700 21743
rect 28640 21707 28661 21725
rect 28679 21707 28700 21725
rect 28640 21680 28700 21707
rect 28760 20213 28820 20240
rect 28760 20195 28781 20213
rect 28799 20195 28820 20213
rect 28760 20177 28820 20195
rect 28760 20159 28781 20177
rect 28799 20159 28820 20177
rect 28760 20141 28820 20159
rect 28760 20123 28781 20141
rect 28799 20140 28820 20141
rect 28799 20123 29180 20140
rect 28760 20105 29180 20123
rect 28760 20087 28781 20105
rect 28799 20087 29180 20105
rect 28760 20060 29180 20087
rect 28520 19815 28541 19833
rect 28559 19815 28580 19833
rect 28520 19797 28580 19815
rect 28520 19779 28541 19797
rect 28559 19779 28580 19797
rect 28520 19761 28580 19779
rect 28520 19743 28541 19761
rect 28559 19743 28580 19761
rect 28520 19725 28580 19743
rect 28520 19707 28541 19725
rect 28559 19707 28580 19725
rect 28520 19680 28580 19707
rect 9420 18023 9441 18041
rect 9459 18023 9480 18041
rect 9420 18005 9480 18023
rect 9420 17987 9441 18005
rect 9459 17987 9480 18005
rect 9420 17969 9480 17987
rect 9420 17951 9441 17969
rect 9459 17951 9480 17969
rect 9420 17933 9480 17951
rect 9420 17915 9441 17933
rect 9459 17915 9480 17933
rect 9420 17897 9480 17915
rect 9420 17879 9441 17897
rect 9459 17879 9480 17897
rect 9420 17860 9480 17879
rect 28640 19453 28700 19480
rect 28640 19435 28661 19453
rect 28679 19435 28700 19453
rect 28640 19417 28700 19435
rect 28640 19399 28661 19417
rect 28679 19399 28700 19417
rect 28640 19381 28700 19399
rect 28640 19363 28661 19381
rect 28679 19363 28700 19381
rect 28640 19345 28700 19363
rect 28640 19327 28661 19345
rect 28679 19327 28700 19345
rect 28640 17440 28700 19327
rect 8820 17320 9140 17400
rect 28640 17360 29180 17440
rect 9080 16401 9140 17320
rect 9080 16383 9101 16401
rect 9119 16383 9140 16401
rect 9080 16365 9140 16383
rect 9080 16347 9101 16365
rect 9119 16347 9140 16365
rect 9080 16329 9140 16347
rect 9080 16311 9101 16329
rect 9119 16311 9140 16329
rect 9080 16293 9140 16311
rect 9080 16275 9101 16293
rect 9119 16275 9140 16293
rect 9080 16257 9140 16275
rect 9080 16239 9101 16257
rect 9119 16239 9140 16257
rect 9080 16220 9140 16239
rect 28520 16653 28580 16680
rect 28520 16635 28541 16653
rect 28559 16635 28580 16653
rect 28520 16617 28580 16635
rect 28520 16599 28541 16617
rect 28559 16599 28580 16617
rect 28520 16581 28580 16599
rect 28520 16563 28541 16581
rect 28559 16563 28580 16581
rect 28520 16545 28580 16563
rect 28520 16527 28541 16545
rect 28559 16527 28580 16545
rect 28520 14740 28580 16527
rect 8820 14620 9120 14700
rect 28520 14660 29180 14740
rect 9060 13293 9120 14620
rect 9060 13275 9081 13293
rect 9099 13275 9120 13293
rect 9060 13257 9120 13275
rect 9060 13239 9081 13257
rect 9099 13239 9120 13257
rect 9060 13221 9120 13239
rect 9060 13203 9081 13221
rect 9099 13203 9120 13221
rect 9060 13185 9120 13203
rect 9060 13167 9081 13185
rect 9099 13167 9120 13185
rect 9060 13140 9120 13167
rect 28660 12103 28720 12120
rect 28660 12085 28681 12103
rect 28699 12085 28720 12103
rect 28660 12067 28720 12085
rect 28660 12049 28681 12067
rect 28699 12049 28720 12067
rect 28660 12040 28720 12049
rect 28660 12031 29180 12040
rect 28660 12013 28681 12031
rect 28699 12013 29180 12031
rect 28660 11995 29180 12013
rect 28660 11977 28681 11995
rect 28699 11977 29180 11995
rect 28660 11960 29180 11977
rect 8820 11539 9080 11560
rect 8820 11521 8861 11539
rect 8879 11521 8897 11539
rect 8915 11521 8933 11539
rect 8951 11521 8969 11539
rect 8987 11521 9005 11539
rect 9023 11521 9041 11539
rect 9059 11521 9080 11539
rect 8820 11503 9080 11521
rect 8820 11485 8861 11503
rect 8879 11485 8897 11503
rect 8915 11485 8933 11503
rect 8951 11485 8969 11503
rect 8987 11485 9005 11503
rect 9023 11485 9041 11503
rect 9059 11485 9080 11503
rect 8820 11467 9080 11485
rect 8820 11449 8861 11467
rect 8879 11449 8897 11467
rect 8915 11449 8933 11467
rect 8951 11449 8969 11467
rect 8987 11449 9005 11467
rect 9023 11449 9041 11467
rect 9059 11449 9080 11467
rect 8820 11431 9080 11449
rect 8820 11413 8861 11431
rect 8879 11413 8897 11431
rect 8915 11413 8933 11431
rect 8951 11413 8969 11431
rect 8987 11413 9005 11431
rect 9023 11413 9041 11431
rect 9059 11413 9080 11431
rect 8820 11395 9080 11413
rect 8820 11377 8861 11395
rect 8879 11377 8897 11395
rect 8915 11377 8933 11395
rect 8951 11377 8969 11395
rect 8987 11377 9005 11395
rect 9023 11377 9041 11395
rect 9059 11377 9080 11395
rect 8820 11359 9080 11377
rect 8820 11341 8861 11359
rect 8879 11341 8897 11359
rect 8915 11341 8933 11359
rect 8951 11341 8969 11359
rect 8987 11341 9005 11359
rect 9023 11341 9041 11359
rect 9059 11341 9080 11359
rect 8820 11323 9080 11341
rect 8820 11305 8861 11323
rect 8879 11305 8897 11323
rect 8915 11305 8933 11323
rect 8951 11305 8969 11323
rect 8987 11305 9005 11323
rect 9023 11305 9041 11323
rect 9059 11305 9080 11323
rect 8820 11287 9080 11305
rect 8820 11269 8861 11287
rect 8879 11269 8897 11287
rect 8915 11269 8933 11287
rect 8951 11269 8969 11287
rect 8987 11269 9005 11287
rect 9023 11269 9041 11287
rect 9059 11269 9080 11287
rect 8820 11251 9080 11269
rect 8820 11233 8861 11251
rect 8879 11233 8897 11251
rect 8915 11233 8933 11251
rect 8951 11233 8969 11251
rect 8987 11233 9005 11251
rect 9023 11233 9041 11251
rect 9059 11233 9080 11251
rect 8820 11215 9080 11233
rect 8820 11197 8861 11215
rect 8879 11197 8897 11215
rect 8915 11197 8933 11215
rect 8951 11197 8969 11215
rect 8987 11197 9005 11215
rect 9023 11197 9041 11215
rect 9059 11197 9080 11215
rect 8820 11179 9080 11197
rect 8820 11161 8861 11179
rect 8879 11161 8897 11179
rect 8915 11161 8933 11179
rect 8951 11161 8969 11179
rect 8987 11161 9005 11179
rect 9023 11161 9041 11179
rect 9059 11161 9080 11179
rect 8820 11143 9080 11161
rect 8820 11125 8861 11143
rect 8879 11125 8897 11143
rect 8915 11125 8933 11143
rect 8951 11125 8969 11143
rect 8987 11125 9005 11143
rect 9023 11125 9041 11143
rect 9059 11125 9080 11143
rect 8820 11107 9080 11125
rect 8820 11089 8861 11107
rect 8879 11089 8897 11107
rect 8915 11089 8933 11107
rect 8951 11089 8969 11107
rect 8987 11089 9005 11107
rect 9023 11089 9041 11107
rect 9059 11089 9080 11107
rect 8820 11071 9080 11089
rect 8820 11053 8861 11071
rect 8879 11053 8897 11071
rect 8915 11053 8933 11071
rect 8951 11053 8969 11071
rect 8987 11053 9005 11071
rect 9023 11053 9041 11071
rect 9059 11053 9080 11071
rect 8820 11035 9080 11053
rect 8820 11017 8861 11035
rect 8879 11017 8897 11035
rect 8915 11017 8933 11035
rect 8951 11017 8969 11035
rect 8987 11017 9005 11035
rect 9023 11017 9041 11035
rect 9059 11017 9080 11035
rect 8820 10999 9080 11017
rect 8820 10981 8861 10999
rect 8879 10981 8897 10999
rect 8915 10981 8933 10999
rect 8951 10981 8969 10999
rect 8987 10981 9005 10999
rect 9023 10981 9041 10999
rect 9059 10981 9080 10999
rect 8820 10963 9080 10981
rect 8820 10945 8861 10963
rect 8879 10945 8897 10963
rect 8915 10945 8933 10963
rect 8951 10945 8969 10963
rect 8987 10945 9005 10963
rect 9023 10945 9041 10963
rect 9059 10945 9080 10963
rect 8820 10927 9080 10945
rect 8820 10909 8861 10927
rect 8879 10909 8897 10927
rect 8915 10909 8933 10927
rect 8951 10909 8969 10927
rect 8987 10909 9005 10927
rect 9023 10909 9041 10927
rect 9059 10909 9080 10927
rect 8820 10891 9080 10909
rect 8820 10873 8861 10891
rect 8879 10873 8897 10891
rect 8915 10873 8933 10891
rect 8951 10873 8969 10891
rect 8987 10873 9005 10891
rect 9023 10873 9041 10891
rect 9059 10873 9080 10891
rect 8820 10855 9080 10873
rect 8820 10837 8861 10855
rect 8879 10837 8897 10855
rect 8915 10837 8933 10855
rect 8951 10837 8969 10855
rect 8987 10837 9005 10855
rect 9023 10837 9041 10855
rect 9059 10837 9080 10855
rect 8820 10819 9080 10837
rect 8820 10801 8861 10819
rect 8879 10801 8897 10819
rect 8915 10801 8933 10819
rect 8951 10801 8969 10819
rect 8987 10801 9005 10819
rect 9023 10801 9041 10819
rect 9059 10801 9080 10819
rect 8820 10783 9080 10801
rect 8820 10765 8861 10783
rect 8879 10765 8897 10783
rect 8915 10765 8933 10783
rect 8951 10765 8969 10783
rect 8987 10765 9005 10783
rect 9023 10765 9041 10783
rect 9059 10765 9080 10783
rect 8820 10747 9080 10765
rect 8820 10729 8861 10747
rect 8879 10729 8897 10747
rect 8915 10729 8933 10747
rect 8951 10729 8969 10747
rect 8987 10729 9005 10747
rect 9023 10729 9041 10747
rect 9059 10729 9080 10747
rect 8820 10711 9080 10729
rect 8820 10693 8861 10711
rect 8879 10693 8897 10711
rect 8915 10693 8933 10711
rect 8951 10693 8969 10711
rect 8987 10693 9005 10711
rect 9023 10693 9041 10711
rect 9059 10693 9080 10711
rect 8820 10675 9080 10693
rect 8820 10657 8861 10675
rect 8879 10657 8897 10675
rect 8915 10657 8933 10675
rect 8951 10657 8969 10675
rect 8987 10657 9005 10675
rect 9023 10657 9041 10675
rect 9059 10657 9080 10675
rect 8820 10639 9080 10657
rect 8820 10621 8861 10639
rect 8879 10621 8897 10639
rect 8915 10621 8933 10639
rect 8951 10621 8969 10639
rect 8987 10621 9005 10639
rect 9023 10621 9041 10639
rect 9059 10621 9080 10639
rect 8820 10603 9080 10621
rect 8820 10585 8861 10603
rect 8879 10585 8897 10603
rect 8915 10585 8933 10603
rect 8951 10585 8969 10603
rect 8987 10585 9005 10603
rect 9023 10585 9041 10603
rect 9059 10585 9080 10603
rect 8820 10567 9080 10585
rect 8820 10549 8861 10567
rect 8879 10549 8897 10567
rect 8915 10549 8933 10567
rect 8951 10549 8969 10567
rect 8987 10549 9005 10567
rect 9023 10549 9041 10567
rect 9059 10549 9080 10567
rect 8820 10531 9080 10549
rect 8820 10513 8861 10531
rect 8879 10513 8897 10531
rect 8915 10513 8933 10531
rect 8951 10513 8969 10531
rect 8987 10513 9005 10531
rect 9023 10513 9041 10531
rect 9059 10513 9080 10531
rect 8820 10495 9080 10513
rect 8820 10477 8861 10495
rect 8879 10477 8897 10495
rect 8915 10477 8933 10495
rect 8951 10477 8969 10495
rect 8987 10477 9005 10495
rect 9023 10477 9041 10495
rect 9059 10477 9080 10495
rect 8820 10459 9080 10477
rect 8820 10441 8861 10459
rect 8879 10441 8897 10459
rect 8915 10441 8933 10459
rect 8951 10441 8969 10459
rect 8987 10441 9005 10459
rect 9023 10441 9041 10459
rect 9059 10441 9080 10459
rect 8820 10423 9080 10441
rect 8820 10405 8861 10423
rect 8879 10405 8897 10423
rect 8915 10405 8933 10423
rect 8951 10405 8969 10423
rect 8987 10405 9005 10423
rect 9023 10405 9041 10423
rect 9059 10405 9080 10423
rect 8820 10387 9080 10405
rect 8820 10369 8861 10387
rect 8879 10369 8897 10387
rect 8915 10369 8933 10387
rect 8951 10369 8969 10387
rect 8987 10369 9005 10387
rect 9023 10369 9041 10387
rect 9059 10369 9080 10387
rect 8820 10351 9080 10369
rect 8820 10333 8861 10351
rect 8879 10333 8897 10351
rect 8915 10333 8933 10351
rect 8951 10333 8969 10351
rect 8987 10333 9005 10351
rect 9023 10333 9041 10351
rect 9059 10333 9080 10351
rect 8820 10315 9080 10333
rect 8820 10297 8861 10315
rect 8879 10297 8897 10315
rect 8915 10297 8933 10315
rect 8951 10297 8969 10315
rect 8987 10297 9005 10315
rect 9023 10297 9041 10315
rect 9059 10297 9080 10315
rect 8820 10279 9080 10297
rect 8820 10261 8861 10279
rect 8879 10261 8897 10279
rect 8915 10261 8933 10279
rect 8951 10261 8969 10279
rect 8987 10261 9005 10279
rect 9023 10261 9041 10279
rect 9059 10261 9080 10279
rect 8820 10240 9080 10261
rect 28540 11143 28600 11160
rect 28540 11125 28561 11143
rect 28579 11125 28600 11143
rect 28540 11107 28600 11125
rect 28540 11089 28561 11107
rect 28579 11089 28600 11107
rect 28540 11071 28600 11089
rect 28540 11053 28561 11071
rect 28579 11053 28600 11071
rect 28540 11035 28600 11053
rect 28540 11017 28561 11035
rect 28579 11017 28600 11035
rect 9800 9579 9980 9600
rect 9800 9561 9827 9579
rect 9845 9561 9863 9579
rect 9881 9561 9899 9579
rect 9917 9561 9935 9579
rect 9953 9561 9980 9579
rect 9800 9540 9980 9561
rect 12720 9579 15640 9600
rect 12720 9561 12747 9579
rect 12765 9561 12783 9579
rect 12801 9561 12819 9579
rect 12837 9561 12855 9579
rect 12873 9561 15487 9579
rect 15505 9561 15523 9579
rect 15541 9561 15559 9579
rect 15577 9561 15595 9579
rect 15613 9561 15640 9579
rect 12720 9540 15640 9561
rect 18480 9579 21100 9600
rect 18480 9561 18507 9579
rect 18525 9561 18543 9579
rect 18561 9561 18579 9579
rect 18597 9561 18615 9579
rect 18633 9561 20947 9579
rect 20965 9561 20983 9579
rect 21001 9561 21019 9579
rect 21037 9561 21055 9579
rect 21073 9561 21100 9579
rect 18480 9540 21100 9561
rect 23780 9579 23940 9600
rect 23780 9561 23797 9579
rect 23815 9561 23833 9579
rect 23851 9561 23869 9579
rect 23887 9561 23905 9579
rect 23923 9561 23940 9579
rect 23780 9540 23940 9561
rect 9800 8820 9880 9540
rect 25000 9480 25080 9580
rect 12500 9459 15560 9480
rect 12500 9441 12527 9459
rect 12545 9441 12563 9459
rect 12581 9441 12599 9459
rect 12617 9441 12635 9459
rect 12653 9441 15407 9459
rect 15425 9441 15443 9459
rect 15461 9441 15479 9459
rect 15497 9441 15515 9459
rect 15533 9441 15560 9459
rect 12500 9420 15560 9441
rect 18280 9459 21340 9480
rect 18280 9441 18307 9459
rect 18325 9441 18343 9459
rect 18361 9441 18379 9459
rect 18397 9441 18415 9459
rect 18433 9441 21187 9459
rect 21205 9441 21223 9459
rect 21241 9441 21259 9459
rect 21277 9441 21295 9459
rect 21313 9441 21340 9459
rect 18280 9420 21340 9441
rect 23400 9459 25080 9480
rect 23400 9441 23427 9459
rect 23445 9441 23463 9459
rect 23481 9441 23499 9459
rect 23517 9441 23535 9459
rect 23553 9441 25080 9459
rect 23400 9420 25080 9441
rect 12500 8820 12580 9420
rect 26080 9360 26160 9600
rect 15200 9339 21160 9360
rect 15200 9321 15227 9339
rect 15245 9321 15263 9339
rect 15281 9321 15299 9339
rect 15317 9321 15335 9339
rect 15353 9321 18107 9339
rect 18125 9321 18143 9339
rect 18161 9321 18179 9339
rect 18197 9321 18215 9339
rect 18233 9321 21007 9339
rect 21025 9321 21043 9339
rect 21061 9321 21079 9339
rect 21097 9321 21115 9339
rect 21133 9321 21160 9339
rect 15200 9300 21160 9321
rect 23580 9339 26160 9360
rect 23580 9321 23607 9339
rect 23625 9321 23643 9339
rect 23661 9321 23679 9339
rect 23697 9321 23715 9339
rect 23733 9321 26160 9339
rect 23580 9300 26160 9321
rect 15200 8820 15280 9300
rect 26500 9240 26560 9600
rect 17900 9219 20960 9240
rect 17900 9201 17927 9219
rect 17945 9201 17963 9219
rect 17981 9201 17999 9219
rect 18017 9201 18035 9219
rect 18053 9201 20807 9219
rect 20825 9201 20843 9219
rect 20861 9201 20879 9219
rect 20897 9201 20915 9219
rect 20933 9201 20960 9219
rect 17900 9180 20960 9201
rect 23860 9219 26560 9240
rect 23860 9201 23887 9219
rect 23905 9201 23923 9219
rect 23941 9201 23959 9219
rect 23977 9201 23995 9219
rect 24013 9201 26560 9219
rect 23860 9180 26560 9201
rect 17900 8820 17980 9180
rect 26900 9120 26960 9600
rect 20600 9099 23240 9120
rect 20600 9081 20627 9099
rect 20645 9081 20663 9099
rect 20681 9081 20699 9099
rect 20717 9081 20735 9099
rect 20753 9081 23087 9099
rect 23105 9081 23123 9099
rect 23141 9081 23159 9099
rect 23177 9081 23195 9099
rect 23213 9081 23240 9099
rect 20600 9060 23240 9081
rect 26280 9099 26960 9120
rect 26280 9081 26307 9099
rect 26325 9081 26343 9099
rect 26361 9081 26379 9099
rect 26397 9081 26415 9099
rect 26433 9081 26960 9099
rect 26280 9060 26960 9081
rect 20600 8820 20680 9060
rect 27260 9000 27320 9600
rect 28540 9373 28600 11017
rect 28540 9355 28561 9373
rect 28579 9355 28600 9373
rect 28540 9337 28600 9355
rect 23300 8979 27320 9000
rect 23300 8961 24747 8979
rect 24765 8961 24783 8979
rect 24801 8961 24819 8979
rect 24837 8961 24855 8979
rect 24873 8961 27167 8979
rect 27185 8961 27203 8979
rect 27221 8961 27239 8979
rect 27257 8961 27275 8979
rect 27293 8961 27320 8979
rect 23300 8940 27320 8961
rect 28160 9297 28340 9320
rect 28160 9279 28187 9297
rect 28205 9279 28223 9297
rect 28241 9279 28259 9297
rect 28277 9279 28295 9297
rect 28313 9279 28340 9297
rect 28160 9261 28340 9279
rect 28160 9243 28187 9261
rect 28205 9243 28223 9261
rect 28241 9243 28259 9261
rect 28277 9243 28295 9261
rect 28313 9243 28340 9261
rect 28160 9220 28340 9243
rect 28540 9319 28561 9337
rect 28579 9319 28600 9337
rect 28540 9301 28600 9319
rect 28540 9283 28561 9301
rect 28579 9283 28600 9301
rect 28540 9265 28600 9283
rect 28540 9247 28561 9265
rect 28579 9247 28600 9265
rect 28540 9220 28600 9247
rect 23300 8820 23380 8940
rect 28160 8820 28260 9220
<< m3contact >>
rect 25477 29041 25495 29059
rect 25513 29041 25531 29059
rect 25549 29041 25567 29059
rect 25585 29041 25603 29059
rect 27257 29041 27275 29059
rect 27293 29041 27311 29059
rect 27329 29041 27347 29059
rect 27365 29041 27383 29059
rect 22787 28921 22805 28939
rect 22823 28921 22841 28939
rect 22859 28921 22877 28939
rect 22895 28921 22913 28939
rect 25157 28921 25175 28939
rect 25193 28921 25211 28939
rect 25229 28921 25247 28939
rect 25265 28921 25283 28939
rect 21527 28801 21545 28819
rect 21563 28801 21581 28819
rect 21599 28801 21617 28819
rect 21635 28801 21653 28819
rect 23467 28801 23485 28819
rect 23503 28801 23521 28819
rect 23539 28801 23557 28819
rect 23575 28801 23593 28819
rect 17387 28681 17405 28699
rect 17423 28681 17441 28699
rect 17459 28681 17477 28699
rect 17495 28681 17513 28699
rect 19147 28681 19165 28699
rect 19183 28681 19201 28699
rect 19219 28681 19237 28699
rect 19255 28681 19273 28699
rect 21047 28681 21065 28699
rect 21083 28681 21101 28699
rect 21119 28681 21137 28699
rect 21155 28681 21173 28699
rect 23207 28681 23225 28699
rect 23243 28681 23261 28699
rect 23279 28681 23297 28699
rect 23315 28681 23333 28699
rect 14687 28561 14705 28579
rect 14723 28561 14741 28579
rect 14759 28561 14777 28579
rect 14795 28561 14813 28579
rect 16247 28561 16265 28579
rect 16283 28561 16301 28579
rect 16319 28561 16337 28579
rect 16355 28561 16373 28579
rect 18407 28561 18425 28579
rect 18443 28561 18461 28579
rect 18479 28561 18497 28579
rect 18515 28561 18533 28579
rect 28801 28795 28819 28813
rect 28801 28759 28819 28777
rect 28801 28723 28819 28741
rect 28681 28655 28699 28673
rect 28801 28687 28819 28705
rect 28681 28619 28699 28637
rect 28681 28583 28699 28601
rect 28681 28547 28699 28565
rect 28801 26261 28819 26279
rect 28837 26261 28855 26279
rect 28873 26261 28891 26279
rect 28909 26261 28927 26279
rect 28945 26261 28963 26279
rect 28981 26261 28999 26279
rect 28681 26141 28699 26159
rect 28717 26141 28735 26159
rect 28753 26141 28771 26159
rect 28789 26141 28807 26159
rect 28825 26141 28843 26159
rect 28861 26141 28879 26159
rect 28781 24375 28799 24393
rect 28781 24339 28799 24357
rect 28781 24303 28799 24321
rect 28781 24267 28799 24285
rect 28661 24075 28679 24093
rect 28661 24039 28679 24057
rect 28661 24003 28679 24021
rect 28661 23967 28679 23985
rect 28541 22775 28559 22793
rect 28541 22739 28559 22757
rect 28541 22703 28559 22721
rect 28541 22667 28559 22685
rect 28781 22135 28799 22153
rect 28781 22099 28799 22117
rect 28781 22063 28799 22081
rect 28781 22027 28799 22045
rect 28661 21815 28679 21833
rect 28661 21779 28679 21797
rect 28661 21743 28679 21761
rect 28661 21707 28679 21725
rect 28781 20195 28799 20213
rect 28781 20159 28799 20177
rect 28781 20123 28799 20141
rect 28781 20087 28799 20105
rect 28541 19815 28559 19833
rect 28541 19779 28559 19797
rect 28541 19743 28559 19761
rect 28541 19707 28559 19725
rect 9441 18023 9459 18041
rect 9441 17987 9459 18005
rect 9441 17951 9459 17969
rect 9441 17915 9459 17933
rect 9441 17879 9459 17897
rect 28661 19435 28679 19453
rect 28661 19399 28679 19417
rect 28661 19363 28679 19381
rect 28661 19327 28679 19345
rect 9101 16383 9119 16401
rect 9101 16347 9119 16365
rect 9101 16311 9119 16329
rect 9101 16275 9119 16293
rect 9101 16239 9119 16257
rect 28541 16635 28559 16653
rect 28541 16599 28559 16617
rect 28541 16563 28559 16581
rect 28541 16527 28559 16545
rect 9081 13275 9099 13293
rect 9081 13239 9099 13257
rect 9081 13203 9099 13221
rect 9081 13167 9099 13185
rect 28681 12085 28699 12103
rect 28681 12049 28699 12067
rect 28681 12013 28699 12031
rect 28681 11977 28699 11995
rect 28561 11125 28579 11143
rect 28561 11089 28579 11107
rect 28561 11053 28579 11071
rect 28561 11017 28579 11035
rect 9827 9561 9845 9579
rect 9863 9561 9881 9579
rect 9899 9561 9917 9579
rect 9935 9561 9953 9579
rect 12747 9561 12765 9579
rect 12783 9561 12801 9579
rect 12819 9561 12837 9579
rect 12855 9561 12873 9579
rect 15487 9561 15505 9579
rect 15523 9561 15541 9579
rect 15559 9561 15577 9579
rect 15595 9561 15613 9579
rect 18507 9561 18525 9579
rect 18543 9561 18561 9579
rect 18579 9561 18597 9579
rect 18615 9561 18633 9579
rect 20947 9561 20965 9579
rect 20983 9561 21001 9579
rect 21019 9561 21037 9579
rect 21055 9561 21073 9579
rect 23797 9561 23815 9579
rect 23833 9561 23851 9579
rect 23869 9561 23887 9579
rect 23905 9561 23923 9579
rect 12527 9441 12545 9459
rect 12563 9441 12581 9459
rect 12599 9441 12617 9459
rect 12635 9441 12653 9459
rect 15407 9441 15425 9459
rect 15443 9441 15461 9459
rect 15479 9441 15497 9459
rect 15515 9441 15533 9459
rect 18307 9441 18325 9459
rect 18343 9441 18361 9459
rect 18379 9441 18397 9459
rect 18415 9441 18433 9459
rect 21187 9441 21205 9459
rect 21223 9441 21241 9459
rect 21259 9441 21277 9459
rect 21295 9441 21313 9459
rect 23427 9441 23445 9459
rect 23463 9441 23481 9459
rect 23499 9441 23517 9459
rect 23535 9441 23553 9459
rect 15227 9321 15245 9339
rect 15263 9321 15281 9339
rect 15299 9321 15317 9339
rect 15335 9321 15353 9339
rect 18107 9321 18125 9339
rect 18143 9321 18161 9339
rect 18179 9321 18197 9339
rect 18215 9321 18233 9339
rect 21007 9321 21025 9339
rect 21043 9321 21061 9339
rect 21079 9321 21097 9339
rect 21115 9321 21133 9339
rect 23607 9321 23625 9339
rect 23643 9321 23661 9339
rect 23679 9321 23697 9339
rect 23715 9321 23733 9339
rect 17927 9201 17945 9219
rect 17963 9201 17981 9219
rect 17999 9201 18017 9219
rect 18035 9201 18053 9219
rect 20807 9201 20825 9219
rect 20843 9201 20861 9219
rect 20879 9201 20897 9219
rect 20915 9201 20933 9219
rect 23887 9201 23905 9219
rect 23923 9201 23941 9219
rect 23959 9201 23977 9219
rect 23995 9201 24013 9219
rect 20627 9081 20645 9099
rect 20663 9081 20681 9099
rect 20699 9081 20717 9099
rect 20735 9081 20753 9099
rect 23087 9081 23105 9099
rect 23123 9081 23141 9099
rect 23159 9081 23177 9099
rect 23195 9081 23213 9099
rect 26307 9081 26325 9099
rect 26343 9081 26361 9099
rect 26379 9081 26397 9099
rect 26415 9081 26433 9099
rect 28561 9355 28579 9373
rect 24747 8961 24765 8979
rect 24783 8961 24801 8979
rect 24819 8961 24837 8979
rect 24855 8961 24873 8979
rect 27167 8961 27185 8979
rect 27203 8961 27221 8979
rect 27239 8961 27257 8979
rect 27275 8961 27293 8979
rect 28187 9279 28205 9297
rect 28223 9279 28241 9297
rect 28259 9279 28277 9297
rect 28295 9279 28313 9297
rect 28187 9243 28205 9261
rect 28223 9243 28241 9261
rect 28259 9243 28277 9261
rect 28295 9243 28313 9261
rect 28561 9319 28579 9337
rect 28561 9283 28579 9301
rect 28561 9247 28579 9265
<< metal3 >>
rect 25460 29059 27400 29080
rect 25460 29041 25477 29059
rect 25495 29041 25513 29059
rect 25531 29041 25549 29059
rect 25567 29041 25585 29059
rect 25603 29041 27257 29059
rect 27275 29041 27293 29059
rect 27311 29041 27329 29059
rect 27347 29041 27365 29059
rect 27383 29041 27400 29059
rect 25460 29020 27400 29041
rect 22760 28939 25300 28960
rect 22760 28921 22787 28939
rect 22805 28921 22823 28939
rect 22841 28921 22859 28939
rect 22877 28921 22895 28939
rect 22913 28921 25157 28939
rect 25175 28921 25193 28939
rect 25211 28921 25229 28939
rect 25247 28921 25265 28939
rect 25283 28921 25300 28939
rect 22760 28900 25300 28921
rect 21500 28819 23620 28840
rect 21500 28801 21527 28819
rect 21545 28801 21563 28819
rect 21581 28801 21599 28819
rect 21617 28801 21635 28819
rect 21653 28801 23467 28819
rect 23485 28801 23503 28819
rect 23521 28801 23539 28819
rect 23557 28801 23575 28819
rect 23593 28801 23620 28819
rect 21500 28780 23620 28801
rect 28780 28813 28840 28840
rect 28780 28795 28801 28813
rect 28819 28795 28840 28813
rect 28780 28777 28840 28795
rect 28780 28759 28801 28777
rect 28819 28759 28840 28777
rect 28780 28741 28840 28759
rect 28780 28723 28801 28741
rect 28819 28723 28840 28741
rect 17360 28699 19300 28720
rect 17360 28681 17387 28699
rect 17405 28681 17423 28699
rect 17441 28681 17459 28699
rect 17477 28681 17495 28699
rect 17513 28681 19147 28699
rect 19165 28681 19183 28699
rect 19201 28681 19219 28699
rect 19237 28681 19255 28699
rect 19273 28681 19300 28699
rect 17360 28660 19300 28681
rect 21020 28699 23360 28720
rect 28780 28705 28840 28723
rect 21020 28681 21047 28699
rect 21065 28681 21083 28699
rect 21101 28681 21119 28699
rect 21137 28681 21155 28699
rect 21173 28681 23207 28699
rect 23225 28681 23243 28699
rect 23261 28681 23279 28699
rect 23297 28681 23315 28699
rect 23333 28681 23360 28699
rect 21020 28660 23360 28681
rect 28660 28673 28720 28700
rect 28660 28655 28681 28673
rect 28699 28655 28720 28673
rect 28660 28637 28720 28655
rect 28660 28619 28681 28637
rect 28699 28619 28720 28637
rect 28660 28601 28720 28619
rect 14660 28579 14840 28600
rect 14660 28561 14687 28579
rect 14705 28561 14723 28579
rect 14741 28561 14759 28579
rect 14777 28561 14795 28579
rect 14813 28561 14840 28579
rect 14660 28540 14840 28561
rect 16220 28579 18560 28600
rect 16220 28561 16247 28579
rect 16265 28561 16283 28579
rect 16301 28561 16319 28579
rect 16337 28561 16355 28579
rect 16373 28561 18407 28579
rect 18425 28561 18443 28579
rect 18461 28561 18479 28579
rect 18497 28561 18515 28579
rect 18533 28561 18560 28579
rect 16220 28540 18560 28561
rect 28660 28583 28681 28601
rect 28699 28583 28720 28601
rect 28660 28565 28720 28583
rect 28660 28547 28681 28565
rect 28699 28547 28720 28565
rect 28660 26180 28720 28547
rect 28780 28687 28801 28705
rect 28819 28687 28840 28705
rect 28780 26300 28840 28687
rect 28780 26279 29020 26300
rect 28780 26261 28801 26279
rect 28819 26261 28837 26279
rect 28855 26261 28873 26279
rect 28891 26261 28909 26279
rect 28927 26261 28945 26279
rect 28963 26261 28981 26279
rect 28999 26261 29020 26279
rect 28780 26240 29020 26261
rect 28660 26159 28900 26180
rect 28660 26141 28681 26159
rect 28699 26141 28717 26159
rect 28735 26141 28753 26159
rect 28771 26141 28789 26159
rect 28807 26141 28825 26159
rect 28843 26141 28861 26159
rect 28879 26141 28900 26159
rect 28660 26120 28900 26141
rect 28420 25920 28820 26000
rect 28500 25460 28700 25520
rect 28520 22793 28580 25220
rect 28640 24093 28700 25460
rect 28760 24393 28820 25920
rect 28760 24375 28781 24393
rect 28799 24375 28820 24393
rect 28760 24357 28820 24375
rect 28760 24339 28781 24357
rect 28799 24339 28820 24357
rect 28760 24321 28820 24339
rect 28760 24303 28781 24321
rect 28799 24303 28820 24321
rect 28760 24285 28820 24303
rect 28760 24267 28781 24285
rect 28799 24267 28820 24285
rect 28760 24240 28820 24267
rect 28640 24075 28661 24093
rect 28679 24075 28700 24093
rect 28640 24057 28700 24075
rect 28640 24039 28661 24057
rect 28679 24039 28700 24057
rect 28640 24021 28700 24039
rect 28640 24003 28661 24021
rect 28679 24003 28700 24021
rect 28640 23985 28700 24003
rect 28640 23967 28661 23985
rect 28679 23967 28700 23985
rect 28640 23940 28700 23967
rect 28520 22775 28541 22793
rect 28559 22775 28580 22793
rect 28520 22757 28580 22775
rect 28520 22739 28541 22757
rect 28559 22739 28580 22757
rect 28520 22721 28580 22739
rect 28520 22703 28541 22721
rect 28559 22703 28580 22721
rect 28520 22685 28580 22703
rect 28520 22667 28541 22685
rect 28559 22667 28580 22685
rect 28520 22640 28580 22667
rect 28760 22153 28820 22180
rect 28760 22135 28781 22153
rect 28799 22135 28820 22153
rect 28760 22117 28820 22135
rect 28760 22099 28781 22117
rect 28799 22099 28820 22117
rect 28760 22081 28820 22099
rect 28760 22063 28781 22081
rect 28799 22063 28820 22081
rect 28760 22045 28820 22063
rect 28760 22027 28781 22045
rect 28799 22027 28820 22045
rect 28640 21833 28700 21860
rect 28640 21815 28661 21833
rect 28679 21815 28700 21833
rect 28640 21797 28700 21815
rect 28640 21779 28661 21797
rect 28679 21779 28700 21797
rect 28640 21761 28700 21779
rect 28640 21743 28661 21761
rect 28679 21743 28700 21761
rect 28640 21725 28700 21743
rect 28640 21707 28661 21725
rect 28679 21707 28700 21725
rect 28520 19833 28580 19860
rect 28520 19815 28541 19833
rect 28559 19815 28580 19833
rect 28520 19797 28580 19815
rect 28520 19779 28541 19797
rect 28559 19779 28580 19797
rect 28520 19761 28580 19779
rect 28520 19743 28541 19761
rect 28559 19743 28580 19761
rect 28520 19725 28580 19743
rect 28520 19707 28541 19725
rect 28559 19707 28580 19725
rect 9420 18041 9480 18060
rect 9420 18023 9441 18041
rect 9459 18023 9480 18041
rect 9420 18005 9480 18023
rect 9420 17987 9441 18005
rect 9459 17987 9480 18005
rect 9420 17969 9480 17987
rect 9420 17951 9441 17969
rect 9459 17951 9480 17969
rect 9420 17933 9480 17951
rect 9420 17915 9441 17933
rect 9459 17915 9480 17933
rect 9420 17897 9480 17915
rect 9420 17879 9441 17897
rect 9459 17879 9480 17897
rect 9420 16480 9480 17879
rect 28520 16653 28580 19707
rect 28640 19453 28700 21707
rect 28760 20213 28820 22027
rect 28760 20195 28781 20213
rect 28799 20195 28820 20213
rect 28760 20177 28820 20195
rect 28760 20159 28781 20177
rect 28799 20159 28820 20177
rect 28760 20141 28820 20159
rect 28760 20123 28781 20141
rect 28799 20123 28820 20141
rect 28760 20105 28820 20123
rect 28760 20087 28781 20105
rect 28799 20087 28820 20105
rect 28760 20060 28820 20087
rect 28640 19435 28661 19453
rect 28679 19435 28700 19453
rect 28640 19417 28700 19435
rect 28640 19399 28661 19417
rect 28679 19399 28700 19417
rect 28640 19381 28700 19399
rect 28640 19363 28661 19381
rect 28679 19363 28700 19381
rect 28640 19345 28700 19363
rect 28640 19327 28661 19345
rect 28679 19327 28700 19345
rect 28640 19300 28700 19327
rect 28520 16635 28541 16653
rect 28559 16635 28580 16653
rect 28520 16617 28580 16635
rect 28520 16599 28541 16617
rect 28559 16599 28580 16617
rect 28520 16581 28580 16599
rect 28520 16563 28541 16581
rect 28559 16563 28580 16581
rect 28520 16545 28580 16563
rect 28520 16527 28541 16545
rect 28559 16527 28580 16545
rect 28520 16500 28580 16527
rect 9080 16401 9140 16420
rect 9080 16383 9101 16401
rect 9119 16383 9140 16401
rect 9420 16400 9840 16480
rect 9080 16365 9140 16383
rect 9080 16347 9101 16365
rect 9119 16347 9140 16365
rect 9080 16329 9140 16347
rect 9080 16311 9101 16329
rect 9119 16311 9140 16329
rect 9080 16300 9140 16311
rect 9080 16293 9840 16300
rect 9080 16275 9101 16293
rect 9119 16275 9840 16293
rect 9080 16257 9840 16275
rect 9080 16239 9101 16257
rect 9119 16239 9840 16257
rect 9080 16220 9840 16239
rect 28500 13820 28720 13880
rect 9060 13293 9120 13320
rect 9060 13275 9081 13293
rect 9099 13275 9120 13293
rect 9060 13257 9120 13275
rect 9060 13239 9081 13257
rect 9099 13239 9120 13257
rect 9060 13221 9120 13239
rect 9060 13203 9081 13221
rect 9099 13220 9120 13221
rect 9099 13203 9840 13220
rect 9060 13185 9840 13203
rect 9060 13167 9081 13185
rect 9099 13167 9840 13185
rect 9060 13140 9840 13167
rect 28420 12380 28600 12440
rect 28540 11143 28600 12380
rect 28660 12103 28720 13820
rect 28660 12085 28681 12103
rect 28699 12085 28720 12103
rect 28660 12067 28720 12085
rect 28660 12049 28681 12067
rect 28699 12049 28720 12067
rect 28660 12031 28720 12049
rect 28660 12013 28681 12031
rect 28699 12013 28720 12031
rect 28660 11995 28720 12013
rect 28660 11977 28681 11995
rect 28699 11977 28720 11995
rect 28660 11960 28720 11977
rect 28540 11125 28561 11143
rect 28579 11125 28600 11143
rect 28540 11107 28600 11125
rect 28540 11089 28561 11107
rect 28579 11089 28600 11107
rect 28540 11071 28600 11089
rect 28540 11053 28561 11071
rect 28579 11053 28600 11071
rect 28540 11035 28600 11053
rect 28540 11017 28561 11035
rect 28579 11017 28600 11035
rect 28540 11000 28600 11017
rect 9800 9579 12900 9600
rect 9800 9561 9827 9579
rect 9845 9561 9863 9579
rect 9881 9561 9899 9579
rect 9917 9561 9935 9579
rect 9953 9561 12747 9579
rect 12765 9561 12783 9579
rect 12801 9561 12819 9579
rect 12837 9561 12855 9579
rect 12873 9561 12900 9579
rect 9800 9540 12900 9561
rect 15460 9579 18660 9600
rect 15460 9561 15487 9579
rect 15505 9561 15523 9579
rect 15541 9561 15559 9579
rect 15577 9561 15595 9579
rect 15613 9561 18507 9579
rect 18525 9561 18543 9579
rect 18561 9561 18579 9579
rect 18597 9561 18615 9579
rect 18633 9561 18660 9579
rect 15460 9540 18660 9561
rect 20920 9579 23940 9600
rect 20920 9561 20947 9579
rect 20965 9561 20983 9579
rect 21001 9561 21019 9579
rect 21037 9561 21055 9579
rect 21073 9561 23797 9579
rect 23815 9561 23833 9579
rect 23851 9561 23869 9579
rect 23887 9561 23905 9579
rect 23923 9561 23940 9579
rect 20920 9540 23940 9561
rect 12500 9459 12680 9480
rect 12500 9441 12527 9459
rect 12545 9441 12563 9459
rect 12581 9441 12599 9459
rect 12617 9441 12635 9459
rect 12653 9441 12680 9459
rect 12500 9420 12680 9441
rect 15380 9459 18460 9480
rect 15380 9441 15407 9459
rect 15425 9441 15443 9459
rect 15461 9441 15479 9459
rect 15497 9441 15515 9459
rect 15533 9441 18307 9459
rect 18325 9441 18343 9459
rect 18361 9441 18379 9459
rect 18397 9441 18415 9459
rect 18433 9441 18460 9459
rect 15380 9420 18460 9441
rect 21160 9459 23580 9480
rect 21160 9441 21187 9459
rect 21205 9441 21223 9459
rect 21241 9441 21259 9459
rect 21277 9441 21295 9459
rect 21313 9441 23427 9459
rect 23445 9441 23463 9459
rect 23481 9441 23499 9459
rect 23517 9441 23535 9459
rect 23553 9441 23580 9459
rect 21160 9420 23580 9441
rect 28540 9373 28600 9400
rect 15200 9339 15380 9360
rect 15200 9321 15227 9339
rect 15245 9321 15263 9339
rect 15281 9321 15299 9339
rect 15317 9321 15335 9339
rect 15353 9321 15380 9339
rect 15200 9300 15380 9321
rect 18080 9339 18260 9360
rect 18080 9321 18107 9339
rect 18125 9321 18143 9339
rect 18161 9321 18179 9339
rect 18197 9321 18215 9339
rect 18233 9321 18260 9339
rect 18080 9300 18260 9321
rect 20980 9339 23760 9360
rect 20980 9321 21007 9339
rect 21025 9321 21043 9339
rect 21061 9321 21079 9339
rect 21097 9321 21115 9339
rect 21133 9321 23607 9339
rect 23625 9321 23643 9339
rect 23661 9321 23679 9339
rect 23697 9321 23715 9339
rect 23733 9321 23760 9339
rect 20980 9300 23760 9321
rect 28540 9355 28561 9373
rect 28579 9355 28600 9373
rect 28540 9337 28600 9355
rect 28540 9320 28561 9337
rect 28160 9319 28561 9320
rect 28579 9319 28600 9337
rect 28160 9301 28600 9319
rect 28160 9297 28561 9301
rect 28160 9279 28187 9297
rect 28205 9279 28223 9297
rect 28241 9279 28259 9297
rect 28277 9279 28295 9297
rect 28313 9283 28561 9297
rect 28579 9283 28600 9301
rect 28313 9279 28600 9283
rect 28160 9265 28600 9279
rect 28160 9261 28561 9265
rect 28160 9243 28187 9261
rect 28205 9243 28223 9261
rect 28241 9243 28259 9261
rect 28277 9243 28295 9261
rect 28313 9247 28561 9261
rect 28579 9247 28600 9265
rect 28313 9243 28600 9247
rect 17900 9219 18080 9240
rect 17900 9201 17927 9219
rect 17945 9201 17963 9219
rect 17981 9201 17999 9219
rect 18017 9201 18035 9219
rect 18053 9201 18080 9219
rect 17900 9180 18080 9201
rect 20780 9219 24040 9240
rect 28160 9220 28600 9243
rect 20780 9201 20807 9219
rect 20825 9201 20843 9219
rect 20861 9201 20879 9219
rect 20897 9201 20915 9219
rect 20933 9201 23887 9219
rect 23905 9201 23923 9219
rect 23941 9201 23959 9219
rect 23977 9201 23995 9219
rect 24013 9201 24040 9219
rect 20780 9180 24040 9201
rect 20600 9099 20780 9120
rect 20600 9081 20627 9099
rect 20645 9081 20663 9099
rect 20681 9081 20699 9099
rect 20717 9081 20735 9099
rect 20753 9081 20780 9099
rect 20600 9060 20780 9081
rect 23060 9099 26460 9120
rect 23060 9081 23087 9099
rect 23105 9081 23123 9099
rect 23141 9081 23159 9099
rect 23177 9081 23195 9099
rect 23213 9081 26307 9099
rect 26325 9081 26343 9099
rect 26361 9081 26379 9099
rect 26397 9081 26415 9099
rect 26433 9081 26460 9099
rect 23060 9060 26460 9081
rect 24720 8979 24900 9000
rect 24720 8961 24747 8979
rect 24765 8961 24783 8979
rect 24801 8961 24819 8979
rect 24837 8961 24855 8979
rect 24873 8961 24900 8979
rect 24720 8940 24900 8961
rect 27140 8979 27320 9000
rect 27140 8961 27167 8979
rect 27185 8961 27203 8979
rect 27221 8961 27239 8979
rect 27257 8961 27275 8979
rect 27293 8961 27320 8979
rect 27140 8940 27320 8961
<< end >>
