magic
tech scmos
magscale 1 2
timestamp 1727495947
<< nwell >>
rect -6 154 106 272
<< ntransistor >>
rect 20 14 24 34
rect 40 14 44 34
rect 60 14 64 34
<< ptransistor >>
rect 20 166 24 246
rect 30 166 34 246
rect 54 206 58 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 46 34
rect 58 14 60 34
rect 64 14 66 34
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 30 246
rect 34 166 36 246
rect 48 206 54 246
rect 58 206 60 246
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
rect 46 14 58 34
rect 66 14 78 34
<< pdcontact >>
rect 6 166 18 246
rect 36 166 48 246
rect 60 206 72 246
<< psubstratepcontact >>
rect 0 -6 100 6
<< nsubstratencontact >>
rect 0 254 100 266
<< polysilicon >>
rect 20 246 24 250
rect 30 246 34 250
rect 54 246 58 250
rect 20 142 24 166
rect 12 138 24 142
rect 30 142 34 166
rect 54 160 58 206
rect 30 138 40 142
rect 12 109 16 138
rect 12 45 16 97
rect 36 45 40 138
rect 12 40 24 45
rect 36 40 44 45
rect 20 34 24 40
rect 40 34 44 40
rect 60 34 64 44
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 52 148 64 160
rect 4 97 16 109
rect 24 91 36 103
rect 52 44 64 56
<< metal1 >>
rect 0 266 100 268
rect 0 252 100 254
rect 36 246 48 252
rect 62 200 76 206
rect 6 160 18 166
rect 6 154 52 160
rect 51 148 52 154
rect 51 56 57 148
rect 70 117 76 200
rect 51 50 52 56
rect 28 44 52 50
rect 28 34 34 44
rect 70 34 76 103
rect 6 8 18 14
rect 46 8 58 14
rect 0 6 100 8
rect 0 -8 100 -6
<< m2contact >>
rect 23 103 37 117
rect 3 83 17 97
rect 63 103 77 117
<< metal2 >>
rect 23 117 37 137
rect 63 83 77 103
rect 3 63 17 83
<< m2p >>
rect 23 123 37 137
rect 63 83 77 97
rect 3 63 17 77
<< labels >>
rlabel metal2 3 63 17 77 0 A
port 0 nsew signal input
rlabel metal2 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal2 63 83 77 97 0 Y
port 2 nsew signal output
rlabel metal1 0 266 100 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 254 100 266 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 252 100 254 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 6 100 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -6 100 6 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -8 100 -6 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
