/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module fir_pe(
    inout vdd,
    inout gnd,
    input [5:0] Cin,
    input Rdy,
    output Vld,
    input [3:0] Xin,
    output [3:0] Xout,
    input [3:0] Yin,
    output [3:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [4:0] LoadCtl ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [3:0] XinHL ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire [3:0] _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire Cin_1_bF$buf0 ;
wire Cin_1_bF$buf1 ;
wire Cin_1_bF$buf2 ;
wire Cin_1_bF$buf3 ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire LoadCtl_0_bF$buf4 ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [3:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire [3:0] Yin0 ;
wire [3:0] Yin1 ;
wire [3:0] Yin2 ;
wire [3:0] Yin3 ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire [3:0] XinH ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [3:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [3:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire LoadCtl_4_bF$buf0 ;
wire LoadCtl_4_bF$buf1 ;
wire LoadCtl_4_bF$buf2 ;
wire LoadCtl_4_bF$buf3 ;
wire LoadCtl_4_bF$buf4 ;
wire LoadCtl_4_bF$buf5 ;
wire LoadCtl_4_bF$buf6 ;
wire LoadCtl_4_bF$buf7 ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [5:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _470__bF$buf0 ;
wire _470__bF$buf1 ;
wire _470__bF$buf2 ;
wire _470__bF$buf3 ;
wire _470__bF$buf4 ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [3:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire [3:0] _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire [13:0] mul ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire [15:0] rYin ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

NAND2X1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_527_),
    .Y(_529_)
);

OAI21X1 _800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_75_),
    .C(_99_),
    .Y(_2_)
);

INVX1 _1486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[2]),
    .Y(_736_)
);

NOR2X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_341_),
    .Y(_342_)
);

INVX1 _1295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[12]),
    .Y(_565_)
);

NAND2X1 _1389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_645_),
    .Y(_650_)
);

BUFX2 _1601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .Y(Vld)
);

AOI21X1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_208_),
    .C(_207_),
    .Y(_210_)
);

INVX1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .Y(_471_)
);

NOR2X1 _1410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_469_),
    .Y(_669_)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .Y(Cin_1_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .Y(Cin_1_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .Y(Cin_1_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[1]),
    .Y(Cin_1_bF$buf0)
);

AOI21X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_201_),
    .C(_204_),
    .Y(_247_)
);

OAI21X1 _1504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .C(Yin1[1]),
    .Y(_747_)
);

OAI21X1 _835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_121_),
    .C(_122_),
    .Y(_14_)
);

OR2X2 _1313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_577_),
    .Y(_582_)
);

DFFPOSX1 _1542_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .CLK(clk_bF$buf2),
    .Q(rYin[12])
);

AOI21X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_392_),
    .C(_348_),
    .Y(_397_)
);

INVX1 _873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .Y(_153_)
);

AOI21X1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_171_),
    .C(_165_),
    .Y(_207_)
);

OAI21X1 _1351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf4),
    .B(_614_),
    .C(_615_),
    .Y(_37_)
);

OAI21X1 _1407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(_664_),
    .C(_653_),
    .Y(_42_)
);

DFFPOSX1 _1580_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_54_),
    .CLK(clk_bF$buf5),
    .Q(Yin2[0])
);

NAND2X1 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[2]),
    .Y(_434_)
);

OAI21X1 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_434_),
    .C(_488_),
    .Y(_489_)
);

OAI21X1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_239_),
    .C(_211_),
    .Y(_244_)
);

OR2X2 _1445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_698_),
    .Y(_701_)
);

NOR2X1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_251_),
    .Y(_301_)
);

AOI22X1 _776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(y[2]),
    .C(_75_),
    .D(y[6]),
    .Y(_84_)
);

OAI21X1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_525_),
    .C(_524_),
    .Y(_526_)
);

INVX1 _1483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[1]),
    .Y(_734_)
);

AOI21X1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_330_),
    .C(_287_),
    .Y(_339_)
);

DFFPOSX1 _1539_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .CLK(clk_bF$buf5),
    .Q(rYin[9])
);

NAND3X1 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_385_),
    .C(_388_),
    .Y(_394_)
);

NAND2X1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_562_),
    .Y(_563_)
);

NAND3X1 _1348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_612_),
    .C(_610_),
    .Y(_613_)
);

DFFPOSX1 _1577_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_51_),
    .CLK(clk_bF$buf6),
    .Q(Yin3[1])
);

AND2X2 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_1_bF$buf0),
    .Y(_431_)
);

NOR2X1 _1386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_345_),
    .Y(_647_)
);

OAI22X1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(LoadCtl_4_bF$buf6),
    .C(_466_),
    .D(_468_),
    .Y(_28_)
);

INVX1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .Y(_560_)
);

INVX1 _1501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .Y(_745_)
);

OAI21X1 _832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_119_),
    .C(_120_),
    .Y(_13_)
);

INVX1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .Y(_373_)
);

OAI21X1 _1310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_572_),
    .C(LoadCtl_4_bF$buf5),
    .Y(_580_)
);

INVX1 _870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .Y(_150_)
);

NOR2X1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_203_),
    .Y(_204_)
);

NOR2X1 _1404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_660_),
    .Y(_664_)
);

OAI21X1 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_480_),
    .C(_483_),
    .Y(_486_)
);

NAND3X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_238_),
    .C(_240_),
    .Y(_241_)
);

NAND2X1 _1442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_697_),
    .Y(_698_)
);

OAI21X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_239_),
    .C(_285_),
    .Y(_298_)
);

OAI21X1 _773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_80_),
    .C(_81_),
    .Y(_759_[1])
);

OAI21X1 _829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_117_),
    .C(_118_),
    .Y(_12_)
);

NAND2X1 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[3]),
    .Y(_523_)
);

NAND2X1 _1307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(_574_),
    .Y(_577_)
);

NAND3X1 _1480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[3]),
    .B(_71_),
    .C(_72_),
    .Y(_732_)
);

INVX1 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .Y(_336_)
);

DFFPOSX1 _1536_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .CLK(clk_bF$buf3),
    .Q(rYin[6])
);

OAI21X1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_391_)
);

NOR2X1 _867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_146_),
    .Y(_147_)
);

INVX1 _1345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .Y(_610_)
);

DFFPOSX1 _1574_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_48_),
    .CLK(clk_bF$buf1),
    .Q(y[14])
);

NOR2X1 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_427_),
    .Y(_428_)
);

INVX1 _1383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_639_),
    .Y(_644_)
);

AOI21X1 _1439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .B(_680_),
    .C(_689_),
    .Y(_695_)
);

NAND3X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_292_),
    .C(_294_),
    .Y(_295_)
);

NOR2X1 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .B(_413_),
    .Y(_466_)
);

INVX1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_519_),
    .Y(_520_)
);

NAND2X1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_275_),
    .Y(_276_)
);

NAND2X1 _1477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .B(_729_),
    .Y(_730_)
);

OAI21X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .C(_289_),
    .Y(_333_)
);

NOR2X1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .B(_556_),
    .Y(_557_)
);

INVX1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .Y(_370_)
);

FILL FILL71250x7350 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .Y(_201_)
);

OAI21X1 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_462_),
    .C(_460_),
    .Y(_463_)
);

NOR2X1 _1401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[8]),
    .B(mul[8]),
    .Y(_661_)
);

FILL FILL71250x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_239_),
    .C(_427_),
    .Y(_483_)
);

FILL FILL70950x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_212_),
    .C(_237_),
    .Y(_238_)
);

NAND2X1 _770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_78_),
    .Y(_79_)
);

OAI21X1 _826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(_115_),
    .C(_116_),
    .Y(_11_)
);

NAND3X1 _1304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_552_),
    .C(_573_),
    .Y(_574_)
);

DFFPOSX1 _1533_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .CLK(clk_bF$buf0),
    .Q(rYin[3])
);

AOI21X1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_323_),
    .C(_387_),
    .Y(_388_)
);

INVX1 _864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[2]),
    .Y(_144_)
);

NOR2X1 _1342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[3]),
    .B(mul[3]),
    .Y(_607_)
);

DFFPOSX1 _1571_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_45_),
    .CLK(clk_bF$buf6),
    .Q(y[11])
);

INVX1 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .Y(_425_)
);

NAND2X1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[4]),
    .Y(_480_)
);

NAND2X1 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[5]),
    .Y(_235_)
);

AND2X2 _1380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_641_),
    .Y(_642_)
);

AOI21X1 _1436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_691_),
    .C(_470__bF$buf3),
    .Y(_693_)
);

OAI21X1 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_212_),
    .C(_291_),
    .Y(_292_)
);

OAI21X1 _767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_73_),
    .C(_76_),
    .Y(_759_[0])
);

AOI21X1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_515_),
    .C(_516_),
    .Y(_517_)
);

NAND3X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_273_)
);

NAND2X1 _1474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[15]),
    .B(_470__bF$buf0),
    .Y(_727_)
);

OAI21X1 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .C(_327_),
    .Y(_330_)
);

OR2X2 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_553_),
    .Y(_554_)
);

NAND2X1 _1339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[2]),
    .B(_470__bF$buf2),
    .Y(_605_)
);

OAI21X1 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_141_),
    .C(_366_),
    .Y(_367_)
);

DFFPOSX1 _1568_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_42_),
    .CLK(clk_bF$buf6),
    .Q(y[8])
);

AND2X2 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_422_)
);

INVX2 _899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .Y(_178_)
);

NOR2X1 _1377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_282_),
    .Y(_639_)
);

AOI22X1 _920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_0_bF$buf0),
    .C(XinHL[3]),
    .D(Cin_1_bF$buf1),
    .Y(_198_)
);

INVX1 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .Y(_460_)
);

FILL FILL70950x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf6),
    .B(_113_),
    .C(_114_),
    .Y(_10_)
);

AOI22X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_310_),
    .C(_312_),
    .D(_309_),
    .Y(_364_)
);

OAI21X1 _1301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_568_),
    .C(_570_),
    .Y(_571_)
);

DFFPOSX1 _1530_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .CLK(clk_bF$buf2),
    .Q(rYin[0])
);

NAND3X1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_382_),
    .C(_384_),
    .Y(_385_)
);

OAI21X1 _861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_141_),
    .C(_137_),
    .Y(_142_)
);

OAI21X1 _917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_166_),
    .C(_170_),
    .Y(_195_)
);

NAND2X1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_439_),
    .Y(_477_)
);

NAND2X1 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_184_),
    .Y(_232_)
);

NOR2X1 _1433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_689_),
    .Y(_690_)
);

AOI21X1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_266_),
    .C(_288_),
    .Y(_289_)
);

INVX2 _764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[1]),
    .Y(_74_)
);

NAND2X1 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(_512_),
    .Y(_514_)
);

NAND2X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .Y(_270_)
);

AOI21X1 _1471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_720_),
    .C(_724_),
    .Y(_725_)
);

OAI21X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_326_),
    .C(_265_),
    .Y(_327_)
);

DFFPOSX1 _1527_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1_),
    .CLK(clk_bF$buf7),
    .Q(XinH[1])
);

AND2X2 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_357_),
    .B(_362_),
    .Y(_382_)
);

INVX1 _858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .Y(_139_)
);

NOR2X1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_420_),
    .Y(_551_)
);

NAND2X1 _1336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_598_),
    .Y(_602_)
);

DFFPOSX1 _1565_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_39_),
    .CLK(clk_bF$buf4),
    .Q(y[5])
);

AOI21X1 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_384_),
    .C(_418_),
    .Y(_419_)
);

AOI21X1 _896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_171_),
    .C(_168_),
    .Y(_175_)
);

AND2X2 _1374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_629_),
    .Y(_636_)
);

OAI21X1 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_452_),
    .C(_419_),
    .Y(_457_)
);

NAND2X1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_502_),
    .Y(_511_)
);

OAI21X1 _1468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_706_),
    .C(_719_),
    .Y(_722_)
);

NAND3X1 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_321_),
    .C(_323_),
    .Y(_324_)
);

NAND2X1 _799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[2]),
    .B(_75_),
    .Y(_99_)
);

AOI21X1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_519_),
    .B(_531_),
    .C(_530_),
    .Y(_548_)
);

OAI21X1 _820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_111_),
    .C(_112_),
    .Y(_9_)
);

OAI21X1 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_212_),
    .C(_360_),
    .Y(_361_)
);

INVX1 _914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .Y(_192_)
);

FILL FILL71250x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL70950x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_473_),
    .C(_456_),
    .Y(_474_)
);

OAI22X1 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(LoadCtl_4_bF$buf7),
    .C(_227_),
    .D(_229_),
    .Y(_24_)
);

NOR2X1 _1430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_687_)
);

OAI21X1 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .B(_285_),
    .C(_245_),
    .Y(_286_)
);

INVX1 _761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .Y(_71_)
);

OAI21X1 _817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .B(_109_),
    .C(_110_),
    .Y(_8_)
);

NAND3X1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_264_),
    .C(_266_),
    .Y(_267_)
);

NAND2X1 _1524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(Xin[3]),
    .Y(_757_)
);

AOI21X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_368_),
    .C(_365_),
    .Y(_379_)
);

NAND2X1 _855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin_1_bF$buf3),
    .Y(_136_)
);

NOR2X1 _1333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[2]),
    .B(mul[2]),
    .Y(_599_)
);

DFFPOSX1 _1562_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .CLK(clk_bF$buf2),
    .Q(y[2])
);

NAND2X1 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(_362_),
    .Y(_416_)
);

NAND3X1 _893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_171_),
    .C(_170_),
    .Y(_172_)
);

AOI21X1 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_226_),
    .C(_192_),
    .Y(_227_)
);

NAND2X1 _1371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[6]),
    .B(_470__bF$buf1),
    .Y(_633_)
);

OAI21X1 _1427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_683_),
    .C(_674_),
    .Y(_44_)
);

AOI21X1 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_283_)
);

OAI21X1 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_452_),
    .C(_451_),
    .Y(_454_)
);

AOI21X1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_507_),
    .C(_470__bF$buf1),
    .Y(_509_)
);

AND2X2 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_245_),
    .Y(_264_)
);

AOI21X1 _1465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_703_),
    .C(_713_),
    .Y(_719_)
);

AND2X2 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_299_),
    .Y(_321_)
);

OAI21X1 _796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_75_),
    .C(_97_),
    .Y(_0_)
);

NAND3X1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf6),
    .B(_540_),
    .C(_545_),
    .Y(_546_)
);

INVX1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .Y(_358_)
);

DFFPOSX1 _1559_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .CLK(clk_bF$buf4),
    .Q(mul[13])
);

OAI21X1 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_346_),
    .C(_412_),
    .Y(_413_)
);

NOR2X1 _1368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(_626_),
    .Y(_631_)
);

NAND2X1 _911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf7),
    .B(_189_),
    .Y(_190_)
);

DFFPOSX1 _1597_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl_0_bF$buf1),
    .CLK(clk_bF$buf6),
    .Q(LoadCtl[1])
);

OAI21X1 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_450_),
    .C(_383_),
    .Y(_451_)
);

OAI21X1 _814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .B(_107_),
    .C(_108_),
    .Y(_7_)
);

OAI21X1 _1521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_236_),
    .C(_755_),
    .Y(_67_)
);

AOI22X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_1_bF$buf2),
    .C(XinH[2]),
    .D(Cin_0_bF$buf3),
    .Y(_376_)
);

NAND3X1 _852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin_0_bF$buf1),
    .C(LoadCtl_4_bF$buf7),
    .Y(_134_)
);

FILL FILL71250x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_185_),
    .C(_186_),
    .Y(_187_)
);

NAND2X1 _1330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[1]),
    .B(_470__bF$buf0),
    .Y(_597_)
);

AND2X2 _890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf0),
    .Y(_169_)
);

AOI21X1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_218_),
    .C(_219_),
    .Y(_224_)
);

INVX1 _1424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .Y(_682_)
);

NAND3X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(_280_),
    .C(_278_),
    .Y(_281_)
);

AOI22X1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_505_),
    .C(_458_),
    .D(_456_),
    .Y(_506_)
);

AOI21X1 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_252_),
    .C(_248_),
    .Y(_261_)
);

AOI21X1 _1462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_715_),
    .C(_470__bF$buf0),
    .Y(_717_)
);

AOI21X1 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .B(_307_),
    .C(_303_),
    .Y(_318_)
);

NAND2X1 _793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(XinHL[3]),
    .Y(_96_)
);

NAND2X1 _1518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[0]),
    .Y(_754_)
);

NAND2X1 _849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(Yin3[3]),
    .Y(_132_)
);

AOI21X1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_412_),
    .C(_542_),
    .Y(_543_)
);

NAND2X1 _1327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_593_),
    .Y(_594_)
);

AND2X2 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[4]),
    .Y(_355_)
);

DFFPOSX1 _1556_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .CLK(clk_bF$buf3),
    .Q(mul[10])
);

INVX1 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[8]),
    .Y(_410_)
);

AOI22X1 _887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin_1_bF$buf3),
    .C(XinHL[3]),
    .D(Cin_0_bF$buf0),
    .Y(_166_)
);

NOR2X1 _1365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_230_),
    .Y(_628_)
);

DFFPOSX1 _1594_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_68_),
    .CLK(clk_bF$buf7),
    .Q(XinHL[2])
);

NAND2X1 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_447_),
    .Y(_448_)
);

NOR2X1 _1459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_713_),
    .Y(_714_)
);

AOI22X1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .C(XinH[1]),
    .D(Cin_0_bF$buf2),
    .Y(_315_)
);

NAND2X1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_517_),
    .Y(_540_)
);

OAI21X1 _811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_105_),
    .C(_106_),
    .Y(_6_)
);

NOR2X1 _1497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[2]),
    .B(_740_),
    .Y(_743_)
);

NAND2X1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[5]),
    .Y(_352_)
);

INVX1 _905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .Y(_184_)
);

FILL FILL70950x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_194_),
    .C(_216_),
    .Y(_221_)
);

NOR2X1 _1421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[10]),
    .B(mul[10]),
    .Y(_679_)
);

OR2X2 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_276_),
    .Y(_278_)
);

OAI21X1 _808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_103_),
    .C(_104_),
    .Y(_5_)
);

AOI21X1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_502_),
    .C(_474_),
    .Y(_503_)
);

NAND3X1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(_257_),
    .C(_247_),
    .Y(_258_)
);

NAND2X1 _790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(XinHL[2]),
    .Y(_94_)
);

AOI21X1 _1515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_736_),
    .C(_752_),
    .Y(_64_)
);

NAND2X1 _846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(Yin3[2]),
    .Y(_130_)
);

NOR2X1 _1324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(_135_),
    .Y(_591_)
);

DFFPOSX1 _1553_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .CLK(clk_bF$buf4),
    .Q(mul[7])
);

NOR2X1 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_403_),
    .Y(_408_)
);

NAND2X1 _884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[2]),
    .Y(_163_)
);

BUFX2 _1609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_[3]),
    .Y(Yout[3])
);

INVX1 _1362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[5]),
    .Y(_625_)
);

OAI21X1 _1418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[9]),
    .B(mul[9]),
    .C(_662_),
    .Y(_676_)
);

DFFPOSX1 _1591_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_65_),
    .CLK(clk_bF$buf0),
    .Q(Yin0[3])
);

NAND2X1 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_432_),
    .Y(_445_)
);

NAND3X1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_492_),
    .C(_495_),
    .Y(_500_)
);

NAND2X1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_249_),
    .Y(_255_)
);

OAI21X1 _1456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_706_),
    .C(_710_),
    .Y(_711_)
);

OAI21X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_141_),
    .C(_306_),
    .Y(_312_)
);

NAND2X1 _787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[1]),
    .Y(_92_)
);

NAND2X1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_535_),
    .Y(_537_)
);

AOI21X1 _1494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_740_),
    .C(_741_),
    .Y(_54_)
);

NAND2X1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_299_),
    .Y(_349_)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf7)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf6)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf5)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf4)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf0)
);

NAND2X1 _1359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_619_),
    .Y(_623_)
);

AOI21X1 _902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_180_),
    .C(_163_),
    .Y(_181_)
);

DFFPOSX1 _1588_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_62_),
    .CLK(clk_bF$buf1),
    .Q(Yin0[0])
);

NOR2X1 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_439_),
    .Y(_442_)
);

AOI21X1 _1397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(_656_),
    .C(_655_),
    .Y(_657_)
);

NAND3X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_202_),
    .C(_205_),
    .Y(_218_)
);

OAI21X1 _805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_101_),
    .C(_102_),
    .Y(_4_)
);

NOR2X1 _1512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(Yin0[1]),
    .Y(_751_)
);

NAND2X1 _843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(Yin3[1]),
    .Y(_128_)
);

NAND2X1 _1321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_587_),
    .Y(_589_)
);

DFFPOSX1 _1550_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .CLK(clk_bF$buf0),
    .Q(mul[4])
);

NAND3X1 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_399_),
    .C(_404_),
    .Y(_405_)
);

INVX1 _881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[3]),
    .Y(_160_)
);

BUFX2 _1606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_[0]),
    .Y(Yout[0])
);

OAI21X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_211_),
    .C(_214_),
    .Y(_215_)
);

OAI21X1 _1415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(LoadCtl_4_bF$buf2),
    .C(_673_),
    .Y(_43_)
);

INVX1 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .Y(_497_)
);

NAND2X1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_196_),
    .Y(_252_)
);

OAI21X1 _1453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_705_),
    .C(_694_),
    .Y(_46_)
);

INVX1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .Y(_309_)
);

NAND2X1 _784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[0]),
    .Y(_90_)
);

OAI21X1 _1509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_745_),
    .C(_749_),
    .Y(_61_)
);

INVX1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .Y(_534_)
);

NOR2X1 _1318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_133_),
    .Y(_586_)
);

OAI21X1 _1491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_732_),
    .C(_739_),
    .Y(_53_)
);

NAND3X1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_279_),
    .C(_340_),
    .Y(_346_)
);

DFFPOSX1 _1547_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .CLK(clk_bF$buf2),
    .Q(mul[1])
);

AOI21X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_335_),
    .C(_401_),
    .Y(_402_)
);

NOR2X1 _878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_156_),
    .Y(_158_)
);

INVX1 _1356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .Y(_620_)
);

DFFPOSX1 _1585_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_59_),
    .CLK(clk_bF$buf4),
    .Q(Yin1[1])
);

OAI21X1 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_372_),
    .C(_371_),
    .Y(_439_)
);

INVX1 _1394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .Y(_654_)
);

NAND3X1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_492_),
    .C(_529_),
    .Y(_531_)
);

OAI21X1 _802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_75_),
    .C(_100_),
    .Y(_3_)
);

OAI21X1 _1488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_732_),
    .C(_737_),
    .Y(_52_)
);

OAI21X1 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_343_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_344_)
);

NOR2X1 _1297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_542_),
    .Y(_567_)
);

NAND2X1 _840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(Yin3[0]),
    .Y(_126_)
);

BUFX2 _1603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_[1]),
    .Y(Xout[1])
);

INVX2 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[4]),
    .Y(_212_)
);

AND2X2 _1412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_667_),
    .B(_670_),
    .Y(_671_)
);

NAND2X1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_432_),
    .Y(_494_)
);

AND2X2 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf2),
    .Y(_249_)
);

NOR2X1 _1450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_700_),
    .Y(_706_)
);

NAND2X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .Y(_306_)
);

AOI22X1 _781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(y[3]),
    .C(_75_),
    .D(y[7]),
    .Y(_88_)
);

OAI21X1 _1506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_74_),
    .C(Yin1[2]),
    .Y(_748_)
);

NAND2X1 _837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(Yin2[3]),
    .Y(_124_)
);

OAI21X1 _1315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_575_),
    .C(LoadCtl_4_bF$buf6),
    .Y(_584_)
);

DFFPOSX1 _1544_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .CLK(clk_bF$buf2),
    .Q(rYin[14])
);

NAND3X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_386_),
    .C(_391_),
    .Y(_399_)
);

NAND3X1 _875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_154_),
    .C(_149_),
    .Y(_155_)
);

NOR2X1 _1353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[4]),
    .B(mul[4]),
    .Y(_617_)
);

NOR2X1 _1409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[9]),
    .B(mul[9]),
    .Y(_668_)
);

DFFPOSX1 _1582_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_56_),
    .CLK(clk_bF$buf5),
    .Q(Yin2[2])
);

INVX1 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .Y(_436_)
);

INVX1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_491_)
);

NAND2X1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_241_),
    .Y(_246_)
);

NAND2X1 _1391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[7]),
    .B(_470__bF$buf3),
    .Y(_652_)
);

NOR2X1 _1447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(_565_),
    .Y(_703_)
);

NAND2X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[2]),
    .Y(_303_)
);

INVX1 _778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[11]),
    .Y(_85_)
);

OAI21X1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_420_),
    .C(_526_),
    .Y(_528_)
);

OAI21X1 _1485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_732_),
    .C(_735_),
    .Y(_51_)
);

AND2X2 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_335_),
    .Y(_341_)
);

NAND2X1 _1294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_564_),
    .Y(_31_)
);

DFFPOSX1 _1579_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_53_),
    .CLK(clk_bF$buf1),
    .Q(Yin3[3])
);

NAND2X1 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_1_bF$buf0),
    .Y(_433_)
);

OR2X2 _1388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_648_),
    .Y(_649_)
);

DFFPOSX1 _1600_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[3]),
    .CLK(clk_bF$buf6),
    .Q(LoadCtl[4])
);

OAI21X1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_204_),
    .C(_201_),
    .Y(_209_)
);

INVX8 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .Y(_470_)
);

FILL FILL70650x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_470__bF$buf0)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

OAI21X1 _1503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_745_),
    .C(_746_),
    .Y(_58_)
);

FILL FILL70950x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(Yin2[2]),
    .Y(_122_)
);

INVX1 _1312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[13]),
    .Y(_581_)
);

DFFPOSX1 _1541_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .CLK(clk_bF$buf5),
    .Q(rYin[11])
);

NAND3X1 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_395_),
    .C(_394_),
    .Y(_396_)
);

NAND3X1 _872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf1),
    .C(_151_),
    .Y(_152_)
);

AOI21X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_202_),
    .C(_195_),
    .Y(_206_)
);

NAND2X1 _1350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[3]),
    .B(_470__bF$buf4),
    .Y(_615_)
);

OAI21X1 _1406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_659_),
    .C(LoadCtl_4_bF$buf4),
    .Y(_666_)
);

NAND2X1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_487_),
    .Y(_488_)
);

NAND2X1 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_237_),
    .Y(_243_)
);

NOR2X1 _1444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_659_),
    .Y(_700_)
);

NAND2X1 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_295_),
    .Y(_300_)
);

OAI21X1 _775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(y[10]),
    .C(_72_),
    .Y(_83_)
);

NAND2X1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin[4]),
    .Y(_525_)
);

INVX1 _1309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .Y(_579_)
);

OAI21X1 _1482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_732_),
    .C(_733_),
    .Y(_50_)
);

AOI21X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_332_),
    .C(_286_),
    .Y(_338_)
);

DFFPOSX1 _1538_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .CLK(clk_bF$buf5),
    .Q(rYin[8])
);

INVX1 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .Y(_393_)
);

OAI21X1 _869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_147_),
    .C(_145_),
    .Y(_149_)
);

OAI21X1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_517_),
    .C(_536_),
    .Y(_562_)
);

INVX1 _1347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_608_),
    .Y(_612_)
);

DFFPOSX1 _1576_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_50_),
    .CLK(clk_bF$buf1),
    .Q(Yin3[0])
);

NAND2X1 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(_429_),
    .Y(_430_)
);

NOR2X1 _1385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[7]),
    .B(mul[7]),
    .Y(_646_)
);

OAI21X1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_467_),
    .C(LoadCtl_4_bF$buf6),
    .Y(_468_)
);

INVX1 _1479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[0]),
    .Y(_731_)
);

NAND3X1 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_284_),
    .C(_331_),
    .Y(_335_)
);

NOR2X1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_558_),
    .Y(_559_)
);

AOI21X1 _1500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_740_),
    .C(_744_),
    .Y(_57_)
);

NAND2X1 _831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(Yin2[1]),
    .Y(_120_)
);

AOI22X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_1_bF$buf0),
    .C(XinH[3]),
    .D(Cin_0_bF$buf3),
    .Y(_372_)
);

NAND2X1 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .Y(_203_)
);

NOR2X1 _1403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_661_),
    .B(_662_),
    .Y(_663_)
);

NAND2X1 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_485_)
);

OAI21X1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_239_),
    .C(_231_),
    .Y(_240_)
);

NAND2X1 _1441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_696_),
    .Y(_697_)
);

NAND2X1 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_291_),
    .Y(_297_)
);

AOI22X1 _772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(y[1]),
    .C(_75_),
    .D(y[5]),
    .Y(_81_)
);

NAND2X1 _828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(Yin2[0]),
    .Y(_118_)
);

NAND2X1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[5]),
    .Y(_522_)
);

OAI21X1 _1306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(_575_),
    .C(_555_),
    .Y(_576_)
);

DFFPOSX1 _1535_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .CLK(clk_bF$buf4),
    .Q(rYin[5])
);

AOI21X1 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_375_),
    .C(_363_),
    .Y(_390_)
);

NAND2X1 _866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin_1_bF$buf3),
    .Y(_146_)
);

FILL FILL71250x36150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_608_),
    .C(_606_),
    .Y(_609_)
);

DFFPOSX1 _1573_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_47_),
    .CLK(clk_bF$buf1),
    .Q(y[13])
);

NAND2X1 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_427_)
);

NAND2X1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(_481_),
    .Y(_482_)
);

OAI21X1 _1382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_642_),
    .C(_633_),
    .Y(_40_)
);

NAND2X1 _1438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[12]),
    .B(_470__bF$buf4),
    .Y(_694_)
);

OAI21X1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_239_),
    .C(_293_),
    .Y(_294_)
);

INVX1 _769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[9]),
    .Y(_78_)
);

INVX1 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .Y(_465_)
);

OAI21X1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_480_),
    .C(_484_),
    .Y(_519_)
);

NAND3X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_273_),
    .C(_274_),
    .Y(_275_)
);

OAI21X1 _1476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_725_),
    .C(_131_),
    .Y(_729_)
);

NAND3X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .C(_327_),
    .Y(_332_)
);

NAND2X1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_554_),
    .Y(_556_)
);

NAND3X1 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_367_),
    .C(_368_),
    .Y(_369_)
);

INVX1 _1379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .Y(_641_)
);

NAND2X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[2]),
    .Y(_200_)
);

AOI21X1 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_449_),
    .C(_417_),
    .Y(_462_)
);

INVX1 _1400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .Y(_660_)
);

AND2X2 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[3]),
    .Y(_237_)
);

NAND2X1 _825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf4),
    .B(Yin1[3]),
    .Y(_116_)
);

INVX1 _1303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .Y(_573_)
);

DFFPOSX1 _1532_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .CLK(clk_bF$buf0),
    .Q(rYin[2])
);

INVX1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .Y(_387_)
);

OAI21X1 _863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(LoadCtl_4_bF$buf3),
    .C(_143_),
    .Y(_21_)
);

NAND2X1 _919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_196_),
    .Y(_197_)
);

AOI21X1 _1341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_601_),
    .C(_600_),
    .Y(_606_)
);

FILL FILL71250x57750 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _1570_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_44_),
    .CLK(clk_bF$buf6),
    .Q(y[10])
);

AOI22X1 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[4]),
    .C(XinH[1]),
    .D(Cin[3]),
    .Y(_424_)
);

FILL FILL70950x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_420_),
    .Y(_479_)
);

AOI21X1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_219_),
    .C(_210_),
    .Y(_234_)
);

OR2X2 _1435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_691_),
    .Y(_692_)
);

AND2X2 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[3]),
    .Y(_291_)
);

AOI22X1 _766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(y[0]),
    .C(_75_),
    .D(y[4]),
    .Y(_76_)
);

OAI21X1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_503_),
    .C(_513_),
    .Y(_516_)
);

NAND3X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_268_),
    .C(_271_),
    .Y(_272_)
);

OAI21X1 _1473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_726_),
    .C(_718_),
    .Y(_48_)
);

AOI21X1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_314_),
    .C(_300_),
    .Y(_329_)
);

DFFPOSX1 _1529_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .CLK(clk_bF$buf7),
    .Q(XinH[3])
);

OAI21X1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_379_),
    .C(_364_),
    .Y(_384_)
);

AND2X2 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_550_),
    .Y(_553_)
);

NAND2X1 _1338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

AND2X2 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .B(Cin_0_bF$buf3),
    .Y(_366_)
);

DFFPOSX1 _1567_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_41_),
    .CLK(clk_bF$buf3),
    .Q(y[7])
);

NOR2X1 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_420_),
    .Y(_421_)
);

OAI21X1 _898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_141_),
    .C(_169_),
    .Y(_177_)
);

NOR2X1 _1376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[6]),
    .B(mul[6]),
    .Y(_638_)
);

NAND3X1 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_458_),
    .C(_455_),
    .Y(_459_)
);

OAI21X1 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_420_),
    .C(_525_),
    .Y(_550_)
);

NAND2X1 _822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf6),
    .B(Yin1[2]),
    .Y(_114_)
);

NAND2X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_357_),
    .Y(_363_)
);

NOR2X1 _1300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_569_),
    .Y(_570_)
);

INVX2 _860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_1_bF$buf2),
    .Y(_141_)
);

OAI21X1 _916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_193_),
    .C(_185_),
    .Y(_194_)
);

INVX1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .Y(_476_)
);

AND2X2 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_231_)
);

INVX1 _1432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .Y(_689_)
);

INVX1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .Y(_288_)
);

OAI21X1 _763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(y[8]),
    .C(_72_),
    .Y(_73_)
);

NAND2X1 _819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf0),
    .B(Yin1[1]),
    .Y(_112_)
);

NAND3X1 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_502_),
    .C(_474_),
    .Y(_513_)
);

OAI21X1 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_206_),
    .C(_218_),
    .Y(_269_)
);

INVX1 _1470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .Y(_724_)
);

AOI21X1 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(_257_),
    .C(_259_),
    .Y(_326_)
);

DFFPOSX1 _1526_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .CLK(clk_bF$buf7),
    .Q(XinH[0])
);

NAND3X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(_375_),
    .C(_380_),
    .Y(_381_)
);

FILL FILL71250x43350 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_137_),
    .Y(_138_)
);

NOR2X1 _1335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_600_),
    .Y(_601_)
);

DFFPOSX1 _1564_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .CLK(clk_bF$buf1),
    .Q(y[4])
);

INVX1 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .Y(_418_)
);

OAI21X1 _895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .B(_148_),
    .C(_152_),
    .Y(_174_)
);

OAI21X1 _1373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_111_),
    .B(_230_),
    .C(_634_),
    .Y(_635_)
);

OAI21X1 _1429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_679_),
    .B(_678_),
    .C(_685_),
    .Y(_686_)
);

NAND2X1 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_285_)
);

NAND3X1 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .B(_443_),
    .C(_448_),
    .Y(_456_)
);

INVX1 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[10]),
    .Y(_510_)
);

OAI21X1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_260_),
    .C(_247_),
    .Y(_266_)
);

INVX1 _1467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .Y(_721_)
);

OAI21X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_318_),
    .C(_302_),
    .Y(_323_)
);

OAI21X1 _798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_75_),
    .C(_98_),
    .Y(_1_)
);

NAND2X1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[11]),
    .B(_470__bF$buf1),
    .Y(_547_)
);

NAND2X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_360_)
);

INVX1 _913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[4]),
    .Y(_191_)
);

DFFPOSX1 _1599_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[2]),
    .CLK(clk_bF$buf6),
    .Q(LoadCtl[3])
);

AOI21X1 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_446_),
    .C(_430_),
    .Y(_453_)
);

AOI21X1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_448_),
    .B(_443_),
    .C(_451_),
    .Y(_473_)
);

NAND2X1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf7),
    .B(_228_),
    .Y(_229_)
);

NOR2X1 _760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[12]),
    .Y(_70_)
);

NAND2X1 _816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .B(Yin1[0]),
    .Y(_110_)
);

OAI21X1 _1523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_176_),
    .C(_756_),
    .Y(_68_)
);

AOI21X1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_373_),
    .C(_370_),
    .Y(_378_)
);

INVX1 _854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[1]),
    .Y(_135_)
);

OAI21X1 _1332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(_135_),
    .C(_594_),
    .Y(_598_)
);

DFFPOSX1 _1561_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .CLK(clk_bF$buf2),
    .Q(y[1])
);

OAI21X1 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_414_),
    .C(_386_),
    .Y(_415_)
);

INVX1 _892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .Y(_171_)
);

OAI21X1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_225_),
    .C(_223_),
    .Y(_226_)
);

OAI21X1 _1370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(LoadCtl_4_bF$buf5),
    .C(_632_),
    .Y(_39_)
);

OAI21X1 _1426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_678_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_684_)
);

INVX1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[6]),
    .Y(_282_)
);

OR2X2 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_507_),
    .Y(_508_)
);

NAND3X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_258_),
    .C(_262_),
    .Y(_263_)
);

NAND2X1 _1464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[14]),
    .B(_470__bF$buf0),
    .Y(_718_)
);

NAND3X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_314_),
    .C(_319_),
    .Y(_320_)
);

NAND2X1 _795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[0]),
    .B(_75_),
    .Y(_97_)
);

OAI21X1 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_543_),
    .C(_544_),
    .Y(_545_)
);

NAND2X1 _1329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .B(_594_),
    .Y(_596_)
);

NAND3X1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_354_),
    .C(_356_),
    .Y(_357_)
);

DFFPOSX1 _1558_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .CLK(clk_bF$buf0),
    .Q(mul[12])
);

NAND2X1 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_411_),
    .Y(_412_)
);

INVX1 _889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .Y(_168_)
);

AND2X2 _1367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_629_),
    .Y(_630_)
);

NAND3X1 _910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_183_),
    .C(_187_),
    .Y(_189_)
);

DFFPOSX1 _1596_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(Rdy),
    .CLK(clk_bF$buf7),
    .Q(LoadCtl[0])
);

AOI21X1 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_374_),
    .C(_377_),
    .Y(_450_)
);

NAND2X1 _813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .B(Yin0[3]),
    .Y(_108_)
);

NOR2X1 _1499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[3]),
    .B(_740_),
    .Y(_744_)
);

OAI21X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_212_),
    .C(_353_),
    .Y(_354_)
);

NAND2X1 _1520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(Xin[1]),
    .Y(_755_)
);

NAND3X1 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_374_),
    .B(_364_),
    .C(_369_),
    .Y(_375_)
);

INVX1 _851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[0]),
    .Y(_133_)
);

OAI21X1 _907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_181_),
    .C(_162_),
    .Y(_186_)
);

AOI21X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_186_),
    .C(_222_),
    .Y(_223_)
);

NOR2X1 _1423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_679_),
    .B(_680_),
    .Y(_681_)
);

INVX1 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .Y(_280_)
);

NAND3X1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_493_),
    .C(_498_),
    .Y(_505_)
);

AOI21X1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_256_),
    .C(_254_),
    .Y(_260_)
);

OR2X2 _1461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_715_),
    .Y(_716_)
);

AOI21X1 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_312_),
    .C(_309_),
    .Y(_317_)
);

INVX2 _792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[3]),
    .Y(_95_)
);

FILL FILL71250x50550 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_738_),
    .C(_753_),
    .Y(_65_)
);

INVX1 _848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[15]),
    .Y(_131_)
);

NAND3X1 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_463_),
    .C(_507_),
    .Y(_542_)
);

FILL FILL70950x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_591_),
    .Y(_593_)
);

DFFPOSX1 _1555_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .CLK(clk_bF$buf5),
    .Q(mul[9])
);

OAI21X1 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(LoadCtl_4_bF$buf0),
    .C(_409_),
    .Y(_27_)
);

NOR2X1 _886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_164_),
    .Y(_165_)
);

NOR2X1 _1364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[5]),
    .B(mul[5]),
    .Y(_627_)
);

DFFPOSX1 _1593_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_67_),
    .CLK(clk_bF$buf7),
    .Q(XinHL[1])
);

NAND2X1 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_445_),
    .Y(_447_)
);

NAND3X1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_501_),
    .C(_500_),
    .Y(_502_)
);

NOR2X1 _1458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(_581_),
    .Y(_713_)
);

NAND3X1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_313_),
    .C(_302_),
    .Y(_314_)
);

INVX2 _789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .Y(_93_)
);

NAND2X1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_538_),
    .Y(_539_)
);

NAND2X1 _810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf5),
    .B(Yin0[2]),
    .Y(_106_)
);

AOI21X1 _1496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_740_),
    .C(_742_),
    .Y(_55_)
);

OAI21X1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_350_),
    .C(_322_),
    .Y(_351_)
);

NAND3X1 _904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_173_),
    .C(_182_),
    .Y(_183_)
);

AND2X2 _1399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

NAND3X1 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_218_),
    .C(_217_),
    .Y(_220_)
);

CLKBUF1 CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

AOI21X1 _1420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_675_),
    .C(_677_),
    .Y(_678_)
);

NAND2X1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_228_),
    .Y(_277_)
);

NAND2X1 _807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(Yin0[1]),
    .Y(_104_)
);

NAND3X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_254_),
    .C(_255_),
    .Y(_257_)
);

NOR2X1 _1514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(Yin0[2]),
    .Y(_752_)
);

INVX1 _845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[14]),
    .Y(_129_)
);

OAI21X1 _1323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf2),
    .B(_589_),
    .C(_590_),
    .Y(_34_)
);

DFFPOSX1 _1552_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .CLK(clk_bF$buf7),
    .Q(mul[6])
);

NAND2X1 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_405_),
    .Y(_407_)
);

AOI21X1 _883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_153_),
    .C(_147_),
    .Y(_162_)
);

BUFX2 _1608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_[2]),
    .Y(Yout[2])
);

NAND3X1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_209_),
    .C(_207_),
    .Y(_217_)
);

OAI21X1 _1361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf4),
    .B(_624_),
    .C(_616_),
    .Y(_38_)
);

AND2X2 _1417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_670_),
    .Y(_675_)
);

DFFPOSX1 _1590_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_64_),
    .CLK(clk_bF$buf3),
    .Q(Yin0[2])
);

AND2X2 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_426_),
    .Y(_444_)
);

NAND3X1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_493_),
    .C(_498_),
    .Y(_499_)
);

INVX1 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .Y(_254_)
);

INVX1 _1455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .Y(_710_)
);

NAND2X1 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_310_),
    .Y(_311_)
);

INVX2 _786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .Y(_91_)
);

NAND3X1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_535_),
    .C(_518_),
    .Y(_536_)
);

NOR2X1 _1493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[0]),
    .B(_740_),
    .Y(_741_)
);

OAI21X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_347_),
    .C(_332_),
    .Y(_348_)
);

DFFPOSX1 _1549_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .CLK(clk_bF$buf0),
    .Q(mul[3])
);

INVX1 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .Y(_404_)
);

NOR2X1 _1358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_618_),
    .Y(_622_)
);

OAI21X1 _901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_179_),
    .C(_151_),
    .Y(_180_)
);

DFFPOSX1 _1587_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_61_),
    .CLK(clk_bF$buf3),
    .Q(Yin1[3])
);

AOI21X1 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_310_),
    .C(_435_),
    .Y(_441_)
);

AND2X2 _1396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_648_),
    .Y(_656_)
);

NAND2X1 _804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin0[0]),
    .B(LoadCtl_4_bF$buf3),
    .Y(_102_)
);

NOR2X1 _1299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_558_),
    .B(_536_),
    .Y(_569_)
);

AOI21X1 _1511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(_731_),
    .C(_750_),
    .Y(_62_)
);

INVX1 _842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[13]),
    .Y(_127_)
);

NAND2X1 _1320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_133_),
    .Y(_588_)
);

OAI21X1 _880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(LoadCtl_4_bF$buf7),
    .C(_159_),
    .Y(_22_)
);

BUFX2 _1605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_[3]),
    .Y(Xout[3])
);

OAI21X1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_212_),
    .C(_213_),
    .Y(_214_)
);

OAI21X1 _1414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_672_),
    .B(_671_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_673_)
);

AOI21X1 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_484_),
    .C(_491_),
    .Y(_496_)
);

NAND2X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_0_bF$buf2),
    .Y(_251_)
);

OAI21X1 _1452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_706_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_708_)
);

NAND3X1 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_307_),
    .C(_305_),
    .Y(_308_)
);

INVX2 _783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .Y(_89_)
);

OAI21X1 _1508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_74_),
    .C(Yin1[3]),
    .Y(_749_)
);

INVX1 _839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[12]),
    .Y(_125_)
);

OAI21X1 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_532_),
    .C(_520_),
    .Y(_533_)
);

AOI22X1 _1317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_470__bF$buf4),
    .C(_582_),
    .D(_585_),
    .Y(_33_)
);

NAND2X1 _1490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[3]),
    .B(_732_),
    .Y(_739_)
);

INVX1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[7]),
    .Y(_345_)
);

DFFPOSX1 _1546_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .CLK(clk_bF$buf0),
    .Q(mul[0])
);

NOR2X1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_400_),
    .Y(_401_)
);

AOI21X1 _877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_154_),
    .C(_138_),
    .Y(_157_)
);

OAI21X1 _1355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_606_),
    .C(_612_),
    .Y(_619_)
);

DFFPOSX1 _1584_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_58_),
    .CLK(clk_bF$buf4),
    .Q(Yin1[0])
);

NOR2X1 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_432_),
    .Y(_438_)
);

NAND2X1 _1393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[8]),
    .B(_470__bF$buf3),
    .Y(_653_)
);

NOR2X1 _1449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .B(_701_),
    .Y(_705_)
);

OAI21X1 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_141_),
    .C(_304_),
    .Y(_305_)
);

AOI21X1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_492_),
    .C(_529_),
    .Y(_530_)
);

NAND2X1 _801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[3]),
    .B(_75_),
    .Y(_100_)
);

NAND2X1 _1487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[2]),
    .B(_732_),
    .Y(_737_)
);

INVX1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .Y(_343_)
);

NAND3X1 _1296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_538_),
    .C(_559_),
    .Y(_566_)
);

BUFX2 _1602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_[0]),
    .Y(Xout[0])
);

NAND2X1 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_211_)
);

AOI21X1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_465_),
    .C(_471_),
    .Y(_472_)
);

NOR2X1 _1411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(_669_),
    .Y(_670_)
);

NAND3X1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(_492_),
    .C(_489_),
    .Y(_493_)
);

NAND2X1 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin[2]),
    .Y(_248_)
);

OAI21X1 _780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[15]),
    .C(_86_),
    .Y(_87_)
);

OAI21X1 _1505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_745_),
    .C(_747_),
    .Y(_59_)
);

INVX1 _836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[11]),
    .Y(_123_)
);

INVX1 _1314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .Y(_583_)
);

DFFPOSX1 _1543_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .CLK(clk_bF$buf1),
    .Q(rYin[13])
);

NAND3X1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_395_),
    .C(_394_),
    .Y(_398_)
);

FILL FILL70650x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_153_),
    .C(_152_),
    .Y(_154_)
);

NAND2X1 _1352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[4]),
    .B(_470__bF$buf3),
    .Y(_616_)
);

AOI21X1 _1408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_663_),
    .C(_662_),
    .Y(_667_)
);

DFFPOSX1 _1581_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_55_),
    .CLK(clk_bF$buf5),
    .Q(Yin2[1])
);

AOI22X1 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin[2]),
    .C(XinH[3]),
    .D(Cin_1_bF$buf0),
    .Y(_435_)
);

FILL FILL71250x10950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_141_),
    .C(_440_),
    .Y(_490_)
);

NAND3X1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_242_),
    .C(_243_),
    .Y(_245_)
);

NAND2X1 _1390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_649_),
    .Y(_651_)
);

NOR2X1 _1446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[12]),
    .B(mul[12]),
    .Y(_702_)
);

AOI21X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_256_),
    .C(_301_),
    .Y(_302_)
);

OAI21X1 _777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_83_),
    .C(_84_),
    .Y(_759_[2])
);

OR2X2 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(_522_),
    .Y(_527_)
);

NAND2X1 _1484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[1]),
    .B(_732_),
    .Y(_735_)
);

OAI21X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_339_),
    .C(_337_),
    .Y(_340_)
);

NAND3X1 _1293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf6),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

NAND2X1 _1349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .B(_613_),
    .Y(_614_)
);

DFFPOSX1 _1578_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_52_),
    .CLK(clk_bF$buf6),
    .Q(Yin3[2])
);

AOI22X1 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_431_),
    .C(_373_),
    .D(_370_),
    .Y(_432_)
);

NOR2X1 _1387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .B(_647_),
    .Y(_648_)
);

NAND3X1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_199_),
    .C(_197_),
    .Y(_208_)
);

INVX1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[9]),
    .Y(_469_)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_470__bF$buf4)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_470__bF$buf3)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_470__bF$buf2)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_470__bF$buf1)
);

OAI21X1 _1502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .C(Yin1[0]),
    .Y(_746_)
);

INVX1 _833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[10]),
    .Y(_121_)
);

NAND3X1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_373_),
    .C(_371_),
    .Y(_374_)
);

OAI22X1 _1311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(LoadCtl_4_bF$buf5),
    .C(_580_),
    .D(_579_),
    .Y(_32_)
);

DFFPOSX1 _1540_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .CLK(clk_bF$buf3),
    .Q(rYin[10])
);

OAI21X1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .C(_351_),
    .Y(_395_)
);

AND2X2 _871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin_1_bF$buf3),
    .Y(_151_)
);

OAI21X1 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_204_),
    .C(_200_),
    .Y(_205_)
);

INVX1 _1405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .Y(_665_)
);

OAI21X1 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_420_),
    .C(_486_),
    .Y(_487_)
);

INVX1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_242_)
);

NAND2X1 _1443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_675_),
    .B(_696_),
    .Y(_699_)
);

NAND3X1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_296_),
    .C(_297_),
    .Y(_299_)
);

NOR2X1 _774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[14]),
    .Y(_82_)
);

OAI21X1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_239_),
    .C(_480_),
    .Y(_524_)
);

NAND2X1 _1308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_572_),
    .Y(_578_)
);

NAND2X1 _1481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin3[0]),
    .B(_732_),
    .Y(_733_)
);

AOI21X1 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_274_),
    .C(_336_),
    .Y(_337_)
);

DFFPOSX1 _1537_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .CLK(clk_bF$buf3),
    .Q(rYin[7])
);

NAND3X1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_386_),
    .C(_391_),
    .Y(_392_)
);

AOI22X1 _868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin_1_bF$buf3),
    .C(XinHL[2]),
    .D(Cin_0_bF$buf1),
    .Y(_148_)
);

NAND3X1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_560_),
    .C(_545_),
    .Y(_561_)
);

INVX1 _1346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .Y(_611_)
);

DFFPOSX1 _1575_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_49_),
    .CLK(clk_bF$buf2),
    .Q(y[15])
);

OAI22X1 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_420_),
    .C(_424_),
    .D(_428_),
    .Y(_429_)
);

OAI21X1 _1384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_637_),
    .C(_644_),
    .Y(_645_)
);

INVX1 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .Y(_467_)
);

NAND2X1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_440_),
    .Y(_521_)
);

OAI21X1 _1478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf0),
    .B(_730_),
    .C(_727_),
    .Y(_49_)
);

NAND3X1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_332_),
    .C(_333_),
    .Y(_334_)
);

AND2X2 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_548_),
    .Y(_558_)
);

INVX1 _830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[9]),
    .Y(_119_)
);

NAND2X1 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_366_),
    .Y(_371_)
);

NAND3X1 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_201_),
    .B(_199_),
    .C(_197_),
    .Y(_202_)
);

NOR2X1 _1402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_410_),
    .Y(_662_)
);

NAND3X1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_479_),
    .C(_482_),
    .Y(_484_)
);

INVX2 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[3]),
    .Y(_239_)
);

NOR2X1 _1440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_682_),
    .Y(_696_)
);

INVX1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .Y(_296_)
);

OAI21X1 _771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(y[13]),
    .C(_79_),
    .Y(_80_)
);

INVX1 _827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[8]),
    .Y(_117_)
);

INVX1 _1305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .Y(_575_)
);

DFFPOSX1 _1534_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .CLK(clk_bF$buf4),
    .Q(rYin[4])
);

AOI21X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_383_),
    .C(_382_),
    .Y(_389_)
);

NAND2X1 _865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[2]),
    .Y(_145_)
);

NOR2X1 _1343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_160_),
    .Y(_608_)
);

DFFPOSX1 _1572_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_46_),
    .CLK(clk_bF$buf1),
    .Q(y[12])
);

NAND3X1 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_421_),
    .C(_423_),
    .Y(_426_)
);

INVX1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .Y(_481_)
);

INVX1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .Y(_236_)
);

OAI21X1 _1381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_637_),
    .C(LoadCtl_4_bF$buf6),
    .Y(_643_)
);

AOI22X1 _1437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_470__bF$buf3),
    .C(_692_),
    .D(_693_),
    .Y(_45_)
);

AND2X2 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_293_)
);

INVX1 _768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .Y(_77_)
);

NAND2X1 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_463_),
    .Y(_464_)
);

NAND2X1 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_499_),
    .Y(_518_)
);

NAND2X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_270_),
    .Y(_274_)
);

NAND3X1 _1475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[14]),
    .B(rYin[15]),
    .C(_722_),
    .Y(_728_)
);

NAND3X1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_330_),
    .C(_325_),
    .Y(_331_)
);

FILL FILL71250x39750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_553_),
    .B(_549_),
    .Y(_555_)
);

FILL FILL70950x54150 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_179_),
    .C(_310_),
    .Y(_368_)
);

DFFPOSX1 _1569_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_43_),
    .CLK(clk_bF$buf5),
    .Q(y[9])
);

NAND3X1 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[4]),
    .C(_422_),
    .Y(_423_)
);

NOR2X1 _1378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_639_),
    .Y(_640_)
);

INVX1 _921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .Y(_199_)
);

AOI21X1 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_457_),
    .B(_456_),
    .C(_416_),
    .Y(_461_)
);

INVX1 _824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[7]),
    .Y(_115_)
);

AOI21X1 _1302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_413_),
    .C(_571_),
    .Y(_572_)
);

DFFPOSX1 _1531_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .CLK(clk_bF$buf0),
    .Q(rYin[1])
);

NAND3X1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_381_),
    .C(_385_),
    .Y(_386_)
);

NAND3X1 _862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf7),
    .B(_142_),
    .C(_139_),
    .Y(_143_)
);

AND2X2 _918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .Y(_196_)
);

OAI21X1 _1340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf2),
    .B(_604_),
    .C(_605_),
    .Y(_36_)
);

OAI21X1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_442_),
    .C(_477_),
    .Y(_478_)
);

INVX1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .Y(_233_)
);

INVX1 _1434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .Y(_691_)
);

NAND2X1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[5]),
    .Y(_290_)
);

NOR2X1 _765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_74_),
    .Y(_75_)
);

NOR2X1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_464_),
    .Y(_515_)
);

NAND2X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_270_),
    .Y(_271_)
);

OAI21X1 _1472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_725_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_726_)
);

AOI21X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_322_),
    .C(_321_),
    .Y(_328_)
);

DFFPOSX1 _1528_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .CLK(clk_bF$buf7),
    .Q(XinH[2])
);

NAND3X1 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_374_),
    .C(_369_),
    .Y(_383_)
);

INVX1 _859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .Y(_140_)
);

NAND2X1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(_551_),
    .Y(_552_)
);

OR2X2 _1337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_601_),
    .Y(_603_)
);

NAND2X1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_365_)
);

DFFPOSX1 _1566_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_40_),
    .CLK(clk_bF$buf3),
    .Q(y[6])
);

INVX2 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin[5]),
    .Y(_420_)
);

INVX2 _897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[2]),
    .Y(_176_)
);

AOI21X1 _1375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_636_),
    .C(_635_),
    .Y(_637_)
);

NAND3X1 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_456_),
    .C(_457_),
    .Y(_458_)
);

FILL FILL71250x25350 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[14]),
    .B(_722_),
    .Y(_723_)
);

NAND3X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .C(_289_),
    .Y(_325_)
);

OAI21X1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_525_),
    .C(_527_),
    .Y(_549_)
);

INVX1 _821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[6]),
    .Y(_113_)
);

NAND3X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_358_),
    .C(_359_),
    .Y(_362_)
);

AOI21X1 _915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_172_),
    .C(_174_),
    .Y(_193_)
);

AOI21X1 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_425_),
    .C(_428_),
    .Y(_475_)
);

INVX1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mul[5]),
    .Y(_230_)
);

NAND2X1 _1431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_688_)
);

INVX1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .Y(_287_)
);

NOR2X1 _762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[1]),
    .B(LoadCtl_0_bF$buf1),
    .Y(_72_)
);

INVX1 _818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[5]),
    .Y(_111_)
);

NAND3X1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_458_),
    .C(_511_),
    .Y(_512_)
);

NAND3X1 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .C(_234_),
    .Y(_268_)
);

OAI21X1 _1525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_178_),
    .C(_757_),
    .Y(_69_)
);

OAI21X1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_379_),
    .C(_377_),
    .Y(_380_)
);

NAND2X1 _856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin_0_bF$buf1),
    .Y(_137_)
);

NOR2X1 _1334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_144_),
    .Y(_600_)
);

DFFPOSX1 _1563_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .CLK(clk_bF$buf1),
    .Q(y[3])
);

INVX1 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .Y(_417_)
);

NAND3X1 _894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_167_),
    .C(_162_),
    .Y(_173_)
);

NAND2X1 _1372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_629_),
    .Y(_634_)
);

INVX1 _1428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .Y(_685_)
);

OAI21X1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_283_),
    .C(_273_),
    .Y(_284_)
);

NAND3X1 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_417_),
    .B(_449_),
    .C(_454_),
    .Y(_455_)
);

AOI22X1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(_470__bF$buf1),
    .C(_508_),
    .D(_509_),
    .Y(_29_)
);

NAND3X1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_257_),
    .C(_253_),
    .Y(_265_)
);

NOR2X1 _1466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_715_),
    .Y(_720_)
);

NAND3X1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_313_),
    .C(_308_),
    .Y(_322_)
);

NAND2X1 _797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Xin[1]),
    .B(_75_),
    .Y(_98_)
);

FILL FILL70950x61350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(LoadCtl_4_bF$buf4),
    .C(_546_),
    .Y(_30_)
);

NAND2X1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_353_),
    .Y(_359_)
);

OAI21X1 _1369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_630_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_632_)
);

OAI22X1 _912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(LoadCtl_4_bF$buf7),
    .C(_188_),
    .D(_190_),
    .Y(_23_)
);

DFFPOSX1 _1598_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(LoadCtl[1]),
    .CLK(clk_bF$buf6),
    .Q(LoadCtl[2])
);

NOR2X1 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_447_),
    .Y(_452_)
);

NAND3X1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_226_),
    .C(_192_),
    .Y(_228_)
);

INVX1 _815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[4]),
    .Y(_109_)
);

NAND2X1 _1522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(Xin[2]),
    .Y(_756_)
);

OAI21X1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_376_),
    .C(_311_),
    .Y(_377_)
);

OAI21X1 _853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(LoadCtl_4_bF$buf7),
    .C(_134_),
    .Y(_20_)
);

AOI21X1 _909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_187_),
    .C(_156_),
    .Y(_188_)
);

OAI21X1 _1331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf2),
    .B(_596_),
    .C(_597_),
    .Y(_35_)
);

DFFPOSX1 _1560_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .CLK(clk_bF$buf2),
    .Q(y[0])
);

AOI21X1 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_385_),
    .C(_351_),
    .Y(_414_)
);

NAND2X1 _891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_169_),
    .Y(_170_)
);

INVX1 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .Y(_225_)
);

AND2X2 _1425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_682_),
    .Y(_683_)
);

OAI21X1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(LoadCtl_4_bF$buf0),
    .C(_281_),
    .Y(_25_)
);

NOR2X1 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_506_),
    .Y(_507_)
);

OAI21X1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_260_),
    .C(_259_),
    .Y(_262_)
);

AOI22X1 _1463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_709_),
    .B(_470__bF$buf4),
    .C(_716_),
    .D(_717_),
    .Y(_47_)
);

OAI21X1 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_318_),
    .C(_316_),
    .Y(_319_)
);

OAI21X1 _794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_95_),
    .C(_96_),
    .Y(_758_[3])
);

OAI21X1 _1519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_140_),
    .C(_754_),
    .Y(_66_)
);

INVX1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .Y(_544_)
);

OAI21X1 _1328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_592_),
    .C(_587_),
    .Y(_595_)
);

OAI21X1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_239_),
    .C(_355_),
    .Y(_356_)
);

DFFPOSX1 _1557_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .CLK(clk_bF$buf5),
    .Q(mul[11])
);

NAND2X1 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_335_),
    .Y(_411_)
);

OAI21X1 _888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_165_),
    .C(_163_),
    .Y(_167_)
);

NOR2X1 _1366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_628_),
    .Y(_629_)
);

DFFPOSX1 _1595_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_69_),
    .CLK(clk_bF$buf7),
    .Q(XinHL[3])
);

NAND3X1 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_448_),
    .C(_419_),
    .Y(_449_)
);

FILL FILL71250x32550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL70950x14550 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_401_),
    .C(_341_),
    .Y(_541_)
);

INVX1 _812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[3]),
    .Y(_107_)
);

AOI21X1 _1498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_740_),
    .C(_743_),
    .Y(_56_)
);

AND2X2 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_353_)
);

OAI21X1 _850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_131_),
    .C(_132_),
    .Y(_19_)
);

NAND3X1 _906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(_172_),
    .C(_167_),
    .Y(_185_)
);

INVX1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .Y(_222_)
);

NOR2X1 _1422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_510_),
    .Y(_680_)
);

AOI22X1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_275_),
    .C(_221_),
    .D(_228_),
    .Y(_279_)
);

INVX1 _809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[2]),
    .Y(_105_)
);

NAND3X1 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_501_),
    .C(_500_),
    .Y(_504_)
);

OAI21X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_200_),
    .C(_197_),
    .Y(_259_)
);

INVX1 _1460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .Y(_715_)
);

OAI21X1 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_315_),
    .C(_255_),
    .Y(_316_)
);

OAI21X1 _791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf3),
    .B(_93_),
    .C(_94_),
    .Y(_758_[2])
);

NOR2X1 _1516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(Yin0[3]),
    .Y(_753_)
);

OAI21X1 _847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_129_),
    .C(_130_),
    .Y(_18_)
);

NOR2X1 _1325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[1]),
    .B(mul[1]),
    .Y(_592_)
);

DFFPOSX1 _1554_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .CLK(clk_bF$buf5),
    .Q(mul[8])
);

OAI21X1 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_408_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_409_)
);

NAND2X1 _885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[3]),
    .B(Cin_0_bF$buf0),
    .Y(_164_)
);

AOI21X1 _1363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_622_),
    .C(_618_),
    .Y(_626_)
);

OAI21X1 _1419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_469_),
    .C(_676_),
    .Y(_677_)
);

DFFPOSX1 _1592_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_66_),
    .CLK(clk_bF$buf7),
    .Q(XinHL[0])
);

NAND2X1 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_439_),
    .Y(_446_)
);

OAI21X1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_497_),
    .C(_478_),
    .Y(_501_)
);

OAI21X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_179_),
    .C(_203_),
    .Y(_256_)
);

NOR2X1 _1457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[13]),
    .B(mul[13]),
    .Y(_712_)
);

NAND3X1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_309_),
    .C(_311_),
    .Y(_313_)
);

OAI21X1 _788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf0),
    .B(_91_),
    .C(_92_),
    .Y(_758_[1])
);

NAND3X1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_499_),
    .C(_537_),
    .Y(_538_)
);

NOR2X1 _1495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin2[1]),
    .B(_740_),
    .Y(_742_)
);

AOI21X1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_313_),
    .C(_316_),
    .Y(_350_)
);

OAI21X1 _903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_181_),
    .C(_174_),
    .Y(_182_)
);

DFFPOSX1 _1589_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_63_),
    .CLK(clk_bF$buf4),
    .Q(Yin0[1])
);

OAI21X1 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_438_),
    .C(_430_),
    .Y(_443_)
);

NAND3X1 _1398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_656_),
    .C(_619_),
    .Y(_658_)
);

INVX1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .Y(_219_)
);

INVX1 _806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[1]),
    .Y(_103_)
);

AOI21X1 _1513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf2),
    .B(_734_),
    .C(_751_),
    .Y(_63_)
);

OAI21X1 _844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf1),
    .B(_127_),
    .C(_128_),
    .Y(_17_)
);

NAND2X1 _1322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[0]),
    .B(_470__bF$buf2),
    .Y(_590_)
);

DFFPOSX1 _1551_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .CLK(clk_bF$buf4),
    .Q(mul[5])
);

NAND3X1 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_392_),
    .C(_396_),
    .Y(_406_)
);

NAND2X1 _882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[0]),
    .B(Cin[3]),
    .Y(_161_)
);

BUFX2 _1607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_[1]),
    .Y(Yout[1])
);

OAI21X1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_210_),
    .C(_215_),
    .Y(_216_)
);

NAND2X1 _1360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_621_),
    .Y(_624_)
);

NAND2X1 _1416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[10]),
    .B(_470__bF$buf3),
    .Y(_674_)
);

OAI21X1 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_497_),
    .C(_495_),
    .Y(_498_)
);

NAND3X1 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_250_),
    .C(_252_),
    .Y(_253_)
);

INVX1 _1454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(y[13]),
    .Y(_709_)
);

AND2X2 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_1_bF$buf2),
    .Y(_310_)
);

OAI21X1 _785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf4),
    .B(_89_),
    .C(_90_),
    .Y(_758_[0])
);

NAND3X1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_519_),
    .B(_531_),
    .C(_534_),
    .Y(_535_)
);

INVX1 _1319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .Y(_587_)
);

NOR2X1 _1492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_77_),
    .Y(_740_)
);

AOI21X1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_320_),
    .C(_327_),
    .Y(_347_)
);

DFFPOSX1 _1548_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .CLK(clk_bF$buf0),
    .Q(mul[2])
);

OAI21X1 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_343_),
    .C(_335_),
    .Y(_403_)
);

NAND2X1 _879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf7),
    .B(_158_),
    .Y(_159_)
);

OAI21X1 _1357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_618_),
    .C(_620_),
    .Y(_621_)
);

INVX1 _900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Cin_0_bF$buf2),
    .Y(_179_)
);

DFFPOSX1 _1586_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_60_),
    .CLK(clk_bF$buf3),
    .Q(Yin1[2])
);

INVX1 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .Y(_440_)
);

CLKBUF1 CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

OAI21X1 _1395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .B(_644_),
    .C(_654_),
    .Y(_655_)
);

INVX1 _803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rYin[0]),
    .Y(_101_)
);

INVX1 _1489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Yin[3]),
    .Y(_738_)
);

OAI22X1 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(LoadCtl_4_bF$buf6),
    .C(_342_),
    .D(_344_),
    .Y(_26_)
);

INVX1 _1298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .Y(_568_)
);

NOR2X1 _1510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_0_bF$buf1),
    .B(Yin0[0]),
    .Y(_750_)
);

OAI21X1 _841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf3),
    .B(_125_),
    .C(_126_),
    .Y(_16_)
);

BUFX2 _1604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_[2]),
    .Y(Xout[2])
);

NAND2X1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_213_)
);

NOR2X1 _1413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_667_),
    .Y(_672_)
);

AOI21X1 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_494_),
    .C(_438_),
    .Y(_495_)
);

NAND2X1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_249_),
    .Y(_250_)
);

INVX1 _1451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .Y(_707_)
);

NAND3X1 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[1]),
    .B(Cin_1_bF$buf2),
    .C(_306_),
    .Y(_307_)
);

OAI21X1 _782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_87_),
    .C(_88_),
    .Y(_759_[3])
);

OAI21X1 _1507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_745_),
    .C(_748_),
    .Y(_60_)
);

OAI21X1 _838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl_4_bF$buf2),
    .B(_123_),
    .C(_124_),
    .Y(_15_)
);

INVX1 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .Y(_532_)
);

NOR2X1 _1316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(_583_),
    .Y(_585_)
);

DFFPOSX1 _1545_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .CLK(clk_bF$buf2),
    .Q(rYin[15])
);

AOI22X1 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_332_),
    .C(_398_),
    .D(_399_),
    .Y(_400_)
);

INVX1 _876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .Y(_156_)
);

NOR2X1 _1354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_191_),
    .Y(_618_)
);

DFFPOSX1 _1583_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_57_),
    .CLK(clk_bF$buf6),
    .Q(Yin2[3])
);

OAI21X1 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_434_),
    .C(_436_),
    .Y(_437_)
);

NAND3X1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_491_),
    .C(_487_),
    .Y(_492_)
);

OAI21X1 _1392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470__bF$buf1),
    .B(_651_),
    .C(_652_),
    .Y(_41_)
);

NOR2X1 _1448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_703_),
    .Y(_704_)
);

AND2X2 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .Y(_304_)
);

NAND2X1 _779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(LoadCtl[2]),
    .B(_85_),
    .Y(_86_)
);

endmodule
