/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module cpu(
    inout vdd,
    inout gnd,
    output [15:0] AB,
    input [7:0] DI,
    output [7:0] DO,
    input IRQ,
    input NMI,
    input RDY,
    output WE,
    input clk,
    input reset
);

wire C ;
wire D ;
wire I ;
wire N ;
wire V ;
wire Z ;
wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire [5:0] _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire IRQ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1__bF$buf10 ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire WE ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire php ;
wire _1192_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire RDY ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire adc_sbc ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _887__bF$buf0 ;
wire _887__bF$buf1 ;
wire _887__bF$buf2 ;
wire _887__bF$buf3 ;
wire _887__bF$buf4 ;
wire _1283_ ;
wire _194_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire write_back ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire index_y ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire clc ;
wire cld ;
wire cli ;
wire clk ;
wire clv ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _830__bF$buf0 ;
wire _830__bF$buf1 ;
wire _830__bF$buf2 ;
wire _830__bF$buf3 ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1271_ ;
wire _182_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire IRHOLD_valid_bF$buf0 ;
wire IRHOLD_valid_bF$buf1 ;
wire IRHOLD_valid_bF$buf2 ;
wire IRHOLD_valid_bF$buf3 ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire HC ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire _1268_ ;
wire _691__bF$buf0 ;
wire _691__bF$buf1 ;
wire _691__bF$buf2 ;
wire _691__bF$buf3 ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire [6:0] ADD ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire RDY_bF$buf0 ;
wire RDY_bF$buf1 ;
wire RDY_bF$buf2 ;
wire RDY_bF$buf3 ;
wire RDY_bF$buf4 ;
wire RDY_bF$buf5 ;
wire RDY_bF$buf6 ;
wire RDY_bF$buf7 ;
wire RDY_bF$buf8 ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire res ;
wire _787_ ;
wire _367_ ;
wire rotate ;
wire [15:0] _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire [3:0] alu_op ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire [1:0] dst_reg ;
wire \u_ALU8.BI7  ;
wire [7:0] DIHOLD ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _1453_ ;
wire _1033_ ;
wire _918__bF$buf0 ;
wire _918__bF$buf1 ;
wire _918__bF$buf2 ;
wire _918__bF$buf3 ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire \u_ALU8.BCD  ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire [7:0] \AXYS[1]  ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _1129__bF$buf0 ;
wire _1129__bF$buf1 ;
wire _1129__bF$buf2 ;
wire _1129__bF$buf3 ;
wire _1129__bF$buf4 ;
wire _853__bF$buf0 ;
wire _853__bF$buf1 ;
wire _853__bF$buf2 ;
wire _853__bF$buf3 ;
wire _853__bF$buf4 ;
wire _853__bF$buf5 ;
wire _853__bF$buf6 ;
wire _853__bF$buf7 ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire store ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire IRHOLD_valid ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _1002__bF$buf0 ;
wire _1002__bF$buf1 ;
wire _1002__bF$buf2 ;
wire _1002__bF$buf3 ;
wire _1002__bF$buf4 ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _1__bF$buf0 ;
wire _1__bF$buf1 ;
wire _1__bF$buf2 ;
wire _1__bF$buf3 ;
wire _1__bF$buf4 ;
wire _1__bF$buf5 ;
wire _1__bF$buf6 ;
wire _1__bF$buf7 ;
wire _1__bF$buf8 ;
wire _1__bF$buf9 ;
wire _919_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire backwards ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _44_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _926__bF$buf0 ;
wire _926__bF$buf1 ;
wire _926__bF$buf2 ;
wire _926__bF$buf3 ;
wire _725_ ;
wire _305_ ;
wire [15:0] PC ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _882__bF$buf0 ;
wire _882__bF$buf1 ;
wire _882__bF$buf2 ;
wire _882__bF$buf3 ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire adj_bcd ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire [7:0] \AXYS[3]  ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire compare ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire load_only ;
wire clk_bF$buf10 ;
wire shift ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire [1:0] src_reg ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _1273_ ;
wire _184_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _869__bF$buf0 ;
wire _869__bF$buf1 ;
wire _869__bF$buf2 ;
wire _869__bF$buf3 ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1270_ ;
wire _181_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _1593_ ;
wire _1173_ ;
wire _1649_ ;
wire _1229_ ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire [2:0] cond_code ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [5:0] state ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire bit_ins ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire [7:0] DI ;
wire [7:0] DO ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire [15:0] AB ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _886__bF$buf0 ;
wire _886__bF$buf1 ;
wire _886__bF$buf2 ;
wire _886__bF$buf3 ;
wire _704_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _1051__bF$buf0 ;
wire _1051__bF$buf1 ;
wire _1051__bF$buf2 ;
wire _1051__bF$buf3 ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire NMI ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire plp ;
wire _1196_ ;
wire _55_ ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1669_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire [7:0] \AXYS[0]  ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire shift_right ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire [7:0] DIMUX ;
wire _1278_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire [3:0] op ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire sec ;
wire sed ;
wire sei ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire [7:0] IRHOLD ;
wire _1275_ ;
wire _186_ ;
wire alu_shift_right ;
wire _1084_ ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _1519_ ;
wire _1272_ ;
wire _183_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire _1269_ ;
wire NMI_1 ;
wire _812_ ;
wire _72_ ;
wire _1649__bF$buf0 ;
wire _1649__bF$buf1 ;
wire _1498_ ;
wire _1649__bF$buf2 ;
wire _1078_ ;
wire _1649__bF$buf3 ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _1219__bF$buf0 ;
wire _1219__bF$buf1 ;
wire _1219__bF$buf2 ;
wire _1219__bF$buf3 ;
wire adc_bcd ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire [7:0] _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _903_ ;
wire [7:0] \AXYS[2]  ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire [7:0] ABH ;
wire [7:0] ABL ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire NMI_edge ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire load_reg ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire inc ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _612_ ;
wire _1298_ ;
wire reset ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

FILL FILL_8__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[6]),
    .B(_1674_),
    .C(_1676_),
    .Y(_1677_)
);

FILL FILL_1__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[6]),
    .Y(_838_)
);

FILL FILL_3__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_586_),
    .C(_588_),
    .Y(_589_)
);

FILL FILL_1__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1526_),
    .B(_1522_),
    .C(_1520_),
    .Y(_1527_)
);

FILL FILL_6__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(DI[7]),
    .Y(_686_)
);

FILL FILL_2__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[10]),
    .B(_853__bF$buf5),
    .Y(_433_)
);

FILL FILL_0__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3250_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_13_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[11])
);

FILL FILL_2__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181350x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[0]),
    .Y(_621_)
);

FILL FILL_6__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_240_),
    .C(_1057_),
    .Y(_264_)
);

OAI21X1 _2101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1235_),
    .C(_1236_),
    .Y(_1237_)
);

FILL FILL_5__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3306_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_60_),
    .CLK(clk_bF$buf10),
    .Q(IRHOLD[7])
);

FILL FILL_1__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[5]),
    .B(_446_),
    .C(_467_),
    .Y(_468_)
);

AND2X2 _2330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(_1279_),
    .Y(_1462_)
);

FILL FILL_4__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1602_),
    .C(_1617_),
    .Y(_1621_)
);

OAI21X1 _3115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf1),
    .B(_758_),
    .C(\AXYS[2] [2]),
    .Y(_761_)
);

FILL FILL_1__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_1323_),
    .Y(_513_)
);

FILL FILL_1__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3344_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_97_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[3] [4])
);

FILL FILL_6__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[7]),
    .Y(_975_)
);

FILL FILL_0__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(res),
    .B(_1051__bF$buf1),
    .C(_344_),
    .Y(_345_)
);

FILL FILL_1__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(_887__bF$buf4)
);

FILL FILL_3__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3573_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1491_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf3),
    .Q(ADD[3])
);

FILL FILL_6__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(_784_),
    .C(_783_),
    .Y(_785_)
);

FILL FILL_2__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_542_),
    .Y(_543_)
);

FILL FILL_6__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[15]),
    .Y(_176_)
);

INVX1 _2004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD[3]),
    .Y(_1140_)
);

FILL FILL_9__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_237_),
    .C(_836_),
    .Y(_105_)
);

FILL FILL_1__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .Y(_1657_)
);

FILL FILL_6__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_373_),
    .C(_378_),
    .Y(_379_)
);

NOR2X1 _2233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .B(_1366_),
    .Y(_1367_)
);

FILL FILL_2__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[2]),
    .Y(_1524_)
);

NAND2X1 _3018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(C),
    .B(_678_),
    .Y(_684_)
);

FILL FILL_1__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(_822_),
    .Y(_823_)
);

FILL FILL_2__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .Y(_1067_)
);

FILL FILL_0__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .Y(_431_)
);

FILL FILL_7__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf2),
    .B(_572_),
    .C(_570_),
    .Y(_42_)
);

FILL FILL_6__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1025_),
    .B(_182_),
    .C(_212_),
    .Y(_213_)
);

INVX1 _2042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .Y(_1178_)
);

FILL FILL_2__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3247_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_10_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[8])
);

FILL FILL_7__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_881_),
    .Y(_886_)
);

FILL FILL_4__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1043_),
    .B(_1044_),
    .C(RDY_bF$buf1),
    .Y(_618_)
);

NOR2X1 _2518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_208_),
    .Y(_261_)
);

FILL FILL_1__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1075_),
    .B(_1264_),
    .C(_413_),
    .Y(_414_)
);

NAND3X1 _2271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1317_),
    .B(_1403_),
    .C(_1404_),
    .Y(_1405_)
);

FILL FILL_2__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(_1560_),
    .C(_1538_),
    .Y(_1562_)
);

FILL FILL_6__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_697_),
    .C(_716_),
    .Y(_717_)
);

FILL FILL_2__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_944_),
    .C(_1100_),
    .Y(_1101_)
);

AOI21X1 _2747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[5]),
    .B(_325_),
    .C(_1284_),
    .Y(_465_)
);

NAND2X1 _2327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1349_),
    .B(_1431_),
    .Y(_1459_)
);

FILL FILL_7__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1155_),
    .Y(_1216_)
);

FILL FILL_5_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3285_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_47_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(src_reg[0])
);

FILL FILL_6__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_911_),
    .B(_913_),
    .C(_923_),
    .Y(_924_)
);

FILL FILL_2__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(ADD[3]),
    .Y(_646_)
);

FILL FILL_6__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_195_),
    .C(DIMUX[5]),
    .Y(_294_)
);

OAI21X1 _2136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_1032_),
    .C(RDY_bF$buf0),
    .Y(_1272_)
);

FILL FILL_7__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_747_),
    .C(_749_),
    .Y(_77_)
);

FILL FILL_2__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_933_),
    .C(_861_),
    .D(_967_),
    .Y(BI[5])
);

FILL FILL_7__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_498_),
    .Y(_499_)
);

OAI21X1 _2365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf3),
    .B(_946_),
    .C(_126_),
    .Y(_127_)
);

FILL FILL_8__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_867_),
    .C(_918__bF$buf0),
    .Y(_325_)
);

OAI21X1 _2174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf2),
    .B(_946_),
    .C(_978_),
    .Y(_1309_)
);

FILL FILL_2__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(BI[7]),
    .Y(_1654_)
);

FILL FILL_0__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(dst_reg[0]),
    .B(_1008_),
    .Y(_1009_)
);

FILL FILL_6__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .Y(_820_)
);

FILL FILL_0__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf1),
    .C(inc),
    .Y(_570_)
);

AOI22X1 _2459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[0]),
    .B(_204_),
    .C(_202_),
    .D(ABL[0]),
    .Y(_210_)
);

NOR2X1 _2039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .B(_1174_),
    .Y(_1175_)
);

FILL FILL_7__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(_1660_),
    .Y(_1674_)
);

FILL FILL_3__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_410_),
    .Y(_411_)
);

NOR2X1 _2268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1315_),
    .Y(_1402_)
);

FILL FILL_7__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1095_),
    .B(_1097_),
    .C(_1096_),
    .Y(_1098_)
);

FILL FILL_2__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_585_),
    .C(_544_),
    .Y(_586_)
);

FILL FILL_3__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_242_),
    .Y(_243_)
);

NAND3X1 _2077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(_1181_),
    .C(_1212_),
    .Y(_1213_)
);

FILL FILL_0__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(C),
    .B(_912_),
    .Y(_921_)
);

FILL FILL_4__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(I),
    .B(_1131_),
    .C(_1132_),
    .Y(_1133_)
);

FILL FILL_8__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3303_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_57_),
    .CLK(clk_bF$buf10),
    .Q(IRHOLD[4])
);

FILL FILL_1__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1597_),
    .B(_1594_),
    .Y(_1618_)
);

OAI21X1 _3112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_757_),
    .C(_759_),
    .Y(_85_)
);

FILL FILL_2__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_1129__bF$buf0),
    .C(_510_),
    .D(_507_),
    .Y(_25_)
);

FILL FILL_1__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3341_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_94_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[3] [1])
);

FILL FILL_6__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_931_),
    .C(_332_),
    .D(_342_),
    .Y(_2_)
);

FILL FILL_0__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3570_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1488_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf3),
    .Q(ADD[0])
);

FILL FILL_8__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_780_),
    .C(_778_),
    .Y(_782_)
);

FILL FILL_2__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_1219__bF$buf1),
    .C(_537_),
    .D(_540_),
    .Y(_33_)
);

FILL FILL_6__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .B(_139_),
    .C(_173_),
    .Y(_174_)
);

AOI21X1 _2001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .B(IRHOLD_valid_bF$buf3),
    .C(_1133_),
    .Y(_1137_)
);

FILL FILL_5__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[3]),
    .Y(_835_)
);

FILL FILL_1__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_376_)
);

OAI21X1 _2230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_927_),
    .B(_1037_),
    .C(_886__bF$buf2),
    .Y(_1364_)
);

FILL FILL_2__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(AI[2]),
    .C(_1653_),
    .Y(_1521_)
);

OAI21X1 _3015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_679_),
    .C(_680_),
    .Y(_681_)
);

FILL FILL_1__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1063_),
    .Y(_1064_)
);

FILL FILL_0__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(_406_),
    .C(_427_),
    .Y(_428_)
);

FILL FILL_7__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3244_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_7_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf2),
    .Q(PC[5])
);

FILL FILL_6__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf0),
    .B(_880_),
    .Y(_883_)
);

FILL FILL_6__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_616_),
    .Y(_617_)
);

AOI21X1 _2515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .B(_182_),
    .C(_258_),
    .Y(_259_)
);

FILL FILL_1__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1546_),
    .B(_1550_),
    .C(_1558_),
    .Y(_1559_)
);

FILL FILL_6__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [2]),
    .B(_693_),
    .Y(_715_)
);

FILL FILL_2__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_283_),
    .C(_462_),
    .Y(_14_)
);

NAND3X1 _2324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1450_),
    .B(_1454_),
    .C(_1456_),
    .Y(_1457_)
);

FILL FILL_5__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1614_),
    .C(_1589_),
    .Y(_1615_)
);

NAND2X1 _3109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_1023_),
    .Y(_757_)
);

FILL FILL_1__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3282_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_44_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(write_back)
);

FILL FILL_6__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_642_),
    .Y(_643_)
);

FILL FILL_6__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[13]),
    .Y(_291_)
);

NAND2X1 _2133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf1),
    .B(_1268_),
    .Y(_1269_)
);

FILL FILL_2__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3338_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_92_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[2] [7])
);

FILL FILL_1__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_1022_),
    .Y(_747_)
);

FILL FILL_2__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[4]),
    .Y(_972_)
);

FILL FILL_4__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_318_),
    .C(_337_),
    .D(_339_),
    .Y(_340_)
);

FILL FILL_1__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(NMI_edge),
    .B(_495_),
    .C(_496_),
    .Y(_18_)
);

INVX1 _2362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(op[2]),
    .Y(_124_)
);

FILL FILL_8__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3567_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1485_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf4),
    .Q(\u_ALU8.BI7 )
);

FILL FILL_6__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf3),
    .B(_880_),
    .C(_1002__bF$buf4),
    .Y(_779_)
);

FILL FILL_7__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1162_),
    .Y(_538_)
);

OAI21X1 _2418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[14]),
    .Y(_171_)
);

FILL FILL_1__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf4),
    .B(_1267_),
    .C(_1051__bF$buf2),
    .Y(_322_)
);

NOR2X1 _2171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1295_),
    .Y(_1306_)
);

FILL FILL_2__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .Y(_1651_)
);

FILL FILL_6__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf0),
    .B(_998_),
    .C(_1005_),
    .Y(_1006_)
);

FILL FILL_6__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_373_),
    .Y(_374_)
);

NAND2X1 _2227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1346_),
    .Y(_1362_)
);

FILL FILL_7__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_809_),
    .C(_816_),
    .Y(_817_)
);

FILL FILL_0__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [1]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [1]),
    .Y(_1061_)
);

FILL FILL_7__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_566_),
    .C(_567_),
    .D(_568_),
    .Y(_40_)
);

FILL FILL_6__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_206_),
    .Y(_207_)
);

NAND2X1 _2036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .B(_1171_),
    .Y(_1172_)
);

FILL FILL_7__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_868_),
    .Y(_880_)
);

FILL FILL_4__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[7]),
    .B(_336_),
    .Y(_408_)
);

OAI21X1 _2265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1159_),
    .C(_1299_),
    .Y(_1399_)
);

FILL FILL_0__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [5]),
    .B(_1022_),
    .Y(_1095_)
);

FILL FILL_7__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .Y(_240_)
);

OR2X2 _2074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_1209_),
    .Y(_1210_)
);

FILL FILL_2__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3279_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_41_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf5),
    .Q(adc_sbc)
);

FILL FILL_0__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_917_),
    .Y(_918_)
);

FILL FILL_4__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _3088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(DIMUX[7]),
    .S(_981_),
    .Y(_745_)
);

FILL FILL_0__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD[1]),
    .Y(_1130_)
);

FILL FILL_8__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(NMI_1),
    .Y(_494_)
);

OAI21X1 _2359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_120_),
    .C(_122_),
    .Y(alu_op[0])
);

FILL FILL_7__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3300_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_54_),
    .CLK(clk_bF$buf5),
    .Q(IRHOLD[1])
);

FILL FILL_3__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_314_),
    .Y(_319_)
);

NAND2X1 _2168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1161_),
    .Y(_1303_)
);

FILL FILL_7__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1001_),
    .B(_1002__bF$buf0),
    .C(_998_),
    .Y(_1003_)
);

FILL FILL_7__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(sec),
    .Y(_508_)
);

FILL FILL_0__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[2]),
    .B(_139_),
    .C(_153_),
    .Y(_154_)
);

FILL FILL_8__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .B(_1040_),
    .Y(_1041_)
);

FILL FILL_8__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_218_),
    .C(_833_),
    .Y(_102_)
);

FILL FILL_1__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1517_),
    .C(_1515_),
    .Y(_1518_)
);

AND2X2 _3012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_676_),
    .Y(_678_)
);

FILL FILL_2__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf2),
    .B(_423_),
    .C(_424_),
    .Y(_425_)
);

FILL FILL_0__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3241_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_4_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(PC[2])
);

FILL FILL_9__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .B(_1168_),
    .C(_603_),
    .Y(_614_)
);

NAND2X1 _2512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_255_),
    .Y(_256_)
);

FILL FILL_9__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1554_),
    .Y(_1556_)
);

FILL FILL_6__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_702_),
    .Y(_712_)
);

FILL FILL_2__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(_410_),
    .C(_367_),
    .Y(_460_)
);

NOR3X1 _2321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .B(_1452_),
    .C(_1451_),
    .Y(_1454_)
);

FILL FILL_9__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .B(_1566_),
    .Y(_1612_)
);

OAI21X1 _3106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_747_),
    .C(_755_),
    .Y(_83_)
);

FILL FILL_1__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(V),
    .B(_636_),
    .Y(_641_)
);

FILL FILL_6__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_268_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _2130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(_1262_),
    .Y(_1266_)
);

FILL FILL_2__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3335_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_89_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[2] [4])
);

FILL FILL_1__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(_933_),
    .C(_855_),
    .D(_967_),
    .Y(BI[2])
);

FILL FILL_0__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[0]),
    .B(_336_),
    .Y(_337_)
);

FILL FILL_1__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .Y(_1640_)
);

FILL FILL_6__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_910_),
    .B(_869__bF$buf2),
    .C(_1224_),
    .Y(_776_)
);

FILL FILL_2__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_526_),
    .Y(_536_)
);

NOR2X1 _2415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_168_),
    .Y(_169_)
);

FILL FILL_1__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _3373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .Y(_1484_)
);

FILL FILL_6__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_371_)
);

NAND3X1 _2224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1357_),
    .C(_1355_),
    .Y(_1359_)
);

FILL FILL_2__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1514_),
    .B(_1512_),
    .Y(_1515_)
);

NAND2X1 _3009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_674_),
    .Y(_675_)
);

FILL FILL_1__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[5]),
    .B(_996_),
    .C(_952_),
    .Y(_814_)
);

FILL FILL_2__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[0]),
    .C(_1058_),
    .Y(_1059_)
);

FILL FILL_1_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .Y(_566_)
);

FILL FILL_6__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf0),
    .B(_1032_),
    .C(_1184_),
    .Y(_204_)
);

INVX1 _2033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf0),
    .Y(_1169_)
);

FILL FILL_2__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3238_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[5]),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf6),
    .Q(state[5])
);

FILL FILL_1__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf0),
    .B(_876_),
    .Y(_877_)
);

FILL FILL_4__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_610_),
    .B(_608_),
    .Y(_611_)
);

INVX1 _2509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[7]),
    .Y(_253_)
);

FILL FILL_1__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_404_),
    .C(_400_),
    .Y(_405_)
);

NAND2X1 _2262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1395_),
    .Y(_1396_)
);

FILL FILL_2__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(_1552_),
    .Y(_1553_)
);

FILL FILL_6__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _3047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(ADD[2]),
    .Y(_709_)
);

FILL FILL_7__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_944_),
    .C(_1092_),
    .Y(_1093_)
);

OR2X2 _2738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_454_),
    .Y(_457_)
);

NAND3X1 _2318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1181_),
    .C(_1211_),
    .Y(_1451_)
);

FILL FILL_1__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_1685_[4])
);

NAND2X1 _2071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1206_),
    .Y(_1207_)
);

FILL FILL_2__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3276_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_38_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(compare)
);

FILL FILL_6__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_888_),
    .Y(_915_)
);

FILL FILL_6__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(ADD[6]),
    .Y(_638_)
);

FILL FILL_6__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_195_),
    .C(DIMUX[4]),
    .Y(_286_)
);

OAI21X1 _2127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf3),
    .B(_891_),
    .C(RDY_bF$buf5),
    .Y(_1263_)
);

FILL FILL_7__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(_698_),
    .Y(_742_)
);

FILL FILL_0__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[1]),
    .Y(_969_)
);

FILL FILL_7__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf0),
    .B(_1124_),
    .C(_1126_),
    .D(_1125_),
    .Y(_1127_)
);

FILL FILL_8__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x160050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_489_),
    .Y(_492_)
);

INVX2 _2356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .Y(_120_)
);

FILL FILL_7__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf4),
    .B(_1133_),
    .C(_315_),
    .Y(_316_)
);

NOR2X1 _2165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(_1295_),
    .Y(_1300_)
);

FILL FILL_0__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_987_),
    .B(_999_),
    .Y(_1000_)
);

FILL FILL_7__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[10]),
    .Y(_151_)
);

FILL FILL_8__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[4]),
    .Y(DO[4])
);

NAND3X1 _3179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_810_),
    .C(_778_),
    .Y(_811_)
);

FILL FILL_0__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .B(_1037_),
    .Y(_1038_)
);

FILL FILL_8__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[0]),
    .B(_869__bF$buf3),
    .C(_905_),
    .Y(_402_)
);

OR2X2 _2259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1392_),
    .B(_1305_),
    .Y(_1393_)
);

FILL FILL182250x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[0]),
    .Y(_832_)
);

FILL FILL_3__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_234_),
    .Y(_235_)
);

OAI21X1 _2068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf0),
    .B(_1029_),
    .C(_1203_),
    .Y(_1204_)
);

FILL FILL_0__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shift),
    .Y(_912_)
);

FILL FILL_4__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1065_),
    .B(_872_),
    .C(_267_),
    .D(_333_),
    .Y(_422_)
);

FILL FILL_0__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1392_),
    .Y(_1430_)
);

FILL FILL_0__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .Y(_1124_)
);

FILL FILL_4__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_893_),
    .Y(_949_)
);

FILL FILL_4__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .B(_1605_),
    .Y(_1609_)
);

OAI21X1 _3103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf3),
    .B(_748_),
    .C(\AXYS[1] [5]),
    .Y(_754_)
);

FILL FILL_1__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3332_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_86_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[2] [1])
);

FILL FILL_2__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf0),
    .B(_1259_),
    .C(_333_),
    .Y(_334_)
);

FILL FILL_1__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .Y(_1638_)
);

FILL FILL_6__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_767_),
    .C(_774_),
    .Y(_99_)
);

FILL FILL_6__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_530_),
    .C(_532_),
    .Y(_533_)
);

OAI21X1 _2412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_1091_),
    .C(_166_),
    .Y(_1686_[4])
);

FILL FILL_0__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.AI7 ),
    .B(CO),
    .Y(_1647_)
);

FILL FILL_6__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_971_),
    .C(_368_),
    .D(_363_),
    .Y(_5_)
);

OAI21X1 _2221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_946_),
    .C(RDY_bF$buf7),
    .Y(_1356_)
);

FILL FILL_2__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(_1510_),
    .C(_1507_),
    .Y(_1512_)
);

NOR2X1 _3006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(write_back),
    .B(_1002__bF$buf3),
    .Y(_672_)
);

FILL FILL_1__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1055_),
    .B(_872_),
    .Y(_1056_)
);

FILL FILL_0__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf0),
    .B(_531_),
    .Y(_564_)
);

FILL FILL_6__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_199_),
    .Y(_201_)
);

NAND3X1 _2030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1127_),
    .B(_1128_),
    .C(_1165_),
    .Y(_1166_)
);

FILL FILL_2__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3235_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[2]),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(state[2])
);

FILL FILL_1__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_866_),
    .Y(_874_)
);

FILL FILL_6__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_523_),
    .C(_547_),
    .Y(_608_)
);

AOI21X1 _2506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .B(_182_),
    .C(_250_),
    .Y(_251_)
);

FILL FILL_1__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(_1542_),
    .C(_1549_),
    .Y(_1550_)
);

FILL FILL_6__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .Y(_707_)
);

FILL FILL_2__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .B(_1089_),
    .C(_1088_),
    .Y(_1090_)
);

OAI21X1 _2735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_333_),
    .C(_1092_),
    .Y(_454_)
);

OAI21X1 _2315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .B(_1447_),
    .C(_1380_),
    .Y(_1448_)
);

FILL FILL_1__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3273_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_35_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(op[3])
);

FILL FILL_6__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .Y(_635_)
);

FILL FILL_6__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[12]),
    .Y(_283_)
);

NOR2X1 _2124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf3),
    .B(_1259_),
    .Y(_1260_)
);

FILL FILL_2__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3329_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_83_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[1] [6])
);

FILL FILL_1__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_738_),
    .C(_739_),
    .Y(_75_)
);

FILL FILL_2__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_958_),
    .B(_966_),
    .C(_948_),
    .Y(_967_)
);

FILL FILL_4__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x121050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_445_),
    .C(_488_),
    .Y(_489_)
);

OR2X2 _2353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_1470_),
    .Y(_1483_[5])
);

FILL FILL_4__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf1),
    .B(_1619_),
    .C(_1636_),
    .Y(_1493_)
);

FILL FILL_6__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [5]),
    .B(_767_),
    .Y(_773_)
);

FILL FILL_7__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .Y(_530_)
);

OAI21X1 _2409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf1),
    .B(_989_),
    .C(_138_),
    .Y(_164_)
);

FILL FILL_1__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_1268_),
    .C(_312_),
    .Y(_313_)
);

NAND2X1 _2162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1154_),
    .Y(_1297_)
);

FILL FILL_2__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(ADD[2]),
    .Y(_1645_)
);

FILL FILL_6__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_996_),
    .C(_992_),
    .Y(_997_)
);

FILL FILL_6__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_364_),
    .B(_355_),
    .C(_365_),
    .D(_361_),
    .Y(_366_)
);

NOR2X1 _2218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf0),
    .B(_1032_),
    .Y(_1353_)
);

FILL FILL_7__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(_139_),
    .C(_148_),
    .Y(_149_)
);

FILL FILL_8__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[1]),
    .Y(DO[1])
);

FILL FILL_6__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .B(_978_),
    .C(_807_),
    .Y(_808_)
);

FILL FILL_0__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .Y(_1053_)
);

FILL FILL_7__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_1178_),
    .Y(_562_)
);

FILL FILL_6__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .Y(_198_)
);

NAND2X1 _2027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1162_),
    .Y(_1163_)
);

FILL FILL_7__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x160050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .B(_870_),
    .Y(_871_)
);

FILL FILL_4__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_945_),
    .Y(_1035_)
);

FILL FILL_8__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_975_),
    .C(_399_),
    .Y(_9_)
);

NOR2X1 _2256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf3),
    .B(_1253_),
    .Y(_1390_)
);

FILL FILL_7__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [4]),
    .B(_1022_),
    .Y(_1087_)
);

FILL FILL_7__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .Y(_1685_[3])
);

NAND3X1 _2065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_1200_),
    .C(_878_),
    .Y(_1201_)
);

FILL FILL_2__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .B(_888_),
    .Y(_909_)
);

FILL FILL_4__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x113250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1424_),
    .C(_1426_),
    .Y(_1427_)
);

FILL FILL_2__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.BCD ),
    .B(_1584_),
    .Y(_1585_)
);

OAI21X1 _3079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_981_),
    .C(_736_),
    .Y(_737_)
);

FILL FILL_0__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(AN),
    .C(_1121_),
    .Y(_1122_)
);

FILL FILL_4__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_915_),
    .B(_945_),
    .Y(_946_)
);

FILL FILL_5__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .B(_629_),
    .C(bit_ins),
    .D(_658_),
    .Y(_666_)
);

NOR2X1 _2579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_120_),
    .Y(alu_shift_right)
);

INVX1 _2159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1294_),
    .Y(_1483_[0])
);

FILL FILL_7__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1605_),
    .B(_1604_),
    .C(_1667_),
    .Y(_1606_)
);

OAI21X1 _3100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_747_),
    .C(_752_),
    .Y(_80_)
);

FILL FILL_4__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[9]),
    .Y(_146_)
);

FILL FILL_6__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_323_),
    .Y(_331_)
);

FILL FILL_9__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1331_),
    .B(_1325_),
    .Y(_1332_)
);

FILL FILL_0__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(_871_),
    .Y(_1032_)
);

FILL FILL_8__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .Y(DIMUX[2])
);

FILL FILL_8__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_1508_),
    .Y(_1509_)
);

MUX2X1 _3003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(AZ),
    .S(_1192_),
    .Y(_670_)
);

FILL FILL_1__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1118_),
    .B(_830__bF$buf2),
    .C(_848_),
    .Y(_116_)
);

FILL FILL_3_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_600_),
    .B(_605_),
    .Y(_606_)
);

OAI21X1 _2503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_226_),
    .C(_247_),
    .Y(_248_)
);

FILL FILL_1__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .B(_1545_),
    .C(_1546_),
    .Y(_1547_)
);

FILL FILL_6__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_703_),
    .Y(_704_)
);

FILL FILL_2__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_450_),
    .C(_430_),
    .Y(_452_)
);

OAI21X1 _2312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1444_),
    .C(_1221_),
    .Y(_1445_)
);

FILL FILL_0__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1602_),
    .Y(_1603_)
);

FILL FILL_1__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3270_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_32_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(op[0])
);

FILL FILL_8__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181350x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(_1002__bF$buf3),
    .Y(_632_)
);

FILL FILL_6__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_196_),
    .C(_280_),
    .Y(_281_)
);

OAI21X1 _2121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf0),
    .B(_959_),
    .C(_1256_),
    .Y(_1257_)
);

FILL FILL_2__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3326_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_80_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[1] [3])
);

FILL FILL_1__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .B(_927_),
    .C(_886__bF$buf3),
    .Y(_964_)
);

FILL FILL_0__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_325_),
    .C(_338_),
    .D(ABH[7]),
    .Y(_486_)
);

NAND3X1 _2350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .B(_1480_),
    .C(_1479_),
    .Y(_1481_)
);

FILL FILL_4__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1614_),
    .C(RDY_bF$buf2),
    .Y(_1635_)
);

FILL FILL_6__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_767_),
    .C(_771_),
    .Y(_96_)
);

FILL FILL_1__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_1219__bF$buf2),
    .C(_527_),
    .Y(_31_)
);

OAI22X1 _2406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_138_),
    .C(_1051__bF$buf3),
    .D(_1144_),
    .Y(_161_)
);

FILL FILL_1__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _3364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[0]),
    .B(ADD[3]),
    .Y(_1642_)
);

FILL FILL_6__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .Y(_994_)
);

FILL FILL_8_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_356_),
    .C(_362_),
    .Y(_363_)
);

INVX1 _2215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .Y(_1350_)
);

FILL FILL_2__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[8]),
    .Y(AB[8])
);

FILL FILL_6__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_916_),
    .C(_794_),
    .Y(_805_)
);

FILL FILL_2__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_1050_)
);

FILL FILL_7__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1314_),
    .C(_509_),
    .Y(_561_)
);

FILL FILL_6__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_121_),
    .C(_884_),
    .Y(_195_)
);

NAND2X1 _2024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf3),
    .B(IRHOLD[6]),
    .Y(_1160_)
);

FILL FILL_2__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[14]),
    .B(_830__bF$buf1),
    .Y(_847_)
);

FILL FILL_1__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .Y(_868_)
);

FILL FILL_4__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181350x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_391_),
    .Y(_397_)
);

NAND2X1 _2253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(_1386_),
    .Y(_1387_)
);

FILL FILL_2__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_1542_),
    .C(_1543_),
    .Y(_1544_)
);

FILL FILL_6__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_698_),
    .Y(_701_)
);

FILL FILL_7__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_944_),
    .C(_1084_),
    .Y(_1085_)
);

FILL FILL_5__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[3]),
    .B(_446_),
    .C(_448_),
    .Y(_449_)
);

OAI21X1 _2309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(_1175_),
    .C(_1142_),
    .Y(_1442_)
);

FILL FILL_7__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(ADD[3]),
    .C(_229_),
    .Y(_230_)
);

NOR2X1 _2062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(write_back),
    .B(_853__bF$buf7),
    .Y(_1198_)
);

FILL FILL_2__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3267_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_29_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf6),
    .Q(sei)
);

FILL FILL_6__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_892_),
    .Y(_906_)
);

FILL FILL_4__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf4),
    .B(_1259_),
    .C(_1002__bF$buf2),
    .Y(_629_)
);

NAND2X1 _2538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[3]),
    .B(_199_),
    .Y(_278_)
);

NOR2X1 _2118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf3),
    .B(_1220_),
    .Y(_1254_)
);

FILL FILL_7__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf2),
    .B(_1037_),
    .Y(_1424_)
);

FILL FILL_2__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .B(_1562_),
    .Y(_1582_)
);

FILL FILL_6__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _3076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(ADD[6]),
    .Y(_734_)
);

FILL FILL_2__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(_945_),
    .Y(_961_)
);

FILL FILL_7__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1118_),
    .B(_872_),
    .Y(_1119_)
);

FILL FILL_8__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_481_),
    .C(_483_),
    .Y(_484_)
);

AOI21X1 _2347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1206_),
    .C(_1289_),
    .Y(_1478_)
);

FILL FILL_7__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_933_),
    .Y(_943_)
);

FILL FILL_5__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .B(_661_),
    .C(_663_),
    .Y(_664_)
);

INVX1 _2576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adc_bcd),
    .Y(_310_)
);

NOR2X1 _2156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1280_),
    .B(_1291_),
    .Y(_1292_)
);

FILL FILL_7__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_989_),
    .C(_990_),
    .Y(_991_)
);

FILL FILL_7__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[0]),
    .B(_139_),
    .C(_143_),
    .Y(_144_)
);

FILL FILL184050x171750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x113250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .Y(_1329_)
);

FILL FILL_2__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_1671_),
    .C(_1668_),
    .Y(_1673_)
);

FILL FILL183450x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_954_),
    .Y(_1029_)
);

FILL FILL_8__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _1694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf1),
    .Y(_853_)
);

FILL FILL_8__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1303_),
    .B(_1314_),
    .Y(_585_)
);

NAND2X1 _2479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_226_),
    .Y(_227_)
);

OAI21X1 _2059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_900_),
    .B(_935_),
    .C(_926__bF$buf0),
    .Y(_1195_)
);

FILL FILL_0__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[4]),
    .B(_1674_),
    .C(_1505_),
    .Y(_1506_)
);

MUX2X1 _3000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(AZ),
    .S(plp),
    .Y(_667_)
);

FILL FILL_4__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1039_),
    .C(_1253_),
    .D(_1352_),
    .Y(_1421_)
);

FILL FILL_0__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1113_),
    .B(_1115_),
    .C(_1114_),
    .Y(_1116_)
);

FILL FILL_2__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .Y(_603_)
);

INVX1 _2500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .Y(_1685_[5])
);

FILL FILL_5__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1232_),
    .Y(_1233_)
);

FILL FILL_0__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_939_),
    .B(_937_),
    .Y(_940_)
);

FILL FILL_4__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1677_),
    .Y(_1600_)
);

FILL FILL_1__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3323_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_77_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[1] [0])
);

FILL FILL_1__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf0),
    .B(_1569_),
    .C(_1632_),
    .Y(_1491_)
);

FILL FILL_6__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [2]),
    .B(_767_),
    .Y(_770_)
);

FILL FILL_2__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(_1296_),
    .C(_1298_),
    .Y(_525_)
);

AOI21X1 _2403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[3]),
    .B(_139_),
    .C(_158_),
    .Y(_159_)
);

FILL FILL_1__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3361_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_114_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(ABH[5])
);

FILL FILL_2__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_359_),
    .C(_1051__bF$buf1),
    .Y(_360_)
);

NOR2X1 _2212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf1),
    .B(_1032_),
    .Y(_1347_)
);

FILL FILL_2__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_1500_),
    .C(_1657_),
    .Y(_1503_)
);

FILL FILL_1__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[5]),
    .Y(AB[5])
);

FILL FILL_6__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_787_),
    .Y(_802_)
);

FILL FILL_2__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1028_),
    .B(_1046_),
    .Y(_1047_)
);

FILL FILL_0__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_1219__bF$buf1),
    .C(_557_),
    .D(_559_),
    .Y(_34_)
);

FILL FILL_6__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_1238_),
    .C(_1363_),
    .Y(_192_)
);

NAND2X1 _2021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf1),
    .B(IRHOLD[7]),
    .Y(_1157_)
);

FILL FILL_8_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_830__bF$buf2),
    .C(_845_),
    .Y(_113_)
);

FILL FILL_1__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .Y(_865_)
);

FILL FILL_0__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_587_),
    .C(_1438_),
    .Y(_601_)
);

FILL FILL_1__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_321_),
    .C(_393_),
    .Y(_394_)
);

NAND2X1 _2250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_1173_),
    .Y(_1384_)
);

FILL FILL_2__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_1540_),
    .C(_1652_),
    .D(_1539_),
    .Y(_1541_)
);

FILL FILL_6__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adj_bcd),
    .B(_310_),
    .Y(_698_)
);

FILL FILL_2__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1079_),
    .B(_1081_),
    .C(_1080_),
    .Y(_1082_)
);

FILL FILL_5__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf3),
    .B(_1259_),
    .C(_320_),
    .Y(_446_)
);

NAND3X1 _2306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(_1438_),
    .C(_1386_),
    .Y(_1439_)
);

FILL FILL_7__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3264_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_26_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf5),
    .Q(cld)
);

FILL FILL_6__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_902_),
    .B(_895_),
    .Y(_903_)
);

FILL FILL_6__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[7]),
    .Y(_628_)
);

FILL FILL_6__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(DIMUX[2]),
    .C(_275_),
    .Y(_276_)
);

OAI21X1 _2115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1250_),
    .B(_1190_),
    .C(RDY_bF$buf6),
    .Y(_1251_)
);

FILL FILL_2__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1535_),
    .B(_1537_),
    .C(_1538_),
    .Y(_1579_)
);

FILL FILL_6__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[5]),
    .B(_1281_),
    .C(_731_),
    .D(_729_),
    .Y(_732_)
);

FILL FILL_2__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(_957_),
    .Y(_958_)
);

FILL FILL_7__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_480_),
    .C(_460_),
    .Y(_481_)
);

NAND3X1 _2344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1421_),
    .B(_1255_),
    .C(_1474_),
    .Y(_1475_)
);

FILL FILL_5__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[2]),
    .B(_1649__bF$buf2),
    .Y(_1631_)
);

OAI21X1 _3129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_767_),
    .C(_768_),
    .Y(_93_)
);

FILL FILL_7__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_1008_),
    .C(_660_),
    .Y(_661_)
);

FILL FILL_6__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .Y(_309_)
);

OAI21X1 _2153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf2),
    .B(_894_),
    .C(_1288_),
    .Y(_1289_)
);

FILL FILL_2__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3358_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_111_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf7),
    .Q(ABH[2])
);

FILL FILL_0__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_914_),
    .Y(_988_)
);

FILL FILL_6__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf5),
    .B(_357_),
    .C(_351_),
    .Y(_4_)
);

NOR2X1 _2209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1343_),
    .Y(_1344_)
);

FILL FILL_7__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_138_),
    .C(_1051__bF$buf3),
    .Y(_141_)
);

FILL FILL_8__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[2]),
    .Y(AB[2])
);

FILL FILL_6__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_797_),
    .B(_315_),
    .C(_798_),
    .Y(_799_)
);

FILL FILL_7__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_556_),
    .Y(_557_)
);

FILL FILL_6__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .B(_188_),
    .Y(_189_)
);

OAI21X1 _2018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf0),
    .B(_861_),
    .C(_1153_),
    .Y(_1154_)
);

FILL FILL_7__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1254_),
    .Y(_1326_)
);

FILL FILL_2__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_1669_),
    .Y(_1670_)
);

FILL FILL_0__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .Y(DIMUX[6])
);

FILL FILL_4__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1025_),
    .Y(_1026_)
);

FILL FILL_8__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_391_),
    .Y(_392_)
);

NAND2X1 _2247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1351_),
    .Y(_1381_)
);

FILL FILL_7__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [3]),
    .B(_1022_),
    .Y(_1079_)
);

FILL FILL_7__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIHOLD[1]),
    .Y(_851_)
);

FILL FILL_8__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1330_),
    .C(_1176_),
    .Y(_583_)
);

FILL FILL_6__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .Y(_224_)
);

INVX1 _2056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .Y(_1192_)
);

FILL FILL_0__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_899_),
    .Y(_900_)
);

FILL FILL_4__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1418_),
    .B(_1271_),
    .Y(_1419_)
);

FILL FILL_2__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [7]),
    .B(_1022_),
    .Y(_1113_)
);

FILL FILL_4__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_1227_),
    .C(_1229_),
    .Y(_1230_)
);

FILL FILL_2__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3299_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_53_),
    .CLK(clk_bF$buf0),
    .Q(IRHOLD[0])
);

FILL FILL_0__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_936_),
    .C(_934_),
    .Y(_937_)
);

FILL FILL_4__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1683_),
    .B(_1596_),
    .C(_1498_),
    .Y(_1597_)
);

FILL FILL_3__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_507_),
    .C(_505_),
    .Y(_24_)
);

NAND2X1 _2379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf3),
    .B(_927_),
    .Y(_138_)
);

FILL FILL_8__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3320_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_74_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[0] [5])
);

FILL FILL_4__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1172_),
    .Y(_1323_)
);

FILL FILL_0__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1018_),
    .B(_1019_),
    .C(_1004_),
    .Y(_1023_)
);

INVX1 _2820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .Y(_523_)
);

OAI21X1 _2400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[11]),
    .Y(_156_)
);

FILL FILL_0__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIHOLD[0]),
    .Y(_849_)
);

FILL FILL_4__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(BI[4]),
    .Y(_1500_)
);

FILL FILL_1__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf2),
    .B(_936_),
    .Y(_1044_)
);

FILL FILL_0__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[11]),
    .B(_830__bF$buf0),
    .Y(_844_)
);

FILL FILL_1__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(dst_reg[0]),
    .Y(_598_)
);

FILL FILL181050x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1663_),
    .B(_1537_),
    .C(_1535_),
    .Y(_1538_)
);

FILL FILL_6__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [0]),
    .B(_693_),
    .Y(_696_)
);

FILL FILL_2__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf5),
    .B(_443_),
    .C(_433_),
    .Y(_12_)
);

NOR2X1 _2303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1429_),
    .B(_1435_),
    .Y(_1436_)
);

FILL FILL_0__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1504_),
    .B(_1506_),
    .C(_1588_),
    .D(_1593_),
    .Y(_1594_)
);

FILL FILL_1__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3261_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_23_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf5),
    .Q(php)
);

FILL FILL_6__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_620_),
    .C(_626_),
    .Y(_58_)
);

FILL FILL_6__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[2]),
    .Y(_273_)
);

AND2X2 _2112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1234_),
    .Y(_1248_)
);

FILL FILL_2__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3317_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_71_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[0] [2])
);

FILL FILL_1__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1575_),
    .Y(_1576_)
);

FILL FILL_6__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_728_),
    .Y(_729_)
);

FILL FILL_2__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_909_),
    .Y(_955_)
);

FILL FILL_4__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .B(_325_),
    .C(_338_),
    .D(ABH[6]),
    .Y(_478_)
);

OAI21X1 _2341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf2),
    .B(_1471_),
    .C(_1376_),
    .Y(_1472_)
);

FILL FILL_5__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1629_),
    .C(_1626_),
    .Y(_1488_)
);

FILL FILL_6__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_757_),
    .C(_766_),
    .Y(_92_)
);

FILL FILL_1__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1162_),
    .Y(_520_)
);

FILL FILL_1__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_1022_),
    .C(_657_),
    .Y(_658_)
);

FILL FILL_6__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_240_),
    .C(_305_),
    .Y(_306_)
);

OAI21X1 _2150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_978_),
    .C(_1285_),
    .Y(_1286_)
);

FILL FILL_2__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3355_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_108_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(ABL[7])
);

FILL FILL_0__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf9)
);

FILL FILL_2__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_984_),
    .B(_964_),
    .Y(_985_)
);

FILL FILL_6__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[2]),
    .B(_321_),
    .C(_354_),
    .Y(_355_)
);

XOR2X1 _2206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1340_),
    .B(cond_code[0]),
    .Y(_1341_)
);

FILL FILL_7__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[13]),
    .Y(AB[13])
);

FILL FILL_6__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_794_),
    .Y(_796_)
);

FILL FILL_2__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_553_),
    .C(_552_),
    .Y(_554_)
);

FILL FILL_6__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(_1052_),
    .Y(_186_)
);

NAND2X1 _2015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf3),
    .B(IRHOLD[4]),
    .Y(_1151_)
);

FILL FILL_2__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1662_),
    .B(_1663_),
    .C(_1659_),
    .Y(_1667_)
);

FILL FILL_2__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .Y(DIMUX[5])
);

FILL FILL_4__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_343_),
    .C(_388_),
    .Y(_389_)
);

NOR2X1 _2244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1377_),
    .B(_1375_),
    .Y(_1378_)
);

FILL FILL_2__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _3449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1524_),
    .B(_1657_),
    .C(_1531_),
    .D(_1534_),
    .Y(_1535_)
);

NAND2X1 _3029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_1020_),
    .Y(_693_)
);

FILL FILL_7__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_944_),
    .C(_1076_),
    .Y(_1077_)
);

FILL FILL_7__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(index_y),
    .Y(_580_)
);

FILL FILL_6__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(_208_),
    .C(_221_),
    .Y(_222_)
);

OAI21X1 _2053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1189_)
);

FILL FILL_2__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3258_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_20_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf6),
    .Q(cond_code[1])
);

FILL FILL_6__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_896_),
    .Y(_897_)
);

FILL FILL_4__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[4]),
    .Y(_625_)
);

AOI21X1 _2529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(DIMUX[1]),
    .C(_270_),
    .Y(_271_)
);

OAI21X1 _2109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_996_),
    .C(RDY_bF$buf7),
    .Y(_1245_)
);

FILL FILL_7__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .Y(_1416_)
);

FILL FILL_2__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1570_),
    .B(_1547_),
    .Y(_1573_)
);

FILL FILL_6__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adj_bcd),
    .B(adc_bcd),
    .C(CO),
    .Y(_726_)
);

FILL FILL_0__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_944_),
    .C(_1110_),
    .Y(_1111_)
);

FILL FILL_4__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_445_),
    .Y(_475_)
);

AND2X2 _2338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(_1128_),
    .Y(_1469_)
);

FILL FILL_7__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf1),
    .B(_955_),
    .Y(_1227_)
);

FILL FILL_2__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3296_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[6]),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf9),
    .Q(DIHOLD[6])
);

FILL FILL_6__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf1),
    .B(_928_),
    .Y(_934_)
);

FILL FILL_5__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(I),
    .B(_651_),
    .Y(_656_)
);

FILL FILL_6__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[15]),
    .Y(_303_)
);

OAI21X1 _2147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf2),
    .B(_1281_),
    .C(_1282_),
    .Y(_1283_)
);

FILL FILL_7__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_938_),
    .C(_981_),
    .Y(_982_)
);

FILL FILL_7__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf0),
    .C(clc),
    .Y(_505_)
);

NAND2X1 _2376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_133_),
    .Y(_1687_)
);

FILL FILL_8__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .Y(_1320_)
);

FILL FILL_0__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(_1018_),
    .C(_1016_),
    .Y(_1020_)
);

FILL FILL_0__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[7]),
    .Y(DO[7])
);

FILL FILL_3__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830__bF$buf1),
    .Y(_831_)
);

FILL FILL_0__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[5]),
    .B(_1674_),
    .C(_1684_),
    .Y(_1497_)
);

FILL FILL_3__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_191_),
    .C(_969_),
    .Y(_421_)
);

AOI21X1 _2279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_878_),
    .B(_1409_),
    .C(_1412_),
    .Y(_1413_)
);

FILL FILL_0__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[10]),
    .B(_830__bF$buf0),
    .Y(_842_)
);

FILL FILL_2__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1400_),
    .B(_595_),
    .C(_594_),
    .Y(_596_)
);

FILL FILL_3__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .Y(_926__bF$buf3)
);

FILL FILL_9__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .Y(_926__bF$buf2)
);

FILL FILL_3__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .Y(_926__bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926_),
    .Y(_926__bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf8)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf7)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf6)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf5)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf4)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf3)
);

FILL FILL_3__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf1),
    .B(_1035_),
    .Y(_1224_)
);

FILL FILL_0__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[0]),
    .Y(_931_)
);

FILL FILL_4__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_440_),
    .C(_439_),
    .Y(_441_)
);

OAI21X1 _2300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf2),
    .B(_1260_),
    .C(_1432_),
    .Y(_1433_)
);

FILL FILL_0__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .Y(_1591_)
);

FILL FILL_1__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3314_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_68_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf9),
    .Q(backwards)
);

FILL FILL_1__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .Y(_952_)
);

FILL FILL_0__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1571_),
    .B(_1559_),
    .C(_1553_),
    .Y(_1627_)
);

FILL FILL_6__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf3),
    .B(_758_),
    .C(\AXYS[2] [6]),
    .Y(_765_)
);

FILL FILL_1__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_1002__bF$buf3),
    .C(sei),
    .Y(_518_)
);

FILL FILL_1__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3352_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_105_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(ABL[4])
);

FILL FILL_2__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(res),
    .B(_1132_),
    .Y(_352_)
);

OAI21X1 _2203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1337_),
    .C(cond_code[1]),
    .Y(_1338_)
);

FILL FILL_9__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_1679_),
    .C(_1657_),
    .Y(_1682_)
);

FILL FILL_1__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[10]),
    .Y(AB[10])
);

FILL FILL_6__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_941_),
    .C(_792_),
    .Y(_793_)
);

FILL FILL_2__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_550_),
    .Y(_551_)
);

FILL FILL_6__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf1),
    .B(_953_),
    .Y(_183_)
);

NAND2X1 _2012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1147_),
    .Y(_1148_)
);

FILL FILL_2__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1055_),
    .B(_830__bF$buf3),
    .C(_840_),
    .Y(_109_)
);

FILL FILL_1__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.BI7 ),
    .B(_1649__bF$buf0),
    .Y(_1665_)
);

FILL FILL_8__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .Y(DIMUX[4])
);

FILL FILL_4__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .B(_1384_),
    .C(_1129__bF$buf3),
    .Y(_593_)
);

FILL FILL_1__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[6]),
    .Y(_386_)
);

INVX1 _2241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1374_),
    .Y(_1375_)
);

FILL FILL_2__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .Y(_1532_)
);

FILL FILL_6__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .Y(_690_)
);

FILL FILL_7__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1073_),
    .Y(_1074_)
);

FILL FILL_0__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_1267_),
    .C(_1051__bF$buf3),
    .Y(_438_)
);

FILL FILL_7__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .B(_1382_),
    .Y(_578_)
);

FILL FILL_8__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .C(ADD[2]),
    .Y(_219_)
);

NAND2X1 _2050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf0),
    .B(_910_),
    .Y(_1186_)
);

FILL FILL_2__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3255_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(NMI),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(NMI_1)
);

FILL FILL183450x171750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf3),
    .B(_893_),
    .Y(_894_)
);

FILL FILL_6__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_620_),
    .C(_623_),
    .Y(_55_)
);

FILL FILL_6__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .Y(_268_)
);

OAI21X1 _2106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1238_),
    .C(_1241_),
    .Y(_1242_)
);

FILL FILL_7__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1548_),
    .Y(_1570_)
);

FILL FILL_6__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[4]),
    .B(_981_),
    .C(_723_),
    .Y(_724_)
);

FILL FILL_2__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[6]),
    .Y(_1108_)
);

NAND2X1 _2755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[12]),
    .B(_323_),
    .Y(_472_)
);

AND2X2 _2335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1466_),
    .B(_1301_),
    .Y(_1467_)
);

FILL FILL_5__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3293_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[3]),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf9),
    .Q(DIHOLD[3])
);

FILL FILL_2__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_951_),
    .C(_649_),
    .Y(_653_)
);

FILL FILL_6__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1108_),
    .B(_268_),
    .C(_300_),
    .Y(_301_)
);

NAND3X1 _2144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1276_),
    .B(_1273_),
    .C(_1279_),
    .Y(_1280_)
);

FILL FILL_2__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3349_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_102_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(ABL[1])
);

FILL FILL_0__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(_977_),
    .C(_978_),
    .Y(_979_)
);

FILL FILL_6__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf0)
);

BUFX2 BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .Y(_1002__bF$buf4)
);

BUFX2 BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .Y(_1002__bF$buf3)
);

BUFX2 BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .Y(_1002__bF$buf2)
);

BUFX2 BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .Y(_1002__bF$buf1)
);

BUFX2 BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .Y(_1002__bF$buf0)
);

BUFX2 BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .Y(_882__bF$buf3)
);

FILL FILL183150x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .Y(_882__bF$buf2)
);

BUFX2 BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .Y(_882__bF$buf1)
);

BUFX2 BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .Y(_882__bF$buf0)
);

FILL FILL_3__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .Y(_503_)
);

NOR2X1 _2373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .B(_130_),
    .Y(_133_)
);

FILL FILL_8__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3578_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1496_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf9),
    .Q(\u_ALU8.AI7 )
);

FILL FILL_6__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1049_),
    .B(_990_),
    .C(_789_),
    .Y(_790_)
);

FILL FILL_7__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_547_),
    .Y(_548_)
);

INVX1 _2429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .Y(_180_)
);

OAI21X1 _2009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1143_),
    .B(NMI_edge),
    .C(_1144_),
    .Y(_1145_)
);

FILL FILL_7__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1316_),
    .Y(_1317_)
);

FILL FILL_2__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[7]),
    .C(_1661_),
    .Y(_1662_)
);

FILL FILL_0__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1005_),
    .B(_1009_),
    .Y(_1017_)
);

FILL FILL_2__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_367_),
    .C(RDY_bF$buf4),
    .Y(_384_)
);

NAND2X1 _2238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1370_),
    .B(_1371_),
    .Y(_1372_)
);

FILL FILL_7__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_827_),
    .C(_825_),
    .D(_818_),
    .Y(_828_)
);

FILL FILL_6__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [2]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [2]),
    .Y(_1071_)
);

FILL FILL_7__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf0),
    .B(_1178_),
    .Y(_575_)
);

FILL FILL_6__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_208_),
    .C(_216_),
    .Y(_217_)
);

INVX1 _2047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1182_),
    .Y(_1183_)
);

FILL FILL_7__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .Y(_891_)
);

FILL FILL_4__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_418_),
    .B(_412_),
    .C(RDY_bF$buf8),
    .Y(_419_)
);

OAI21X1 _2276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf2),
    .B(_880_),
    .C(_853__bF$buf2),
    .Y(_1410_)
);

FILL FILL_2__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [6]),
    .B(_1020_),
    .Y(_1105_)
);

FILL FILL_7__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1150_),
    .Y(_1221_)
);

FILL FILL_5_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_928_),
    .B(_927_),
    .C(_926__bF$buf1),
    .Y(_929_)
);

FILL FILL_4__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_1569_),
    .C(_1587_),
    .Y(_1588_)
);

FILL FILL_3__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf0),
    .B(_748_),
    .C(\AXYS[1] [3]),
    .Y(_752_)
);

FILL FILL_0__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3311_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_65_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf5),
    .Q(N)
);

FILL FILL_3__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x78150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_329_),
    .C(_324_),
    .Y(_330_)
);

AND2X2 _2179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1147_),
    .B(_1145_),
    .Y(_1314_)
);

FILL FILL_0__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_1649__bF$buf3),
    .Y(_1625_)
);

FILL FILL_6__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_757_),
    .C(_763_),
    .Y(_89_)
);

FILL FILL_2__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1163_),
    .Y(_516_)
);

FILL FILL_0__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_349_),
    .Y(_350_)
);

AND2X2 _2200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[2]),
    .B(Z),
    .Y(_1335_)
);

FILL FILL_4__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(BI[5]),
    .Y(_1679_)
);

FILL FILL_1__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[7]),
    .Y(_839_)
);

FILL FILL_1__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x31350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .Y(DIMUX[3])
);

FILL FILL_0__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .Y(_591_)
);

FILL FILL_1__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1675_),
    .Y(_1529_)
);

FILL FILL_6__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_633_),
    .Y(_687_)
);

FILL FILL_2__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_1002__bF$buf4),
    .C(_1145_),
    .Y(_435_)
);

FILL FILL_5__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3252_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_15_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(PC[13])
);

FILL FILL_2__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[1]),
    .Y(_622_)
);

FILL FILL_6__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_262_),
    .C(_265_),
    .Y(_266_)
);

NAND2X1 _2103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf0),
    .B(_1037_),
    .Y(_1239_)
);

FILL FILL184050x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3308_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_62_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf9),
    .Q(V)
);

FILL FILL_1__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .Y(_1567_)
);

FILL FILL_6__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [3]),
    .B(_693_),
    .Y(_722_)
);

FILL FILL_2__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_460_),
    .Y(_470_)
);

NAND3X1 _2332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1276_),
    .C(_1243_),
    .Y(_1464_)
);

FILL FILL_5__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .B(_1619_),
    .C(_1610_),
    .Y(_1623_)
);

OAI21X1 _3117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf3),
    .B(_758_),
    .C(\AXYS[2] [3]),
    .Y(_762_)
);

FILL FILL_1__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3290_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[0]),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(DIHOLD[0])
);

FILL FILL_2__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(sed),
    .Y(_514_)
);

FILL FILL_1__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_978_),
    .C(_632_),
    .Y(_650_)
);

FILL FILL_6__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_208_),
    .C(_298_),
    .Y(_1685_[13])
);

INVX1 _2141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_990_),
    .Y(_1277_)
);

FILL FILL_2__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3346_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_99_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[3] [6])
);

FILL FILL_6__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x171750 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf0),
    .B(_926__bF$buf1),
    .C(_953_),
    .Y(_976_)
);

FILL FILL_0__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_343_),
    .C(_346_),
    .Y(_347_)
);

FILL FILL_1__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf1)
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf0)
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .Y(_886__bF$buf3)
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .Y(_886__bF$buf2)
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .Y(_886__bF$buf1)
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .Y(_886__bF$buf0)
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .Y(_1649__bF$buf3)
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .Y(_1649__bF$buf2)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .Y(_1649__bF$buf1)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .Y(_1649__bF$buf0)
);

FILL FILL_3__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_1159_),
    .C(_501_),
    .Y(_21_)
);

OAI21X1 _2370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_120_),
    .C(_131_),
    .Y(alu_op[2])
);

FILL FILL_8__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3575_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1493_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf4),
    .Q(ADD[5])
);

FILL FILL_6__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .Y(_787_)
);

FILL FILL_2__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_544_),
    .C(_543_),
    .Y(_545_)
);

FILL FILL_6__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_128_),
    .C(_177_),
    .Y(_178_)
);

OAI21X1 _2006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf2),
    .B(DIMUX[3]),
    .C(_1141_),
    .Y(_1142_)
);

FILL FILL_7__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1658_),
    .B(_1656_),
    .C(_1650_),
    .Y(_1659_)
);

FILL FILL_6__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(src_reg[1]),
    .Y(_1014_)
);

FILL FILL_2__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[5]),
    .B(_336_),
    .Y(_381_)
);

NAND3X1 _2235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_943_),
    .C(_1341_),
    .Y(_1369_)
);

FILL FILL_3_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_824_),
    .Y(_825_)
);

FILL FILL_2__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[1]),
    .C(_1068_),
    .Y(_1069_)
);

FILL FILL_7__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf0),
    .B(_521_),
    .C(_573_),
    .Y(_43_)
);

FILL FILL_6__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .C(ADD[1]),
    .Y(_214_)
);

OAI21X1 _2044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1177_),
    .B(_1179_),
    .C(_1176_),
    .Y(_1180_)
);

FILL FILL_2__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3249_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_12_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[10])
);

FILL FILL_7__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .Y(_888_)
);

FILL FILL_4__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[8]),
    .B(_415_),
    .C(_414_),
    .Y(_416_)
);

NAND3X1 _2273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1406_),
    .C(_1398_),
    .Y(_1407_)
);

FILL FILL_2__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(_1529_),
    .Y(_1564_)
);

FILL FILL_6__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_717_),
    .B(_718_),
    .Y(_719_)
);

FILL FILL_0__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1099_),
    .C(_1102_),
    .Y(AI[5])
);

FILL FILL_4__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_464_),
    .Y(_467_)
);

NAND3X1 _2329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1374_),
    .B(_1204_),
    .C(_1411_),
    .Y(_1461_)
);

FILL FILL_7__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1044_),
    .C(_1217_),
    .D(_1129__bF$buf4),
    .Y(_1218_)
);

FILL FILL_5_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3287_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_49_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf1),
    .Q(dst_reg[0])
);

FILL FILL_6__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[5]),
    .B(_917_),
    .Y(_926_)
);

FILL FILL_4__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _2978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[3]),
    .B(_647_),
    .S(_1260_),
    .Y(_648_)
);

FILL FILL_6__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[5]),
    .B(_1075_),
    .C(_295_),
    .Y(_296_)
);

INVX1 _2138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_1274_)
);

FILL FILL_7__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_747_),
    .C(_750_),
    .Y(_78_)
);

FILL FILL_2__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_933_),
    .C(_863_),
    .D(_967_),
    .Y(BI[6])
);

FILL FILL_7__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[1]),
    .B(_853__bF$buf7),
    .Y(_500_)
);

NOR2X1 _2367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1353_),
    .Y(_129_)
);

FILL FILL_7__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(ABL[0]),
    .Y(_327_)
);

NOR2X1 _2176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1310_),
    .Y(_1311_)
);

FILL FILL_2__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .B(src_reg[0]),
    .S(_1006_),
    .Y(_1011_)
);

FILL FILL_7__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .B(BI[6]),
    .C(_1675_),
    .Y(_1676_)
);

FILL FILL_3__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_245_),
    .C(_837_),
    .Y(_106_)
);

FILL FILL_3__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_587_),
    .C(_549_),
    .Y(_588_)
);

FILL FILL_3__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1098_),
    .B(_182_),
    .C(_244_),
    .Y(_245_)
);

NAND2X1 _2079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_1173_),
    .Y(_1215_)
);

FILL FILL_0__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1525_),
    .Y(_1526_)
);

FILL FILL_6__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(backwards),
    .Y(_685_)
);

FILL FILL_2__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_267_),
    .C(_432_),
    .D(_428_),
    .Y(_11_)
);

FILL FILL_0__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf2),
    .B(DIMUX[1]),
    .C(_1134_),
    .Y(_1135_)
);

FILL FILL_2__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .Y(_620_)
);

FILL FILL_8__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[0]),
    .Y(_263_)
);

NAND2X1 _2100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1039_),
    .Y(_1236_)
);

FILL FILL_9__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3305_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_59_),
    .CLK(clk_bF$buf5),
    .Q(IRHOLD[6])
);

FILL FILL_1__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1598_),
    .Y(_1620_)
);

OAI21X1 _3114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_757_),
    .C(_760_),
    .Y(_86_)
);

FILL FILL_1__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1303_),
    .Y(_512_)
);

FILL FILL_1__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3343_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_96_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[3] [3])
);

FILL FILL_6__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[1]),
    .B(_338_),
    .Y(_344_)
);

FILL FILL_1__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf7)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf6)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf5)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf4)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf3)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf2)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf1)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf0)
);

FILL FILL_3__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3572_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1490_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf3),
    .Q(ADD[2])
);

FILL FILL_6__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_917_),
    .C(_893_),
    .Y(_784_)
);

FILL FILL_2__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_541_),
    .C(_1350_),
    .Y(_542_)
);

FILL FILL_6__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1116_),
    .Y(_175_)
);

NAND2X1 _2003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .B(_1138_),
    .Y(_1139_)
);

FILL FILL_5__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[4]),
    .Y(_836_)
);

FILL FILL_1__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[7]),
    .C(_1655_),
    .D(_1652_),
    .Y(_1656_)
);

FILL FILL_6__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_343_),
    .C(_377_),
    .Y(_378_)
);

OAI21X1 _2232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_918__bF$buf0),
    .C(_1365_),
    .Y(_1366_)
);

FILL FILL_2__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .Y(_1523_)
);

OAI21X1 _3017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1260_),
    .B(_681_),
    .C(_682_),
    .Y(_683_)
);

FILL FILL_1__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _3190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_935_),
    .Y(_822_)
);

FILL FILL_2__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1065_),
    .B(_872_),
    .Y(_1066_)
);

FILL FILL_0__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_416_),
    .C(_426_),
    .D(_429_),
    .Y(_430_)
);

FILL FILL_7__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1323_),
    .B(_551_),
    .C(_571_),
    .D(_498_),
    .Y(_572_)
);

FILL FILL_6__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_208_),
    .C(_211_),
    .Y(_212_)
);

NAND2X1 _2041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .B(_1148_),
    .Y(_1177_)
);

FILL FILL_2__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3246_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_9_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf7),
    .Q(PC[7])
);

FILL FILL_7__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_872_),
    .Y(_885_)
);

FILL FILL_6__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf4),
    .B(res),
    .Y(_52_)
);

INVX1 _2517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[8]),
    .Y(_260_)
);

FILL FILL_1__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf1),
    .B(_882__bF$buf3),
    .C(_946_),
    .D(_916_),
    .Y(_413_)
);

AOI21X1 _2270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1164_),
    .C(_1217_),
    .Y(_1404_)
);

FILL FILL_2__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(_1535_),
    .Y(_1561_)
);

FILL FILL_6__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .Y(_716_)
);

FILL FILL_2__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[5]),
    .B(_1075_),
    .Y(_1100_)
);

OAI21X1 _2746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_333_),
    .C(_1100_),
    .Y(_464_)
);

OAI21X1 _2326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1437_),
    .C(_1458_),
    .Y(_1483_[3])
);

FILL FILL_7__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3284_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_46_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf6),
    .Q(index_y)
);

FILL FILL_6__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rotate),
    .B(_922_),
    .C(_919_),
    .Y(_923_)
);

FILL FILL184350x19650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(D),
    .B(_644_),
    .Y(_645_)
);

FILL FILL_6__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[5]),
    .Y(_293_)
);

NOR3X1 _2135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1270_),
    .C(_1258_),
    .Y(_1271_)
);

FILL FILL_0__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf2),
    .B(_748_),
    .C(\AXYS[1] [0]),
    .Y(_749_)
);

FILL FILL_2__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[5]),
    .Y(_973_)
);

FILL FILL_7__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .Y(_498_)
);

INVX1 _2364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .Y(_126_)
);

FILL FILL_8__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3569_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1487_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf0),
    .Q(HC)
);

OAI21X1 _3149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_917_),
    .C(_927_),
    .Y(_781_)
);

FILL FILL_7__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x160050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .Y(_324_)
);

NAND2X1 _2173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1307_),
    .B(_1301_),
    .Y(_1308_)
);

FILL FILL_2__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .Y(_1653_)
);

FILL FILL_6__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf2),
    .Y(_1008_)
);

FILL FILL_6__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .Y(_375_)
);

INVX1 _2229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1228_),
    .Y(_1363_)
);

FILL FILL_7__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .Y(_819_)
);

FILL FILL_0__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_566_),
    .C(_568_),
    .Y(_41_)
);

FILL FILL_6__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .C(ADD[0]),
    .Y(_209_)
);

INVX1 _2038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .Y(_1174_)
);

FILL FILL_7__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_881_),
    .Y(_882_)
);

FILL FILL_4__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_409_),
    .Y(_410_)
);

NAND2X1 _2267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1400_),
    .Y(_1401_)
);

FILL FILL_7__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [5]),
    .B(_1020_),
    .Y(_1097_)
);

FILL FILL_7__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[5]),
    .B(_199_),
    .C(_241_),
    .Y(_242_)
);

AND2X2 _2076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1211_),
    .B(_1197_),
    .Y(_1212_)
);

FILL FILL_2__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(compare),
    .Y(_920_)
);

FILL FILL_4__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x152250 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(NMI_edge),
    .Y(_1132_)
);

FILL FILL_8__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3302_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_56_),
    .CLK(clk_bF$buf10),
    .Q(IRHOLD[3])
);

FILL FILL_3__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(_1615_),
    .Y(_1617_)
);

OAI21X1 _3111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf2),
    .B(_758_),
    .C(\AXYS[2] [0]),
    .Y(_759_)
);

FILL FILL_2__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_509_),
    .Y(_510_)
);

FILL FILL_0__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1082_),
    .Y(_155_)
);

FILL FILL_8__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3340_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_93_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[3] [0])
);

FILL FILL_6__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_341_),
    .Y(_342_)
);

FILL FILL_0__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .Y(_1043_)
);

FILL FILL182250x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_539_),
    .C(_1159_),
    .Y(_540_)
);

FILL FILL_6__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_128_),
    .C(_172_),
    .Y(_173_)
);

INVX1 _2000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD[0]),
    .Y(_1136_)
);

FILL FILL_5__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_223_),
    .C(_834_),
    .Y(_103_)
);

FILL FILL_1__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(alu_shift_right),
    .Y(_1520_)
);

NAND2X1 _3014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(_673_),
    .Y(_680_)
);

FILL FILL_1__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1060_),
    .B(_1062_),
    .C(_1061_),
    .Y(_1063_)
);

FILL FILL_0__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_324_),
    .C(_426_),
    .Y(_427_)
);

FILL FILL_5__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3243_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_6_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(PC[4])
);

FILL FILL_2__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_615_),
    .C(_614_),
    .Y(_616_)
);

OAI21X1 _2514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_208_),
    .C(_257_),
    .Y(_258_)
);

FILL FILL_1__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1556_),
    .Y(_1558_)
);

FILL FILL_6__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[2]),
    .B(_1281_),
    .C(_713_),
    .D(_711_),
    .Y(_714_)
);

FILL FILL_2__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_461_),
    .Y(_462_)
);

NOR2X1 _2323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1308_),
    .B(_1455_),
    .Y(_1456_)
);

FILL FILL_5__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1613_),
    .B(_1611_),
    .C(_1586_),
    .Y(_1614_)
);

OAI21X1 _3108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_747_),
    .C(_756_),
    .Y(_84_)
);

FILL FILL_1__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3281_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_43_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(load_only)
);

FILL FILL_6__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(cld),
    .Y(_642_)
);

FILL FILL_6__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_208_),
    .C(_290_),
    .Y(_1685_[12])
);

XOR2X1 _2132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(backwards),
    .Y(_1268_)
);

FILL FILL_2__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3337_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_91_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[2] [6])
);

FILL FILL_1__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_745_),
    .C(_746_),
    .Y(_76_)
);

FILL FILL_2__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_933_),
    .C(_857_),
    .D(_967_),
    .Y(BI[3])
);

FILL FILL_4__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[0]),
    .B(_338_),
    .C(_321_),
    .D(ADD[0]),
    .Y(_339_)
);

FILL FILL_1__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf0),
    .B(_961_),
    .C(NMI_edge),
    .Y(_496_)
);

OAI21X1 _2361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_120_),
    .C(_122_),
    .Y(alu_op[1])
);

FILL FILL_8__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf2),
    .B(_1640_),
    .C(_1641_),
    .Y(_1496_)
);

FILL FILL_6__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(_777_),
    .Y(_778_)
);

FILL FILL_7__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_1219__bF$buf1),
    .C(_534_),
    .D(_537_),
    .Y(_32_)
);

NAND2X1 _2417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1106_),
    .Y(_170_)
);

FILL FILL_1__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_191_),
    .C(_320_),
    .Y(_321_)
);

NAND2X1 _2170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1304_),
    .Y(_1305_)
);

FILL FILL_2__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(CI),
    .Y(_1650_)
);

FILL FILL_6__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(_982_),
    .C(_985_),
    .Y(_1005_)
);

FILL FILL_6__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .B(_343_),
    .C(_372_),
    .Y(_373_)
);

AND2X2 _2226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1349_),
    .B(_1360_),
    .Y(_1361_)
);

FILL FILL_7__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_815_),
    .B(_814_),
    .Y(_816_)
);

FILL FILL_2__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [1]),
    .B(_1022_),
    .Y(_1060_)
);

FILL FILL_7__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1304_),
    .B(_566_),
    .C(_1175_),
    .Y(_568_)
);

FILL FILL_6__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_203_),
    .Y(_206_)
);

AOI21X1 _2035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(_857_),
    .C(_1170_),
    .Y(_1171_)
);

FILL FILL_0__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(state[0]),
    .Y(_879_)
);

FILL FILL_4__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[6]),
    .B(_336_),
    .Y(_407_)
);

NOR2X1 _2264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1391_),
    .B(_1397_),
    .Y(_1398_)
);

FILL FILL_2__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_1540_),
    .Y(_1555_)
);

NAND2X1 _3049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_702_),
    .Y(_711_)
);

FILL FILL_7__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1091_),
    .C(_1094_),
    .Y(AI[4])
);

FILL FILL_1__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[5]),
    .Y(_239_)
);

NAND3X1 _2073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1207_),
    .C(_1204_),
    .Y(_1209_)
);

FILL FILL_2__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3278_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_40_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf5),
    .Q(adc_bcd)
);

FILL FILL_6__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _1764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .Y(_917_)
);

FILL FILL_4__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(AV),
    .C(_639_),
    .Y(_640_)
);

AOI21X1 _2549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[4]),
    .B(_1075_),
    .C(_287_),
    .Y(_288_)
);

OAI21X1 _2129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(_1264_),
    .C(_1263_),
    .Y(_1265_)
);

FILL FILL_7__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .B(_743_),
    .Y(_744_)
);

FILL FILL_0__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf1),
    .Y(_1129_)
);

FILL FILL_8__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf5),
    .B(_492_),
    .C(_493_),
    .Y(_17_)
);

NAND3X1 _2358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf2),
    .B(_121_),
    .C(_120_),
    .Y(_122_)
);

FILL FILL_7__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

INVX1 _2167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_894_),
    .Y(_1302_)
);

FILL FILL_7__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_914_),
    .C(_869__bF$buf1),
    .Y(_1002_)
);

FILL FILL_7__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(_128_),
    .C(_152_),
    .Y(_153_)
);

FILL FILL_8__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x152250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1039_),
    .Y(_1040_)
);

FILL FILL_8__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[1]),
    .Y(_833_)
);

FILL FILL_9__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1514_),
    .B(_1516_),
    .Y(_1517_)
);

AOI21X1 _3011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shift),
    .B(_1191_),
    .C(_1260_),
    .Y(_677_)
);

FILL FILL_2__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[1]),
    .B(_1133_),
    .C(_1008_),
    .Y(_424_)
);

FILL FILL_0__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf0),
    .B(_1035_),
    .C(_853__bF$buf2),
    .Y(_1432_)
);

FILL FILL_0__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3240_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_3_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(PC[1])
);

FILL FILL_2__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1173_),
    .B(_520_),
    .C(_612_),
    .Y(_613_)
);

AOI21X1 _2511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(AN),
    .C(_254_),
    .Y(_255_)
);

FILL FILL_7__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf0),
    .B(_880_),
    .Y(_951_)
);

OAI21X1 _2740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_324_),
    .C(_458_),
    .Y(_459_)
);

NAND3X1 _2320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1276_),
    .B(_1357_),
    .C(_1234_),
    .Y(_1453_)
);

FILL FILL_4__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(_1518_),
    .Y(_1611_)
);

OAI21X1 _3105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf2),
    .B(_748_),
    .C(\AXYS[1] [6]),
    .Y(_755_)
);

FILL FILL_1__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3334_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_88_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[2] [3])
);

FILL FILL_1__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[2]),
    .Y(_970_)
);

FILL FILL_0__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_321_),
    .C(_335_),
    .Y(_336_)
);

FILL FILL_1__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1638_),
    .B(RDY_bF$buf2),
    .C(_1639_),
    .Y(_1495_)
);

FILL FILL_6__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_767_),
    .C(_775_),
    .Y(_100_)
);

FILL FILL_6__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .Y(_535_)
);

OAI21X1 _2414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_128_),
    .C(_167_),
    .Y(_168_)
);

FILL FILL_1__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _3372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(_1648_),
    .Y(AV)
);

FILL FILL_6__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[4]),
    .Y(_370_)
);

NAND3X1 _2223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf2),
    .B(_927_),
    .C(_1356_),
    .Y(_1358_)
);

FILL FILL_2__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[3]),
    .B(_1674_),
    .C(_1513_),
    .Y(_1514_)
);

NOR2X1 _3008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(clc),
    .Y(_674_)
);

FILL FILL_1__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .B(_812_),
    .Y(_813_)
);

FILL FILL_2__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(_944_),
    .C(_1057_),
    .Y(_1058_)
);

FILL FILL_0__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1036_),
    .C(RDY_bF$buf1),
    .Y(_565_)
);

FILL FILL_6__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .Y(_203_)
);

NAND2X1 _2032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1152_),
    .Y(_1168_)
);

FILL FILL_2__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3237_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[4]),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf6),
    .Q(state[4])
);

FILL FILL_1__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_874_),
    .Y(_876_)
);

FILL FILL_4__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1320_),
    .B(_1384_),
    .C(_609_),
    .Y(_610_)
);

NAND2X1 _2508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_190_),
    .Y(_252_)
);

FILL FILL_1__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf2),
    .B(_402_),
    .C(_403_),
    .Y(_404_)
);

NOR2X1 _2261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1394_),
    .B(_1156_),
    .Y(_1395_)
);

FILL FILL_2__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x179550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(_1675_),
    .C(CI),
    .Y(_1552_)
);

FILL FILL_6__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_707_),
    .C(_708_),
    .Y(_70_)
);

FILL FILL_7__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[4]),
    .B(_1075_),
    .Y(_1092_)
);

OAI21X1 _2737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_359_),
    .C(_455_),
    .Y(_456_)
);

INVX1 _2317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .Y(_1450_)
);

FILL FILL_1__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1090_),
    .B(_182_),
    .C(_236_),
    .Y(_237_)
);

OAI21X1 _2070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf4),
    .B(_916_),
    .C(_853__bF$buf0),
    .Y(_1206_)
);

FILL FILL_2__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3275_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_37_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(shift_right)
);

FILL FILL_6__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(state[3]),
    .Y(_914_)
);

FILL FILL_6__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf3),
    .B(_988_),
    .C(DIMUX[6]),
    .Y(_637_)
);

INVX1 _2546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[4]),
    .Y(_285_)
);

OAI21X1 _2126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1260_),
    .C(_1261_),
    .Y(_1262_)
);

FILL FILL_7__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_726_),
    .C(_740_),
    .Y(_741_)
);

FILL FILL_2__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[1]),
    .Y(_968_)
);

FILL FILL_7__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .B(RDY_bF$buf1),
    .Y(_1126_)
);

FILL FILL_8__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_490_),
    .C(_460_),
    .Y(_491_)
);

OAI21X1 _2355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_918__bF$buf3),
    .C(_911_),
    .Y(_119_)
);

FILL FILL184050x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf0),
    .B(_926__bF$buf3),
    .C(_193_),
    .Y(_315_)
);

NAND2X1 _2164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1298_),
    .Y(_1299_)
);

FILL FILL_2__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1646_),
    .Y(AZ)
);

FILL FILL184050x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf3),
    .B(_988_),
    .C(_998_),
    .Y(_999_)
);

FILL FILL_6__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1073_),
    .Y(_150_)
);

FILL FILL_8__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[3]),
    .Y(DO[3])
);

FILL FILL_6__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_992_),
    .Y(_810_)
);

FILL FILL_0__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .B(_1129__bF$buf3),
    .C(_563_),
    .Y(_38_)
);

NAND3X1 _2449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1123_),
    .C(_1186_),
    .Y(_200_)
);

NAND3X1 _2029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf2),
    .B(_1150_),
    .C(_1164_),
    .Y(_1165_)
);

FILL FILL_7__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181350x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_1037_)
);

FILL FILL_8__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1055_),
    .B(_872_),
    .C(_260_),
    .D(_333_),
    .Y(_401_)
);

INVX1 _2258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .Y(_1392_)
);

FILL FILL_7__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [4]),
    .B(_1020_),
    .Y(_1089_)
);

FILL FILL_2__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[4]),
    .B(_204_),
    .C(_202_),
    .D(ABL[4]),
    .Y(_234_)
);

OAI21X1 _2067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf2),
    .B(_916_),
    .C(_853__bF$buf0),
    .Y(_1203_)
);

FILL FILL_0__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_910_),
    .C(_886__bF$buf1),
    .Y(_911_)
);

FILL FILL_4__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1428_),
    .B(_1361_),
    .Y(_1429_)
);

FILL FILL_2__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf1),
    .B(_900_),
    .Y(_1123_)
);

FILL FILL_4__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_940_),
    .B(_947_),
    .Y(_948_)
);

FILL FILL_5__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(_1607_),
    .Y(_1608_)
);

OAI21X1 _3102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_747_),
    .C(_753_),
    .Y(_81_)
);

FILL FILL_8__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3331_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_85_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[2] [0])
);

FILL FILL_2__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf1),
    .B(_953_),
    .C(_1145_),
    .Y(_333_)
);

FILL FILL_0__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_938_),
    .C(_1333_),
    .Y(_1334_)
);

FILL FILL_0__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf1),
    .B(_1622_),
    .C(_1637_),
    .Y(_1494_)
);

FILL FILL_6__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [6]),
    .B(_767_),
    .Y(_774_)
);

FILL FILL_8__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_526_),
    .Y(_532_)
);

AND2X2 _2411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_165_),
    .Y(_166_)
);

FILL FILL_0__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(DI[3]),
    .C(_856_),
    .Y(_857_)
);

FILL FILL_8__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_367_),
    .Y(_368_)
);

OAI21X1 _2220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1353_),
    .C(_1354_),
    .Y(_1355_)
);

FILL FILL_2__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[3]),
    .B(_1508_),
    .C(_1657_),
    .Y(_1511_)
);

OAI21X1 _3005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(_670_),
    .C(_671_),
    .Y(_66_)
);

FILL FILL_1__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[0]),
    .Y(_1055_)
);

FILL FILL_0__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3234_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[1]),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(state[1])
);

FILL FILL_1__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .Y(_873_)
);

FILL FILL_6__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(load_reg),
    .Y(_607_)
);

OAI21X1 _2505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_208_),
    .C(_249_),
    .Y(_250_)
);

FILL FILL_1__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1548_),
    .Y(_1549_)
);

FILL FILL_6__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_981_),
    .C(_705_),
    .Y(_706_)
);

FILL FILL_2__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_277_),
    .C(_453_),
    .D(_451_),
    .Y(_13_)
);

NAND3X1 _2314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1446_),
    .C(_1441_),
    .Y(_1447_)
);

FILL FILL_1__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1662_),
    .C(_1667_),
    .Y(_1605_)
);

FILL FILL_1__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3272_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_34_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf1),
    .Q(op[2])
);

FILL FILL_6__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(clv),
    .B(_633_),
    .Y(_634_)
);

FILL FILL_6__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_208_),
    .C(_282_),
    .Y(_1685_[11])
);

NAND2X1 _2123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(_868_),
    .Y(_1259_)
);

FILL FILL_2__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3328_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_82_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[1] [5])
);

FILL FILL_1__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [6]),
    .B(_693_),
    .Y(_739_)
);

FILL FILL_2__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_963_),
    .Y(_966_)
);

FILL FILL_4__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[7]),
    .B(_446_),
    .C(_487_),
    .Y(_488_)
);

NAND3X1 _2352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1252_),
    .B(_1408_),
    .C(_1482_),
    .Y(_117_)
);

FILL FILL_4__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[5]),
    .B(_1649__bF$buf1),
    .Y(_1636_)
);

FILL FILL_6__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_767_),
    .C(_772_),
    .Y(_97_)
);

FILL FILL_7__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x179550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_1175_),
    .Y(_529_)
);

OAI21X1 _2408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf3),
    .B(_1035_),
    .C(_981_),
    .Y(_163_)
);

FILL FILL_1__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_900_),
    .B(_1037_),
    .C(_869__bF$buf3),
    .Y(_312_)
);

OAI21X1 _2161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1152_),
    .C(_1145_),
    .Y(_1296_)
);

FILL FILL_2__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(ADD[6]),
    .Y(_1644_)
);

FILL FILL_2__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(_879_),
    .Y(_996_)
);

FILL FILL_6__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[3]),
    .B(_336_),
    .Y(_365_)
);

NOR2X1 _2217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf2),
    .B(_1168_),
    .Y(_1352_)
);

FILL FILL_7__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_128_),
    .C(_147_),
    .Y(_148_)
);

FILL FILL_8__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[0]),
    .Y(DO[0])
);

FILL FILL_6__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_804_),
    .Y(_807_)
);

FILL FILL_0__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf1),
    .B(_891_),
    .C(_1051__bF$buf3),
    .Y(_1052_)
);

FILL FILL_7__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_1219__bF$buf1),
    .C(_558_),
    .Y(_37_)
);

FILL FILL_6__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf3),
    .B(_891_),
    .C(_196_),
    .Y(_197_)
);

AND2X2 _2026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1161_),
    .B(_1145_),
    .Y(_1162_)
);

FILL FILL_7__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .Y(_870_)
);

FILL FILL_4__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf1),
    .B(_926__bF$buf2),
    .C(_893_),
    .Y(_1034_)
);

FILL FILL_8__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_398_),
    .C(_397_),
    .Y(_399_)
);

OAI21X1 _2255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1323_),
    .C(_1321_),
    .Y(_1389_)
);

FILL FILL_2__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1083_),
    .C(_1086_),
    .Y(AI[3])
);

FILL FILL_7__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(_182_),
    .C(_231_),
    .Y(_232_)
);

NOR2X1 _2064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(write_back),
    .B(_1125_),
    .Y(_1200_)
);

FILL FILL_2__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3269_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_31_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf5),
    .Q(bit_ins)
);

FILL FILL_7__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(rotate),
    .Y(_908_)
);

FILL FILL_4__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_1274_),
    .C(_1425_),
    .Y(_1426_)
);

FILL FILL_2__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1581_),
    .C(_1583_),
    .Y(_1584_)
);

FILL FILL_6__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_734_),
    .C(_735_),
    .Y(_736_)
);

FILL FILL_0__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_944_),
    .C(_1120_),
    .Y(_1121_)
);

FILL FILL_4__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_485_),
    .Y(_16_)
);

NOR2X1 _2349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1237_),
    .Y(_1480_)
);

FILL FILL_7__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(_866_),
    .Y(_945_)
);

FILL FILL_5__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_664_),
    .C(_665_),
    .Y(_65_)
);

INVX1 _2578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(shift_right),
    .Y(_311_)
);

NOR3X1 _2158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1249_),
    .C(_1213_),
    .Y(_1294_)
);

FILL FILL_7__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_917_),
    .Y(_993_)
);

FILL FILL_7__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1063_),
    .Y(_145_)
);

FILL FILL_8__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .B(_1326_),
    .C(_1328_),
    .Y(_1331_)
);

FILL FILL_0__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_),
    .Y(_1031_)
);

FILL FILL_8__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(DI[2]),
    .C(_854_),
    .Y(_855_)
);

FILL FILL_8__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(BI[3]),
    .Y(_1508_)
);

OAI21X1 _3002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1260_),
    .B(_667_),
    .C(_668_),
    .Y(_669_)
);

FILL FILL_5__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[15]),
    .B(_830__bF$buf2),
    .Y(_848_)
);

FILL FILL_3_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1172_),
    .B(_594_),
    .C(_604_),
    .Y(_605_)
);

AOI22X1 _2502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[6]),
    .B(_204_),
    .C(_202_),
    .D(ABL[6]),
    .Y(_247_)
);

FILL FILL_5__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .B(_935_),
    .Y(_1235_)
);

FILL FILL_0__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[1]),
    .Y(_1546_)
);

FILL FILL_8__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .Y(_703_)
);

FILL FILL_2__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_441_),
    .C(_450_),
    .Y(_451_)
);

INVX1 _2311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .Y(_1444_)
);

FILL FILL_0__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1601_),
    .C(_1599_),
    .Y(_1602_)
);

FILL FILL_1__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_1031_),
    .C(_630_),
    .Y(_631_)
);

FILL FILL_6__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_278_),
    .Y(_280_)
);

OAI21X1 _2120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_989_),
    .C(RDY_bF$buf0),
    .Y(_1256_)
);

FILL FILL_2__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3325_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_79_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[1] [2])
);

FILL FILL_1__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(_959_),
    .Y(_963_)
);

FILL FILL_0__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x160050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1593_),
    .B(_1588_),
    .Y(_1634_)
);

FILL FILL_6__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [3]),
    .B(_767_),
    .Y(_771_)
);

FILL FILL_1__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf2),
    .B(_526_),
    .Y(_527_)
);

INVX1 _2405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .Y(_160_)
);

FILL FILL_1__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3363_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_116_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(ABH[7])
);

FILL FILL_2__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_343_),
    .C(_361_),
    .Y(_362_)
);

AOI22X1 _2214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1347_),
    .C(_1348_),
    .D(_1129__bF$buf4),
    .Y(_1349_)
);

FILL FILL_2__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .B(BI[4]),
    .C(_1675_),
    .Y(_1505_)
);

FILL FILL_1__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[7]),
    .Y(AB[7])
);

FILL FILL_6__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_798_),
    .Y(_804_)
);

FILL FILL_2__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .Y(_1049_)
);

FILL FILL_0__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_1129__bF$buf3),
    .C(_560_),
    .Y(_35_)
);

FILL FILL_6__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf3),
    .B(_193_),
    .Y(_194_)
);

NAND2X1 _2023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1158_),
    .Y(_1159_)
);

FILL FILL_2__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_830__bF$buf3),
    .C(_846_),
    .Y(_114_)
);

FILL FILL_1__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(_866_),
    .Y(_867_)
);

FILL FILL_4__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_1219__bF$buf1),
    .C(_602_),
    .Y(_49_)
);

FILL FILL_1__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_395_),
    .Y(_396_)
);

AOI21X1 _2252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1180_),
    .C(_1385_),
    .Y(_1386_)
);

FILL FILL_2__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[0]),
    .Y(_1543_)
);

FILL FILL_6__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .Y(_700_)
);

FILL FILL_7__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[3]),
    .B(_1075_),
    .Y(_1084_)
);

FILL FILL_5__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf1),
    .B(_1084_),
    .C(_447_),
    .Y(_448_)
);

NOR2X1 _2308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1430_),
    .Y(_1441_)
);

FILL FILL_7__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_205_),
    .C(_228_),
    .D(_201_),
    .Y(_229_)
);

NAND3X1 _2061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_1196_),
    .C(_1190_),
    .Y(_1197_)
);

FILL FILL_2__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3266_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_28_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf5),
    .Q(cli)
);

FILL FILL_6__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_867_),
    .Y(_905_)
);

FILL FILL_6__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(_1129__bF$buf3),
    .C(_618_),
    .Y(_61_)
);

FILL FILL_6__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[11]),
    .Y(_277_)
);

NOR2X1 _2117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .B(_1171_),
    .Y(_1253_)
);

FILL FILL_7__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1422_),
    .B(_1421_),
    .Y(_1423_)
);

FILL FILL_2__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(_1578_),
    .Y(_1581_)
);

FILL FILL_6__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_732_),
    .C(_733_),
    .Y(_74_)
);

FILL FILL_0__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .Y(_960_)
);

FILL FILL_7__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[7]),
    .Y(_1118_)
);

FILL FILL_8__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_479_),
    .C(_482_),
    .Y(_483_)
);

NOR2X1 _2346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1476_),
    .Y(_1477_)
);

FILL FILL_7__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf2),
    .B(_941_),
    .Y(_942_)
);

FILL FILL_5__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_1191_),
    .C(_662_),
    .Y(_663_)
);

FILL FILL_6__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adc_sbc),
    .B(D),
    .Y(_0_)
);

NAND2X1 _2155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(_1290_),
    .Y(_1291_)
);

FILL FILL_0__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf2),
    .B(_876_),
    .Y(_990_)
);

FILL FILL_7__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_128_),
    .C(_142_),
    .Y(_143_)
);

FILL FILL_8__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[4]),
    .Y(AB[4])
);

NAND3X1 _3169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_800_),
    .C(_791_),
    .Y(_801_)
);

FILL FILL_7__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _2193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_1327_),
    .S(RDY_bF$buf0),
    .Y(_1328_)
);

FILL FILL_2__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[6]),
    .B(_1669_),
    .C(_1657_),
    .Y(_1672_)
);

FILL FILL_0__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf3),
    .B(_901_),
    .C(_1027_),
    .Y(_1028_)
);

FILL FILL_8__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_393_)
);

NOR2X1 _2249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .B(_1382_),
    .Y(_1383_)
);

FILL FILL_7__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_851_),
    .C(_852_),
    .Y(DIMUX[1])
);

FILL FILL_8__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(_1129__bF$buf1),
    .C(_584_),
    .Y(_46_)
);

FILL FILL_6__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1075_),
    .B(_225_),
    .Y(_226_)
);

OAI21X1 _2058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf2),
    .B(_926__bF$buf2),
    .C(_1193_),
    .Y(_1194_)
);

FILL FILL_0__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf3),
    .B(_901_),
    .C(_898_),
    .Y(_902_)
);

FILL FILL_4__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1420_),
    .Y(_1483_[2])
);

FILL FILL_0__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [7]),
    .B(_1020_),
    .Y(_1115_)
);

FILL FILL_4__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1049_),
    .C(_1231_),
    .Y(_1232_)
);

FILL FILL_0__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf2),
    .B(_936_),
    .C(_938_),
    .Y(_939_)
);

FILL FILL_4__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(_1673_),
    .Y(_1599_)
);

FILL FILL_1__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3322_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_76_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[0] [7])
);

FILL FILL_5__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[3]),
    .B(_1649__bF$buf0),
    .Y(_1632_)
);

FILL FILL_6__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_767_),
    .C(_769_),
    .Y(_94_)
);

FILL FILL_2__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bit_ins),
    .Y(_524_)
);

OAI21X1 _2402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_128_),
    .C(_157_),
    .Y(_158_)
);

FILL FILL_0__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3360_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_113_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(ABH[4])
);

FILL FILL_2__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .Y(_359_)
);

NOR3X1 _2211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1308_),
    .C(_1345_),
    .Y(_1346_)
);

FILL FILL_9__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[4]),
    .C(_1501_),
    .D(_1652_),
    .Y(_1502_)
);

FILL FILL_1__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1030_),
    .B(_1045_),
    .C(_1042_),
    .Y(_1046_)
);

FILL FILL_0__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_558_),
    .Y(_559_)
);

FILL FILL_8__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf3),
    .B(_905_),
    .Y(_191_)
);

INVX1 _2020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1155_),
    .Y(_1156_)
);

FILL FILL_2__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[12]),
    .B(_830__bF$buf2),
    .Y(_845_)
);

FILL FILL_1__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .Y(DIMUX[7])
);

FILL FILL_0__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_599_),
    .C(_549_),
    .Y(_600_)
);

FILL FILL_1__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .B(AI[0]),
    .Y(_1540_)
);

FILL FILL_6__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adj_bcd),
    .B(adc_bcd),
    .C(HC),
    .Y(_697_)
);

FILL FILL_2__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [3]),
    .B(_1020_),
    .Y(_1081_)
);

FILL FILL_5__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1145_),
    .C(_414_),
    .D(_415_),
    .Y(_445_)
);

NOR2X1 _2305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf3),
    .B(_1217_),
    .Y(_1438_)
);

FILL FILL_5__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3263_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_25_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf5),
    .Q(sec)
);

FILL FILL_6__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_620_),
    .C(_627_),
    .Y(_59_)
);

FILL FILL_6__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_268_),
    .C(_274_),
    .Y(_275_)
);

INVX1 _2114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(write_back),
    .Y(_1250_)
);

FILL FILL_9__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3319_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_73_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [4])
);

FILL FILL_1__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1577_),
    .B(_1574_),
    .Y(_1578_)
);

FILL FILL_6__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_730_),
    .Y(_731_)
);

FILL FILL_2__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .B(_954_),
    .C(_956_),
    .Y(_957_)
);

FILL FILL_4__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_475_),
    .Y(_480_)
);

NOR2X1 _2343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1472_),
    .Y(_1474_)
);

FILL FILL_9__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf2),
    .B(_1581_),
    .C(_1630_),
    .Y(_1489_)
);

FILL FILL_6__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [0]),
    .B(_767_),
    .Y(_768_)
);

FILL FILL_7__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_521_),
    .Y(_522_)
);

FILL FILL_1__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(AN),
    .C(_1008_),
    .Y(_660_)
);

FILL FILL_6__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1118_),
    .B(_268_),
    .C(_307_),
    .Y(_308_)
);

NAND2X1 _2152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf0),
    .B(_1287_),
    .Y(_1288_)
);

FILL FILL_2__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3357_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_110_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(ABH[1])
);

FILL FILL_0__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_980_),
    .B(_983_),
    .C(_986_),
    .Y(_987_)
);

FILL FILL_6__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_356_),
    .Y(_357_)
);

OAI22X1 _2208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_872_),
    .C(_1342_),
    .D(_1341_),
    .Y(_1343_)
);

FILL FILL_7__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(php),
    .Y(_140_)
);

FILL FILL_8__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[15]),
    .Y(AB[15])
);

FILL FILL_6__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1193_),
    .B(_926__bF$buf3),
    .C(_881_),
    .D(_905_),
    .Y(_798_)
);

FILL FILL_7__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1162_),
    .B(_549_),
    .C(_555_),
    .Y(_556_)
);

FILL FILL_6__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .B(_990_),
    .C(_1235_),
    .Y(_188_)
);

NAND2X1 _2017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf0),
    .B(IRHOLD[5]),
    .Y(_1153_)
);

FILL FILL_7__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_934_),
    .C(_1324_),
    .D(_1322_),
    .Y(_1325_)
);

FILL FILL_2__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(BI[6]),
    .Y(_1669_)
);

FILL FILL_0__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(DI[6]),
    .C(_862_),
    .Y(_863_)
);

FILL FILL_4__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1013_),
    .B(_1021_),
    .C(_1024_),
    .Y(_1025_)
);

FILL FILL_8__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_385_),
    .Y(_391_)
);

AOI21X1 _2246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1368_),
    .C(_1379_),
    .Y(_1380_)
);

FILL FILL_7__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1074_),
    .C(_1078_),
    .Y(AI[2])
);

FILL FILL_7__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_849_),
    .C(_850_),
    .Y(DIMUX[0])
);

FILL FILL_8__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_581_),
    .Y(_582_)
);

FILL FILL_6__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .Y(_1685_[2])
);

FILL FILL183450x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf4),
    .B(_989_),
    .Y(_1191_)
);

FILL FILL_0__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[0]),
    .B(_870_),
    .Y(_899_)
);

FILL FILL_4__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1223_),
    .B(_1276_),
    .Y(_1418_)
);

FILL FILL_2__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .Y(_1575_)
);

INVX1 _3069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .Y(_728_)
);

FILL FILL_0__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1107_),
    .C(_1112_),
    .Y(AI[6])
);

FILL FILL_4__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_1228_),
    .Y(_1229_)
);

FILL FILL_2__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3298_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_52_),
    .S(_1__bF$buf8),
    .R(vdd),
    .CLK(clk_bF$buf7),
    .Q(res)
);

FILL FILL_6__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .Y(_936_)
);

FILL FILL_4__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(compare),
    .B(_633_),
    .Y(_657_)
);

OAI21X1 _2569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_195_),
    .C(DIMUX[7]),
    .Y(_305_)
);

NAND2X1 _2149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1284_),
    .Y(_1285_)
);

FILL FILL_7__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1595_),
    .Y(_1596_)
);

FILL FILL_3__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x54750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_1394_),
    .Y(_507_)
);

OAI21X1 _2378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1281_),
    .C(PC[8]),
    .Y(_137_)
);

FILL FILL_6__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .Y(_1322_)
);

FILL FILL_0__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1016_),
    .B(_1011_),
    .Y(_1022_)
);

FILL FILL_0__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[5]),
    .Y(_1499_)
);

FILL FILL_1__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[3]),
    .Y(_843_)
);

FILL FILL_2__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1219__bF$buf0),
    .C(_589_),
    .D(_597_),
    .Y(_48_)
);

FILL FILL_1__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1536_),
    .Y(_1537_)
);

FILL FILL_6__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[0]),
    .B(_981_),
    .C(_694_),
    .Y(_695_)
);

FILL FILL_2__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_441_),
    .Y(_443_)
);

NAND3X1 _2302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1431_),
    .C(_1434_),
    .Y(_1435_)
);

FILL FILL_0__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .Y(_1593_)
);

FILL FILL_1__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3260_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_22_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(plp)
);

FILL FILL_8__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[5]),
    .Y(_626_)
);

FILL FILL_6__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[10]),
    .Y(_272_)
);

AND2X2 _2111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(_1246_),
    .Y(_1247_)
);

FILL FILL_2__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3316_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_70_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [1])
);

FILL FILL_1__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x175650 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf2),
    .B(_953_),
    .Y(_954_)
);

FILL FILL_0__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1284_),
    .B(_1109_),
    .Y(_477_)
);

INVX1 _2340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .Y(_1471_)
);

FILL FILL_4__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1572_),
    .B(_1628_),
    .C(RDY_bF$buf2),
    .Y(_1629_)
);

FILL FILL_6__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf3),
    .B(_758_),
    .C(\AXYS[2] [7]),
    .Y(_766_)
);

FILL FILL_1__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf1),
    .C(clv),
    .Y(_519_)
);

FILL FILL_1__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3354_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_107_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf9),
    .Q(ABL[6])
);

FILL FILL_2__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_955_),
    .Y(_984_)
);

FILL FILL_6__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf1),
    .B(_352_),
    .C(_353_),
    .Y(_354_)
);

OAI21X1 _2205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[1]),
    .B(_1339_),
    .C(_1338_),
    .Y(_1340_)
);

FILL FILL_5__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[12]),
    .Y(AB[12])
);

FILL FILL_6__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_943_),
    .B(_937_),
    .Y(_795_)
);

FILL FILL_2__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1168_),
    .C(_1214_),
    .Y(_553_)
);

FILL FILL_6__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_1227_),
    .C(_184_),
    .Y(_185_)
);

NOR2X1 _2014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1149_),
    .Y(_1150_)
);

FILL FILL_2__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1065_),
    .B(_830__bF$buf3),
    .C(_841_),
    .Y(_110_)
);

FILL FILL_1__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .Y(_1666_)
);

FILL FILL_2__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(DI[5]),
    .C(_860_),
    .Y(_861_)
);

FILL FILL_4__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .B(_321_),
    .C(_387_),
    .Y(_388_)
);

OAI21X1 _2243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf1),
    .B(_1002__bF$buf2),
    .C(_1376_),
    .Y(_1377_)
);

FILL FILL_2__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[1]),
    .B(_1533_),
    .C(_1657_),
    .Y(_1534_)
);

FILL FILL_6__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf2),
    .Y(_692_)
);

FILL FILL_7__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[2]),
    .B(_1075_),
    .Y(_1076_)
);

NAND3X1 _2719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[10]),
    .B(_415_),
    .C(_414_),
    .Y(_440_)
);

FILL FILL_7__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_579_),
    .C(_576_),
    .Y(_45_)
);

FILL FILL_6__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_220_),
    .Y(_221_)
);

NOR2X1 _2052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1187_),
    .Y(_1188_)
);

FILL FILL_2__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3257_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_19_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(cond_code[0])
);

FILL FILL_7__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(state[3]),
    .Y(_896_)
);

FILL FILL_4__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_620_),
    .C(_624_),
    .Y(_56_)
);

FILL FILL_6__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1065_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

NOR2X1 _2108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_936_),
    .Y(_1244_)
);

FILL FILL_7__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1380_),
    .B(_1414_),
    .C(_1407_),
    .Y(_1415_)
);

FILL FILL_2__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .Y(_1572_)
);

FILL FILL_6__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_724_),
    .C(_725_),
    .Y(_73_)
);

FILL FILL_2__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .Y(_1110_)
);

AOI22X1 _2757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_472_),
    .C(_468_),
    .D(_473_),
    .Y(_474_)
);

NAND3X1 _2337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1468_),
    .C(_1467_),
    .Y(_1483_[4])
);

FILL FILL_7__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1224_),
    .C(_1225_),
    .Y(_1226_)
);

FILL FILL_2__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3295_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[5]),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf2),
    .Q(DIHOLD[5])
);

FILL FILL_0__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf2),
    .B(_900_),
    .Y(_933_)
);

FILL FILL_5__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_653_),
    .B(_652_),
    .C(_654_),
    .Y(_655_)
);

FILL FILL_6__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_208_),
    .C(_302_),
    .Y(_1685_[14])
);

OAI21X1 _2146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf2),
    .B(_961_),
    .C(_853__bF$buf2),
    .Y(_1282_)
);

FILL FILL_7__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf1),
    .B(_893_),
    .Y(_981_)
);

FILL FILL_7__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x58650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_1129__bF$buf1),
    .C(_504_),
    .Y(_23_)
);

OAI21X1 _2375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1182_),
    .B(_134_),
    .C(store),
    .Y(_135_)
);

FILL FILL_8__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(_1313_),
    .C(_1318_),
    .Y(_1319_)
);

FILL FILL_2__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1663_),
    .C(_1662_),
    .Y(_1664_)
);

FILL FILL_0__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1006_),
    .B(src_reg[0]),
    .Y(_1019_)
);

FILL FILL_0__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[6]),
    .Y(DO[6])
);

FILL FILL_3__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .Y(_830_)
);

FILL FILL_0__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x97650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1161_),
    .C(_1145_),
    .Y(_577_)
);

INVX1 _2469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .Y(_1685_[1])
);

INVX1 _2049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .Y(_1185_)
);

FILL FILL_7__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .B(BI[5]),
    .C(_1675_),
    .Y(_1684_)
);

FILL FILL_3__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .Y(_420_)
);

OAI21X1 _2278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1186_),
    .C(_1411_),
    .Y(_1412_)
);

FILL FILL_0__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .Y(_1107_)
);

FILL FILL_2__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1297_),
    .C(_520_),
    .Y(_595_)
);

FILL FILL_3__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_943_),
    .C(_1222_),
    .Y(_1223_)
);

FILL FILL_0__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_904_),
    .B(_930_),
    .Y(CI)
);

FILL FILL_4__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1506_),
    .Y(_1590_)
);

FILL FILL_1__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3313_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_67_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf5),
    .Q(C)
);

FILL FILL_1__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[0]),
    .B(_1649__bF$buf2),
    .Y(_1626_)
);

FILL FILL_6__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_757_),
    .C(_764_),
    .Y(_90_)
);

FILL FILL_2__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_1129__bF$buf1),
    .C(_506_),
    .D(_517_),
    .Y(_28_)
);

FILL FILL_1__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3351_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_104_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf2),
    .Q(ABL[3])
);

FILL FILL_2__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[2]),
    .B(_853__bF$buf5),
    .Y(_351_)
);

NOR2X1 _2202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[2]),
    .B(_1336_),
    .Y(_1337_)
);

FILL FILL_5__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[5]),
    .C(_1680_),
    .D(_1652_),
    .Y(_1681_)
);

FILL FILL_1__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[1]),
    .Y(AB[1])
);

FILL FILL_6__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf2),
    .B(_926__bF$buf0),
    .C(_900_),
    .Y(_792_)
);

FILL FILL_2__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .Y(_550_)
);

FILL FILL_6__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_181_),
    .Y(_182_)
);

OAI21X1 _2011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf1),
    .B(_855_),
    .C(_1146_),
    .Y(_1147_)
);

FILL FILL_9__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_266_),
    .C(_830__bF$buf3),
    .Y(_840_)
);

FILL FILL_1__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(DI[4]),
    .C(_858_),
    .Y(_859_)
);

FILL FILL_9__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf0),
    .B(_591_),
    .C(_592_),
    .Y(_47_)
);

FILL FILL_1__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_367_),
    .Y(_385_)
);

OAI21X1 _2240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1029_),
    .C(_1373_),
    .Y(_1374_)
);

FILL FILL_9__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[1]),
    .C(_1530_),
    .D(_1652_),
    .Y(_1531_)
);

NOR2X1 _3025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(_688_),
    .Y(_689_)
);

FILL FILL_0__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1070_),
    .B(_1072_),
    .C(_1071_),
    .Y(_1073_)
);

FILL FILL_0__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[2]),
    .Y(_437_)
);

FILL FILL_7__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3254_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_17_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[15])
);

FILL FILL_2__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(_892_),
    .Y(_893_)
);

FILL FILL_6__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[2]),
    .Y(_623_)
);

FILL FILL_6__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[9]),
    .Y(_267_)
);

NAND2X1 _2105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1240_),
    .Y(_1241_)
);

FILL FILL_5__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(_1519_),
    .Y(_1569_)
);

FILL FILL_6__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_949_),
    .C(_285_),
    .Y(_723_)
);

FILL FILL_2__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf5),
    .B(_471_),
    .C(_463_),
    .Y(_15_)
);

NOR2X1 _2334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1461_),
    .B(_1465_),
    .Y(_1466_)
);

FILL FILL_5__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1666_),
    .B(_1649__bF$buf3),
    .C(_1624_),
    .D(_1608_),
    .Y(_1486_)
);

OAI21X1 _3119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf0),
    .B(_758_),
    .C(\AXYS[2] [4]),
    .Y(_763_)
);

FILL FILL_1__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3292_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[2]),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf9),
    .Q(DIHOLD[2])
);

FILL FILL_6__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1260_),
    .Y(_652_)
);

FILL FILL_6__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(ADD[6]),
    .C(_1109_),
    .Y(_300_)
);

OAI21X1 _2143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf0),
    .B(_1277_),
    .C(_1278_),
    .Y(_1279_)
);

FILL FILL_2__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3348_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_101_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf8),
    .Q(ABL[0])
);

FILL FILL_0__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf1),
    .B(_906_),
    .Y(_978_)
);

FILL FILL_6__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_340_),
    .Y(_349_)
);

FILL FILL_4_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .Y(_918__bF$buf2)
);

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .Y(_918__bF$buf1)
);

BUFX2 BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .Y(_918__bF$buf0)
);

BUFX2 BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf7)
);

BUFX2 BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf6)
);

BUFX2 BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf5)
);

BUFX2 BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf4)
);

BUFX2 BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf3)
);

BUFX2 BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf2)
);

BUFX2 BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .Y(_853__bF$buf1)
);

FILL FILL_3__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_1129__bF$buf1),
    .C(_1299_),
    .D(_1324_),
    .Y(_22_)
);

NOR2X1 _2372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_120_),
    .Y(alu_op[3])
);

FILL FILL_8__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3577_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1495_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf0),
    .Q(AN)
);

FILL FILL_6__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf0),
    .B(_906_),
    .C(_1044_),
    .Y(_789_)
);

FILL FILL_7__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1323_),
    .Y(_547_)
);

FILL FILL_6__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_179_),
    .C(_175_),
    .Y(_1686_[7])
);

NAND2X1 _2008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1131_),
    .B(_1132_),
    .Y(_1144_)
);

FILL FILL_7__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1315_),
    .Y(_1316_)
);

FILL FILL_2__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[7]),
    .C(_1660_),
    .Y(_1661_)
);

FILL FILL_6__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1006_),
    .C(_1015_),
    .Y(_1016_)
);

FILL FILL_2__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .Y(_383_)
);

NOR2X1 _2237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1268_),
    .B(_872_),
    .Y(_1371_)
);

FILL FILL_7__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _3195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_826_),
    .B(_1183_),
    .Y(_827_)
);

FILL FILL_0__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [2]),
    .B(_1022_),
    .Y(_1070_)
);

FILL FILL_7__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1250_),
    .B(_1129__bF$buf2),
    .C(_520_),
    .D(_574_),
    .Y(_44_)
);

FILL FILL_6__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_215_),
    .Y(_216_)
);

NOR2X1 _2046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_936_),
    .Y(_1182_)
);

FILL FILL_7__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_889_),
    .Y(_890_)
);

FILL FILL_4__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_416_),
    .C(_417_),
    .Y(_418_)
);

NOR2X1 _2275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_1200_),
    .Y(_1409_)
);

FILL FILL_2__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x156150 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [6]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [6]),
    .Y(_1104_)
);

FILL FILL_7__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .Y(_1220_)
);

FILL FILL_5_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3289_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_51_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(load_reg)
);

FILL FILL_0__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_889_),
    .Y(_928_)
);

FILL FILL_4__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1586_),
    .Y(_1587_)
);

FILL FILL_3__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_747_),
    .C(_751_),
    .Y(_79_)
);

FILL FILL_0__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[2]),
    .B(_853__bF$buf7),
    .Y(_501_)
);

AOI21X1 _2369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(backwards),
    .B(_1075_),
    .C(_130_),
    .Y(_131_)
);

FILL FILL_7__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3310_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_64_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf9),
    .Q(I)
);

FILL FILL_3__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_327_),
    .C(_1008_),
    .Y(_329_)
);

NAND3X1 _2178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_926__bF$buf0),
    .C(_890_),
    .Y(_1313_)
);

FILL FILL_0__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [0]),
    .B(_1012_),
    .Y(_1013_)
);

FILL FILL_7__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cli),
    .Y(_515_)
);

FILL FILL_0__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[6]),
    .Y(_1678_)
);

FILL FILL_1__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_251_),
    .C(_838_),
    .Y(_107_)
);

FILL FILL_1__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_523_),
    .C(_589_),
    .Y(_590_)
);

FILL FILL_1__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(alu_op[3]),
    .Y(_1528_)
);

FILL FILL_6__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf1),
    .B(_685_),
    .C(_686_),
    .Y(_68_)
);

FILL FILL_2__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1264_),
    .B(_413_),
    .C(DIMUX[2]),
    .Y(_434_)
);

FILL FILL_0__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3251_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_14_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf7),
    .Q(PC[12])
);

FILL FILL_2__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x144450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(_620_),
    .C(_621_),
    .Y(_53_)
);

FILL FILL_6__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(DIMUX[0]),
    .C(_264_),
    .Y(_265_)
);

NAND2X1 _2102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf0),
    .B(_935_),
    .Y(_1238_)
);

FILL FILL_5__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3307_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_61_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf1),
    .Q(IRHOLD_valid)
);

FILL FILL_1__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1565_),
    .C(_1563_),
    .Y(_1566_)
);

FILL FILL_8__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _3060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[3]),
    .B(_981_),
    .C(_720_),
    .D(_719_),
    .Y(_721_)
);

FILL FILL_2__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_324_),
    .C(_468_),
    .Y(_469_)
);

NAND3X1 _2331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(_1127_),
    .C(_1462_),
    .Y(_1463_)
);

FILL FILL_5__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1621_),
    .B(_1620_),
    .Y(_1622_)
);

OAI21X1 _3116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_757_),
    .C(_761_),
    .Y(_87_)
);

FILL FILL_1__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_513_),
    .C(_511_),
    .Y(_26_)
);

FILL FILL_1__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_951_),
    .Y(_649_)
);

FILL FILL_6__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_298_)
);

OAI21X1 _2140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf0),
    .B(_1274_),
    .C(_1275_),
    .Y(_1276_)
);

FILL FILL_2__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3345_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_98_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[3] [5])
);

FILL FILL_6__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_933_),
    .C(_864_),
    .D(_967_),
    .Y(BI[7])
);

FILL FILL_0__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(_321_),
    .C(_345_),
    .Y(_346_)
);

FILL FILL_1__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(_887__bF$buf3)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(_887__bF$buf2)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(_887__bF$buf1)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .Y(_887__bF$buf0)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .Y(_869__bF$buf3)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .Y(_869__bF$buf2)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .Y(_869__bF$buf1)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .Y(_869__bF$buf0)
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf3)
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid),
    .Y(IRHOLD_valid_bF$buf2)
);

FILL FILL_3__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3574_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1492_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf0),
    .Q(ADD[4])
);

FILL FILL_6__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_785_),
    .B(_782_),
    .Y(_786_)
);

FILL FILL_2__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1155_),
    .B(_512_),
    .Y(_544_)
);

FILL FILL_6__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(N),
    .B(_141_),
    .Y(_177_)
);

AOI21X1 _2005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf2),
    .B(_1140_),
    .C(_1133_),
    .Y(_1141_)
);

FILL FILL_5__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[7]),
    .B(_1654_),
    .C(_1657_),
    .Y(_1658_)
);

FILL FILL_6__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[4]),
    .B(_336_),
    .Y(_380_)
);

NAND3X1 _2234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1364_),
    .C(_1367_),
    .Y(_1368_)
);

FILL FILL_2__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_1523_),
    .C(_1524_),
    .Y(_1525_)
);

OAI21X1 _3019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_683_),
    .C(_684_),
    .Y(_67_)
);

FILL FILL_1__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_783_),
    .C(_823_),
    .Y(_824_)
);

FILL FILL_2__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_944_),
    .C(_1067_),
    .Y(_1068_)
);

FILL FILL_0__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf0),
    .C(load_only),
    .Y(_573_)
);

FILL FILL_6__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_213_),
    .Y(_1685_[0])
);

NAND2X1 _2043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1178_),
    .Y(_1179_)
);

FILL FILL_2__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3248_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_11_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[9])
);

FILL FILL_7__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _1734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf3),
    .Y(_887_)
);

FILL FILL_4__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .Y(_619_)
);

AOI21X1 _2519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[0]),
    .B(_199_),
    .C(_182_),
    .Y(_262_)
);

FILL FILL_1__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .Y(_415_)
);

INVX1 _2272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .Y(_1406_)
);

FILL FILL_2__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_1527_),
    .Y(_1563_)
);

FILL FILL_6__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _3057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(ADD[3]),
    .Y(_718_)
);

FILL FILL_0__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[5]),
    .C(_1101_),
    .Y(_1102_)
);

FILL FILL_4__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_359_),
    .C(_465_),
    .Y(_466_)
);

NOR2X1 _2328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1459_),
    .Y(_1460_)
);

FILL FILL_7__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1216_),
    .B(_1215_),
    .Y(_1217_)
);

FILL FILL_5_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3286_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_48_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(src_reg[1])
);

FILL FILL_6__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(C),
    .B(_908_),
    .C(_924_),
    .Y(_925_)
);

FILL FILL_2__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(cld),
    .C(_646_),
    .Y(_647_)
);

FILL FILL_6__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_240_),
    .C(_294_),
    .Y(_295_)
);

OAI21X1 _2137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf0),
    .B(_878_),
    .C(_1272_),
    .Y(_1273_)
);

FILL FILL_7__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf1),
    .B(_748_),
    .C(\AXYS[1] [1]),
    .Y(_750_)
);

FILL FILL_2__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[6]),
    .Y(_974_)
);

FILL FILL_7__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_497_),
    .C(_499_),
    .Y(_19_)
);

INVX2 _2366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .Y(_128_)
);

FILL FILL_7__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x156150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[0]),
    .B(_325_),
    .C(_321_),
    .D(ADD[0]),
    .Y(_326_)
);

NAND3X1 _2175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf3),
    .B(_1235_),
    .C(_1188_),
    .Y(_1310_)
);

FILL FILL_2__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .B(_1009_),
    .C(_1005_),
    .Y(_1010_)
);

FILL FILL_7__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .B(_993_),
    .C(_933_),
    .Y(_821_)
);

FILL FILL_0__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .Y(_1675_)
);

FILL FILL_3__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_411_),
    .Y(_412_)
);

AOI22X1 _2269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1401_),
    .B(_1402_),
    .C(_1399_),
    .D(_1316_),
    .Y(_1403_)
);

FILL FILL_7__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[5]),
    .Y(_837_)
);

FILL FILL_3__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_498_),
    .Y(_587_)
);

FILL FILL_3__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_208_),
    .C(_243_),
    .Y(_244_)
);

INVX1 _2078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .Y(_1214_)
);

FILL FILL_0__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(load_only),
    .B(_921_),
    .C(_920_),
    .Y(_922_)
);

FILL FILL_4__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_398_),
    .C(RDY_bF$buf8),
    .Y(_432_)
);

FILL FILL_0__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf2),
    .B(_1130_),
    .C(_1133_),
    .Y(_1134_)
);

FILL FILL_8__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3304_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_58_),
    .CLK(clk_bF$buf10),
    .Q(IRHOLD[5])
);

FILL FILL_1__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1617_),
    .Y(_1619_)
);

OAI21X1 _3113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf0),
    .B(_758_),
    .C(\AXYS[2] [1]),
    .Y(_760_)
);

FILL FILL_1__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf3),
    .C(cld),
    .Y(_511_)
);

FILL FILL_1__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3342_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_95_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[3] [2])
);

FILL FILL_6__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2615_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .Y(_343_)
);

FILL FILL_1__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x144450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf2)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf1)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY),
    .Y(RDY_bF$buf0)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1051__bF$buf3)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1051__bF$buf2)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1051__bF$buf1)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1051__bF$buf0)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf10)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf9)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_),
    .Y(_1__bF$buf8)
);

FILL FILL_3__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3571_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1489_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf3),
    .Q(ADD[1])
);

FILL FILL_6__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_1327_),
    .C(_994_),
    .Y(_783_)
);

FILL FILL_2__2844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3382_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(_1383_),
    .Y(_541_)
);

FILL FILL_6__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_174_),
    .C(_170_),
    .Y(_1686_[6])
);

OAI21X1 _2002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf3),
    .B(DIMUX[0]),
    .C(_1137_),
    .Y(_1138_)
);

FILL FILL_5__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_232_),
    .C(_835_),
    .Y(_104_)
);

FILL FILL_1__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[7]),
    .B(_1654_),
    .Y(_1655_)
);

FILL FILL_6__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2653_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2233_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[5]),
    .B(_321_),
    .C(_376_),
    .Y(_377_)
);

NAND2X1 _2231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_905_),
    .Y(_1365_)
);

FILL FILL_2__1924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[2]),
    .B(_1651_),
    .C(_1521_),
    .D(_1652_),
    .Y(_1522_)
);

NAND2X1 _3016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(_1260_),
    .Y(_682_)
);

FILL FILL_1__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[1]),
    .Y(_1065_)
);

FILL FILL_0__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[9]),
    .B(_415_),
    .C(_414_),
    .Y(_429_)
);

FILL FILL_7__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_550_),
    .B(_541_),
    .Y(_571_)
);

FILL FILL_8__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_210_),
    .Y(_211_)
);

NAND2X1 _2040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1173_),
    .Y(_1176_)
);

FILL FILL_2__1733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3245_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_8_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf7),
    .Q(PC[6])
);

FILL FILL_0__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2271_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .B(_878_),
    .Y(_884_)
);

FILL FILL_6__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3056_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_1219__bF$buf0),
    .C(_611_),
    .D(_617_),
    .Y(_51_)
);

INVX1 _2516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .Y(_1685_[7])
);

FILL FILL_1__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1551_),
    .C(_1559_),
    .D(_1553_),
    .Y(_1560_)
);

FILL FILL_6__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_714_),
    .C(_715_),
    .Y(_71_)
);

FILL FILL_2__2747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2327_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1098_),
    .Y(_1099_)
);

NAND2X1 _2745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[13]),
    .B(_853__bF$buf5),
    .Y(_463_)
);

NOR2X1 _2325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1457_),
    .Y(_1458_)
);

FILL FILL_5__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3283_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_45_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(store)
);

FILL FILL_6__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3094_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf3),
    .B(_643_),
    .C(_629_),
    .Y(_644_)
);

FILL FILL_6__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[5]),
    .Y(_292_)
);

OAI22X1 _2134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_1269_),
    .C(RDY_bF$buf1),
    .D(_1267_),
    .Y(_1270_)
);

FILL FILL_2__1827_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3339_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_0_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(adj_bcd)
);

FILL FILL_1__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1022_),
    .Y(_748_)
);

FILL FILL_2__2785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2365_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .B(_933_),
    .C(_859_),
    .D(_967_),
    .Y(BI[4])
);

FILL FILL_4__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(cond_code[0]),
    .Y(_497_)
);

NOR2X1 _2363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf0),
    .B(_961_),
    .Y(_125_)
);

FILL FILL_8__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3568_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1486_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf0),
    .Q(CO)
);

FILL FILL_6__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_951_),
    .Y(_780_)
);

FILL FILL_7__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_538_),
    .B(_1350_),
    .Y(_539_)
);

NAND2X1 _2419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(V),
    .B(_141_),
    .Y(_172_)
);

FILL FILL_1__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_321_),
    .Y(_323_)
);

AOI22X1 _2172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_1302_),
    .C(_1306_),
    .D(_1129__bF$buf4),
    .Y(_1307_)
);

FILL FILL_2__1865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_1651_),
    .Y(_1652_)
);

FILL FILL_6__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .B(_997_),
    .C(index_y),
    .Y(_1007_)
);

FILL FILL_6__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x132750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(_374_),
    .C(_369_),
    .Y(_6_)
);

OR2X2 _2228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1293_),
    .Y(_1483_[1])
);

FILL FILL_7__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_813_),
    .B(_817_),
    .C(_811_),
    .Y(_818_)
);

FILL FILL_0__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3400_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [1]),
    .B(_1020_),
    .Y(_1062_)
);

FILL FILL_7__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adc_sbc),
    .Y(_569_)
);

FILL FILL_6__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_207_),
    .Y(_208_)
);

INVX1 _2037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1172_),
    .Y(_1173_)
);

FILL FILL_7__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2268_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[5]),
    .Y(_881_)
);

FILL FILL_4__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_388_),
    .C(_408_),
    .D(_394_),
    .Y(_409_)
);

INVX1 _2266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .Y(_1400_)
);

FILL FILL_7__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [5]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [5]),
    .Y(_1096_)
);

FILL FILL_7__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_205_),
    .C(_239_),
    .D(_240_),
    .Y(_241_)
);

AOI21X1 _2075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1189_),
    .B(_1198_),
    .C(_1210_),
    .Y(_1211_)
);

FILL FILL_2__1768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_916_),
    .Y(_919_)
);

FILL FILL_7__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [7]),
    .B(_693_),
    .Y(_746_)
);

FILL FILL_0__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRQ),
    .Y(_1131_)
);

FILL FILL184050x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _3301_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_55_),
    .CLK(clk_bF$buf10),
    .Q(IRHOLD[2])
);

FILL FILL_3__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf0),
    .B(_926__bF$buf3),
    .C(_1193_),
    .D(_193_),
    .Y(_320_)
);

NOR2X1 _2169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1303_),
    .Y(_1304_)
);

FILL FILL_7__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1597_),
    .Y(_1616_)
);

FILL FILL_8__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _3110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .Y(_758_)
);

FILL FILL_2__2803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf1),
    .B(_499_),
    .Y(_509_)
);

FILL FILL_0__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_154_),
    .C(_150_),
    .Y(_1686_[2])
);

FILL FILL183150x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2612_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .Y(_341_)
);

FILL FILL_0__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(_1041_),
    .Y(_1042_)
);

FILL FILL_6__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_829_),
    .C(ABL[2]),
    .Y(_834_)
);

FILL FILL_1__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2650_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .Y(_1519_)
);

AOI21X1 _3013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .B(ADD[0]),
    .C(_674_),
    .Y(_679_)
);

FILL FILL_1__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(_425_),
    .C(_421_),
    .Y(_426_)
);

FILL FILL_9__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3242_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_5_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(PC[3])
);

FILL FILL_2__2935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_1159_),
    .C(_1175_),
    .Y(_615_)
);

INVX1 _2513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .Y(_257_)
);

FILL FILL_1__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .B(_1543_),
    .C(alu_shift_right),
    .Y(_1557_)
);

FILL FILL_6__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_712_),
    .Y(_713_)
);

FILL FILL_2__2744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2324_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_459_),
    .Y(_461_)
);

INVX1 _2322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1332_),
    .Y(_1455_)
);

FILL FILL_5__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1581_),
    .C(_1610_),
    .Y(_1613_)
);

OAI21X1 _3107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf3),
    .B(_748_),
    .C(\AXYS[1] [7]),
    .Y(_756_)
);

FILL FILL_1__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3280_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_42_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(inc)
);

FILL FILL_6__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_640_),
    .C(_641_),
    .Y(_62_)
);

FILL FILL_6__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .Y(_290_)
);

NAND2X1 _2131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf1),
    .B(_905_),
    .Y(_1267_)
);

FILL FILL_2__1824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3336_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_90_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[2] [5])
);

FILL FILL_1__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2609_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2362_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _1822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[3]),
    .Y(_971_)
);

FILL FILL_0__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf4),
    .B(_1145_),
    .Y(_338_)
);

FILL FILL_1__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(NMI),
    .B(_494_),
    .Y(_495_)
);

INVX1 _2360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(op[1]),
    .Y(_123_)
);

FILL FILL_8__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[7]),
    .B(RDY_bF$buf2),
    .Y(_1641_)
);

FILL FILL_6__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_1035_),
    .C(_776_),
    .Y(_777_)
);

FILL FILL_0__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_535_),
    .C(_1219__bF$buf1),
    .Y(_537_)
);

OAI21X1 _2416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_1099_),
    .C(_169_),
    .Y(_1686_[5])
);

FILL FILL_1__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _3374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf2),
    .Y(_1649_)
);

FILL FILL_6__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2647_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1000_),
    .B(src_reg[1]),
    .C(_1003_),
    .Y(_1004_)
);

FILL FILL_6__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[4]),
    .B(_321_),
    .C(_371_),
    .Y(_372_)
);

AOI21X1 _2225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1351_),
    .B(_1352_),
    .C(_1359_),
    .Y(_1360_)
);

FILL FILL_9__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_1032_),
    .C(_1227_),
    .Y(_815_)
);

FILL FILL_2__2876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1026_),
    .C(_1059_),
    .Y(AI[0])
);

FILL FILL_7__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(D),
    .B(_1159_),
    .Y(_567_)
);

FILL FILL_6__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .Y(_205_)
);

OAI21X1 _2034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(IRHOLD[3]),
    .C(_1145_),
    .Y(_1170_)
);

FILL FILL_2__1727_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3239_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_2_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf8),
    .Q(PC[0])
);

FILL FILL_1__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2685_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2265_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .Y(_878_)
);

FILL FILL_4__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_324_),
    .C(_405_),
    .Y(_406_)
);

NAND3X1 _2263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .B(_1396_),
    .C(_1393_),
    .Y(_1397_)
);

FILL FILL_2__1956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _3468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[1]),
    .B(_1542_),
    .S(alu_op[0]),
    .Y(_1554_)
);

FILL FILL_6__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_709_),
    .Y(_710_)
);

FILL FILL_7__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[4]),
    .C(_1093_),
    .Y(_1094_)
);

AOI21X1 _2739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[4]),
    .B(_446_),
    .C(_457_),
    .Y(_458_)
);

OR2X2 _2319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1258_),
    .B(_1291_),
    .Y(_1452_)
);

FILL FILL_1__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .C(ADD[5]),
    .Y(_238_)
);

NAND2X1 _2072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf0),
    .B(_919_),
    .Y(_1208_)
);

FILL FILL_2__1765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3277_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_39_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(shift)
);

FILL FILL_6__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_915_),
    .Y(_916_)
);

FILL FILL_4__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002__bF$buf2),
    .B(_638_),
    .C(_637_),
    .Y(_639_)
);

OAI21X1 _2548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_240_),
    .C(_286_),
    .Y(_287_)
);

NOR3X1 _2128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_867_),
    .C(_882__bF$buf3),
    .Y(_1264_)
);

FILL FILL_7__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _3086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(AN),
    .Y(_743_)
);

FILL FILL_0__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2359_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_933_),
    .C(_969_),
    .D(_967_),
    .Y(BI[1])
);

FILL FILL_7__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_938_),
    .B(RDY_bF$buf6),
    .Y(_1128_)
);

FILL FILL_8__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[15]),
    .B(_853__bF$buf5),
    .Y(_493_)
);

INVX1 _2357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1244_),
    .Y(_121_)
);

FILL FILL_7__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_978_),
    .B(_1365_),
    .C(_992_),
    .Y(_317_)
);

AOI22X1 _2166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1281_),
    .C(_1300_),
    .D(_1129__bF$buf4),
    .Y(_1301_)
);

FILL FILL_7__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(dst_reg[1]),
    .Y(_1001_)
);

FILL FILL_7__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(I),
    .B(_141_),
    .Y(_152_)
);

FILL FILL_8__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x82050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1038_),
    .Y(_1039_)
);

FILL FILL_8__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_213_),
    .C(_832_),
    .Y(_101_)
);

FILL FILL_3__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .B(_208_),
    .C(_235_),
    .Y(_236_)
);

OAI21X1 _2069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_887__bF$buf4),
    .C(RDY_bF$buf1),
    .Y(_1205_)
);

FILL FILL_0__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1663_),
    .Y(_1516_)
);

FILL FILL_8__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_675_),
    .C(_672_),
    .Y(_676_)
);

FILL FILL_2__2703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(_869__bF$buf3),
    .C(_905_),
    .Y(_423_)
);

FILL FILL_0__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181350x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1224_),
    .C(_1430_),
    .D(_1129__bF$buf4),
    .Y(_1431_)
);

FILL FILL_0__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3050_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(store),
    .Y(_1125_)
);

FILL FILL_4__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1382_),
    .B(_498_),
    .Y(_612_)
);

FILL FILL_8__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_205_),
    .C(_253_),
    .D(_201_),
    .Y(_254_)
);

FILL FILL_4__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2321_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .Y(_950_)
);

FILL FILL_4__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\u_ALU8.BCD ),
    .Y(_1610_)
);

OAI21X1 _3104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_747_),
    .C(_754_),
    .Y(_82_)
);

FILL FILL_1__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181650x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3333_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_87_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[2] [2])
);

FILL FILL_1__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2606_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3144_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .Y(_335_)
);

FILL FILL_1__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf2),
    .B(_1609_),
    .Y(_1639_)
);

FILL FILL_6__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [7]),
    .B(_767_),
    .Y(_775_)
);

FILL FILL_6__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .Y(_534_)
);

AOI22X1 _2413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(ADD[5]),
    .C(PC[13]),
    .D(_163_),
    .Y(_167_)
);

FILL FILL_1__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _3371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(\u_ALU8.BI7 ),
    .Y(_1648_)
);

FILL FILL_6__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2644_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[4]),
    .B(_853__bF$buf4),
    .Y(_369_)
);

OAI21X1 _2222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1284_),
    .C(_1356_),
    .Y(_1357_)
);

FILL FILL_2__1915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .B(BI[3]),
    .C(_1675_),
    .Y(_1513_)
);

NAND3X1 _3007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_912_),
    .C(_920_),
    .Y(_673_)
);

FILL FILL_1__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x70350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .Y(_812_)
);

FILL FILL_2__2873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .Y(_1057_)
);

FILL FILL_0__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_912_),
    .B(_1129__bF$buf1),
    .C(_1329_),
    .D(_564_),
    .Y(_39_)
);

FILL FILL_6__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _2451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_201_),
    .Y(_202_)
);

INVX1 _2031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .Y(_1167_)
);

FILL FILL_2__1724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3236_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[3]),
    .S(_1__bF$buf10),
    .R(vdd),
    .CLK(clk_bF$buf8),
    .Q(state[3])
);

FILL FILL_7__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2682_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2262_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(state[0]),
    .Y(_875_)
);

FILL FILL_6__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_522_),
    .Y(_609_)
);

INVX1 _2507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .Y(_1685_[6])
);

FILL FILL_1__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[0]),
    .B(_1133_),
    .C(_1008_),
    .Y(_403_)
);

NAND2X1 _2260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1303_),
    .Y(_1394_)
);

FILL FILL_2__1953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1550_),
    .Y(_1551_)
);

FILL FILL_6__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [1]),
    .B(_693_),
    .Y(_708_)
);

FILL FILL_2__2738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2318_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1090_),
    .Y(_1091_)
);

AOI21X1 _2736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[4]),
    .B(_325_),
    .C(_1284_),
    .Y(_455_)
);

NAND2X1 _2316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1431_),
    .Y(_1449_)
);

FILL FILL_1__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3274_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_36_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(rotate)
);

FILL FILL_6__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_912_),
    .B(inc),
    .C(rotate),
    .Y(_913_)
);

FILL FILL_6__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(adc_sbc),
    .B(_635_),
    .C(_631_),
    .Y(_636_)
);

FILL FILL_6__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[4]),
    .Y(_284_)
);

OAI21X1 _2125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf0),
    .B(_891_),
    .C(RDY_bF$buf3),
    .Y(_1261_)
);

FILL FILL_2__1818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_730_),
    .Y(_740_)
);

FILL FILL_2__2776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2356_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_933_),
    .C(_932_),
    .D(_967_),
    .Y(BI[0])
);

FILL FILL_7__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183150x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .Y(_490_)
);

INVX1 _2354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(op[0]),
    .Y(_118_)
);

FILL FILL_4__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .B(_1649__bF$buf1),
    .Y(_1637_)
);

OAI21X1 _3139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_767_),
    .C(_773_),
    .Y(_98_)
);

FILL FILL_7__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_1193_),
    .C(_313_),
    .Y(_314_)
);

NOR2X1 _2163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1162_),
    .Y(_1298_)
);

FILL FILL_2__1856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1644_),
    .C(_1645_),
    .Y(_1646_)
);

FILL FILL_6__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2394_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .B(_997_),
    .Y(_998_)
);

FILL FILL_6__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3179_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_340_),
    .C(_366_),
    .Y(_367_)
);

OAI21X1 _2219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf0),
    .B(_936_),
    .C(RDY_bF$buf3),
    .Y(_1354_)
);

FILL FILL_7__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_149_),
    .C(_145_),
    .Y(_1686_[1])
);

FILL FILL_8__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[2]),
    .Y(DO[2])
);

FILL FILL_6__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1347_),
    .B(_1284_),
    .Y(_809_)
);

FILL FILL_0__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_554_),
    .C(_1129__bF$buf3),
    .Y(_563_)
);

FILL FILL_6__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf1),
    .B(_989_),
    .C(_911_),
    .Y(_199_)
);

NOR2X1 _2028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1156_),
    .B(_1163_),
    .Y(_1164_)
);

FILL FILL_7__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2679_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2259_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3200_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf1),
    .B(_871_),
    .C(_868_),
    .Y(_872_)
);

FILL FILL_4__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_1035_),
    .Y(_1036_)
);

FILL FILL_8__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_191_),
    .C(_932_),
    .Y(_400_)
);

NAND3X1 _2257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .B(_1390_),
    .C(_1389_),
    .Y(_1391_)
);

FILL FILL_7__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [4]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [4]),
    .Y(_1088_)
);

FILL FILL_7__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_197_),
    .C(ADD[4]),
    .Y(_233_)
);

OAI21X1 _2066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1199_),
    .C(_1201_),
    .Y(_1202_)
);

FILL FILL_2__1759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2297_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_909_),
    .Y(_910_)
);

FILL FILL_4__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1427_),
    .B(_1423_),
    .Y(_1428_)
);

FILL FILL_2__1988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1117_),
    .C(_1122_),
    .Y(AI[7])
);

FILL FILL_5_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_946_),
    .C(_944_),
    .Y(_947_)
);

FILL FILL_5__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[0]),
    .Y(_1607_)
);

OAI21X1 _3101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf1),
    .B(_748_),
    .C(\AXYS[1] [4]),
    .Y(_753_)
);

FILL FILL_3__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x140550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Z),
    .B(_141_),
    .Y(_147_)
);

FILL FILL_6__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3330_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_84_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf4),
    .Q(\AXYS[1] [7])
);

FILL FILL_8__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_330_),
    .B(_331_),
    .C(_319_),
    .Y(_332_)
);

FILL FILL_0__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf3),
    .B(_886__bF$buf2),
    .C(_890_),
    .Y(_1333_)
);

FILL FILL_0__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3370_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _1889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_1032_),
    .C(load_only),
    .D(_1031_),
    .Y(_1033_)
);

NOR2X1 _2830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1400_),
    .Y(_531_)
);

FILL FILL_8__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(ADD[4]),
    .C(PC[12]),
    .D(_163_),
    .Y(_165_)
);

FILL FILL_0__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2641_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf5),
    .B(DIHOLD[3]),
    .Y(_856_)
);

FILL FILL_8__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[3]),
    .C(_1509_),
    .D(_1652_),
    .Y(_1510_)
);

NAND2X1 _3004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(Z),
    .B(_666_),
    .Y(_671_)
);

FILL FILL_1__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1049_),
    .B(_1053_),
    .C(_1050_),
    .Y(_1054_)
);

FILL FILL_0__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3233_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1483_[0]),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(state[0])
);

FILL FILL_1__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3044_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1001_),
    .B(_1219__bF$buf0),
    .C(_606_),
    .Y(_50_)
);

AOI21X1 _2504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .B(_190_),
    .C(_248_),
    .Y(_249_)
);

FILL FILL_1__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x117150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[0]),
    .C(_1660_),
    .Y(_1548_)
);

FILL FILL_6__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(_699_),
    .C(_704_),
    .Y(_705_)
);

FILL FILL_2__2735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2315_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(_398_),
    .C(RDY_bF$buf8),
    .Y(_453_)
);

NOR2X1 _2313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1443_),
    .B(_1445_),
    .Y(_1446_)
);

FILL FILL_1__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1677_),
    .C(_1598_),
    .D(_1603_),
    .Y(_1604_)
);

FILL FILL_1__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3271_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_33_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(op[1])
);

FILL FILL_6__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3082_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .Y(_633_)
);

FILL FILL_6__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .Y(_282_)
);

NAND2X1 _2122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_1255_),
    .Y(_1258_)
);

FILL FILL_2__1815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3327_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_81_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[1] [4])
);

FILL FILL_1__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .Y(_738_)
);

FILL FILL_2__2773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2353_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_891_),
    .C(_964_),
    .Y(_965_)
);

FILL FILL_4__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf2),
    .B(_486_),
    .C(_1120_),
    .Y(_487_)
);

NOR2X1 _2351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1475_),
    .B(_1481_),
    .Y(_1482_)
);

FILL FILL_4__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1634_),
    .B(_1635_),
    .C(_1633_),
    .Y(_1492_)
);

FILL FILL_6__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [4]),
    .B(_767_),
    .Y(_772_)
);

FILL FILL_7__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1304_),
    .Y(_528_)
);

AOI21X1 _2407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_127_),
    .B(PC[4]),
    .C(_161_),
    .Y(_162_)
);

FILL FILL_1__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _2580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .Y(_1_)
);

INVX1 _2160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .Y(_1295_)
);

FILL FILL_2__1853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x23550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[5]),
    .B(ADD[4]),
    .Y(_1643_)
);

FILL FILL_2__2638_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[2]),
    .B(state[3]),
    .Y(_995_)
);

FILL FILL_6__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[2]),
    .B(_336_),
    .Y(_364_)
);

OAI21X1 _2216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1172_),
    .B(_1350_),
    .C(_1315_),
    .Y(_1351_)
);

FILL FILL_7__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[9]),
    .Y(AB[9])
);

FILL FILL_6__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .B(_805_),
    .Y(_806_)
);

FILL FILL_2__2867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf3),
    .B(_893_),
    .Y(_1051_)
);

FILL FILL_7__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_1129__bF$buf0),
    .C(_561_),
    .D(_535_),
    .Y(_36_)
);

FILL FILL_6__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_195_),
    .Y(_196_)
);

OAI21X1 _2025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf3),
    .B(_863_),
    .C(_1160_),
    .Y(_1161_)
);

FILL FILL_0__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2676_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2256_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[5]),
    .B(state[4]),
    .Y(_869_)
);

FILL FILL_4__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_395_),
    .C(_385_),
    .Y(_398_)
);

INVX1 _2254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .Y(_1388_)
);

FILL FILL_2__1947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x62550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1544_),
    .Y(_1545_)
);

OAI21X1 _3039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_701_),
    .C(ADD[1]),
    .Y(_702_)
);

FILL FILL_7__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[3]),
    .C(_1085_),
    .Y(_1086_)
);

FILL FILL_5__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_208_),
    .C(_230_),
    .Y(_231_)
);

NAND2X1 _2063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf1),
    .B(_883_),
    .Y(_1199_)
);

FILL FILL_2__1756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3268_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_30_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(clv)
);

FILL FILL_6__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2294_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_906_),
    .C(_886__bF$buf0),
    .Y(_907_)
);

FILL FILL_4__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x105450 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .Y(_630_)
);

AOI22X1 _2539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[3]),
    .B(_1075_),
    .C(_200_),
    .D(ADD[3]),
    .Y(_279_)
);

AOI22X1 _2119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf6),
    .B(_1185_),
    .C(_1254_),
    .D(_1253_),
    .Y(_1255_)
);

FILL FILL_7__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .B(_887__bF$buf2),
    .C(_853__bF$buf3),
    .Y(_1425_)
);

FILL FILL_2__1985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1538_),
    .B(_1567_),
    .C(_1578_),
    .Y(_1583_)
);

FILL FILL_6__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_734_),
    .C(_1281_),
    .Y(_735_)
);

FILL FILL_0__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .Y(_1120_)
);

FILL FILL_4__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf4),
    .B(_299_),
    .Y(_485_)
);

AND2X2 _2348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(_1262_),
    .Y(_1479_)
);

FILL FILL_7__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2302_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_943_),
    .B(_942_),
    .Y(_944_)
);

FILL FILL_5__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(N),
    .B(_659_),
    .Y(_665_)
);

FILL FILL_6__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_1031_),
    .Y(\u_ALU8.BCD )
);

NAND3X1 _2157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1252_),
    .B(_1292_),
    .C(_1271_),
    .Y(_1293_)
);

FILL FILL_7__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2388_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf2),
    .B(_927_),
    .Y(_992_)
);

FILL FILL_7__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_144_),
    .C(_136_),
    .Y(_1686_[0])
);

FILL FILL_8__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x39150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x97650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2340_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x11850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1329_),
    .Y(_1330_)
);

FILL FILL_0__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2816_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1029_),
    .B(_951_),
    .Y(_1030_)
);

FILL FILL_8__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2625_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2205_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf2),
    .B(DIHOLD[2]),
    .Y(_854_)
);

FILL FILL_8__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[4]),
    .Y(_1507_)
);

NAND2X1 _3001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[1]),
    .B(_1260_),
    .Y(_668_)
);

FILL FILL_5__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3219_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _2289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .B(_959_),
    .S(_853__bF$buf3),
    .Y(_1422_)
);

FILL FILL_0__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1108_),
    .B(_830__bF$buf1),
    .C(_847_),
    .Y(_115_)
);

FILL FILL_3_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_603_),
    .C(_593_),
    .Y(_604_)
);

INVX1 _2501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[6]),
    .Y(_246_)
);

FILL FILL_5__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2663_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2243_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1233_),
    .B(_1226_),
    .Y(_1234_)
);

FILL FILL_0__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2312_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2719_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .Y(_941_)
);

FILL FILL_4__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_445_),
    .C(_449_),
    .Y(_450_)
);

NAND2X1 _2310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(_1389_),
    .Y(_1443_)
);

FILL FILL_0__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1600_),
    .Y(_1601_)
);

FILL FILL_1__2892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3324_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_78_),
    .S(vdd),
    .R(_1__bF$buf4),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[1] [1])
);

FILL FILL_1__2281_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7_BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2350_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf0),
    .B(_961_),
    .C(_907_),
    .Y(_962_)
);

FILL FILL_0__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2337_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[4]),
    .B(_1649__bF$buf3),
    .Y(_1633_)
);

FILL FILL_6__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_767_),
    .C(_770_),
    .Y(_95_)
);

FILL FILL_1__2090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3364_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_525_),
    .Y(_526_)
);

NAND3X1 _2404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_159_),
    .C(_155_),
    .Y(_1686_[3])
);

FILL FILL_1__1781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x27450 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3362_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_115_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf7),
    .Q(ABH[6])
);

FILL FILL_2__2635_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x85950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[3]),
    .B(_321_),
    .C(_360_),
    .Y(_361_)
);

NOR2X1 _2213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1330_),
    .Y(_1348_)
);

FILL FILL_2__1906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .B(_1502_),
    .C(_1499_),
    .Y(_1504_)
);

FILL FILL_1__2795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[6]),
    .Y(AB[6])
);

FILL FILL_6__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1277_),
    .Y(_803_)
);

FILL FILL_2__2864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2024_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf1),
    .B(_946_),
    .Y(_1048_)
);

FILL FILL_0__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_537_),
    .Y(_560_)
);

FILL FILL_6__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_899_),
    .B(_892_),
    .Y(_193_)
);

OAI21X1 _2022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf1),
    .B(_864_),
    .C(_1157_),
    .Y(_1158_)
);

FILL FILL_8_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[13]),
    .B(_830__bF$buf0),
    .Y(_846_)
);

FILL FILL_1__2184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2673_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2253_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[3]),
    .Y(_866_)
);

FILL FILL_4__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_600_),
    .B(_601_),
    .Y(_602_)
);

FILL FILL_1__1875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_343_),
    .C(_394_),
    .Y(_395_)
);

OAI21X1 _2251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1215_),
    .C(_1384_),
    .Y(_1385_)
);

FILL FILL_2__1944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .Y(_1542_)
);

FILL FILL_6__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(HC),
    .B(_698_),
    .C(_697_),
    .Y(_699_)
);

FILL FILL_7__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2309_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2062_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .Y(_1083_)
);

FILL FILL_5__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[3]),
    .B(_325_),
    .C(_338_),
    .D(ABH[3]),
    .Y(_447_)
);

NAND2X1 _2307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1396_),
    .B(_1317_),
    .Y(_1440_)
);

FILL FILL_7__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[3]),
    .Y(_228_)
);

NAND3X1 _2060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(_1195_),
    .C(_1192_),
    .Y(_1196_)
);

FILL FILL_2__1753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3265_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_27_),
    .S(vdd),
    .R(_1__bF$buf6),
    .CLK(clk_bF$buf6),
    .Q(sed)
);

FILL FILL_6__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2291_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(_885_),
    .C(_903_),
    .Y(_904_)
);

FILL FILL_6__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3076_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_620_),
    .C(_628_),
    .Y(_60_)
);

FILL FILL_6__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_208_),
    .C(_276_),
    .Y(_1685_[10])
);

OAI21X1 _2116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_942_),
    .C(_1251_),
    .Y(_1252_)
);

FILL FILL_7__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2286_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2278_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x121050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x167850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .B(_1579_),
    .Y(_1580_)
);

FILL FILL_6__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [5]),
    .B(_693_),
    .Y(_733_)
);

FILL FILL_2__2767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2347_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .Y(_959_)
);

FILL FILL_7__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .Y(_1117_)
);

FILL FILL_8__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_460_),
    .Y(_482_)
);

NAND2X1 _2345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1355_),
    .Y(_1476_)
);

FILL FILL_5__2095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2576_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3512_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3504_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .Y(_662_)
);

FILL FILL_6__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_208_),
    .C(_309_),
    .Y(_1685_[15])
);

NOR2X1 _2154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1289_),
    .B(_1286_),
    .Y(_1290_)
);

FILL FILL_2__1847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3359_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_112_),
    .S(vdd),
    .R(_1__bF$buf8),
    .CLK(clk_bF$buf7),
    .Q(ABH[3])
);

FILL FILL_0__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2385_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_871_),
    .Y(_989_)
);

FILL FILL_6__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(C),
    .B(_141_),
    .Y(_142_)
);

FILL FILL_8__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[3]),
    .Y(AB[3])
);

FILL FILL_6__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_963_),
    .Y(_800_)
);

FILL FILL_7__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3399_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_1383_),
    .C(_1219__bF$buf2),
    .Y(_558_)
);

NAND2X1 _2439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_187_),
    .Y(_190_)
);

OAI21X1 _2019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1154_),
    .C(_1145_),
    .Y(_1155_)
);

FILL FILL_7__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x15750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3550_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3130_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[4]),
    .B(_989_),
    .Y(_1327_)
);

FILL FILL_2__1885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(BI[6]),
    .C(_1670_),
    .D(_1652_),
    .Y(_1671_)
);

FILL FILL_0__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2821_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2401_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .Y(_1027_)
);

FILL FILL_8__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_974_),
    .C(_390_),
    .D(_392_),
    .Y(_8_)
);

INVX1 _2248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .Y(_1382_)
);

FILL FILL_7__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3420_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [3]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [3]),
    .Y(_1080_)
);

FILL FILL_2__3000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2630_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2622_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(DI[1]),
    .Y(_852_)
);

FILL FILL_8__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3415_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_583_),
    .B(_582_),
    .C(_1129__bF$buf2),
    .Y(_584_)
);

FILL FILL_6__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_192_),
    .Y(_225_)
);

NOR2X1 _2057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_899_),
    .Y(_1193_)
);

FILL FILL_0__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2288_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_900_),
    .Y(_901_)
);

FILL FILL_4__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1417_),
    .C(_1419_),
    .Y(_1420_)
);

FILL FILL_2__1979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2915_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2907_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [7]),
    .B(_1023_),
    .C(_1012_),
    .D(\AXYS[3] [7]),
    .Y(_1114_)
);

FILL FILL_4__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2660_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2240_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3453_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3033_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1036_),
    .Y(_1231_)
);

FILL FILL_0__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2724_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2304_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2716_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf2),
    .B(_900_),
    .Y(_938_)
);

FILL FILL_4__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3509_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1597_),
    .B(_1594_),
    .C(_1498_),
    .Y(_1598_)
);

FILL FILL_3__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2953_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3321_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_75_),
    .S(vdd),
    .R(_1__bF$buf9),
    .CLK(clk_bF$buf10),
    .Q(\AXYS[0] [6])
);

FILL FILL_5__3491_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3071_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1804_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL181950x7950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2762_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2342_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2334_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3547_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3127_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf2),
    .B(_1323_),
    .Y(_1324_)
);

FILL FILL_0__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf2),
    .B(_1612_),
    .C(_1631_),
    .Y(_1490_)
);

FILL FILL_8__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[3] [1]),
    .B(_767_),
    .Y(_769_)
);

FILL FILL_8__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2818_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(_523_),
    .C(_519_),
    .Y(_30_)
);

NAND2X1 _2401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(D),
    .B(_141_),
    .Y(_157_)
);

FILL FILL_0__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2991_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2571_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2632_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x89850 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2627_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2619_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3170_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DI[0]),
    .B(RDY_bF$buf4),
    .Y(_850_)
);

FILL FILL_4__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .Y(_358_)
);

NAND2X1 _2210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1344_),
    .B(_1332_),
    .Y(_1345_)
);

FILL FILL_2__1903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[4]),
    .B(_1500_),
    .Y(_1501_)
);

FILL FILL_1__2792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3585_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1043_),
    .B(_1044_),
    .Y(_1045_)
);

FILL FILL_0__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_830__bF$buf1),
    .C(_844_),
    .Y(_112_)
);

FILL FILL_1__2181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3394_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2670_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2250_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _1710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DI[7]),
    .B(DIHOLD[7]),
    .S(RDY_bF$buf5),
    .Y(_864_)
);

FILL FILL_0__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(_1168_),
    .C(_1214_),
    .Y(_599_)
);

FILL FILL_1__1872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2665_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2245_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2657_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2237_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[0]),
    .B(_1653_),
    .Y(_1539_)
);

FILL FILL_6__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_695_),
    .C(_696_),
    .Y(_69_)
);

FILL FILL_2__2726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2306_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1928_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_398_),
    .Y(_444_)
);

NAND3X1 _2304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1346_),
    .B(_1436_),
    .C(_1294_),
    .Y(_1437_)
);

FILL FILL_5__2894_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2054_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(alu_op[2]),
    .C(_1497_),
    .Y(_1595_)
);

FILL FILL_1__2886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3262_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_24_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(clc)
);

FILL FILL_6__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182250x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3073_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[6]),
    .Y(_627_)
);

FILL FILL_6__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABH[2]),
    .B(_1075_),
    .C(_200_),
    .D(ADD[2]),
    .Y(_274_)
);

NAND3X1 _2113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(_1223_),
    .C(_1248_),
    .Y(_1249_)
);

FILL FILL_2__1806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2283_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3318_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_72_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[0] [3])
);

FILL FILL_1__2695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2275_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3488_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3068_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

MUX2X1 _3491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(_1575_),
    .S(_1535_),
    .Y(_1577_)
);

FILL FILL_6__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_293_),
    .B(_728_),
    .Y(_730_)
);

FILL FILL_2__2764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2344_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_953_),
    .B(_955_),
    .C(_869__bF$buf3),
    .Y(_956_)
);

FILL FILL_4__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2759_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2339_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_478_),
    .C(_477_),
    .Y(_479_)
);

OAI21X1 _2342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf0),
    .B(_1192_),
    .C(_1426_),
    .Y(_1473_)
);

FILL FILL_5__2092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ADD[1]),
    .B(_1649__bF$buf2),
    .Y(_1630_)
);

FILL FILL_6__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_1012_),
    .Y(_767_)
);

FILL FILL_7__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2573_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2153_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1783_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_520_),
    .Y(_521_)
);

FILL FILL_1__1775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2568_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .B(_631_),
    .C(_658_),
    .Y(_659_)
);

FILL FILL_6__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(_306_),
    .Y(_307_)
);

NOR2X1 _2151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf4),
    .B(_961_),
    .Y(_1287_)
);

FILL FILL_2__1844_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3356_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_109_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(ABH[0])
);

FILL FILL_0__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2629_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2209_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182550x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

CLKBUF1 CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL FILL_2__2382_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .Y(_986_)
);

FILL FILL_6__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(_343_),
    .C(_355_),
    .Y(_356_)
);

NAND2X1 _2207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf6),
    .B(_943_),
    .Y(_1342_)
);

FILL FILL_7__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2369_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(php),
    .B(_138_),
    .C(_1192_),
    .Y(_139_)
);

FILL FILL_8__2620_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2200_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2446_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[14]),
    .Y(AB[14])
);

FILL FILL_6__2026_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_1193_),
    .Y(_797_)
);

FILL FILL_0__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2438_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2018_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3405_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x121050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1822_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2607_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2191_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3396_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .Y(_555_)
);

FILL FILL_6__1717_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_186_),
    .Y(_187_)
);

OAI21X1 _2016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf0),
    .B(_859_),
    .C(_1151_),
    .Y(_1152_)
);

FILL FILL_7__2780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2360_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1709_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1882_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2675_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2255_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_shift_right),
    .B(AI[7]),
    .Y(_1668_)
);

FILL FILL_2__2667_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2247_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3214_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf2),
    .B(DIHOLD[6]),
    .Y(_862_)
);

FILL FILL_4__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _1880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[2] [0]),
    .B(_1023_),
    .C(_1022_),
    .D(\AXYS[1] [0]),
    .Y(_1024_)
);

FILL FILL_8__1700_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3603_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1946_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_385_),
    .Y(_390_)
);

NAND3X1 _2245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1372_),
    .C(_1378_),
    .Y(_1379_)
);

FILL FILL_2__1938_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2905_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3374_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1691_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2476_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3443_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2056_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3023_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[2]),
    .C(_1077_),
    .Y(_1078_)
);

FILL FILL_7__1860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2645_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3412_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3404_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_520_),
    .Y(_581_)
);

FILL FILL_6__1755_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1073_),
    .B(_182_),
    .C(_222_),
    .Y(_223_)
);

INVX1 _2054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1189_),
    .Y(_1190_)
);

FILL FILL_2__1747_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2714_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3259_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_21_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf5),
    .Q(cond_code[2])
);

FILL FILL_7__3183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1916_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2293_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2285_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869__bF$buf0),
    .B(_897_),
    .Y(_898_)
);

FILL FILL_4__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2874_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3221_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1984_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1345_),
    .Y(_1417_)
);

FILL FILL_2__1976_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2943_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2523_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2103_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2769_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1572_),
    .B(_1573_),
    .C(_1571_),
    .Y(_1574_)
);

FILL FILL_6__2349_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CO),
    .B(_698_),
    .C(_726_),
    .Y(_727_)
);

FILL FILL_0__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2912_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2094_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2904_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _1974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(ADD[6]),
    .C(_1111_),
    .Y(_1112_)
);

FILL FILL_4__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1264_),
    .B(_413_),
    .C(DIMUX[6]),
    .Y(_476_)
);

NAND3X1 _2339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1218_),
    .C(_1307_),
    .Y(_1470_)
);

FILL FILL_7__2683_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2263_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3450_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3030_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1793_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf2),
    .B(_946_),
    .Y(_1228_)
);

FILL FILL_2__1785_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2752_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2332_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2578_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2158_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3297_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[7]),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf9),
    .Q(DIHOLD[7])
);

FILL FILL184050x156150 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3117_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2721_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2301_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2319_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_899_),
    .B(_874_),
    .Y(_935_)
);

FILL FILL_4__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3506_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(_655_),
    .C(_656_),
    .Y(_64_)
);

FILL FILL_6__1849_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .Y(_304_)
);

INVX2 _2148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051__bF$buf3),
    .Y(_1284_)
);

FILL FILL_7__2492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2808_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2981_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2561_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2141_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x171750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2387_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2379_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_983_)
);

FILL FILL_7__1763_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2950_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1832_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1352_),
    .Y(_506_)
);

NAND2X1 _2377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_1025_),
    .Y(_136_)
);

FILL FILL_8__2617_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1819_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2370_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2188_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3155_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2357_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2331_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3224_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3544_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3124_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1887_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1320_),
    .Y(_1321_)
);

FILL FILL_2__1879_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2846_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2426_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2006_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2400_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2815_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2807_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [0]),
    .B(_1020_),
    .Y(_1021_)
);

FILL FILL_0__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .Y(WE)
);

FILL FILL_1__2980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1870_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1688_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2655_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2235_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1857_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2624_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8_BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2616_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1926_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3409_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1900_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .B(_1683_),
    .Y(_1498_)
);

FILL FILL_3__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3582_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3162_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2884_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2464_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2044_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2853_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1735_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3218_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2502_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_830__bF$buf0),
    .C(_842_),
    .Y(_111_)
);

FILL FILL_2__2914_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3391_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1704_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2273_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2909_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3058_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_596_),
    .Y(_597_)
);

FILL FILL_3__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2662_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2242_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2654_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2234_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1964_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3447_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3027_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf1),
    .B(_946_),
    .C(_853__bF$buf6),
    .Y(_1225_)
);

FILL FILL_0__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2749_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2731_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(BI[1]),
    .C(_1660_),
    .Y(_1536_)
);

FILL FILL_6__2311_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2329_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_949_),
    .C(_263_),
    .Y(_694_)
);

FILL FILL_2__2723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2303_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2082_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2718_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_417_),
    .Y(_442_)
);

OR2X2 _2301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1219__bF$buf3),
    .Y(_1434_)
);

FILL FILL_0__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2891_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2051_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1504_),
    .B(_1591_),
    .C(_1589_),
    .Y(_1592_)
);

FILL FILL_1__2883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1773_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2978_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2558_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2138_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2532_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2112_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2947_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3070_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_620_),
    .C(_625_),
    .Y(_57_)
);

FILL FILL_8__1829_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1811_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_208_),
    .C(_271_),
    .Y(_1685_[9])
);

OAI21X1 _2110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf7),
    .B(_1244_),
    .C(_1245_),
    .Y(_1246_)
);

FILL FILL_2__1803_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2298_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2280_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3315_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_69_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf0),
    .Q(\AXYS[0] [0])
);

FILL FILL_1__2692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2272_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__3165_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3485_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3065_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2787_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2367_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2341_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _1801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_879_),
    .Y(_953_)
);

FILL FILL_0__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2856_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2756_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2336_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2748_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2328_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2825_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1570_),
    .C(_1571_),
    .Y(_1628_)
);

FILL FILL_6__2405_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_757_),
    .C(_765_),
    .Y(_91_)
);

FILL FILL_1__2081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2817_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__1707_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2596_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2176_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2570_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2150_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1780_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1798_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(_510_),
    .C(_518_),
    .Y(_29_)
);

FILL FILL_1__1772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2985_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2565_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2145_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2977_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1867_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1841_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2634_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2214_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3353_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_106_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf9),
    .Q(ABL[5])
);

FILL FILL_2__2626_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2206_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3095_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1836_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1905_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(ABL[2]),
    .B(_338_),
    .Y(_353_)
);

MUX2X1 _2204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(C),
    .B(N),
    .S(cond_code[2]),
    .Y(_1339_)
);

FILL FILL182550x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2794_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2374_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1682_),
    .B(_1681_),
    .C(_1678_),
    .Y(_1683_)
);

FILL FILL_1__2786_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3579_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3159_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2443_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[11]),
    .Y(AB[11])
);

FILL FILL_6__2023_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .Y(_794_)
);

FILL FILL_2__2855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2435_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3402_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2015_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2604_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3393_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_551_),
    .Y(_552_)
);

FILL FILL_6__1714_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1274_),
    .B(_1048_),
    .Y(_184_)
);

NAND2X1 _2013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1148_),
    .Y(_1149_)
);

FILL FILL_2__1706_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2183_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2919_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[9]),
    .B(_830__bF$buf3),
    .Y(_841_)
);

FILL FILL_1__2595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3388_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2672_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf0),
    .B(_1664_),
    .C(_1665_),
    .Y(_1485_)
);

FILL FILL_6__2252_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2664_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2244_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3211_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(DIHOLD[5]),
    .Y(_860_)
);

FILL FILL_4__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1874_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _2909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_498_),
    .C(_551_),
    .Y(_594_)
);

FILL FILL_1__1866_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2413_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2659_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2239_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3600_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1943_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_359_),
    .C(_1051__bF$buf0),
    .Y(_387_)
);

OAI21X1 _2242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf0),
    .B(_1287_),
    .C(_1370_),
    .Y(_1376_)
);

FILL FILL_2__1935_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2902_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2728_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[0]),
    .B(_1532_),
    .Y(_1533_)
);

FILL FILL_6__2308_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_690_),
    .C(RDY_bF$buf2),
    .Y(_691_)
);

FILL FILL_7__3371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3197_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3189_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2499_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2481_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2079_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2061_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2473_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2053_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _1933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_918__bF$buf0),
    .C(_889_),
    .Y(_1075_)
);

FILL FILL_0__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x101550 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _2718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_438_),
    .C(_436_),
    .Y(_439_)
);

FILL FILL_7__2642_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2222_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2988_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2888_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2468_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2048_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3401_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_578_),
    .C(_577_),
    .Y(_579_)
);

FILL FILL_6__1752_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[2]),
    .B(_204_),
    .C(_202_),
    .D(ABL[2]),
    .Y(_220_)
);

OAI21X1 _2051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918__bF$buf2),
    .B(_936_),
    .C(_1186_),
    .Y(_1187_)
);

FILL FILL_2__1744_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2537_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2117_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3256_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_18_),
    .S(vdd),
    .R(_1__bF$buf2),
    .CLK(clk_bF$buf8),
    .Q(NMI_edge)
);

FILL FILL_7__3180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2529_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2109_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1913_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x136650 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1739_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2290_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2282_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf3),
    .B(_891_),
    .C(_894_),
    .Y(_895_)
);

FILL FILL_6__3495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(reset),
    .B(_618_),
    .C(IRHOLD[3]),
    .Y(_624_)
);

FILL FILL_6__1808_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(ADD[1]),
    .C(_1066_),
    .Y(_269_)
);

NOR2X1 _2107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1237_),
    .B(_1242_),
    .Y(_1243_)
);

FILL FILL_7__2871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2451_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2031_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9__2797_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2697_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2277_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2689_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2269_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3210_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1999_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1981_ (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _2280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1413_),
    .Y(_1414_)
);

FILL FILL_2__1973_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2520_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2100_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2766_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1663_),
    .B(_1570_),
    .C(_1547_),
    .Y(_1571_)
);

FILL FILL_6__2346_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [4]),
    .B(_693_),
    .Y(_725_)
);

FILL FILL_0__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2338_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1722_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1968_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2507_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2091_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2901_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1108_),
    .B(_872_),
    .Y(_1109_)
);

NAND2X1 _2756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[13]),
    .B(_323_),
    .Y(_473_)
);

NOR2X1 _2336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1423_),
    .B(_1325_),
    .Y(_1468_)
);

FILL FILL_7__2680_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2260_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2086_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2498_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2078_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1790_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1782_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2575_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2155_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3294_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[4]),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf9),
    .Q(DIHOLD[4])
);

FILL FILL_2__2987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2567_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2147_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3114_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1951_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1777_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1769_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2316_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2710_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[0]),
    .Y(_932_)
);

FILL FILL_5__3503_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_652_),
    .C(_978_),
    .Y(_654_)
);

FILL FILL_6__1846_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(DIMUX[6]),
    .C(_301_),
    .Y(_302_)
);

INVX4 _2145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_981_),
    .Y(_1281_)
);

FILL FILL_2__1838_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2805_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2384_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2376_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_980_)
);

FILL FILL_7__1760_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1998_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2545_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2125_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .Y(_691__bF$buf3)
);

BUFX2 BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .Y(_691__bF$buf2)
);

BUFX2 BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .Y(_691__bF$buf1)
);

BUFX2 BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .Y(_691__bF$buf0)
);

BUFX2 BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1219__bF$buf3)
);

BUFX2 BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1219__bF$buf2)
);

BUFX2 BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1219__bF$buf1)
);

BUFX2 BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1219__bF$buf0)
);

NAND2X1 _2794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .B(_503_),
    .Y(_504_)
);

OAI21X1 _2374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf0),
    .B(_901_),
    .C(_1188_),
    .Y(_134_)
);

FILL FILL_8__2614_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_[0]),
    .Y(AB[0])
);

NOR2X1 _3159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_790_),
    .Y(_791_)
);

FILL FILL_7__3083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1816_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183450x35250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2193_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2185_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3152_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2774_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2354_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3541_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3121_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3533_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3113_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1884_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1317_),
    .B(_1219__bF$buf3),
    .Y(_1318_)
);

FILL FILL_2__1876_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2843_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2423_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2003_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2669_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _3388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[2]),
    .B(_1660_),
    .Y(_1663_)
);

FILL FILL_6__2249_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2812_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2804_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1006_),
    .B(_1007_),
    .C(_1017_),
    .Y(_1018_)
);

FILL FILL_2__3199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(_973_),
    .C(_384_),
    .D(_379_),
    .Y(_7_)
);

OAI21X1 _2239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf2),
    .B(_961_),
    .C(RDY_bF$buf3),
    .Y(_1373_)
);

FILL FILL_7__2583_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2163_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _3600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_[5]),
    .Y(DO[5])
);

FILL FILL_3__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3368_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1693_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2652_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2232_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2478_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2058_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(_828_),
    .C(RDY_bF$buf5),
    .Y(_829_)
);

FILL FILL_0__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3017_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1854_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2639_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2621_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2201_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2219_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2613_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x171750 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1923_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3406_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf1),
    .C(store),
    .Y(_576_)
);

FILL FILL_6__1749_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1063_),
    .B(_182_),
    .C(_217_),
    .Y(_218_)
);

NAND2X1 _2048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886__bF$buf3),
    .B(_897_),
    .Y(_1184_)
);

FILL FILL_7__2392_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2708_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3151_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2461_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2041_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL183750x74250 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2287_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2279_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3220_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[3]),
    .B(_873_),
    .Y(_892_)
);

FILL FILL_4__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2850_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2430_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2448_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2028_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2010_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2842_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2422_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2002_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1732_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3215_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3207_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1978_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_260_),
    .C(_419_),
    .Y(_10_)
);

OAI21X1 _2277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf2),
    .B(_1277_),
    .C(_1410_),
    .Y(_1411_)
);

FILL FILL_0__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2937_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2517_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184050x109350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3380_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1701_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1719_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2270_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2096_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2906_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2088_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3055_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1103_),
    .B(_1105_),
    .C(_1104_),
    .Y(_1106_)
);

FILL FILL_7__1892_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2677_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2257_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2651_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2231_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1961_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3444_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3024_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3436_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3016_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1787_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219__bF$buf3),
    .B(_1221_),
    .Y(_1222_)
);

FILL FILL_2__1779_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2746_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2326_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2300_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2646_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2226_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184350x124950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2966_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2546_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2126_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1948_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1930_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1922_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1848_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2715_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2707_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _1777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_929_),
    .C(_925_),
    .Y(_930_)
);

FILL FILL_4__3184_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3084_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1917_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2486_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2066_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1817_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1506_),
    .B(_1504_),
    .Y(_1589_)
);

FILL FILL_1__2880_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2460_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2040_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2386_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1770_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1990_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2975_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2555_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2135_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2875_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2455_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2035_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6_BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2775_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2355_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1757_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1731_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2944_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2524_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2104_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2936_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2516_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1826_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1800_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1726_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2295_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3312_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_66_),
    .S(vdd),
    .R(_1__bF$buf10),
    .CLK(clk_bF$buf9),
    .Q(Z)
);

FILL FILL_3__2195_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3482_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3062_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3474_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3054_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2784_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2364_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert28 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_CLKBUF1_insert29 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2684_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2264_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2584_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2164_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1986_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3469_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3049_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1960_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1886_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3369_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2753_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2333_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x148350 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2745_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2325_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3538_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3118_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1955_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1855_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2822_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649__bF$buf3),
    .B(_1614_),
    .C(_1625_),
    .Y(_1487_)
);

FILL FILL_6__2402_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf0),
    .B(_758_),
    .C(\AXYS[2] [5]),
    .Y(_764_)
);

FILL FILL_9_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2814_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2593_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2173_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2493_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2073_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2809_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2393_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3378_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1795_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_1323_),
    .Y(_517_)
);

FILL FILL_3__1695_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3598_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3178_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2982_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2562_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2142_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2974_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2554_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2134_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3421_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3001_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1864_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1764_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2649_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2631_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2211_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3350_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_103_),
    .S(vdd),
    .R(_1__bF$buf5),
    .CLK(clk_bF$buf9),
    .Q(ABL[2])
);

FILL FILL_8__2229_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2623_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2203_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2969_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2549_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2129_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2869_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2449_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2029_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3416_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3092_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1833_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1825_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2618_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3087_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1902_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf8),
    .B(_968_),
    .C(_348_),
    .D(_350_),
    .Y(_3_)
);

INVX1 _2201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(V),
    .Y(_1336_)
);

FILL FILL_5__2791_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2371_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2389_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _3406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AI[5]),
    .B(_1679_),
    .Y(_1680_)
);

FILL FILL_1__2783_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2363_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2289_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3230_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3156_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3148_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1993_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1893_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2860_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2878_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2458_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2440_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2038_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2020_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2432_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2012_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2778_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2358_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2678_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2258_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3225_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2601_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2921_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2501_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2847_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2427_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2007_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2839_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2419_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3390_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .Y(_549_)
);

FILL FILL_6__1711_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1729_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf3),
    .B(_901_),
    .C(_1034_),
    .Y(_181_)
);

NAND2X1 _2010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IRHOLD_valid_bF$buf1),
    .B(IRHOLD[2]),
    .Y(_1146_)
);

FILL FILL_2__1703_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2180_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2198_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1949_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2916_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_259_),
    .C(_839_),
    .Y(_108_)
);

FILL FILL_1__2592_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2172_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2098_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3385_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3377_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2687_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2267_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2661_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2241_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2587_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2167_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _1701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(RDY_bF$buf4),
    .B(DIHOLD[4]),
    .Y(_858_)
);

FILL FILL_0__2487_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3454_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2067_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3034_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3446_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3026_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1871_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1889_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf1),
    .B(_1002__bF$buf0),
    .C(src_reg[0]),
    .Y(_592_)
);

FILL FILL_1__1863_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2830_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2410_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1789_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2730_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2310_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2656_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2236_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2648_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2228_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3515_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1940_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1958_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1932_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1858_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1758_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2725_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2305_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _3444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(BI[1]),
    .B(AI[1]),
    .C(_1653_),
    .Y(_1530_)
);

OAI21X1 _3024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887__bF$buf1),
    .B(_1035_),
    .C(_981_),
    .Y(_688_)
);

FILL FILL_2__2717_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3194_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3186_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1927_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2496_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2076_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1919_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2890_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2470_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2050_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2396_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[0] [2]),
    .B(_1020_),
    .Y(_1072_)
);

FILL FILL_0__2296_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1698_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_333_),
    .C(_1076_),
    .Y(_436_)
);

FILL FILL_5__2885_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2465_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2045_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2877_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2457_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2037_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3424_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3004_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1767_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1741_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert30 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert31 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert32 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert33 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert34 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert35 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL182850x163950 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert36 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert37 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4_CLKBUF1_insert38 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1987_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2954_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2534_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2114_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3253_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_16_),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf7),
    .Q(PC[14])
);

FILL FILL_2__2946_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2526_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2106_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1910_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1810_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1736_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1728_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3492_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3072_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3484_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3064_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0_BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_620_),
    .C(_622_),
    .Y(_54_)
);

FILL FILL_6__1805_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_266_),
    .Y(_1685_[8])
);

INVX1 _2104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .Y(_1240_)
);

FILL FILL_5__2694_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2274_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3309_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_63_),
    .S(vdd),
    .R(_1__bF$buf3),
    .CLK(clk_bF$buf5),
    .Q(D)
);

FILL FILL_1__2686_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2266_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3553_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3133_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1996_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3479_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3059_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1970_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1896_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1796_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2763_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _3482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1529_),
    .C(_1562_),
    .D(_1567_),
    .Y(_1568_)
);

FILL FILL_6__2343_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_721_),
    .C(_722_),
    .Y(_72_)
);

FILL FILL_2__2755_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2335_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3202_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3548_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3128_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3522_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3102_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1965_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1957_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2924_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2504_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2824_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2404_ (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _2753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(_469_),
    .Y(_471_)
);

OR2X2 _2333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1464_),
    .B(_1463_),
    .Y(_1465_)
);

FILL FILL_5__2083_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2819_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _3538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1609_),
    .B(_1623_),
    .C(_1649__bF$buf3),
    .Y(_1624_)
);

OAI21X1 _3118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_757_),
    .C(_762_),
    .Y(_88_)
);

FILL FILL_1__2495_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3462_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2075_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3042_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2992_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2572_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2152_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3291_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(DIMUX[1]),
    .S(vdd),
    .R(_1__bF$buf0),
    .CLK(clk_bF$buf2),
    .Q(DIHOLD[1])
);

FILL FILL_2__2984_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2564_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3531_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2144_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3111_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3431_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3011_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1774_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_1129__bF$buf0),
    .C(_513_),
    .D(_510_),
    .Y(_27_)
);

FILL FILL_1__1766_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2733_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2313_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2633_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2213_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2979_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2559_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2139_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3500_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3518_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3418_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _2982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(sei),
    .B(_649_),
    .C(_951_),
    .D(_650_),
    .Y(_651_)
);

FILL FILL_6__1843_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(PC[14]),
    .Y(_299_)
);

OAI21X1 _2142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf1),
    .B(_1032_),
    .C(RDY_bF$buf0),
    .Y(_1278_)
);

FILL FILL_2__1835_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2802_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2702_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2628_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3347_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_100_),
    .S(vdd),
    .R(_1__bF$buf1),
    .CLK(clk_bF$buf3),
    .Q(\AXYS[3] [7])
);

FILL FILL_6__2208_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2602_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3591_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3171_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3097_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3089_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1904_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2399_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2381_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2793_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2373_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2299_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_926__bF$buf2),
    .B(_897_),
    .Y(_977_)
);

FILL FILL_0__2199_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3586_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3166_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3560_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3140_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3158_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x136650 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_340_),
    .Y(_348_)
);

FILL FILL_1__1995_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2962_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2542_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2122_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2862_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2442_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2022_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2788_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2368_ (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1129__bF$buf4)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1129__bF$buf3)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1129__bF$buf2)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1129__bF$buf1)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1129__bF$buf0)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .Y(_830__bF$buf3)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .Y(_830__bF$buf2)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .Y(_830__bF$buf1)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .Y(_830__bF$buf0)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .Y(_918__bF$buf3)
);

FILL FILL_3__3227_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _2791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(plp),
    .Y(_502_)
);

INVX1 _2371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(op[3]),
    .Y(_132_)
);

FILL FILL_8__2611_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2931_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2511_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2857_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3576_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_1494_),
    .S(vdd),
    .R(_1484_),
    .CLK(clk_bF$buf4),
    .Q(ADD[6])
);

FILL FILL_6__2437_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2017_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_936_),
    .C(_1184_),
    .Y(_788_)
);

FILL FILL_7__3080_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2849_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2831_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2429_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2411_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2009_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1813_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1713_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2190_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2182_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2918_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3395_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3387_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1178_),
    .Y(_546_)
);

FILL FILL_6__1708_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _2427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(AN),
    .B(_139_),
    .C(_178_),
    .Y(_179_)
);

INVX1 _2007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(I),
    .Y(_1143_)
);

FILL FILL_7__2771_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2351_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2671_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2251_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2597_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2177_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2589_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2169_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3556_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3136_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3530_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3110_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3456_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3036_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1881_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1899_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _2180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1314_),
    .Y(_1315_)
);

FILL FILL_2__1873_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2840_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2420_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2000_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1799_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2740_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2320_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1699_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2666_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX4 _3385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(alu_op[3]),
    .Y(_1660_)
);

FILL FILL_6__2246_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2658_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2640_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2238_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2220_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3205_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3525_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3105_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1942_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3425_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3005_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__1868_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2827_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2407_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2801_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2727_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2307_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _1871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1003_),
    .Y(_1015_)
);

FILL FILL_2__3196_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1937_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_372_),
    .C(_381_),
    .D(_377_),
    .Y(_382_)
);

OAI21X1 _2236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_887__bF$buf4),
    .C(_853__bF$buf0),
    .Y(_1370_)
);

FILL FILL_7__2580_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2160_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1929_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1911_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2480_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2060_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2398_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3365_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1690_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2895_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2475_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2055_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_937_),
    .B(_821_),
    .C(_822_),
    .Y(_826_)
);

FILL FILL_2__2887_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2467_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3434_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2047_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3014_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _1927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1064_),
    .C(_1069_),
    .Y(AI[1])
);

FILL FILL_7__1851_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1751_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2636_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2216_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2610_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2956_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2536_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2116_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1920_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3403_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1820_ (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _2885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_1219__bF$buf2),
    .Y(_574_)
);

FILL FILL_6__1746_ (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _2465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DIMUX[1]),
    .B(_204_),
    .C(_202_),
    .D(ABL[1]),
    .Y(_215_)
);

NAND3X1 _2045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf2),
    .B(_1168_),
    .C(_1180_),
    .Y(_1181_)
);

FILL FILL_2__1738_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1720_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2705_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2605_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3594_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3174_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2925_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2505_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3494_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3074_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1907_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1807_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2284_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2696_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2276_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(state[1]),
    .B(_888_),
    .Y(_889_)
);

FILL FILL_4__3563_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3143_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3489_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3069_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1980_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3463_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3043_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__1898_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2865_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2445_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2025_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2765_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2345_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3212_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3204_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1975_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_367_),
    .Y(_417_)
);

AOI22X1 _2274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_951_),
    .C(_1385_),
    .D(_1129__bF$buf4),
    .Y(_1408_)
);

FILL FILL_2__1967_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2934_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2514_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2834_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2414_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _3479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .Y(_1565_)
);

OAI21X1 _3059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_717_),
    .C(_981_),
    .Y(_720_)
);

FILL FILL_0__2734_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2314_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1716_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3519_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2093_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2903_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3472_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2085_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3052_ (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _1965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\AXYS[1] [6]),
    .B(_1022_),
    .Y(_1103_)
);

FILL FILL_4__3372_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2674_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2254_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2994_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2574_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2154_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3459_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3441_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3039_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3021_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3433_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3013_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1784_ (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _2083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129__bF$buf3),
    .Y(_1219_)
);

FILL FILL_5_BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__1776_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2743_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2323_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5_BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2643_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2223_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2989_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2569_ (
    .gnd(gnd),
    .vdd(vdd)
);

DFFSR _3288_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_50_),
    .S(vdd),
    .R(_1__bF$buf7),
    .CLK(clk_bF$buf1),
    .Q(dst_reg[1])
);

FILL FILL_6__2149_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2963_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2543_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3528_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__3510_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2123_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3108_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3502_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1945_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3428_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3008_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1845_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2712_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2704_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(_874_),
    .Y(_927_)
);

FILL FILL_4__3181_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3081_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3099_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1914_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .B(_648_),
    .C(_645_),
    .Y(_63_)
);

OAI21X1 _2559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_268_),
    .C(_296_),
    .Y(_297_)
);

OAI21X1 _2139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882__bF$buf1),
    .B(_989_),
    .C(RDY_bF$buf0),
    .Y(_1275_)
);

FILL FILL_7__2483_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2063_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1814_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1568_),
    .C(_1515_),
    .Y(_1586_)
);

FILL FILL_3__2383_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3588_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3168_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2972_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2552_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2132_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2872_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2452_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2032_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2798_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2378_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _3097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691__bF$buf1),
    .B(_748_),
    .C(\AXYS[1] [2]),
    .Y(_751_)
);

FILL FILL_0__2772_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2352_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1754_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3557_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3137_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2941_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2959_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2521_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2539_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2119_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2101_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3090_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2933_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2513_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2859_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2439_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2019_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1823_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1723_ (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _2788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853__bF$buf7),
    .B(_1303_),
    .C(_500_),
    .Y(_20_)
);

NAND3X1 _2368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_129_),
    .C(_128_),
    .Y(_130_)
);

FILL FILL_7__2292_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2608_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2192_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2928_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2508_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3497_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__3077_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2828_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2408_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3471_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3051_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__3397_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2781_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2361_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2681_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2261_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__2187_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2581_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2599_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2161_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2179_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3566_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3146_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3540_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__3120_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__1983_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3466_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__3046_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1883_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3366_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2750_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2768_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2330_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2348_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2742_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2322_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2668_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2248_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3535_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__3115_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3527_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__3107_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1952_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_6__1878_ (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _2597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_1133_),
    .Y(_328_)
);

NAND2X1 _2177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1309_),
    .B(_1311_),
    .Y(_1312_)
);

FILL FILL_0__1852_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2837_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2417_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_9_BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_2__2811_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2737_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2317_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2637_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2217_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2590_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__2170_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1939_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2490_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__2070_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_5__2806_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__2390_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__3375_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL184650x124950 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _1868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1004_),
    .B(_1011_),
    .Y(_1012_)
);

FILL FILL_7__1792_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3595_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__1692_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__3175_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2997_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2577_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_7__2157_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_0__1908_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2971_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2551_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_1__2131_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2897_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2477_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_3__2057_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_8__1861_ (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL_4__1761_ (
    .gnd(gnd),
    .vdd(vdd)
);

endmodule
