magic
tech scmos
magscale 1 2
timestamp 1727908185
<< nwell >>
rect -14 134 132 252
<< ntransistor >>
rect 24 14 28 54
rect 32 14 36 54
rect 53 14 57 54
rect 61 14 65 54
<< ptransistor >>
rect 20 146 24 226
rect 40 146 44 226
rect 60 146 64 226
rect 80 146 84 226
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 32 54
rect 36 14 39 54
rect 51 14 53 54
rect 57 14 61 54
rect 65 14 67 54
<< pdiffusion >>
rect 18 148 20 226
rect 6 146 20 148
rect 24 160 26 226
rect 38 160 40 226
rect 24 146 40 160
rect 44 148 46 226
rect 58 148 60 226
rect 44 146 60 148
rect 64 212 80 226
rect 64 146 66 212
rect 78 146 80 212
rect 84 146 86 226
<< ndcontact >>
rect 10 14 22 54
rect 39 14 51 54
rect 67 14 79 54
<< pdcontact >>
rect 6 148 18 226
rect 26 160 38 226
rect 46 148 58 226
rect 66 146 78 212
rect 86 146 98 226
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 234 126 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 80 226 84 230
rect 20 124 24 146
rect 40 124 44 146
rect 11 118 24 124
rect 32 118 44 124
rect 11 109 17 118
rect 32 103 36 118
rect 60 103 64 146
rect 80 124 84 146
rect 80 118 90 124
rect 84 109 90 118
rect 11 83 17 97
rect 60 91 63 103
rect 11 71 28 83
rect 24 54 28 71
rect 32 54 36 91
rect 60 82 64 91
rect 53 71 64 82
rect 53 54 57 71
rect 84 63 90 97
rect 61 59 90 63
rect 61 54 65 59
rect 24 10 28 14
rect 32 10 36 14
rect 53 10 57 14
rect 61 10 65 14
<< polycontact >>
rect 5 97 17 109
rect 25 91 37 103
rect 63 91 75 103
rect 84 97 96 109
<< metal1 >>
rect -6 246 126 248
rect -6 232 126 234
rect 26 226 38 232
rect 18 148 46 154
rect 58 218 86 226
rect 6 146 58 148
rect 66 140 78 146
rect 49 132 78 140
rect 23 103 37 117
rect 3 83 17 97
rect 49 97 57 132
rect 43 83 57 97
rect 63 103 77 117
rect 83 83 97 97
rect 43 54 51 83
rect 10 8 22 14
rect 67 8 79 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m1p >>
rect 23 103 37 117
rect 63 103 77 117
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal1 43 83 57 97 0 Y
port 4 nsew signal output
rlabel metal1 83 83 97 97 0 C
port 2 nsew signal input
rlabel metal1 23 103 37 117 0 B
port 1 nsew signal input
rlabel metal1 63 103 77 117 0 D
port 3 nsew signal input
rlabel metal1 -6 232 126 248 0 vdd
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 120 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
