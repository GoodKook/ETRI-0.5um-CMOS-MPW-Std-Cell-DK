magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect 46 142 134 181
rect 46 139 154 142
rect -14 61 154 139
rect -14 58 74 61
<< nwell >>
rect -12 154 153 272
<< ntransistor >>
rect 22 14 26 54
rect 42 14 46 34
rect 54 14 58 34
rect 82 14 86 34
rect 92 14 96 34
rect 114 14 118 54
<< ptransistor >>
rect 22 166 26 246
rect 44 206 48 246
rect 54 206 58 246
rect 82 226 86 246
rect 92 226 96 246
rect 114 166 118 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 28 54
rect 40 14 42 34
rect 46 14 54 34
rect 58 14 64 34
rect 76 14 82 34
rect 86 14 92 34
rect 96 14 100 34
rect 112 14 114 54
rect 118 14 120 54
<< pdiffusion >>
rect 20 166 22 246
rect 26 166 28 246
rect 40 206 44 246
rect 48 206 54 246
rect 58 206 62 246
rect 75 226 82 246
rect 86 226 92 246
rect 96 226 100 246
rect 112 166 114 246
rect 118 166 120 246
<< ndcontact >>
rect 8 14 20 54
rect 28 14 40 54
rect 64 14 76 34
rect 100 14 112 54
rect 120 14 132 54
<< pdcontact >>
rect 8 166 20 246
rect 28 166 40 246
rect 62 206 75 246
rect 100 166 112 246
rect 120 166 132 246
<< psubstratepcontact >>
rect -6 -6 146 6
<< nsubstratencontact >>
rect -6 254 146 266
<< polysilicon >>
rect 22 246 26 250
rect 44 246 48 250
rect 54 246 58 250
rect 82 246 86 250
rect 92 246 96 250
rect 114 246 118 250
rect 22 83 26 166
rect 44 160 48 206
rect 42 148 48 160
rect 42 129 46 148
rect 22 54 26 71
rect 42 34 46 117
rect 54 142 58 206
rect 82 191 86 226
rect 74 187 86 191
rect 54 79 58 130
rect 74 99 78 187
rect 92 115 96 226
rect 114 160 118 166
rect 116 148 118 160
rect 54 74 86 79
rect 54 54 57 66
rect 54 34 58 54
rect 82 34 86 74
rect 92 34 96 103
rect 114 54 118 148
rect 22 10 26 14
rect 42 10 46 14
rect 54 10 58 14
rect 82 10 86 14
rect 92 10 96 14
rect 114 10 118 14
<< polycontact >>
rect 34 117 46 129
rect 22 71 34 83
rect 54 130 66 142
rect 66 87 78 99
rect 104 148 116 160
rect 92 103 104 115
rect 57 54 69 66
<< metal1 >>
rect -6 266 146 268
rect -6 252 146 254
rect 28 246 40 252
rect 100 246 112 252
rect 8 142 16 166
rect 78 152 104 160
rect 8 136 54 142
rect 8 54 16 136
rect 78 125 83 139
rect 78 123 86 125
rect 46 117 86 123
rect 124 116 132 166
rect 118 102 132 116
rect 36 87 66 97
rect 57 66 64 87
rect 124 54 132 102
rect 62 14 64 34
rect 28 8 40 14
rect 100 8 112 14
rect -6 6 146 8
rect -6 -8 146 -6
<< m2contact >>
rect 64 192 78 206
rect 64 152 78 166
rect 83 125 97 139
rect 104 103 118 117
rect 22 83 36 97
rect 64 34 78 48
<< metal2 >>
rect 64 166 72 192
rect 26 97 34 114
rect 64 48 72 152
rect 86 139 94 154
rect 106 86 114 103
<< m1p >>
rect -6 252 146 268
rect -6 -8 146 8
<< m2p >>
rect 86 141 94 154
rect 26 99 34 114
rect 106 86 114 101
<< labels >>
rlabel metal2 90 152 90 152 1 D
port 1 n signal input
rlabel metal2 30 111 30 111 1 CLK
port 2 n signal input
rlabel metal2 110 89 110 89 3 Q
port 3 n signal output
rlabel metal1 -6 252 146 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 146 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
