* NGSPICE file created from AOI21X1.ext - technology: scmos

.subckt AOI21X1 A B C Y vdd gnd
M1000 Y C a_4_108# vdd pfet w=12u l=0.6u
+  ad=18p pd=27.000002u as=10.8p ps=13.8u
M1001 a_24_12# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=9p ps=15.000001u
M1002 a_4_108# B vdd vdd pfet w=12u l=0.6u
+  ad=10.8p pd=13.8u as=10.8p ps=13.8u
M1003 gnd C Y gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=4.95p ps=7.8u
M1004 Y B a_24_12# gnd nfet w=6u l=0.6u
+  ad=4.95p pd=7.8u as=2.7p ps=6.9u
M1005 vdd A a_4_108# vdd pfet w=12u l=0.6u
+  ad=10.8p pd=13.8u as=18p ps=27.000002u
.ends

