magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -7 71 57 79
rect -17 30 67 71
<< nwell >>
rect -6 77 56 136
<< ntransistor >>
rect 9 7 11 27
rect 19 7 21 27
rect 29 7 31 27
rect 39 7 41 27
<< ptransistor >>
rect 9 83 11 123
rect 14 83 16 123
rect 29 83 31 123
rect 34 83 36 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 22 19 27
rect 11 7 12 22
rect 18 7 19 22
rect 21 7 22 27
rect 28 7 29 27
rect 31 13 32 27
rect 38 13 39 27
rect 31 7 39 13
rect 41 7 42 27
<< pdiffusion >>
rect 8 83 9 123
rect 11 83 14 123
rect 16 83 17 123
rect 28 83 29 123
rect 31 83 34 123
rect 36 83 37 123
<< ndcontact >>
rect 2 7 8 27
rect 12 7 18 22
rect 22 7 28 27
rect 32 13 38 27
rect 42 7 48 27
<< pdcontact >>
rect 2 83 8 123
rect 17 83 28 123
rect 37 83 43 123
<< psubstratepcontact >>
rect -3 -3 53 3
<< nsubstratencontact >>
rect -3 127 53 133
<< polysilicon >>
rect 9 123 11 125
rect 14 123 16 125
rect 29 123 31 125
rect 34 123 36 125
rect 9 82 11 83
rect 5 80 11 82
rect 14 82 16 83
rect 14 80 21 82
rect 5 64 8 80
rect 5 41 8 58
rect 19 51 21 80
rect 18 45 21 51
rect 5 38 11 41
rect 9 27 11 38
rect 19 27 21 45
rect 29 27 31 83
rect 34 82 36 83
rect 34 80 43 82
rect 41 64 43 80
rect 41 41 43 58
rect 39 38 43 41
rect 39 27 41 38
rect 9 5 11 7
rect 19 5 21 7
rect 29 5 31 7
rect 39 5 41 7
<< polycontact >>
rect 2 58 8 64
rect 12 45 18 51
rect 41 58 47 64
rect 31 45 37 51
<< metal1 >>
rect -3 133 53 134
rect -3 126 53 127
rect 2 123 8 126
rect 37 123 43 126
rect 21 58 25 83
rect 21 36 25 51
rect 21 32 36 36
rect 2 27 28 28
rect 33 27 36 32
rect 8 25 22 27
rect 28 7 42 10
rect 12 4 18 7
rect -3 3 53 4
rect -3 -4 53 -3
<< m2contact >>
rect 1 51 8 58
rect 11 51 18 58
rect 21 51 28 58
rect 31 51 38 58
rect 41 51 48 58
<< metal2 >>
rect 13 58 17 67
rect 33 58 37 67
rect 3 43 7 51
rect 23 43 27 51
rect 43 43 47 51
<< m1p >>
rect -3 126 53 134
rect -3 -4 53 4
<< m2p >>
rect 13 59 17 67
rect 33 59 37 67
rect 3 43 7 50
rect 23 43 27 50
rect 43 43 47 50
<< labels >>
rlabel metal2 5 45 5 45 1 A
port 1 n signal input
rlabel metal2 15 65 15 65 1 B
port 2 n signal input
rlabel metal2 45 45 45 45 1 C
port 3 n signal input
rlabel metal2 35 65 35 65 1 D
port 4 n signal input
rlabel metal2 25 44 25 44 5 Y
port 5 n signal output
rlabel metal1 -3 126 53 134 0 vdd
port 6 nsew power bidirectional abutment
rlabel metal1 -3 -4 53 4 0 gnd
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 50 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
