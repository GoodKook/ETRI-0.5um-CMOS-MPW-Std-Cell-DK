magic
tech scmos
magscale 1 2
timestamp 1728305200
<< nwell >>
rect -12 134 132 252
<< ntransistor >>
rect 21 14 25 54
rect 41 14 45 54
rect 61 14 65 54
rect 81 14 85 54
<< ptransistor >>
rect 21 146 25 226
rect 31 146 35 226
rect 61 146 65 226
rect 71 146 75 226
<< ndiffusion >>
rect 19 14 21 54
rect 25 44 41 54
rect 25 14 27 44
rect 39 14 41 44
rect 45 14 47 54
rect 59 14 61 54
rect 65 26 67 54
rect 79 26 81 54
rect 65 14 81 26
rect 85 14 87 54
<< pdiffusion >>
rect 19 146 21 226
rect 25 146 31 226
rect 35 146 37 226
rect 59 146 61 226
rect 65 146 71 226
rect 75 146 77 226
<< ndcontact >>
rect 7 14 19 54
rect 27 14 39 44
rect 47 14 59 54
rect 67 26 79 54
rect 87 14 99 54
<< pdcontact >>
rect 7 146 19 226
rect 37 146 59 226
rect 77 146 89 226
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 234 126 246
<< polysilicon >>
rect 21 226 25 230
rect 31 226 35 230
rect 61 226 65 230
rect 71 226 75 230
rect 21 142 25 146
rect 11 138 25 142
rect 31 142 35 146
rect 31 138 45 142
rect 11 123 16 138
rect 10 65 16 111
rect 39 89 45 138
rect 61 89 65 146
rect 71 142 75 146
rect 71 138 85 142
rect 81 123 85 138
rect 81 111 83 123
rect 36 77 45 89
rect 10 61 25 65
rect 21 54 25 61
rect 41 54 45 77
rect 61 54 65 77
rect 81 54 85 111
rect 21 10 25 14
rect 41 10 45 14
rect 61 10 65 14
rect 81 10 85 14
<< polycontact >>
rect 4 111 16 123
rect 83 111 95 123
rect 24 77 36 89
rect 60 77 72 89
<< metal1 >>
rect -6 246 126 248
rect -6 232 126 234
rect 7 226 19 232
rect 77 226 89 232
rect 47 111 55 146
rect 46 71 54 97
rect 46 64 75 71
rect 7 54 59 56
rect 69 54 75 64
rect 19 50 47 54
rect 59 14 87 20
rect 27 8 39 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 97 17 111
rect 23 89 37 103
rect 43 97 57 111
rect 63 89 77 103
rect 83 97 97 111
<< metal2 >>
rect 3 83 17 97
rect 23 103 37 117
rect 43 83 57 97
rect 63 103 77 117
rect 83 83 97 97
<< m1p >>
rect -6 232 126 248
rect -6 -8 126 8
<< m2p >>
rect 23 103 37 117
rect 63 103 77 117
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 -6 232 126 248 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 23 103 37 117 0 B
port 1 nsew signal input
rlabel metal2 83 83 97 97 0 C
port 2 nsew signal input
rlabel metal2 43 83 57 97 0 Y
port 4 nsew signal output
rlabel metal2 63 103 77 117 0 D
port 3 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
