magic
tech scmos
magscale 1 2
timestamp 1727490190
<< nwell >>
rect -6 154 206 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
rect 100 14 104 54
rect 120 14 124 54
rect 140 14 144 54
rect 160 14 164 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
rect 100 166 104 246
rect 120 166 124 246
rect 140 166 144 246
rect 160 166 164 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
rect 78 14 80 54
rect 84 14 86 54
rect 98 14 100 54
rect 104 14 106 54
rect 118 14 120 54
rect 124 14 126 54
rect 138 14 140 54
rect 144 14 146 54
rect 158 14 160 54
rect 164 14 166 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 26 246
rect 38 166 40 246
rect 44 166 46 246
rect 58 166 60 246
rect 64 166 66 246
rect 78 166 80 246
rect 84 166 86 246
rect 98 166 100 246
rect 104 166 106 246
rect 118 166 120 246
rect 124 166 126 246
rect 138 166 140 246
rect 144 166 146 246
rect 158 166 160 246
rect 164 166 166 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
rect 86 14 98 54
rect 106 14 118 54
rect 126 14 138 54
rect 146 14 158 54
rect 166 14 178 54
<< pdcontact >>
rect 6 166 18 246
rect 26 166 38 246
rect 46 166 58 246
rect 66 166 78 246
rect 86 166 98 246
rect 106 166 118 246
rect 126 166 138 246
rect 146 166 158 246
rect 166 166 178 246
<< psubstratepcontact >>
rect 0 -6 200 6
<< nsubstratencontact >>
rect 0 254 200 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 100 246 104 250
rect 120 246 124 250
rect 140 246 144 250
rect 160 246 164 250
rect 20 54 24 166
rect 40 103 44 166
rect 36 91 44 103
rect 40 54 44 91
rect 60 86 64 166
rect 80 86 84 166
rect 72 74 84 86
rect 60 54 64 74
rect 80 54 84 74
rect 100 86 104 166
rect 120 86 124 166
rect 112 74 124 86
rect 100 54 104 74
rect 120 54 124 74
rect 140 86 144 166
rect 160 86 164 166
rect 152 74 164 86
rect 140 54 144 74
rect 160 54 164 74
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
rect 100 10 104 14
rect 120 10 124 14
rect 140 10 144 14
rect 160 10 164 14
<< polycontact >>
rect 24 91 36 103
rect 60 74 72 86
rect 100 74 112 86
rect 140 74 152 86
<< metal1 >>
rect 0 266 200 268
rect 0 252 200 254
rect 6 246 18 252
rect 46 246 58 252
rect 86 246 98 252
rect 126 246 138 252
rect 166 246 178 252
rect 26 160 38 166
rect 66 160 78 166
rect 106 160 118 166
rect 146 160 158 166
rect 26 152 52 160
rect 66 152 92 160
rect 106 152 132 160
rect 146 152 164 160
rect 44 82 52 152
rect 44 74 60 82
rect 84 82 92 152
rect 84 74 100 82
rect 124 82 132 152
rect 158 117 164 152
rect 158 103 163 117
rect 124 74 140 82
rect 44 68 52 74
rect 84 68 92 74
rect 124 68 132 74
rect 158 68 164 103
rect 26 60 52 68
rect 66 60 92 68
rect 106 60 132 68
rect 146 60 164 68
rect 26 54 38 60
rect 66 54 78 60
rect 106 54 118 60
rect 146 54 158 60
rect 6 8 18 14
rect 46 8 58 14
rect 86 8 98 14
rect 126 8 138 14
rect 166 8 178 14
rect 0 6 200 8
rect 0 -8 200 -6
<< m2contact >>
rect 23 103 37 117
rect 163 103 177 117
<< metal2 >>
rect 23 117 37 137
rect 163 117 177 137
<< m2p >>
rect 23 123 37 137
rect 163 123 177 137
<< labels >>
rlabel metal2 23 123 37 137 0 A
port 0 nsew signal input
rlabel metal2 163 123 177 137 0 Y
port 1 nsew signal output
rlabel metal1 0 266 200 268 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal1 0 254 200 266 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal1 0 252 200 254 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal1 0 6 200 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 0 -6 200 6 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 0 -8 200 -6 0 gnd
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 200 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
