magic
tech scmos
magscale 1 2
timestamp 1727908812
<< nwell >>
rect -12 134 112 252
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
<< ptransistor >>
rect 26 146 30 226
rect 34 146 38 226
rect 56 186 60 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 24 146 26 226
rect 30 146 34 226
rect 38 146 40 226
rect 52 186 56 226
rect 60 186 62 226
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
<< pdcontact >>
rect 12 146 24 226
rect 40 146 52 226
rect 62 186 74 226
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 234 106 246
<< polysilicon >>
rect 26 226 30 230
rect 34 226 38 230
rect 56 226 60 230
rect 26 142 30 146
rect 12 134 30 142
rect 12 109 16 134
rect 34 103 38 146
rect 56 142 60 186
rect 56 134 66 142
rect 60 103 66 134
rect 12 66 16 97
rect 36 91 44 103
rect 12 59 24 66
rect 20 54 24 59
rect 40 54 44 91
rect 60 54 64 103
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 4 97 16 109
rect 24 91 36 103
rect 64 91 76 103
<< metal1 >>
rect -6 246 106 248
rect -6 232 106 234
rect 12 226 24 232
rect 62 226 74 232
rect 23 103 37 117
rect 3 83 17 97
rect 44 97 52 146
rect 63 103 77 117
rect 43 85 57 97
rect 43 77 74 85
rect 10 60 54 68
rect 10 54 18 60
rect 46 54 54 60
rect 66 54 74 77
rect 26 8 38 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 23 103 37 117
rect 63 103 77 117
rect 3 83 17 97
rect 43 83 57 97
<< labels >>
rlabel metal1 -6 -8 106 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal1 43 83 57 97 0 Y
port 3 nsew signal output
rlabel metal1 23 103 37 117 0 B
port 1 nsew signal input
rlabel metal1 63 103 77 117 0 C
port 2 nsew signal input
rlabel metal1 -6 232 106 248 0 vdd
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
