magic
tech scmos
magscale 1 2
timestamp 1700713733
<< checkpaint >>
rect -24 308 79 321
rect -30 306 79 308
rect -46 214 79 306
rect -30 212 79 214
rect -24 114 79 212
rect -30 46 66 48
rect -46 -46 66 46
rect -30 -48 66 -46
<< nwell >>
rect -12 154 22 272
<< psubstratepcontact >>
rect -6 -6 16 6
<< nsubstratencontact >>
rect -6 254 16 266
<< metal1 >>
rect -6 266 16 268
rect -6 252 16 254
rect -6 6 16 8
rect -6 -8 16 -6
<< m1p >>
rect -6 252 16 268
rect -6 -8 16 8
<< labels >>
rlabel metal1 1 267 1 267 0 vdd
port 3 nsew
rlabel metal1 2 -7 2 -7 0 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 10 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
