magic
tech scmos
magscale 1 6
timestamp 1569139307
<< checkpaint >>
rect -140 -1950 2540 5180
<< metal2 >>
rect 522 5032 586 5060
use DOUBLE_GUARD  DOUBLE_GUARD_0
timestamp 1569139307
transform 1 0 0 0 1 1660
box -20 -20 2419 500
use INV24  INV24_0
timestamp 1569139307
transform 1 0 296 0 1 4220
box 0 -88 1488 840
use METAL_RING  METAL_RING_0
timestamp 1569139307
transform 1 0 0 0 1 0
box 0 0 2400 5012
use NDRV  NDRV_0
timestamp 1569139307
transform 1 0 0 0 1 0
box 0 0 2400 1560
use PAD_80  PAD_80_0
timestamp 1569139307
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_POB24  PAD_METAL_POB24_0
timestamp 1569139307
transform 1 0 0 0 1 0
box 0 0 2400 4200
use PDRV  PDRV_0
timestamp 1569139307
transform 1 0 0 0 1 2260
box -20 -20 2420 1580
use SINGLE_GUARD  SINGLE_GUARD_0
timestamp 1569139307
transform 1 0 0 0 1 3920
box 0 0 2400 200
<< labels >>
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 PAD
flabel m3p s 0 3018 0 3018 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4339 0 4339 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4788 0 4788 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 752 0 752 0 FreeSans 1000 0 0 0 VSS
flabel m2p s 557 5060 557 5060 0 FreeSans 400 0 0 0 A
<< end >>
