magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -50 -50 300 300
<< psubstratepdiff >>
rect 10 220 240 240
rect 10 30 30 220
rect 220 30 240 220
rect 10 10 240 30
<< metal1 >>
rect 10 220 240 240
rect 10 30 30 220
rect 220 30 240 220
rect 10 10 240 30
use ptap_CDNS_7230122529122  ptap_CDNS_7230122529122_0
timestamp 1723012252
transform 1 0 216 0 1 26
box 4 4 24 194
use ptap_CDNS_7230122529122  ptap_CDNS_7230122529122_1
timestamp 1723012252
transform 0 1 26 1 0 216
box 4 4 24 194
use ptap_CDNS_7230122529122  ptap_CDNS_7230122529122_2
timestamp 1723012252
transform 0 1 26 1 0 6
box 4 4 24 194
use ptap_CDNS_7230122529122  ptap_CDNS_7230122529122_3
timestamp 1723012252
transform 1 0 6 0 1 26
box 4 4 24 194
<< end >>
