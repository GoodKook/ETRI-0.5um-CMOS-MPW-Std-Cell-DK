magic
tech scmos
magscale 1 2
timestamp 1702306673
<< nwell >>
rect -12 154 72 272
<< ntransistor >>
rect 21 14 25 54
rect 31 14 35 54
<< ptransistor >>
rect 18 206 22 246
rect 38 206 42 246
<< ndiffusion >>
rect 19 14 21 54
rect 25 14 31 54
rect 35 14 41 54
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 206 38 246
rect 42 206 44 246
<< ndcontact >>
rect 7 14 19 54
rect 41 14 53 54
<< pdcontact >>
rect 4 206 16 246
rect 24 206 36 246
rect 44 206 56 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 18 117 22 206
rect 17 105 22 117
rect 18 80 22 105
rect 38 117 42 206
rect 38 105 43 117
rect 38 80 42 105
rect 18 75 25 80
rect 21 54 25 75
rect 31 75 42 80
rect 31 54 35 75
rect 21 10 25 14
rect 31 10 35 14
<< polycontact >>
rect 5 105 17 117
rect 43 105 55 117
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 4 246 16 252
rect 44 246 56 252
rect 3 123 17 137
rect 5 117 17 123
rect 26 117 34 206
rect 43 123 57 137
rect 43 117 55 123
rect 23 103 37 117
rect 26 60 34 103
rect 26 54 53 60
rect 7 8 15 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m1p >>
rect -6 252 66 268
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect -6 -8 66 8
<< labels >>
rlabel nsubstratencontact 30 260 30 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 30 0 30 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 50 127 50 127 0 B
port 2 nsew signal input
rlabel metal1 30 110 30 110 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
