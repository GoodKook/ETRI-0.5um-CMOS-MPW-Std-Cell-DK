magic
tech scmos
magscale 1 3
timestamp 1537935238
<< checkpaint >>
rect -70 -70 1270 850
<< nwell >>
rect -10 -10 1210 790
<< nsubstratendiff >>
rect 0 730 1200 780
rect 0 50 50 730
rect 1150 50 1200 730
rect 0 0 1200 50
<< metal1 >>
rect 0 730 1200 780
rect 0 50 50 730
rect 1150 50 1200 730
rect 0 0 1200 50
<< metal2 >>
rect 0 0 40 780
rect 1150 0 1200 780
<< metal3 >>
rect 0 0 50 780
rect 1150 0 1200 780
<< filln >>
rect 56 56 1144 724
use CONT  CONT_0
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 1175 0 1 12
box -3 -3 3 3
use CONT  CONT_1
array 0 90 12 0 2 12
timestamp 1537935238
transform 1 0 59 0 1 743
box -3 -3 3 3
use CONT  CONT_2
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 25 0 1 12
box -3 -3 3 3
use CONT  CONT_3
array 0 90 12 0 2 12
timestamp 1537935238
transform 1 0 59 0 1 13
box -3 -3 3 3
use PLEAF  PLEAF_0
array 0 7 126 0 0 0
timestamp 1537935238
transform 1 0 83 0 1 90
box -13 -10 165 628
use VIA1  VIA1_0
array 0 1 30 0 42 18
timestamp 1537935238
transform 1 0 1160 0 1 12
box -4 -4 4 4
use VIA1  VIA1_1
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 10 0 1 12
box -4 -4 4 4
use VIA2  VIA2_0
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 1175 0 1 12
box -4 -4 4 4
use VIA2  VIA2_1
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 25 0 1 12
box -4 -4 4 4
<< end >>
