// 256 bytes read from wozmon.bin
// Offset address: FF00
	16'hFF00: 8'hD8;
	16'hFF01: 8'h58;
	16'hFF02: 8'hA0;
	16'hFF03: 8'h7F;
	16'hFF04: 8'h8C;
	16'hFF05: 8'h12;
	16'hFF06: 8'hD0;
	16'hFF07: 8'hA9;
	16'hFF08: 8'hA7;
	16'hFF09: 8'h8D;
	16'hFF0A: 8'h11;
	16'hFF0B: 8'hD0;
	16'hFF0C: 8'h8D;
	16'hFF0D: 8'h13;
	16'hFF0E: 8'hD0;
	16'hFF0F: 8'hC9;
	16'hFF10: 8'hDF;
	16'hFF11: 8'hF0;
	16'hFF12: 8'h13;
	16'hFF13: 8'hC9;
	16'hFF14: 8'h9B;
	16'hFF15: 8'hF0;
	16'hFF16: 8'h03;
	16'hFF17: 8'hC8;
	16'hFF18: 8'h10;
	16'hFF19: 8'h0F;
	16'hFF1A: 8'hA9;
	16'hFF1B: 8'hDC;
	16'hFF1C: 8'h20;
	16'hFF1D: 8'hEF;
	16'hFF1E: 8'hFF;
	16'hFF1F: 8'hA9;
	16'hFF20: 8'h8D;
	16'hFF21: 8'h20;
	16'hFF22: 8'hEF;
	16'hFF23: 8'hFF;
	16'hFF24: 8'hA0;
	16'hFF25: 8'h01;
	16'hFF26: 8'h88;
	16'hFF27: 8'h30;
	16'hFF28: 8'hF6;
	16'hFF29: 8'hAD;
	16'hFF2A: 8'h11;
	16'hFF2B: 8'hD0;
	16'hFF2C: 8'h10;
	16'hFF2D: 8'hFB;
	16'hFF2E: 8'hAD;
	16'hFF2F: 8'h10;
	16'hFF30: 8'hD0;
	16'hFF31: 8'h99;
	16'hFF32: 8'h00;
	16'hFF33: 8'h02;
	16'hFF34: 8'h20;
	16'hFF35: 8'hEF;
	16'hFF36: 8'hFF;
	16'hFF37: 8'hC9;
	16'hFF38: 8'h8D;
	16'hFF39: 8'hD0;
	16'hFF3A: 8'hD4;
	16'hFF3B: 8'hA0;
	16'hFF3C: 8'hFF;
	16'hFF3D: 8'hA9;
	16'hFF3E: 8'h00;
	16'hFF3F: 8'hAA;
	16'hFF40: 8'h0A;
	16'hFF41: 8'h85;
	16'hFF42: 8'h2B;
	16'hFF43: 8'hC8;
	16'hFF44: 8'hB9;
	16'hFF45: 8'h00;
	16'hFF46: 8'h02;
	16'hFF47: 8'hC9;
	16'hFF48: 8'h8D;
	16'hFF49: 8'hF0;
	16'hFF4A: 8'hD4;
	16'hFF4B: 8'hC9;
	16'hFF4C: 8'hAE;
	16'hFF4D: 8'h90;
	16'hFF4E: 8'hF4;
	16'hFF4F: 8'hF0;
	16'hFF50: 8'hF0;
	16'hFF51: 8'hC9;
	16'hFF52: 8'hBA;
	16'hFF53: 8'hF0;
	16'hFF54: 8'hEB;
	16'hFF55: 8'hC9;
	16'hFF56: 8'hD2;
	16'hFF57: 8'hF0;
	16'hFF58: 8'h3B;
	16'hFF59: 8'h86;
	16'hFF5A: 8'h28;
	16'hFF5B: 8'h86;
	16'hFF5C: 8'h29;
	16'hFF5D: 8'h84;
	16'hFF5E: 8'h2A;
	16'hFF5F: 8'hB9;
	16'hFF60: 8'h00;
	16'hFF61: 8'h02;
	16'hFF62: 8'h49;
	16'hFF63: 8'hB0;
	16'hFF64: 8'hC9;
	16'hFF65: 8'h0A;
	16'hFF66: 8'h90;
	16'hFF67: 8'h06;
	16'hFF68: 8'h69;
	16'hFF69: 8'h88;
	16'hFF6A: 8'hC9;
	16'hFF6B: 8'hFA;
	16'hFF6C: 8'h90;
	16'hFF6D: 8'h11;
	16'hFF6E: 8'h0A;
	16'hFF6F: 8'h0A;
	16'hFF70: 8'h0A;
	16'hFF71: 8'h0A;
	16'hFF72: 8'hA2;
	16'hFF73: 8'h04;
	16'hFF74: 8'h0A;
	16'hFF75: 8'h26;
	16'hFF76: 8'h28;
	16'hFF77: 8'h26;
	16'hFF78: 8'h29;
	16'hFF79: 8'hCA;
	16'hFF7A: 8'hD0;
	16'hFF7B: 8'hF8;
	16'hFF7C: 8'hC8;
	16'hFF7D: 8'hD0;
	16'hFF7E: 8'hE0;
	16'hFF7F: 8'hC4;
	16'hFF80: 8'h2A;
	16'hFF81: 8'hF0;
	16'hFF82: 8'h97;
	16'hFF83: 8'h24;
	16'hFF84: 8'h2B;
	16'hFF85: 8'h50;
	16'hFF86: 8'h10;
	16'hFF87: 8'hA5;
	16'hFF88: 8'h28;
	16'hFF89: 8'h81;
	16'hFF8A: 8'h26;
	16'hFF8B: 8'hE6;
	16'hFF8C: 8'h26;
	16'hFF8D: 8'hD0;
	16'hFF8E: 8'hB5;
	16'hFF8F: 8'hE6;
	16'hFF90: 8'h27;
	16'hFF91: 8'h4C;
	16'hFF92: 8'h44;
	16'hFF93: 8'hFF;
	16'hFF94: 8'h6C;
	16'hFF95: 8'h24;
	16'hFF96: 8'h00;
	16'hFF97: 8'h30;
	16'hFF98: 8'h2B;
	16'hFF99: 8'hA2;
	16'hFF9A: 8'h02;
	16'hFF9B: 8'hB5;
	16'hFF9C: 8'h27;
	16'hFF9D: 8'h95;
	16'hFF9E: 8'h25;
	16'hFF9F: 8'h95;
	16'hFFA0: 8'h23;
	16'hFFA1: 8'hCA;
	16'hFFA2: 8'hD0;
	16'hFFA3: 8'hF7;
	16'hFFA4: 8'hD0;
	16'hFFA5: 8'h14;
	16'hFFA6: 8'hA9;
	16'hFFA7: 8'h8D;
	16'hFFA8: 8'h20;
	16'hFFA9: 8'hEF;
	16'hFFAA: 8'hFF;
	16'hFFAB: 8'hA5;
	16'hFFAC: 8'h25;
	16'hFFAD: 8'h20;
	16'hFFAE: 8'hDC;
	16'hFFAF: 8'hFF;
	16'hFFB0: 8'hA5;
	16'hFFB1: 8'h24;
	16'hFFB2: 8'h20;
	16'hFFB3: 8'hDC;
	16'hFFB4: 8'hFF;
	16'hFFB5: 8'hA9;
	16'hFFB6: 8'hBA;
	16'hFFB7: 8'h20;
	16'hFFB8: 8'hEF;
	16'hFFB9: 8'hFF;
	16'hFFBA: 8'hA9;
	16'hFFBB: 8'hA0;
	16'hFFBC: 8'h20;
	16'hFFBD: 8'hEF;
	16'hFFBE: 8'hFF;
	16'hFFBF: 8'hA1;
	16'hFFC0: 8'h24;
	16'hFFC1: 8'h20;
	16'hFFC2: 8'hDC;
	16'hFFC3: 8'hFF;
	16'hFFC4: 8'h86;
	16'hFFC5: 8'h2B;
	16'hFFC6: 8'hA5;
	16'hFFC7: 8'h24;
	16'hFFC8: 8'hC5;
	16'hFFC9: 8'h28;
	16'hFFCA: 8'hA5;
	16'hFFCB: 8'h25;
	16'hFFCC: 8'hE5;
	16'hFFCD: 8'h29;
	16'hFFCE: 8'hB0;
	16'hFFCF: 8'hC1;
	16'hFFD0: 8'hE6;
	16'hFFD1: 8'h24;
	16'hFFD2: 8'hD0;
	16'hFFD3: 8'h02;
	16'hFFD4: 8'hE6;
	16'hFFD5: 8'h25;
	16'hFFD6: 8'hA5;
	16'hFFD7: 8'h24;
	16'hFFD8: 8'h29;
	16'hFFD9: 8'h07;
	16'hFFDA: 8'h10;
	16'hFFDB: 8'hC8;
	16'hFFDC: 8'h48;
	16'hFFDD: 8'h4A;
	16'hFFDE: 8'h4A;
	16'hFFDF: 8'h4A;
	16'hFFE0: 8'h4A;
	16'hFFE1: 8'h20;
	16'hFFE2: 8'hE5;
	16'hFFE3: 8'hFF;
	16'hFFE4: 8'h68;
	16'hFFE5: 8'h29;
	16'hFFE6: 8'h0F;
	16'hFFE7: 8'h09;
	16'hFFE8: 8'hB0;
	16'hFFE9: 8'hC9;
	16'hFFEA: 8'hBA;
	16'hFFEB: 8'h90;
	16'hFFEC: 8'h02;
	16'hFFED: 8'h69;
	16'hFFEE: 8'h06;
	16'hFFEF: 8'h2C;
	16'hFFF0: 8'h12;
	16'hFFF1: 8'hD0;
	16'hFFF2: 8'h30;
	16'hFFF3: 8'hFB;
	16'hFFF4: 8'h8D;
	16'hFFF5: 8'h12;
	16'hFFF6: 8'hD0;
	16'hFFF7: 8'h60;
	16'hFFF8: 8'h00;
	16'hFFF9: 8'h00;
	16'hFFFA: 8'h00;
	16'hFFFB: 8'h0F;
	16'hFFFC: 8'h00;
	16'hFFFD: 8'hFF;
	16'hFFFE: 8'h00;
	16'hFFFF: 8'h00;
