magic
tech scmos
magscale 1 3
timestamp 1537935238
<< checkpaint >>
rect -60 -60 1008 840
<< psubstratepdiff >>
rect 0 730 948 780
rect 0 50 50 730
rect 898 50 948 730
rect 0 0 948 50
<< metal1 >>
rect 0 730 948 780
rect 0 50 50 730
rect 898 50 948 730
rect 0 0 948 50
<< metal2 >>
rect 0 0 50 780
rect 898 0 948 780
<< filln >>
rect 56 56 892 724
use CONT  CONT_0
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 923 0 1 12
box -3 -3 3 3
use CONT  CONT_1
array 0 45 18 0 1 18
timestamp 1537935238
transform 1 0 59 0 1 746
box -3 -3 3 3
use CONT  CONT_2
array 0 0 0 0 42 18
timestamp 1537935238
transform 1 0 25 0 1 12
box -3 -3 3 3
use CONT  CONT_3
array 0 45 18 0 1 18
timestamp 1537935238
transform 1 0 59 0 1 16
box -3 -3 3 3
use NLEAF1  NLEAF1_0
array 0 5 126 0 0 0
timestamp 1537935238
transform 1 0 83 0 1 90
box -13 -10 165 628
use VIA1  VIA1_0
array 0 1 30 0 36 18
timestamp 1537935238
transform 1 0 908 0 1 66
box -4 -4 4 4
use VIA1  VIA1_1
array 0 1 30 0 36 18
timestamp 1537935238
transform 1 0 10 0 1 66
box -4 -4 4 4
<< end >>
