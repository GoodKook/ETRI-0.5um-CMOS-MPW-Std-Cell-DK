magic
tech scmos
magscale 1 6
timestamp 1569139307
<< checkpaint >>
rect -120 -120 2520 320
<< psubstratepdiff >>
rect 0 0 2400 200
<< metal1 >>
rect 0 0 2400 200
use CONT  CONT_0
timestamp 1569139307
transform 1 0 164 0 1 63
box -6 -6 6 6
use CONT  CONT_1
timestamp 1569139307
transform 1 0 128 0 1 63
box -6 -6 6 6
use CONT  CONT_2
timestamp 1569139307
transform 1 0 92 0 1 63
box -6 -6 6 6
use CONT  CONT_3
timestamp 1569139307
transform 1 0 236 0 1 27
box -6 -6 6 6
use CONT  CONT_4
timestamp 1569139307
transform 1 0 200 0 1 27
box -6 -6 6 6
use CONT  CONT_5
timestamp 1569139307
transform 1 0 164 0 1 27
box -6 -6 6 6
use CONT  CONT_6
timestamp 1569139307
transform 1 0 524 0 1 63
box -6 -6 6 6
use CONT  CONT_7
timestamp 1569139307
transform 1 0 488 0 1 63
box -6 -6 6 6
use CONT  CONT_8
timestamp 1569139307
transform 1 0 452 0 1 63
box -6 -6 6 6
use CONT  CONT_9
timestamp 1569139307
transform 1 0 416 0 1 63
box -6 -6 6 6
use CONT  CONT_10
timestamp 1569139307
transform 1 0 380 0 1 63
box -6 -6 6 6
use CONT  CONT_11
timestamp 1569139307
transform 1 0 344 0 1 63
box -6 -6 6 6
use CONT  CONT_12
timestamp 1569139307
transform 1 0 308 0 1 63
box -6 -6 6 6
use CONT  CONT_13
timestamp 1569139307
transform 1 0 272 0 1 63
box -6 -6 6 6
use CONT  CONT_14
timestamp 1569139307
transform 1 0 596 0 1 99
box -6 -6 6 6
use CONT  CONT_15
timestamp 1569139307
transform 1 0 560 0 1 99
box -6 -6 6 6
use CONT  CONT_16
timestamp 1569139307
transform 1 0 524 0 1 99
box -6 -6 6 6
use CONT  CONT_17
timestamp 1569139307
transform 1 0 488 0 1 99
box -6 -6 6 6
use CONT  CONT_18
timestamp 1569139307
transform 1 0 452 0 1 99
box -6 -6 6 6
use CONT  CONT_19
timestamp 1569139307
transform 1 0 416 0 1 99
box -6 -6 6 6
use CONT  CONT_20
timestamp 1569139307
transform 1 0 380 0 1 99
box -6 -6 6 6
use CONT  CONT_21
timestamp 1569139307
transform 1 0 344 0 1 99
box -6 -6 6 6
use CONT  CONT_22
timestamp 1569139307
transform 1 0 308 0 1 99
box -6 -6 6 6
use CONT  CONT_23
timestamp 1569139307
transform 1 0 272 0 1 99
box -6 -6 6 6
use CONT  CONT_24
timestamp 1569139307
transform 1 0 236 0 1 99
box -6 -6 6 6
use CONT  CONT_25
timestamp 1569139307
transform 1 0 200 0 1 99
box -6 -6 6 6
use CONT  CONT_26
timestamp 1569139307
transform 1 0 164 0 1 99
box -6 -6 6 6
use CONT  CONT_27
timestamp 1569139307
transform 1 0 128 0 1 99
box -6 -6 6 6
use CONT  CONT_28
timestamp 1569139307
transform 1 0 236 0 1 63
box -6 -6 6 6
use CONT  CONT_29
timestamp 1569139307
transform 1 0 200 0 1 63
box -6 -6 6 6
use CONT  CONT_30
timestamp 1569139307
transform 1 0 596 0 1 63
box -6 -6 6 6
use CONT  CONT_31
timestamp 1569139307
transform 1 0 596 0 1 135
box -6 -6 6 6
use CONT  CONT_32
timestamp 1569139307
transform 1 0 560 0 1 135
box -6 -6 6 6
use CONT  CONT_33
timestamp 1569139307
transform 1 0 524 0 1 135
box -6 -6 6 6
use CONT  CONT_34
timestamp 1569139307
transform 1 0 488 0 1 135
box -6 -6 6 6
use CONT  CONT_35
timestamp 1569139307
transform 1 0 452 0 1 135
box -6 -6 6 6
use CONT  CONT_36
timestamp 1569139307
transform 1 0 416 0 1 135
box -6 -6 6 6
use CONT  CONT_37
timestamp 1569139307
transform 1 0 380 0 1 135
box -6 -6 6 6
use CONT  CONT_38
timestamp 1569139307
transform 1 0 344 0 1 135
box -6 -6 6 6
use CONT  CONT_39
timestamp 1569139307
transform 1 0 596 0 1 171
box -6 -6 6 6
use CONT  CONT_40
timestamp 1569139307
transform 1 0 560 0 1 171
box -6 -6 6 6
use CONT  CONT_41
timestamp 1569139307
transform 1 0 524 0 1 171
box -6 -6 6 6
use CONT  CONT_42
timestamp 1569139307
transform 1 0 488 0 1 171
box -6 -6 6 6
use CONT  CONT_43
timestamp 1569139307
transform 1 0 452 0 1 171
box -6 -6 6 6
use CONT  CONT_44
timestamp 1569139307
transform 1 0 416 0 1 171
box -6 -6 6 6
use CONT  CONT_45
timestamp 1569139307
transform 1 0 380 0 1 171
box -6 -6 6 6
use CONT  CONT_46
timestamp 1569139307
transform 1 0 344 0 1 171
box -6 -6 6 6
use CONT  CONT_47
timestamp 1569139307
transform 1 0 308 0 1 171
box -6 -6 6 6
use CONT  CONT_48
timestamp 1569139307
transform 1 0 272 0 1 171
box -6 -6 6 6
use CONT  CONT_49
timestamp 1569139307
transform 1 0 236 0 1 171
box -6 -6 6 6
use CONT  CONT_50
timestamp 1569139307
transform 1 0 200 0 1 171
box -6 -6 6 6
use CONT  CONT_51
timestamp 1569139307
transform 1 0 164 0 1 171
box -6 -6 6 6
use CONT  CONT_52
timestamp 1569139307
transform 1 0 128 0 1 171
box -6 -6 6 6
use CONT  CONT_53
timestamp 1569139307
transform 1 0 92 0 1 171
box -6 -6 6 6
use CONT  CONT_54
timestamp 1569139307
transform 1 0 56 0 1 171
box -6 -6 6 6
use CONT  CONT_55
timestamp 1569139307
transform 1 0 92 0 1 99
box -6 -6 6 6
use CONT  CONT_56
timestamp 1569139307
transform 1 0 56 0 1 99
box -6 -6 6 6
use CONT  CONT_57
timestamp 1569139307
transform 1 0 56 0 1 63
box -6 -6 6 6
use CONT  CONT_58
timestamp 1569139307
transform 1 0 56 0 1 27
box -6 -6 6 6
use CONT  CONT_59
timestamp 1569139307
transform 1 0 308 0 1 135
box -6 -6 6 6
use CONT  CONT_60
timestamp 1569139307
transform 1 0 272 0 1 135
box -6 -6 6 6
use CONT  CONT_61
timestamp 1569139307
transform 1 0 236 0 1 135
box -6 -6 6 6
use CONT  CONT_62
timestamp 1569139307
transform 1 0 200 0 1 135
box -6 -6 6 6
use CONT  CONT_63
timestamp 1569139307
transform 1 0 164 0 1 135
box -6 -6 6 6
use CONT  CONT_64
timestamp 1569139307
transform 1 0 128 0 1 135
box -6 -6 6 6
use CONT  CONT_65
timestamp 1569139307
transform 1 0 92 0 1 135
box -6 -6 6 6
use CONT  CONT_66
timestamp 1569139307
transform 1 0 56 0 1 135
box -6 -6 6 6
use CONT  CONT_67
timestamp 1569139307
transform 1 0 128 0 1 27
box -6 -6 6 6
use CONT  CONT_68
timestamp 1569139307
transform 1 0 92 0 1 27
box -6 -6 6 6
use CONT  CONT_69
timestamp 1569139307
transform 1 0 560 0 1 63
box -6 -6 6 6
use CONT  CONT_70
timestamp 1569139307
transform 1 0 596 0 1 27
box -6 -6 6 6
use CONT  CONT_71
timestamp 1569139307
transform 1 0 560 0 1 27
box -6 -6 6 6
use CONT  CONT_72
timestamp 1569139307
transform 1 0 524 0 1 27
box -6 -6 6 6
use CONT  CONT_73
timestamp 1569139307
transform 1 0 488 0 1 27
box -6 -6 6 6
use CONT  CONT_74
timestamp 1569139307
transform 1 0 452 0 1 27
box -6 -6 6 6
use CONT  CONT_75
timestamp 1569139307
transform 1 0 416 0 1 27
box -6 -6 6 6
use CONT  CONT_76
timestamp 1569139307
transform 1 0 380 0 1 27
box -6 -6 6 6
use CONT  CONT_77
timestamp 1569139307
transform 1 0 344 0 1 27
box -6 -6 6 6
use CONT  CONT_78
timestamp 1569139307
transform 1 0 308 0 1 27
box -6 -6 6 6
use CONT  CONT_79
timestamp 1569139307
transform 1 0 272 0 1 27
box -6 -6 6 6
use CONT  CONT_80
timestamp 1569139307
transform 1 0 1172 0 1 99
box -6 -6 6 6
use CONT  CONT_81
timestamp 1569139307
transform 1 0 1136 0 1 99
box -6 -6 6 6
use CONT  CONT_82
timestamp 1569139307
transform 1 0 920 0 1 99
box -6 -6 6 6
use CONT  CONT_83
timestamp 1569139307
transform 1 0 884 0 1 99
box -6 -6 6 6
use CONT  CONT_84
timestamp 1569139307
transform 1 0 848 0 1 99
box -6 -6 6 6
use CONT  CONT_85
timestamp 1569139307
transform 1 0 812 0 1 99
box -6 -6 6 6
use CONT  CONT_86
timestamp 1569139307
transform 1 0 776 0 1 99
box -6 -6 6 6
use CONT  CONT_87
timestamp 1569139307
transform 1 0 740 0 1 99
box -6 -6 6 6
use CONT  CONT_88
timestamp 1569139307
transform 1 0 704 0 1 99
box -6 -6 6 6
use CONT  CONT_89
timestamp 1569139307
transform 1 0 668 0 1 99
box -6 -6 6 6
use CONT  CONT_90
timestamp 1569139307
transform 1 0 776 0 1 63
box -6 -6 6 6
use CONT  CONT_91
timestamp 1569139307
transform 1 0 1172 0 1 171
box -6 -6 6 6
use CONT  CONT_92
timestamp 1569139307
transform 1 0 1136 0 1 171
box -6 -6 6 6
use CONT  CONT_93
timestamp 1569139307
transform 1 0 920 0 1 171
box -6 -6 6 6
use CONT  CONT_94
timestamp 1569139307
transform 1 0 884 0 1 171
box -6 -6 6 6
use CONT  CONT_95
timestamp 1569139307
transform 1 0 848 0 1 171
box -6 -6 6 6
use CONT  CONT_96
timestamp 1569139307
transform 1 0 812 0 1 171
box -6 -6 6 6
use CONT  CONT_97
timestamp 1569139307
transform 1 0 776 0 1 171
box -6 -6 6 6
use CONT  CONT_98
timestamp 1569139307
transform 1 0 740 0 1 171
box -6 -6 6 6
use CONT  CONT_99
timestamp 1569139307
transform 1 0 704 0 1 171
box -6 -6 6 6
use CONT  CONT_100
timestamp 1569139307
transform 1 0 668 0 1 171
box -6 -6 6 6
use CONT  CONT_101
timestamp 1569139307
transform 1 0 740 0 1 63
box -6 -6 6 6
use CONT  CONT_102
timestamp 1569139307
transform 1 0 1172 0 1 27
box -6 -6 6 6
use CONT  CONT_103
timestamp 1569139307
transform 1 0 1136 0 1 27
box -6 -6 6 6
use CONT  CONT_104
timestamp 1569139307
transform 1 0 920 0 1 27
box -6 -6 6 6
use CONT  CONT_105
timestamp 1569139307
transform 1 0 884 0 1 27
box -6 -6 6 6
use CONT  CONT_106
timestamp 1569139307
transform 1 0 848 0 1 27
box -6 -6 6 6
use CONT  CONT_107
timestamp 1569139307
transform 1 0 812 0 1 27
box -6 -6 6 6
use CONT  CONT_108
timestamp 1569139307
transform 1 0 776 0 1 27
box -6 -6 6 6
use CONT  CONT_109
timestamp 1569139307
transform 1 0 740 0 1 27
box -6 -6 6 6
use CONT  CONT_110
timestamp 1569139307
transform 1 0 704 0 1 27
box -6 -6 6 6
use CONT  CONT_111
timestamp 1569139307
transform 1 0 668 0 1 27
box -6 -6 6 6
use CONT  CONT_112
timestamp 1569139307
transform 1 0 704 0 1 63
box -6 -6 6 6
use CONT  CONT_113
timestamp 1569139307
transform 1 0 1172 0 1 135
box -6 -6 6 6
use CONT  CONT_114
timestamp 1569139307
transform 1 0 1136 0 1 135
box -6 -6 6 6
use CONT  CONT_115
timestamp 1569139307
transform 1 0 920 0 1 135
box -6 -6 6 6
use CONT  CONT_116
timestamp 1569139307
transform 1 0 884 0 1 135
box -6 -6 6 6
use CONT  CONT_117
timestamp 1569139307
transform 1 0 848 0 1 135
box -6 -6 6 6
use CONT  CONT_118
timestamp 1569139307
transform 1 0 812 0 1 135
box -6 -6 6 6
use CONT  CONT_119
timestamp 1569139307
transform 1 0 776 0 1 135
box -6 -6 6 6
use CONT  CONT_120
timestamp 1569139307
transform 1 0 740 0 1 135
box -6 -6 6 6
use CONT  CONT_121
timestamp 1569139307
transform 1 0 704 0 1 135
box -6 -6 6 6
use CONT  CONT_122
timestamp 1569139307
transform 1 0 668 0 1 135
box -6 -6 6 6
use CONT  CONT_123
timestamp 1569139307
transform 1 0 668 0 1 63
box -6 -6 6 6
use CONT  CONT_124
timestamp 1569139307
transform 1 0 1172 0 1 63
box -6 -6 6 6
use CONT  CONT_125
timestamp 1569139307
transform 1 0 1136 0 1 63
box -6 -6 6 6
use CONT  CONT_126
timestamp 1569139307
transform 1 0 920 0 1 63
box -6 -6 6 6
use CONT  CONT_127
timestamp 1569139307
transform 1 0 884 0 1 63
box -6 -6 6 6
use CONT  CONT_128
timestamp 1569139307
transform 1 0 848 0 1 63
box -6 -6 6 6
use CONT  CONT_129
timestamp 1569139307
transform 1 0 812 0 1 63
box -6 -6 6 6
use CONT  CONT_130
timestamp 1569139307
transform 1 0 632 0 1 99
box -6 -6 6 6
use CONT  CONT_131
timestamp 1569139307
transform 1 0 632 0 1 171
box -6 -6 6 6
use CONT  CONT_132
timestamp 1569139307
transform 1 0 632 0 1 27
box -6 -6 6 6
use CONT  CONT_133
timestamp 1569139307
transform 1 0 632 0 1 135
box -6 -6 6 6
use CONT  CONT_134
timestamp 1569139307
transform 1 0 632 0 1 63
box -6 -6 6 6
use CONT  CONT_135
timestamp 1569139307
transform 1 0 1388 0 1 135
box -6 -6 6 6
use CONT  CONT_136
timestamp 1569139307
transform 1 0 1352 0 1 135
box -6 -6 6 6
use CONT  CONT_137
timestamp 1569139307
transform 1 0 1316 0 1 135
box -6 -6 6 6
use CONT  CONT_138
timestamp 1569139307
transform 1 0 1280 0 1 135
box -6 -6 6 6
use CONT  CONT_139
timestamp 1569139307
transform 1 0 1244 0 1 135
box -6 -6 6 6
use CONT  CONT_140
timestamp 1569139307
transform 1 0 1316 0 1 27
box -6 -6 6 6
use CONT  CONT_141
timestamp 1569139307
transform 1 0 1748 0 1 63
box -6 -6 6 6
use CONT  CONT_142
timestamp 1569139307
transform 1 0 1532 0 1 63
box -6 -6 6 6
use CONT  CONT_143
timestamp 1569139307
transform 1 0 1496 0 1 63
box -6 -6 6 6
use CONT  CONT_144
timestamp 1569139307
transform 1 0 1460 0 1 63
box -6 -6 6 6
use CONT  CONT_145
timestamp 1569139307
transform 1 0 1424 0 1 63
box -6 -6 6 6
use CONT  CONT_146
timestamp 1569139307
transform 1 0 1388 0 1 63
box -6 -6 6 6
use CONT  CONT_147
timestamp 1569139307
transform 1 0 1352 0 1 63
box -6 -6 6 6
use CONT  CONT_148
timestamp 1569139307
transform 1 0 1316 0 1 63
box -6 -6 6 6
use CONT  CONT_149
timestamp 1569139307
transform 1 0 1280 0 1 63
box -6 -6 6 6
use CONT  CONT_150
timestamp 1569139307
transform 1 0 1244 0 1 63
box -6 -6 6 6
use CONT  CONT_151
timestamp 1569139307
transform 1 0 1244 0 1 27
box -6 -6 6 6
use CONT  CONT_152
timestamp 1569139307
transform 1 0 1748 0 1 171
box -6 -6 6 6
use CONT  CONT_153
timestamp 1569139307
transform 1 0 1532 0 1 171
box -6 -6 6 6
use CONT  CONT_154
timestamp 1569139307
transform 1 0 1496 0 1 171
box -6 -6 6 6
use CONT  CONT_155
timestamp 1569139307
transform 1 0 1460 0 1 171
box -6 -6 6 6
use CONT  CONT_156
timestamp 1569139307
transform 1 0 1424 0 1 171
box -6 -6 6 6
use CONT  CONT_157
timestamp 1569139307
transform 1 0 1388 0 1 171
box -6 -6 6 6
use CONT  CONT_158
timestamp 1569139307
transform 1 0 1352 0 1 171
box -6 -6 6 6
use CONT  CONT_159
timestamp 1569139307
transform 1 0 1316 0 1 171
box -6 -6 6 6
use CONT  CONT_160
timestamp 1569139307
transform 1 0 1280 0 1 171
box -6 -6 6 6
use CONT  CONT_161
timestamp 1569139307
transform 1 0 1244 0 1 171
box -6 -6 6 6
use CONT  CONT_162
timestamp 1569139307
transform 1 0 1352 0 1 27
box -6 -6 6 6
use CONT  CONT_163
timestamp 1569139307
transform 1 0 1532 0 1 27
box -6 -6 6 6
use CONT  CONT_164
timestamp 1569139307
transform 1 0 1496 0 1 27
box -6 -6 6 6
use CONT  CONT_165
timestamp 1569139307
transform 1 0 1460 0 1 27
box -6 -6 6 6
use CONT  CONT_166
timestamp 1569139307
transform 1 0 1424 0 1 27
box -6 -6 6 6
use CONT  CONT_167
timestamp 1569139307
transform 1 0 1388 0 1 27
box -6 -6 6 6
use CONT  CONT_168
timestamp 1569139307
transform 1 0 1748 0 1 27
box -6 -6 6 6
use CONT  CONT_169
timestamp 1569139307
transform 1 0 1748 0 1 99
box -6 -6 6 6
use CONT  CONT_170
timestamp 1569139307
transform 1 0 1532 0 1 99
box -6 -6 6 6
use CONT  CONT_171
timestamp 1569139307
transform 1 0 1496 0 1 99
box -6 -6 6 6
use CONT  CONT_172
timestamp 1569139307
transform 1 0 1460 0 1 99
box -6 -6 6 6
use CONT  CONT_173
timestamp 1569139307
transform 1 0 1424 0 1 99
box -6 -6 6 6
use CONT  CONT_174
timestamp 1569139307
transform 1 0 1388 0 1 99
box -6 -6 6 6
use CONT  CONT_175
timestamp 1569139307
transform 1 0 1352 0 1 99
box -6 -6 6 6
use CONT  CONT_176
timestamp 1569139307
transform 1 0 1316 0 1 99
box -6 -6 6 6
use CONT  CONT_177
timestamp 1569139307
transform 1 0 1280 0 1 99
box -6 -6 6 6
use CONT  CONT_178
timestamp 1569139307
transform 1 0 1244 0 1 99
box -6 -6 6 6
use CONT  CONT_179
timestamp 1569139307
transform 1 0 1280 0 1 27
box -6 -6 6 6
use CONT  CONT_180
timestamp 1569139307
transform 1 0 1748 0 1 135
box -6 -6 6 6
use CONT  CONT_181
timestamp 1569139307
transform 1 0 1532 0 1 135
box -6 -6 6 6
use CONT  CONT_182
timestamp 1569139307
transform 1 0 1496 0 1 135
box -6 -6 6 6
use CONT  CONT_183
timestamp 1569139307
transform 1 0 1460 0 1 135
box -6 -6 6 6
use CONT  CONT_184
timestamp 1569139307
transform 1 0 1424 0 1 135
box -6 -6 6 6
use CONT  CONT_185
timestamp 1569139307
transform 1 0 2360 0 1 171
box -6 -6 6 6
use CONT  CONT_186
timestamp 1569139307
transform 1 0 2324 0 1 171
box -6 -6 6 6
use CONT  CONT_187
timestamp 1569139307
transform 1 0 2288 0 1 171
box -6 -6 6 6
use CONT  CONT_188
timestamp 1569139307
transform 1 0 2252 0 1 171
box -6 -6 6 6
use CONT  CONT_189
timestamp 1569139307
transform 1 0 2216 0 1 171
box -6 -6 6 6
use CONT  CONT_190
timestamp 1569139307
transform 1 0 2180 0 1 171
box -6 -6 6 6
use CONT  CONT_191
timestamp 1569139307
transform 1 0 2144 0 1 171
box -6 -6 6 6
use CONT  CONT_192
timestamp 1569139307
transform 1 0 2108 0 1 171
box -6 -6 6 6
use CONT  CONT_193
timestamp 1569139307
transform 1 0 2072 0 1 171
box -6 -6 6 6
use CONT  CONT_194
timestamp 1569139307
transform 1 0 2036 0 1 171
box -6 -6 6 6
use CONT  CONT_195
timestamp 1569139307
transform 1 0 2000 0 1 171
box -6 -6 6 6
use CONT  CONT_196
timestamp 1569139307
transform 1 0 1964 0 1 171
box -6 -6 6 6
use CONT  CONT_197
timestamp 1569139307
transform 1 0 1928 0 1 171
box -6 -6 6 6
use CONT  CONT_198
timestamp 1569139307
transform 1 0 1892 0 1 171
box -6 -6 6 6
use CONT  CONT_199
timestamp 1569139307
transform 1 0 1856 0 1 171
box -6 -6 6 6
use CONT  CONT_200
timestamp 1569139307
transform 1 0 1820 0 1 171
box -6 -6 6 6
use CONT  CONT_201
timestamp 1569139307
transform 1 0 1928 0 1 27
box -6 -6 6 6
use CONT  CONT_202
timestamp 1569139307
transform 1 0 2360 0 1 135
box -6 -6 6 6
use CONT  CONT_203
timestamp 1569139307
transform 1 0 2324 0 1 135
box -6 -6 6 6
use CONT  CONT_204
timestamp 1569139307
transform 1 0 2288 0 1 135
box -6 -6 6 6
use CONT  CONT_205
timestamp 1569139307
transform 1 0 2252 0 1 135
box -6 -6 6 6
use CONT  CONT_206
timestamp 1569139307
transform 1 0 2216 0 1 135
box -6 -6 6 6
use CONT  CONT_207
timestamp 1569139307
transform 1 0 2180 0 1 135
box -6 -6 6 6
use CONT  CONT_208
timestamp 1569139307
transform 1 0 2144 0 1 135
box -6 -6 6 6
use CONT  CONT_209
timestamp 1569139307
transform 1 0 2108 0 1 135
box -6 -6 6 6
use CONT  CONT_210
timestamp 1569139307
transform 1 0 2072 0 1 135
box -6 -6 6 6
use CONT  CONT_211
timestamp 1569139307
transform 1 0 2036 0 1 135
box -6 -6 6 6
use CONT  CONT_212
timestamp 1569139307
transform 1 0 2000 0 1 135
box -6 -6 6 6
use CONT  CONT_213
timestamp 1569139307
transform 1 0 1964 0 1 135
box -6 -6 6 6
use CONT  CONT_214
timestamp 1569139307
transform 1 0 1928 0 1 135
box -6 -6 6 6
use CONT  CONT_215
timestamp 1569139307
transform 1 0 1892 0 1 135
box -6 -6 6 6
use CONT  CONT_216
timestamp 1569139307
transform 1 0 1856 0 1 135
box -6 -6 6 6
use CONT  CONT_217
timestamp 1569139307
transform 1 0 1820 0 1 135
box -6 -6 6 6
use CONT  CONT_218
timestamp 1569139307
transform 1 0 1892 0 1 27
box -6 -6 6 6
use CONT  CONT_219
timestamp 1569139307
transform 1 0 2360 0 1 99
box -6 -6 6 6
use CONT  CONT_220
timestamp 1569139307
transform 1 0 2324 0 1 99
box -6 -6 6 6
use CONT  CONT_221
timestamp 1569139307
transform 1 0 2288 0 1 99
box -6 -6 6 6
use CONT  CONT_222
timestamp 1569139307
transform 1 0 2252 0 1 99
box -6 -6 6 6
use CONT  CONT_223
timestamp 1569139307
transform 1 0 2216 0 1 99
box -6 -6 6 6
use CONT  CONT_224
timestamp 1569139307
transform 1 0 2180 0 1 99
box -6 -6 6 6
use CONT  CONT_225
timestamp 1569139307
transform 1 0 2144 0 1 99
box -6 -6 6 6
use CONT  CONT_226
timestamp 1569139307
transform 1 0 2108 0 1 99
box -6 -6 6 6
use CONT  CONT_227
timestamp 1569139307
transform 1 0 2072 0 1 99
box -6 -6 6 6
use CONT  CONT_228
timestamp 1569139307
transform 1 0 2036 0 1 99
box -6 -6 6 6
use CONT  CONT_229
timestamp 1569139307
transform 1 0 2000 0 1 99
box -6 -6 6 6
use CONT  CONT_230
timestamp 1569139307
transform 1 0 1964 0 1 99
box -6 -6 6 6
use CONT  CONT_231
timestamp 1569139307
transform 1 0 1928 0 1 99
box -6 -6 6 6
use CONT  CONT_232
timestamp 1569139307
transform 1 0 1892 0 1 99
box -6 -6 6 6
use CONT  CONT_233
timestamp 1569139307
transform 1 0 1856 0 1 99
box -6 -6 6 6
use CONT  CONT_234
timestamp 1569139307
transform 1 0 1820 0 1 99
box -6 -6 6 6
use CONT  CONT_235
timestamp 1569139307
transform 1 0 1856 0 1 27
box -6 -6 6 6
use CONT  CONT_236
timestamp 1569139307
transform 1 0 2360 0 1 63
box -6 -6 6 6
use CONT  CONT_237
timestamp 1569139307
transform 1 0 2324 0 1 63
box -6 -6 6 6
use CONT  CONT_238
timestamp 1569139307
transform 1 0 2288 0 1 63
box -6 -6 6 6
use CONT  CONT_239
timestamp 1569139307
transform 1 0 2252 0 1 63
box -6 -6 6 6
use CONT  CONT_240
timestamp 1569139307
transform 1 0 2216 0 1 63
box -6 -6 6 6
use CONT  CONT_241
timestamp 1569139307
transform 1 0 2180 0 1 63
box -6 -6 6 6
use CONT  CONT_242
timestamp 1569139307
transform 1 0 2144 0 1 63
box -6 -6 6 6
use CONT  CONT_243
timestamp 1569139307
transform 1 0 2108 0 1 63
box -6 -6 6 6
use CONT  CONT_244
timestamp 1569139307
transform 1 0 2072 0 1 63
box -6 -6 6 6
use CONT  CONT_245
timestamp 1569139307
transform 1 0 2036 0 1 63
box -6 -6 6 6
use CONT  CONT_246
timestamp 1569139307
transform 1 0 2000 0 1 63
box -6 -6 6 6
use CONT  CONT_247
timestamp 1569139307
transform 1 0 1964 0 1 63
box -6 -6 6 6
use CONT  CONT_248
timestamp 1569139307
transform 1 0 1928 0 1 63
box -6 -6 6 6
use CONT  CONT_249
timestamp 1569139307
transform 1 0 1892 0 1 63
box -6 -6 6 6
use CONT  CONT_250
timestamp 1569139307
transform 1 0 1856 0 1 63
box -6 -6 6 6
use CONT  CONT_251
timestamp 1569139307
transform 1 0 1820 0 1 63
box -6 -6 6 6
use CONT  CONT_252
timestamp 1569139307
transform 1 0 1820 0 1 27
box -6 -6 6 6
use CONT  CONT_253
timestamp 1569139307
transform 1 0 2360 0 1 27
box -6 -6 6 6
use CONT  CONT_254
timestamp 1569139307
transform 1 0 2324 0 1 27
box -6 -6 6 6
use CONT  CONT_255
timestamp 1569139307
transform 1 0 2288 0 1 27
box -6 -6 6 6
use CONT  CONT_256
timestamp 1569139307
transform 1 0 2252 0 1 27
box -6 -6 6 6
use CONT  CONT_257
timestamp 1569139307
transform 1 0 2216 0 1 27
box -6 -6 6 6
use CONT  CONT_258
timestamp 1569139307
transform 1 0 2180 0 1 27
box -6 -6 6 6
use CONT  CONT_259
timestamp 1569139307
transform 1 0 2144 0 1 27
box -6 -6 6 6
use CONT  CONT_260
timestamp 1569139307
transform 1 0 2108 0 1 27
box -6 -6 6 6
use CONT  CONT_261
timestamp 1569139307
transform 1 0 2072 0 1 27
box -6 -6 6 6
use CONT  CONT_262
timestamp 1569139307
transform 1 0 2036 0 1 27
box -6 -6 6 6
use CONT  CONT_263
timestamp 1569139307
transform 1 0 2000 0 1 27
box -6 -6 6 6
use CONT  CONT_264
timestamp 1569139307
transform 1 0 1964 0 1 27
box -6 -6 6 6
use CONT  CONT_265
timestamp 1569139307
transform 1 0 1784 0 1 171
box -6 -6 6 6
use CONT  CONT_266
timestamp 1569139307
transform 1 0 1784 0 1 135
box -6 -6 6 6
use CONT  CONT_267
timestamp 1569139307
transform 1 0 1784 0 1 99
box -6 -6 6 6
use CONT  CONT_268
timestamp 1569139307
transform 1 0 1784 0 1 63
box -6 -6 6 6
use CONT  CONT_269
timestamp 1569139307
transform 1 0 1784 0 1 27
box -6 -6 6 6
use CONT  CONT_270
timestamp 1569139307
transform 1 0 1208 0 1 171
box -6 -6 6 6
use CONT  CONT_271
timestamp 1569139307
transform 1 0 1208 0 1 135
box -6 -6 6 6
use CONT  CONT_272
timestamp 1569139307
transform 1 0 1208 0 1 99
box -6 -6 6 6
use CONT  CONT_273
timestamp 1569139307
transform 1 0 1208 0 1 63
box -6 -6 6 6
use CONT  CONT_274
timestamp 1569139307
transform 1 0 1208 0 1 27
box -6 -6 6 6
<< end >>
