magic
tech scmos
magscale 1 2
timestamp 1700034436
<< checkpaint >>
rect -50 -46 124 250
<< nwell >>
rect -10 96 84 210
<< ntransistor >>
rect 14 12 18 32
rect 48 12 52 52
rect 58 12 62 52
<< ptransistor >>
rect 14 148 18 188
rect 48 108 52 188
rect 58 108 62 188
<< ndiffusion >>
rect 38 51 48 52
rect 4 31 14 32
rect 12 13 14 31
rect 4 12 14 13
rect 18 31 28 32
rect 18 13 20 31
rect 18 12 28 13
rect 46 13 48 51
rect 38 12 48 13
rect 52 12 58 52
rect 62 51 72 52
rect 62 13 64 51
rect 62 12 72 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 149 14 187
rect 4 148 14 149
rect 18 187 28 188
rect 18 149 20 187
rect 18 148 28 149
rect 38 187 48 188
rect 46 109 48 187
rect 38 108 48 109
rect 52 108 58 188
rect 62 187 72 188
rect 62 109 64 187
rect 62 108 72 109
<< ndcontact >>
rect 4 13 12 31
rect 20 13 28 31
rect 38 13 46 51
rect 64 13 72 51
<< pdcontact >>
rect 4 149 12 187
rect 20 149 28 187
rect 38 109 46 187
rect 64 109 72 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 44 -4 52 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 44 196 52 204
<< polysilicon >>
rect 14 188 18 192
rect 48 188 52 192
rect 58 188 62 192
rect 14 134 18 148
rect 14 58 18 126
rect 48 70 52 108
rect 34 66 52 70
rect 58 74 62 108
rect 58 66 60 74
rect 14 54 52 58
rect 14 32 18 54
rect 48 52 52 54
rect 58 52 62 66
rect 14 8 18 12
rect 48 8 52 12
rect 58 8 62 12
<< polycontact >>
rect 12 126 20 134
rect 26 66 34 74
rect 60 66 68 74
<< metal1 >>
rect -4 204 84 206
rect 4 196 44 204
rect 52 196 84 204
rect -4 194 84 196
rect 4 187 12 194
rect 4 148 12 149
rect 20 187 28 188
rect 38 187 46 188
rect 28 149 32 154
rect 20 148 32 149
rect 4 126 12 134
rect 26 106 32 148
rect 38 108 46 109
rect 64 187 72 194
rect 64 108 72 109
rect 24 100 32 106
rect 24 80 30 100
rect 40 94 46 108
rect 36 86 46 94
rect 24 74 32 80
rect 26 32 32 66
rect 40 52 46 86
rect 68 66 76 74
rect 4 31 12 32
rect 4 6 12 13
rect 20 31 32 32
rect 28 24 32 31
rect 38 51 46 52
rect 20 12 28 13
rect 38 12 46 13
rect 64 51 72 52
rect 64 6 72 13
rect -4 4 84 6
rect 4 -4 44 4
rect 52 -4 84 4
rect -4 -6 84 -4
<< m1p >>
rect 4 126 12 134
rect 36 86 44 94
rect 68 66 76 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
port 4 se
rlabel metal1 8 0 8 0 4 gnd
port 5 se
rlabel metal1 8 130 8 130 4 EN
port 2 se
rlabel metal1 72 70 72 70 4 A
port 1 se
rlabel metal1 40 90 40 90 4 Y
port 3 se
<< end >>
