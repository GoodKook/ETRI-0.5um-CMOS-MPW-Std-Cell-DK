magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -15 -15 455 455
use pnp5_CDNS_7230122529116  pnp5_CDNS_7230122529116_0
timestamp 1555596690
transform 1 0 0 0 1 0
box 45 45 395 395
<< end >>
