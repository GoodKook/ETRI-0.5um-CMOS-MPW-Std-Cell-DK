magic
tech scmos
magscale 1 2
timestamp 1727518396
<< checkpaint >>
rect -97 -84 6617 6604
<< error_p >>
rect 4073 6173 4087 6187
rect 1873 4193 1887 4207
rect 5313 4193 5327 4207
rect 4052 3253 4066 3267
rect 6113 2013 6127 2027
rect 4413 1753 4427 1767
rect 5813 973 5827 987
<< nwell >>
rect 4175 5622 4189 5626
rect 5317 4193 5327 4207
<< metal1 >>
rect -57 6258 3 6518
rect 6490 6502 6577 6518
rect 357 6427 363 6473
rect 806 6423 820 6427
rect 806 6413 823 6423
rect 817 6287 823 6413
rect 1577 6287 1583 6413
rect 2337 6327 2343 6413
rect 2497 6307 2503 6333
rect 2617 6327 2623 6473
rect 3077 6327 3083 6353
rect 4677 6287 4683 6453
rect 5457 6303 5463 6353
rect 5437 6297 5463 6303
rect -57 6242 30 6258
rect -57 5738 3 6242
rect 857 6047 863 6153
rect 1017 6027 1023 6173
rect 2097 6067 2103 6133
rect 2537 6047 2543 6213
rect 3477 6027 3483 6133
rect 4077 6127 4083 6173
rect 6517 5998 6577 6502
rect 6490 5982 6577 5998
rect 1937 5767 1943 5893
rect 2297 5767 2303 5813
rect 2317 5787 2323 5933
rect 2457 5787 2463 5953
rect 2477 5767 2483 5953
rect 2497 5767 2503 5813
rect 2757 5767 2763 5953
rect 3557 5807 3563 5873
rect 4597 5767 4603 5793
rect 5197 5787 5203 5813
rect 5317 5767 5323 5953
rect 5497 5807 5503 5853
rect 5817 5807 5823 5893
rect 6257 5867 6263 5933
rect -57 5722 30 5738
rect -57 5218 3 5722
rect 1360 5703 1373 5707
rect 1357 5693 1373 5703
rect 357 5567 363 5653
rect 1357 5567 1363 5693
rect 1677 5567 1683 5673
rect 1857 5607 1863 5693
rect 3357 5647 3363 5673
rect 2017 5527 2023 5593
rect 3357 5587 3363 5612
rect 3377 5527 3383 5613
rect 3617 5527 3623 5693
rect 3737 5647 3743 5673
rect 3897 5567 3903 5693
rect 4617 5507 4623 5693
rect 4937 5567 4943 5693
rect 5737 5567 5743 5693
rect 4897 5507 4903 5553
rect 6097 5507 6103 5653
rect 6377 5627 6383 5673
rect 6497 5567 6503 5693
rect 4617 5497 4632 5507
rect 4620 5493 4632 5497
rect 6517 5478 6577 5982
rect 6490 5462 6577 5478
rect 1747 5440 1783 5443
rect 1747 5437 1787 5440
rect 817 5267 823 5433
rect 1773 5427 1787 5437
rect 1773 5420 1774 5427
rect 1240 5403 1253 5407
rect 1237 5393 1253 5403
rect 1237 5287 1243 5393
rect 1417 5307 1423 5353
rect 1757 5327 1763 5413
rect 3317 5387 3323 5433
rect 3217 5247 3223 5293
rect 3597 5247 3603 5433
rect 3800 5423 3812 5427
rect 3797 5413 3812 5423
rect 3617 5287 3623 5413
rect 3797 5247 3803 5413
rect 4057 5247 4063 5433
rect 4457 5247 4463 5353
rect 4477 5267 4483 5393
rect 5297 5267 5303 5333
rect 5317 5287 5323 5413
rect 5577 5407 5583 5433
rect 5597 5347 5603 5413
rect 5857 5287 5863 5413
rect 5877 5307 5883 5433
rect -57 5202 30 5218
rect -57 4698 3 5202
rect 197 5007 203 5153
rect 537 4987 543 5173
rect 1117 5047 1123 5173
rect 1457 5027 1463 5173
rect 1477 5047 1483 5153
rect 1617 5047 1623 5133
rect 1797 5047 1803 5173
rect 2297 5007 2303 5153
rect 2637 5147 2643 5173
rect 2637 5067 2643 5133
rect 2757 5127 2763 5173
rect 3057 5107 3063 5153
rect 2917 5027 2923 5073
rect 2957 5007 2963 5093
rect 2948 4997 2963 5007
rect 2948 4993 2960 4997
rect 3257 4987 3263 5173
rect 3377 4987 3383 5133
rect 3397 4987 3403 5173
rect 3897 5063 3903 5133
rect 4437 5087 4443 5153
rect 4457 5127 4463 5173
rect 3897 5057 3923 5063
rect 3917 5047 3923 5057
rect 3917 5037 3934 5047
rect 3920 5033 3934 5037
rect 4597 4987 4603 5153
rect 5697 5127 5703 5153
rect 5817 5127 5823 5173
rect 5257 4987 5263 5093
rect 5457 4987 5463 5033
rect 6517 4958 6577 5462
rect 6490 4942 6577 4958
rect 1177 4847 1183 4893
rect 1497 4867 1503 4893
rect 2237 4887 2243 4913
rect 1177 4837 1193 4847
rect 1180 4833 1193 4837
rect 737 4767 743 4813
rect 1497 4727 1503 4753
rect 1797 4747 1803 4813
rect 2617 4727 2623 4893
rect 2877 4727 2883 4833
rect 2917 4807 2923 4873
rect 3077 4727 3083 4913
rect 3197 4767 3203 4913
rect 3677 4897 3714 4903
rect 3677 4803 3683 4897
rect 3657 4797 3683 4803
rect 3377 4727 3383 4773
rect 3657 4747 3663 4797
rect 3777 4727 3783 4773
rect 4477 4727 4483 4853
rect 4497 4767 4503 4913
rect 4537 4727 4543 4893
rect 4677 4747 4683 4913
rect 4877 4807 4883 4913
rect 5197 4727 5203 4913
rect 5677 4787 5683 4913
rect 2877 4717 2893 4727
rect 2880 4713 2893 4717
rect -57 4682 30 4698
rect -57 4178 3 4682
rect 477 4637 513 4643
rect 17 4547 23 4593
rect 477 4487 483 4637
rect 497 4527 503 4613
rect 1177 4487 1183 4653
rect 1317 4487 1323 4593
rect 1997 4567 2003 4613
rect 2137 4547 2143 4653
rect 2297 4507 2303 4653
rect 2637 4527 2643 4653
rect 3640 4643 3653 4647
rect 3637 4633 3653 4643
rect 5460 4643 5473 4647
rect 5457 4633 5473 4643
rect 2957 4507 2963 4633
rect 3197 4527 3203 4633
rect 3217 4487 3223 4513
rect 3637 4487 3643 4633
rect 4597 4567 4603 4633
rect 5457 4587 5463 4633
rect 4857 4467 4863 4513
rect 6517 4438 6577 4942
rect 6490 4422 6577 4438
rect 1037 4247 1043 4393
rect 1057 4227 1063 4253
rect 1197 4207 1203 4373
rect 1337 4207 1343 4393
rect 1697 4307 1703 4333
rect 1877 4207 1883 4393
rect 2037 4227 2043 4373
rect 2057 4247 2063 4393
rect 2537 4247 2543 4353
rect 2957 4207 2963 4333
rect 3173 4227 3187 4233
rect 3317 4227 3323 4333
rect 3167 4220 3187 4227
rect 3167 4217 3183 4220
rect 3167 4213 3180 4217
rect 3697 4207 3703 4373
rect 3837 4247 3843 4293
rect 4557 4247 4563 4393
rect 5317 4207 5323 4333
rect 5437 4207 5443 4233
rect 5477 4207 5483 4373
rect 5957 4287 5963 4333
rect 2957 4197 2973 4207
rect 2960 4193 2973 4197
rect 5317 4193 5326 4207
rect -57 4162 30 4178
rect -57 3658 3 4162
rect 737 4007 743 4093
rect 897 4047 903 4093
rect 1177 3967 1183 4073
rect 1277 3947 1283 4113
rect 1577 4007 1583 4133
rect 1737 4047 1743 4093
rect 2057 4007 2063 4133
rect 2217 4007 2223 4073
rect 2217 3997 2233 4007
rect 2220 3993 2233 3997
rect 2457 3947 2463 3993
rect 2677 3947 2683 4113
rect 3017 4087 3023 4133
rect 3157 4087 3163 4113
rect 3577 3947 3583 4033
rect 3717 3947 3723 4133
rect 4537 3967 4543 4133
rect 4557 4047 4563 4093
rect 4677 3947 4683 4133
rect 4837 3987 4843 4113
rect 5597 3947 5603 4133
rect 5617 3947 5623 3973
rect 5777 3947 5783 4053
rect 5917 3967 5923 4093
rect 6057 3967 6063 4113
rect 6377 4007 6383 4133
rect 6517 3918 6577 4422
rect 6490 3902 6577 3918
rect 2326 3880 2363 3883
rect 2326 3877 2367 3880
rect 2353 3867 2367 3877
rect 2353 3860 2354 3867
rect 657 3827 663 3853
rect 337 3687 343 3813
rect 497 3707 503 3813
rect 2317 3687 2323 3813
rect 2337 3687 2343 3853
rect 2477 3727 2483 3813
rect 3137 3747 3143 3853
rect 4577 3687 4583 3753
rect 4597 3727 4603 3793
rect 4737 3767 4743 3853
rect 4917 3707 4923 3873
rect 5037 3787 5043 3853
rect 5677 3827 5683 3853
rect 5557 3727 5563 3813
rect 5697 3687 5703 3773
rect 5717 3707 5723 3853
rect 6017 3727 6023 3833
rect 6397 3767 6403 3853
rect -57 3642 30 3658
rect -57 3138 3 3642
rect 837 3487 843 3573
rect 857 3427 863 3613
rect 1617 3487 1623 3573
rect 2117 3487 2123 3613
rect 2497 3467 2503 3553
rect 2517 3447 2523 3593
rect 3237 3547 3243 3613
rect 3357 3427 3363 3473
rect 4777 3447 4783 3573
rect 5597 3427 5603 3573
rect 5737 3427 5743 3593
rect 5757 3447 5763 3533
rect 5957 3447 5963 3573
rect 6297 3427 6303 3533
rect 6517 3398 6577 3902
rect 6490 3382 6577 3398
rect 677 3187 683 3213
rect 957 3167 963 3313
rect 977 3227 983 3333
rect 2177 3267 2183 3353
rect 2197 3207 2203 3353
rect 2337 3187 2343 3353
rect 2357 3207 2363 3293
rect 2537 3207 2543 3293
rect 3777 3207 3783 3353
rect 4057 3281 4063 3353
rect 4177 3167 4183 3353
rect 4528 3263 4540 3267
rect 4528 3253 4543 3263
rect 4537 3207 4543 3253
rect 4637 3227 4643 3353
rect 4837 3307 4843 3333
rect 4627 3217 4643 3227
rect 4627 3213 4640 3217
rect 5057 3187 5063 3353
rect 5077 3167 5083 3353
rect 6400 3363 6413 3367
rect 6397 3353 6413 3363
rect 5237 3207 5243 3333
rect 5857 3167 5863 3293
rect 5897 3187 5903 3352
rect 6197 3167 6203 3293
rect 6397 3267 6403 3353
rect -57 3122 30 3138
rect -57 2618 3 3122
rect 237 2967 243 3093
rect 2197 3027 2203 3073
rect 2217 2967 2223 3093
rect 2517 2907 2523 3093
rect 2537 2907 2543 3013
rect 2717 2907 2723 3033
rect 4517 2907 4523 3093
rect 4657 2927 4663 3013
rect 4697 2927 4703 3093
rect 4837 2927 4843 3013
rect 4997 2967 5003 3093
rect 5477 2967 5483 3073
rect 4857 2907 4863 2953
rect 5157 2907 5163 2953
rect 5797 2927 5803 3073
rect 5977 2907 5983 3053
rect 6137 2907 6143 3073
rect 6157 2907 6163 3053
rect 6297 2907 6303 3073
rect 6457 2907 6463 3093
rect 6497 2987 6503 3093
rect 2537 2897 2553 2907
rect 2540 2893 2553 2897
rect 6127 2897 6143 2907
rect 6127 2893 6140 2897
rect 6517 2878 6577 3382
rect 6490 2862 6577 2878
rect 617 2727 623 2813
rect 757 2747 763 2793
rect 317 2687 323 2713
rect 1177 2667 1183 2773
rect 2257 2727 2263 2833
rect 2397 2687 2403 2773
rect 2697 2667 2703 2833
rect 3517 2687 3523 2813
rect 4477 2787 4483 2833
rect 4137 2667 4143 2733
rect 4737 2727 4743 2813
rect 4437 2687 4443 2713
rect 4857 2687 4863 2733
rect 4437 2677 4454 2687
rect 4440 2673 4454 2677
rect 4877 2647 4883 2773
rect 4897 2687 4903 2813
rect 5017 2783 5023 2833
rect 5017 2777 5043 2783
rect 5037 2667 5043 2777
rect 5397 2747 5403 2813
rect 5577 2647 5583 2813
rect -57 2602 30 2618
rect -57 2098 3 2602
rect 357 2407 363 2433
rect 817 2387 823 2473
rect 977 2447 983 2573
rect 2137 2427 2143 2553
rect 2397 2507 2403 2573
rect 2437 2467 2443 2573
rect 2557 2527 2563 2573
rect 2417 2407 2423 2433
rect 3197 2407 3203 2553
rect 3568 2543 3580 2547
rect 3568 2533 3583 2543
rect 3457 2407 3463 2493
rect 3477 2387 3483 2433
rect 3577 2407 3583 2533
rect 3597 2447 3603 2533
rect 3737 2427 3743 2573
rect 3757 2387 3763 2513
rect 4037 2447 4043 2573
rect 4217 2387 4223 2573
rect 4317 2387 4323 2533
rect 4457 2387 4463 2573
rect 4737 2547 4743 2573
rect 4917 2427 4923 2533
rect 5097 2447 5103 2573
rect 5117 2467 5123 2513
rect 5137 2427 5143 2573
rect 5417 2447 5423 2573
rect 6157 2387 6163 2553
rect 6297 2447 6303 2573
rect 6517 2358 6577 2862
rect 6490 2342 6577 2358
rect 1397 2127 1403 2153
rect 1717 2147 1723 2253
rect 3097 2147 3103 2213
rect 3437 2147 3443 2273
rect 3457 2127 3463 2253
rect 3657 2147 3663 2293
rect 3977 2223 3983 2313
rect 3977 2217 4003 2223
rect 3997 2147 4003 2217
rect 4117 2187 4123 2253
rect 4137 2147 4143 2213
rect 4457 2147 4463 2193
rect 4897 2127 4903 2253
rect 5477 2127 5483 2193
rect 6257 2167 6263 2253
rect -57 2082 30 2098
rect -57 1578 3 2082
rect 197 1887 203 1973
rect 1737 1887 1743 1933
rect 2577 1887 2583 1993
rect 2597 1867 2603 2053
rect 2737 1947 2743 2053
rect 2857 2007 2863 2033
rect 3257 1867 3263 1933
rect 3697 1887 3703 1933
rect 4000 1883 4013 1887
rect 3997 1880 4013 1883
rect 3993 1873 4013 1880
rect 3993 1867 4007 1873
rect 4037 1867 4043 2033
rect 4177 1947 4183 2053
rect 4317 1867 4323 1953
rect 4417 1887 4423 2053
rect 4557 1867 4563 1913
rect 4577 1907 4583 2033
rect 4757 1947 4763 2033
rect 5057 1967 5063 2013
rect 5077 1887 5083 2053
rect 5217 1887 5223 1953
rect 5237 1867 5243 2013
rect 5257 1967 5263 2053
rect 5497 2027 5503 2053
rect 6117 1964 6123 1996
rect 6517 1838 6577 2342
rect 6490 1822 6577 1838
rect 3126 1803 3140 1807
rect 3126 1800 3143 1803
rect 3126 1793 3147 1800
rect 197 1747 203 1793
rect 1337 1607 1343 1653
rect 1377 1647 1383 1773
rect 1557 1607 1563 1773
rect 1697 1687 1703 1793
rect 1717 1627 1723 1773
rect 1857 1627 1863 1773
rect 2057 1607 2063 1793
rect 2177 1647 2183 1793
rect 3133 1787 3147 1793
rect 3267 1777 3293 1783
rect 2217 1687 2223 1773
rect 2637 1607 2643 1773
rect 2837 1687 2843 1733
rect 2857 1627 2863 1693
rect 2877 1607 2883 1633
rect 3397 1607 3403 1753
rect 3577 1627 3583 1773
rect 3737 1607 3743 1733
rect 3757 1627 3763 1793
rect 3877 1747 3883 1773
rect 3917 1627 3923 1773
rect 4037 1627 4043 1673
rect 4257 1667 4263 1773
rect 4540 1763 4553 1767
rect 4537 1760 4553 1763
rect 4533 1753 4553 1760
rect 4533 1747 4547 1753
rect 4277 1647 4283 1733
rect 4417 1667 4423 1739
rect 4546 1740 4547 1747
rect 5077 1667 5083 1793
rect 6197 1747 6203 1793
rect 4037 1617 4053 1627
rect 4040 1613 4053 1617
rect 5557 1607 5563 1733
rect 6497 1647 6503 1773
rect 1547 1597 1563 1607
rect 1547 1593 1560 1597
rect 3397 1597 3413 1607
rect 3400 1593 3413 1597
rect -57 1562 30 1578
rect -57 1058 3 1562
rect 177 1367 183 1473
rect 197 1347 203 1513
rect 377 1407 383 1513
rect 1277 1347 1283 1533
rect 1717 1507 1723 1533
rect 2477 1367 2483 1473
rect 2937 1467 2943 1513
rect 2617 1347 2623 1373
rect 3237 1367 3243 1453
rect 3377 1347 3383 1373
rect 3397 1347 3403 1413
rect 3637 1367 3643 1453
rect 3657 1427 3663 1513
rect 3777 1447 3783 1493
rect 3797 1347 3803 1513
rect 4157 1387 4163 1513
rect 4617 1347 4623 1533
rect 4997 1407 5003 1513
rect 5317 1387 5323 1493
rect 5337 1387 5343 1413
rect 5307 1377 5323 1387
rect 5307 1373 5320 1377
rect 5617 1347 5623 1533
rect 5637 1427 5643 1513
rect 5657 1367 5663 1393
rect 6517 1318 6577 1822
rect 6490 1302 6577 1318
rect 4967 1283 4980 1287
rect 4967 1273 4983 1283
rect 217 1147 223 1253
rect 537 1127 543 1153
rect 526 1117 543 1127
rect 526 1113 540 1117
rect 957 1107 963 1213
rect 2557 1127 2563 1253
rect 2717 1127 2723 1253
rect 2737 1227 2743 1273
rect 2837 1087 2843 1213
rect 3137 1107 3143 1213
rect 4197 1107 4203 1273
rect 4326 1223 4340 1227
rect 4326 1213 4343 1223
rect 4337 1127 4343 1213
rect 4357 1147 4363 1253
rect 4377 1107 4383 1273
rect 4977 1127 4983 1273
rect 5317 1107 5323 1253
rect 5457 1087 5463 1213
rect 5477 1107 5483 1273
rect 5637 1217 5673 1223
rect 5637 1087 5643 1217
rect -57 1042 30 1058
rect -57 538 3 1042
rect 517 847 523 873
rect 657 847 663 973
rect 1277 847 1283 933
rect 1737 867 1743 993
rect 2337 827 2343 993
rect 3097 827 3103 933
rect 3257 887 3263 973
rect 3277 827 3283 993
rect 3297 987 3303 1013
rect 3417 827 3423 873
rect 3437 827 3443 1013
rect 4217 827 4223 993
rect 4357 847 4363 973
rect 4677 847 4683 993
rect 5617 923 5623 973
rect 5617 917 5643 923
rect 4357 837 4373 847
rect 4360 833 4373 837
rect 4697 827 4703 913
rect 5637 887 5643 917
rect 5817 867 5823 959
rect 6517 798 6577 1302
rect 6490 782 6577 798
rect 477 607 483 693
rect 817 627 823 733
rect 957 587 963 753
rect 1977 567 1983 693
rect 2137 567 2143 693
rect 2757 567 2763 733
rect 2937 587 2943 693
rect 3277 627 3283 733
rect 3297 667 3303 753
rect 3317 567 3323 653
rect 3437 627 3443 733
rect 3620 703 3634 707
rect 3617 693 3634 703
rect 3617 567 3623 693
rect 4217 567 4223 753
rect 4917 707 4923 753
rect 5777 707 5783 733
rect 4397 587 4403 693
rect 4577 587 4583 693
rect 5057 567 5063 693
rect 5217 607 5223 693
rect 5417 567 5423 633
rect 5580 583 5593 587
rect 5577 580 5593 583
rect 5573 573 5593 580
rect 5573 567 5587 573
rect -57 522 30 538
rect -57 18 3 522
rect 817 327 823 493
rect 837 387 843 433
rect 977 347 983 453
rect 977 337 993 347
rect 980 333 993 337
rect 1777 327 1783 493
rect 3097 407 3103 473
rect 3317 467 3323 493
rect 3517 367 3523 493
rect 3837 307 3843 493
rect 3857 347 3863 493
rect 4037 347 4043 493
rect 3857 337 3873 347
rect 3860 333 3873 337
rect 4217 307 4223 473
rect 5497 327 5503 453
rect 5617 307 5623 473
rect 5997 327 6003 453
rect 6517 278 6577 782
rect 6490 262 6577 278
rect 217 87 223 173
rect 357 67 363 213
rect 377 147 383 173
rect 677 87 683 133
rect 697 47 703 213
rect 717 87 723 233
rect 857 87 863 213
rect 1037 87 1043 173
rect 1157 47 1163 213
rect 1197 67 1203 173
rect 1337 87 1343 233
rect 2157 47 2163 213
rect 2297 87 2303 233
rect 3037 47 3043 153
rect 3217 87 3223 173
rect 3537 127 3543 213
rect 3697 67 3703 173
rect 3717 147 3723 193
rect 3877 127 3883 233
rect 3897 87 3903 153
rect 4937 67 4943 213
rect 6037 67 6043 173
rect 6197 127 6203 233
rect 6217 87 6223 173
rect -57 2 30 18
rect 6517 2 6577 262
<< m2contact >>
rect 353 6473 367 6487
rect 2613 6473 2627 6487
rect 353 6413 367 6427
rect 792 6413 806 6427
rect 1573 6413 1587 6427
rect 2333 6413 2347 6427
rect 2493 6333 2507 6347
rect 2333 6313 2347 6327
rect 4673 6453 4687 6467
rect 3073 6353 3087 6367
rect 2613 6313 2627 6327
rect 3073 6313 3087 6327
rect 2493 6293 2507 6307
rect 5453 6353 5467 6367
rect 813 6273 827 6287
rect 1573 6273 1587 6287
rect 4672 6273 4686 6287
rect 2534 6213 2548 6227
rect 5170 6213 5184 6227
rect 1013 6173 1027 6187
rect 853 6153 867 6167
rect 853 6033 867 6047
rect 2093 6133 2107 6147
rect 2093 6053 2107 6067
rect 5317 6193 5331 6207
rect 4073 6173 4087 6187
rect 3473 6133 3487 6147
rect 2533 6033 2547 6047
rect 4073 6113 4087 6127
rect 1013 6013 1027 6027
rect 3473 6013 3487 6027
rect 2452 5953 2466 5967
rect 2474 5953 2488 5967
rect 2753 5953 2767 5967
rect 5313 5953 5327 5967
rect 2313 5933 2327 5947
rect 1933 5893 1947 5907
rect 2293 5813 2307 5827
rect 2314 5773 2328 5787
rect 2453 5773 2467 5787
rect 2493 5813 2507 5827
rect 3553 5873 3567 5887
rect 5193 5813 5207 5827
rect 3553 5793 3567 5807
rect 4594 5793 4608 5807
rect 5193 5773 5207 5787
rect 6253 5933 6267 5947
rect 5813 5893 5827 5907
rect 5493 5853 5507 5867
rect 6253 5853 6267 5867
rect 5494 5793 5508 5807
rect 5813 5793 5827 5807
rect 1933 5753 1947 5767
rect 2293 5753 2307 5767
rect 2472 5753 2486 5767
rect 2494 5753 2508 5767
rect 2752 5753 2766 5767
rect 4592 5753 4606 5767
rect 5314 5753 5328 5767
rect 1373 5693 1387 5707
rect 1853 5693 1867 5707
rect 3613 5693 3627 5707
rect 3893 5693 3907 5707
rect 4613 5693 4627 5707
rect 4933 5693 4947 5707
rect 5733 5693 5747 5707
rect 6493 5693 6507 5707
rect 353 5653 367 5667
rect 1673 5673 1687 5687
rect 3353 5673 3367 5687
rect 3353 5633 3367 5647
rect 3352 5612 3366 5626
rect 3374 5613 3388 5627
rect 1853 5593 1867 5607
rect 2013 5593 2027 5607
rect 352 5553 366 5567
rect 1353 5553 1367 5567
rect 1672 5553 1686 5567
rect 3353 5573 3367 5587
rect 3733 5673 3747 5687
rect 3733 5633 3747 5647
rect 3893 5553 3907 5567
rect 2013 5513 2027 5527
rect 3373 5513 3387 5527
rect 3613 5513 3627 5527
rect 6373 5673 6387 5687
rect 6093 5653 6107 5667
rect 4893 5553 4907 5567
rect 4933 5553 4947 5567
rect 5733 5553 5747 5567
rect 6373 5613 6387 5627
rect 6493 5553 6507 5567
rect 4632 5493 4646 5507
rect 4893 5493 4907 5507
rect 6093 5493 6107 5507
rect 813 5433 827 5447
rect 1733 5433 1747 5447
rect 3312 5433 3326 5447
rect 3593 5433 3607 5447
rect 4053 5433 4067 5447
rect 5574 5433 5588 5447
rect 5873 5433 5887 5447
rect 1752 5413 1766 5427
rect 1774 5413 1788 5427
rect 1253 5393 1267 5407
rect 1413 5353 1427 5367
rect 3313 5373 3327 5387
rect 1753 5313 1767 5327
rect 1413 5293 1427 5307
rect 3213 5293 3227 5307
rect 1233 5273 1247 5287
rect 813 5253 827 5267
rect 3613 5413 3627 5427
rect 3812 5413 3826 5427
rect 3613 5273 3627 5287
rect 5313 5413 5327 5427
rect 4473 5393 4487 5407
rect 4453 5353 4467 5367
rect 5293 5333 5307 5347
rect 5593 5413 5607 5427
rect 5853 5413 5867 5427
rect 5573 5393 5587 5407
rect 5593 5333 5607 5347
rect 5873 5293 5887 5307
rect 5313 5273 5327 5287
rect 5853 5273 5867 5287
rect 4473 5253 4487 5267
rect 5293 5253 5307 5267
rect 3213 5233 3227 5247
rect 3593 5233 3607 5247
rect 3793 5233 3807 5247
rect 4053 5233 4067 5247
rect 4453 5233 4467 5247
rect 533 5173 547 5187
rect 1113 5173 1127 5187
rect 1453 5173 1467 5187
rect 1793 5173 1807 5187
rect 2633 5173 2647 5187
rect 2753 5173 2767 5187
rect 3253 5173 3267 5187
rect 3393 5173 3407 5187
rect 4453 5173 4467 5187
rect 5813 5173 5827 5187
rect 193 5153 207 5167
rect 193 4993 207 5007
rect 1113 5033 1127 5047
rect 1473 5153 1487 5167
rect 1613 5133 1627 5147
rect 2293 5153 2307 5167
rect 1473 5033 1487 5047
rect 1613 5033 1627 5047
rect 1793 5033 1807 5047
rect 1453 5013 1467 5027
rect 2634 5133 2648 5147
rect 3053 5153 3067 5167
rect 2752 5113 2766 5127
rect 2953 5093 2967 5107
rect 3053 5093 3067 5107
rect 2913 5073 2927 5087
rect 2633 5053 2647 5067
rect 2914 5013 2928 5027
rect 2293 4993 2307 5007
rect 2934 4993 2948 5007
rect 3373 5133 3387 5147
rect 4433 5153 4447 5167
rect 3892 5133 3906 5147
rect 4593 5153 4607 5167
rect 5693 5153 5707 5167
rect 4453 5113 4467 5127
rect 4433 5073 4447 5087
rect 3934 5033 3948 5047
rect 5692 5113 5706 5127
rect 5813 5113 5827 5127
rect 5253 5093 5267 5107
rect 5453 5033 5467 5047
rect 533 4973 547 4987
rect 3253 4973 3267 4987
rect 3372 4973 3386 4987
rect 3394 4973 3408 4987
rect 4593 4973 4607 4987
rect 5253 4973 5267 4987
rect 5453 4973 5467 4987
rect 2233 4913 2247 4927
rect 3073 4913 3087 4927
rect 3193 4913 3207 4927
rect 4493 4913 4507 4927
rect 4673 4913 4687 4927
rect 4873 4913 4887 4927
rect 5193 4913 5207 4927
rect 5674 4913 5688 4927
rect 1173 4893 1187 4907
rect 1492 4893 1506 4907
rect 2613 4893 2627 4907
rect 2233 4873 2247 4887
rect 1493 4853 1507 4867
rect 1193 4833 1207 4847
rect 733 4813 747 4827
rect 1793 4813 1807 4827
rect 733 4753 747 4767
rect 1493 4753 1507 4767
rect 1793 4733 1807 4747
rect 2913 4873 2927 4887
rect 2873 4833 2887 4847
rect 2913 4793 2927 4807
rect 3714 4893 3728 4907
rect 4473 4853 4487 4867
rect 3373 4773 3387 4787
rect 3193 4753 3207 4767
rect 3773 4773 3787 4787
rect 3652 4733 3666 4747
rect 4533 4893 4547 4907
rect 4493 4753 4507 4767
rect 4873 4793 4887 4807
rect 4673 4733 4687 4747
rect 5673 4773 5687 4787
rect 1493 4713 1507 4727
rect 2613 4713 2627 4727
rect 2893 4713 2907 4727
rect 3073 4713 3087 4727
rect 3374 4713 3388 4727
rect 3773 4713 3787 4727
rect 4473 4713 4487 4727
rect 4533 4713 4547 4727
rect 5193 4713 5207 4727
rect 1173 4653 1187 4667
rect 2133 4653 2147 4667
rect 2293 4653 2307 4667
rect 2633 4653 2647 4667
rect 13 4593 27 4607
rect 13 4533 27 4547
rect 513 4633 527 4647
rect 493 4613 507 4627
rect 493 4513 507 4527
rect 1993 4613 2007 4627
rect 1313 4593 1327 4607
rect 1993 4553 2007 4567
rect 2133 4533 2147 4547
rect 2953 4633 2967 4647
rect 3193 4633 3207 4647
rect 3653 4633 3667 4647
rect 4593 4633 4607 4647
rect 5473 4633 5487 4647
rect 2633 4513 2647 4527
rect 3192 4513 3206 4527
rect 3214 4513 3228 4527
rect 2293 4493 2307 4507
rect 2953 4493 2967 4507
rect 5453 4573 5467 4587
rect 4593 4553 4607 4567
rect 4853 4513 4867 4527
rect 473 4473 487 4487
rect 1174 4473 1188 4487
rect 1313 4473 1327 4487
rect 3213 4473 3227 4487
rect 3633 4473 3647 4487
rect 4853 4453 4867 4467
rect 1033 4393 1047 4407
rect 1333 4393 1347 4407
rect 1873 4393 1887 4407
rect 2053 4393 2067 4407
rect 4553 4393 4567 4407
rect 1193 4373 1207 4387
rect 1053 4253 1067 4267
rect 1033 4233 1047 4247
rect 1053 4213 1067 4227
rect 1693 4333 1707 4347
rect 1693 4293 1707 4307
rect 2033 4373 2047 4387
rect 3693 4373 3707 4387
rect 2533 4353 2547 4367
rect 2953 4333 2967 4347
rect 3313 4333 3327 4347
rect 2053 4233 2067 4247
rect 2533 4233 2547 4247
rect 2033 4213 2047 4227
rect 3173 4233 3187 4247
rect 3153 4213 3167 4227
rect 3313 4213 3327 4227
rect 3833 4293 3847 4307
rect 5473 4373 5487 4387
rect 5314 4333 5328 4347
rect 3833 4233 3847 4247
rect 4553 4233 4567 4247
rect 5433 4233 5447 4247
rect 5954 4333 5968 4347
rect 5953 4273 5967 4287
rect 1193 4193 1207 4207
rect 1333 4193 1347 4207
rect 1873 4193 1887 4207
rect 2973 4193 2987 4207
rect 3692 4193 3706 4207
rect 5326 4193 5340 4207
rect 5432 4193 5446 4207
rect 5472 4193 5486 4207
rect 1573 4133 1587 4147
rect 2053 4133 2067 4147
rect 3013 4133 3027 4147
rect 3713 4133 3727 4147
rect 4533 4133 4547 4147
rect 4673 4133 4687 4147
rect 5593 4133 5607 4147
rect 6373 4133 6387 4147
rect 1273 4113 1287 4127
rect 733 4093 747 4107
rect 893 4093 907 4107
rect 1173 4073 1187 4087
rect 893 4033 907 4047
rect 733 3993 747 4007
rect 1173 3953 1187 3967
rect 1733 4093 1747 4107
rect 1733 4033 1747 4047
rect 2673 4113 2687 4127
rect 2213 4073 2227 4087
rect 1572 3993 1586 4007
rect 2053 3993 2067 4007
rect 2233 3993 2247 4007
rect 2452 3993 2466 4007
rect 3154 4113 3168 4127
rect 3013 4073 3027 4087
rect 3153 4073 3167 4087
rect 3573 4033 3587 4047
rect 4553 4093 4567 4107
rect 4553 4033 4567 4047
rect 4533 3953 4547 3967
rect 4833 4113 4847 4127
rect 4833 3973 4847 3987
rect 6053 4113 6067 4127
rect 5913 4093 5927 4107
rect 5773 4053 5787 4067
rect 5613 3973 5627 3987
rect 6373 3993 6387 4007
rect 5913 3953 5927 3967
rect 6053 3953 6067 3967
rect 1274 3933 1288 3947
rect 2453 3933 2467 3947
rect 2673 3933 2687 3947
rect 3573 3933 3587 3947
rect 3713 3933 3727 3947
rect 4672 3933 4686 3947
rect 5592 3933 5606 3947
rect 5614 3933 5628 3947
rect 5774 3933 5788 3947
rect 2312 3873 2326 3887
rect 4914 3873 4928 3887
rect 653 3853 667 3867
rect 2332 3853 2346 3867
rect 2354 3853 2368 3867
rect 3133 3853 3147 3867
rect 4733 3853 4747 3867
rect 333 3813 347 3827
rect 492 3813 506 3827
rect 653 3813 667 3827
rect 2313 3813 2327 3827
rect 493 3693 507 3707
rect 2473 3813 2487 3827
rect 4593 3793 4607 3807
rect 4573 3753 4587 3767
rect 3133 3733 3147 3747
rect 2473 3713 2487 3727
rect 4734 3753 4748 3767
rect 4592 3713 4606 3727
rect 5033 3853 5047 3867
rect 5674 3853 5688 3867
rect 5713 3853 5727 3867
rect 6393 3853 6407 3867
rect 5553 3813 5567 3827
rect 5673 3813 5687 3827
rect 5033 3773 5047 3787
rect 5693 3773 5707 3787
rect 5553 3713 5567 3727
rect 4913 3693 4927 3707
rect 6013 3833 6027 3847
rect 6393 3753 6407 3767
rect 6013 3713 6027 3727
rect 5713 3693 5727 3707
rect 333 3673 347 3687
rect 2312 3673 2326 3687
rect 2334 3673 2348 3687
rect 4572 3673 4586 3687
rect 5693 3673 5707 3687
rect 853 3613 867 3627
rect 2113 3613 2127 3627
rect 3233 3613 3247 3627
rect 833 3573 847 3587
rect 833 3473 847 3487
rect 1613 3573 1627 3587
rect 2513 3593 2527 3607
rect 2493 3553 2507 3567
rect 1613 3473 1627 3487
rect 2113 3473 2127 3487
rect 2493 3453 2507 3467
rect 5734 3593 5748 3607
rect 4773 3573 4787 3587
rect 5593 3573 5607 3587
rect 3233 3533 3247 3547
rect 3353 3473 3367 3487
rect 2513 3433 2527 3447
rect 4773 3433 4787 3447
rect 5953 3573 5967 3587
rect 5753 3533 5767 3547
rect 6293 3533 6307 3547
rect 5753 3433 5767 3447
rect 5953 3433 5967 3447
rect 853 3413 867 3427
rect 3353 3413 3367 3427
rect 5593 3413 5607 3427
rect 5733 3413 5747 3427
rect 6294 3413 6308 3427
rect 2172 3353 2186 3367
rect 2194 3353 2208 3367
rect 2333 3353 2347 3367
rect 3774 3353 3788 3367
rect 4053 3353 4067 3367
rect 4173 3353 4187 3367
rect 4633 3353 4647 3367
rect 5052 3353 5066 3367
rect 5072 3353 5086 3367
rect 973 3333 987 3347
rect 953 3313 967 3327
rect 673 3213 687 3227
rect 673 3173 687 3187
rect 2173 3253 2187 3267
rect 973 3213 987 3227
rect 2193 3193 2207 3207
rect 2353 3293 2367 3307
rect 2533 3293 2547 3307
rect 4052 3267 4066 3281
rect 2353 3193 2367 3207
rect 2533 3193 2547 3207
rect 3773 3193 3787 3207
rect 2333 3173 2347 3187
rect 4514 3253 4528 3267
rect 4833 3333 4847 3347
rect 4833 3293 4847 3307
rect 4613 3213 4627 3227
rect 4533 3193 4547 3207
rect 5053 3173 5067 3187
rect 5893 3352 5907 3366
rect 6413 3353 6427 3367
rect 5233 3333 5247 3347
rect 5853 3293 5867 3307
rect 5233 3193 5247 3207
rect 6194 3293 6208 3307
rect 5893 3173 5907 3187
rect 6393 3253 6407 3267
rect 953 3153 967 3167
rect 4173 3153 4187 3167
rect 5073 3153 5087 3167
rect 5853 3153 5867 3167
rect 6193 3153 6207 3167
rect 233 3093 247 3107
rect 2213 3093 2227 3107
rect 2512 3093 2526 3107
rect 4513 3093 4527 3107
rect 4693 3093 4707 3107
rect 4993 3093 5007 3107
rect 6453 3093 6467 3107
rect 6494 3093 6508 3107
rect 2193 3073 2207 3087
rect 2193 3013 2207 3027
rect 233 2953 247 2967
rect 2213 2953 2227 2967
rect 2713 3033 2727 3047
rect 2533 3013 2547 3027
rect 4653 3013 4667 3027
rect 4833 3013 4847 3027
rect 5473 3073 5487 3087
rect 5793 3073 5807 3087
rect 6133 3073 6147 3087
rect 6293 3073 6307 3087
rect 4853 2953 4867 2967
rect 4993 2953 5007 2967
rect 5153 2953 5167 2967
rect 5473 2953 5487 2967
rect 4653 2913 4667 2927
rect 4693 2913 4707 2927
rect 4833 2913 4847 2927
rect 5973 3053 5987 3067
rect 5793 2913 5807 2927
rect 6153 3053 6167 3067
rect 6493 2973 6507 2987
rect 2512 2893 2526 2907
rect 2553 2893 2567 2907
rect 2713 2893 2727 2907
rect 4513 2893 4527 2907
rect 4852 2893 4866 2907
rect 5153 2893 5167 2907
rect 5973 2893 5987 2907
rect 6113 2893 6127 2907
rect 6154 2893 6168 2907
rect 6293 2893 6307 2907
rect 6453 2893 6467 2907
rect 2253 2833 2267 2847
rect 2693 2833 2707 2847
rect 4474 2833 4488 2847
rect 5013 2833 5027 2847
rect 613 2813 627 2827
rect 753 2793 767 2807
rect 1172 2773 1186 2787
rect 753 2733 767 2747
rect 313 2713 327 2727
rect 613 2713 627 2727
rect 313 2673 327 2687
rect 2393 2773 2407 2787
rect 2253 2713 2267 2727
rect 2393 2673 2407 2687
rect 3513 2813 3527 2827
rect 4733 2813 4747 2827
rect 4893 2813 4907 2827
rect 4473 2773 4487 2787
rect 4133 2733 4147 2747
rect 3513 2673 3527 2687
rect 4873 2773 4887 2787
rect 4853 2733 4867 2747
rect 4433 2713 4447 2727
rect 4733 2713 4747 2727
rect 4454 2673 4468 2687
rect 4853 2673 4867 2687
rect 1173 2653 1187 2667
rect 2693 2653 2707 2667
rect 4133 2653 4147 2667
rect 5393 2813 5407 2827
rect 5573 2813 5587 2827
rect 4893 2673 4907 2687
rect 5393 2733 5407 2747
rect 5033 2653 5047 2667
rect 4873 2633 4887 2647
rect 5573 2633 5587 2647
rect 973 2573 987 2587
rect 2393 2573 2407 2587
rect 2434 2573 2448 2587
rect 2553 2573 2567 2587
rect 3734 2573 3748 2587
rect 4033 2573 4047 2587
rect 4213 2573 4227 2587
rect 4453 2573 4467 2587
rect 4733 2573 4747 2587
rect 5093 2573 5107 2587
rect 5133 2573 5147 2587
rect 5413 2573 5427 2587
rect 6293 2573 6307 2587
rect 813 2473 827 2487
rect 353 2433 367 2447
rect 352 2393 366 2407
rect 2133 2553 2147 2567
rect 973 2433 987 2447
rect 2393 2493 2407 2507
rect 3193 2553 3207 2567
rect 2553 2513 2567 2527
rect 2433 2453 2447 2467
rect 2413 2433 2427 2447
rect 2133 2413 2147 2427
rect 3554 2533 3568 2547
rect 3594 2533 3608 2547
rect 3454 2493 3468 2507
rect 3473 2433 3487 2447
rect 2413 2393 2427 2407
rect 3193 2393 3207 2407
rect 3453 2393 3467 2407
rect 3592 2433 3606 2447
rect 3753 2513 3767 2527
rect 3733 2413 3747 2427
rect 3572 2393 3586 2407
rect 4033 2433 4047 2447
rect 4313 2533 4327 2547
rect 4734 2533 4748 2547
rect 4913 2533 4927 2547
rect 5113 2513 5127 2527
rect 5113 2453 5127 2467
rect 5093 2433 5107 2447
rect 6153 2553 6167 2567
rect 5413 2433 5427 2447
rect 4914 2413 4928 2427
rect 5133 2413 5147 2427
rect 6293 2433 6307 2447
rect 813 2373 827 2387
rect 3473 2373 3487 2387
rect 3753 2373 3767 2387
rect 4213 2373 4227 2387
rect 4313 2373 4327 2387
rect 4453 2373 4467 2387
rect 6153 2373 6167 2387
rect 3973 2313 3987 2327
rect 3653 2293 3667 2307
rect 3433 2273 3447 2287
rect 1713 2253 1727 2267
rect 1393 2153 1407 2167
rect 3093 2213 3107 2227
rect 3453 2253 3467 2267
rect 1713 2133 1727 2147
rect 3093 2133 3107 2147
rect 3433 2133 3447 2147
rect 4113 2253 4127 2267
rect 4893 2253 4907 2267
rect 6253 2253 6267 2267
rect 4133 2213 4147 2227
rect 4113 2173 4127 2187
rect 4453 2193 4467 2207
rect 3653 2133 3667 2147
rect 3993 2133 4007 2147
rect 4133 2133 4147 2147
rect 4453 2133 4467 2147
rect 5473 2193 5487 2207
rect 6253 2153 6267 2167
rect 1393 2113 1407 2127
rect 3452 2113 3466 2127
rect 4893 2113 4907 2127
rect 5473 2113 5487 2127
rect 2593 2053 2607 2067
rect 2732 2053 2746 2067
rect 4173 2053 4187 2067
rect 4413 2053 4427 2067
rect 5072 2053 5086 2067
rect 5253 2053 5267 2067
rect 5493 2053 5507 2067
rect 2573 1993 2587 2007
rect 193 1973 207 1987
rect 1733 1933 1747 1947
rect 193 1873 207 1887
rect 1733 1873 1747 1887
rect 2573 1873 2587 1887
rect 2853 2033 2867 2047
rect 4033 2033 4047 2047
rect 2853 1993 2867 2007
rect 2733 1933 2747 1947
rect 3253 1933 3267 1947
rect 3693 1933 3707 1947
rect 3693 1873 3707 1887
rect 4013 1873 4027 1887
rect 4313 1953 4327 1967
rect 4173 1933 4187 1947
rect 4573 2033 4587 2047
rect 4752 2033 4766 2047
rect 4553 1913 4567 1927
rect 4413 1873 4427 1887
rect 5053 2013 5067 2027
rect 5053 1953 5067 1967
rect 4753 1933 4767 1947
rect 4573 1893 4587 1907
rect 5233 2013 5247 2027
rect 5213 1953 5227 1967
rect 5073 1873 5087 1887
rect 5213 1873 5227 1887
rect 5494 2013 5508 2027
rect 6113 1996 6127 2010
rect 5253 1953 5267 1967
rect 6113 1950 6127 1964
rect 2593 1853 2607 1867
rect 3253 1853 3267 1867
rect 3993 1853 4007 1867
rect 4033 1853 4047 1867
rect 4314 1853 4328 1867
rect 4553 1853 4567 1867
rect 5233 1853 5247 1867
rect 193 1793 207 1807
rect 1693 1793 1707 1807
rect 2053 1793 2067 1807
rect 2173 1793 2187 1807
rect 3112 1793 3126 1807
rect 3753 1793 3767 1807
rect 5073 1793 5087 1807
rect 6193 1793 6207 1807
rect 1373 1773 1387 1787
rect 1553 1773 1567 1787
rect 193 1733 207 1747
rect 1333 1653 1347 1667
rect 1373 1633 1387 1647
rect 1714 1773 1728 1787
rect 1853 1773 1867 1787
rect 1693 1673 1707 1687
rect 1713 1613 1727 1627
rect 1853 1613 1867 1627
rect 2214 1773 2228 1787
rect 2633 1773 2647 1787
rect 3133 1773 3147 1787
rect 3253 1773 3267 1787
rect 3293 1773 3307 1787
rect 3573 1773 3587 1787
rect 2213 1673 2227 1687
rect 2172 1633 2186 1647
rect 3393 1753 3407 1767
rect 2833 1733 2847 1747
rect 2853 1693 2867 1707
rect 2833 1673 2847 1687
rect 2873 1633 2887 1647
rect 2853 1613 2867 1627
rect 3733 1733 3747 1747
rect 3573 1613 3587 1627
rect 3873 1773 3887 1787
rect 3913 1773 3927 1787
rect 4253 1773 4267 1787
rect 3873 1733 3887 1747
rect 4033 1673 4047 1687
rect 4553 1753 4567 1767
rect 4273 1733 4287 1747
rect 4413 1739 4427 1753
rect 4253 1653 4267 1667
rect 4532 1733 4546 1747
rect 6493 1773 6507 1787
rect 5553 1733 5567 1747
rect 6193 1733 6207 1747
rect 4413 1653 4427 1667
rect 5073 1653 5087 1667
rect 4273 1633 4287 1647
rect 3753 1613 3767 1627
rect 3913 1613 3927 1627
rect 4053 1613 4067 1627
rect 6493 1633 6507 1647
rect 1333 1593 1347 1607
rect 1533 1593 1547 1607
rect 2053 1593 2067 1607
rect 2632 1593 2646 1607
rect 2873 1593 2887 1607
rect 3413 1593 3427 1607
rect 3733 1593 3747 1607
rect 5553 1593 5567 1607
rect 1273 1533 1287 1547
rect 1713 1533 1727 1547
rect 4612 1533 4626 1547
rect 5613 1533 5627 1547
rect 192 1513 206 1527
rect 373 1513 387 1527
rect 173 1473 187 1487
rect 172 1353 186 1367
rect 374 1393 388 1407
rect 2933 1513 2947 1527
rect 3652 1513 3666 1527
rect 3793 1513 3807 1527
rect 4153 1513 4167 1527
rect 1713 1493 1727 1507
rect 2473 1473 2487 1487
rect 2933 1453 2947 1467
rect 3233 1453 3247 1467
rect 3633 1453 3647 1467
rect 2613 1373 2627 1387
rect 2473 1353 2487 1367
rect 3393 1413 3407 1427
rect 3373 1373 3387 1387
rect 3233 1353 3247 1367
rect 3773 1493 3787 1507
rect 3773 1433 3787 1447
rect 3653 1413 3667 1427
rect 3633 1353 3647 1367
rect 4153 1373 4167 1387
rect 4993 1513 5007 1527
rect 5313 1493 5327 1507
rect 4993 1393 5007 1407
rect 5333 1413 5347 1427
rect 5293 1373 5307 1387
rect 5334 1373 5348 1387
rect 5633 1513 5647 1527
rect 5633 1413 5647 1427
rect 5653 1393 5667 1407
rect 5653 1353 5667 1367
rect 194 1333 208 1347
rect 1273 1333 1287 1347
rect 2613 1333 2627 1347
rect 3372 1333 3386 1347
rect 3394 1333 3408 1347
rect 3793 1333 3807 1347
rect 4613 1333 4627 1347
rect 5613 1333 5627 1347
rect 2733 1273 2747 1287
rect 4193 1273 4207 1287
rect 4373 1273 4387 1287
rect 4953 1273 4967 1287
rect 5472 1273 5486 1287
rect 213 1253 227 1267
rect 2553 1253 2567 1267
rect 2713 1253 2727 1267
rect 953 1213 967 1227
rect 533 1153 547 1167
rect 213 1133 227 1147
rect 512 1113 526 1127
rect 2734 1213 2748 1227
rect 2834 1213 2848 1227
rect 3133 1213 3147 1227
rect 2554 1113 2568 1127
rect 2713 1113 2727 1127
rect 953 1093 967 1107
rect 4353 1253 4367 1267
rect 4312 1213 4326 1227
rect 4353 1133 4367 1147
rect 4334 1113 4348 1127
rect 5313 1253 5327 1267
rect 4973 1113 4987 1127
rect 5453 1213 5467 1227
rect 3133 1093 3147 1107
rect 4193 1093 4207 1107
rect 4373 1093 4387 1107
rect 5313 1093 5327 1107
rect 5473 1093 5487 1107
rect 5673 1213 5687 1227
rect 2833 1073 2847 1087
rect 5452 1073 5466 1087
rect 5633 1073 5647 1087
rect 3293 1013 3307 1027
rect 3433 1013 3447 1027
rect 1733 993 1747 1007
rect 2333 993 2347 1007
rect 3273 993 3287 1007
rect 653 973 667 987
rect 512 873 526 887
rect 1273 933 1287 947
rect 1733 853 1747 867
rect 513 833 527 847
rect 653 833 667 847
rect 1273 833 1287 847
rect 3253 973 3267 987
rect 3093 933 3107 947
rect 3254 873 3268 887
rect 3293 973 3307 987
rect 3413 873 3427 887
rect 4212 993 4226 1007
rect 4673 993 4687 1007
rect 4353 973 4367 987
rect 5613 973 5627 987
rect 4693 913 4707 927
rect 5813 959 5827 973
rect 4373 833 4387 847
rect 4673 833 4687 847
rect 5633 873 5647 887
rect 5813 853 5827 867
rect 2333 813 2347 827
rect 3093 813 3107 827
rect 3273 813 3287 827
rect 3412 813 3426 827
rect 3434 813 3448 827
rect 4213 813 4227 827
rect 4694 813 4708 827
rect 953 753 967 767
rect 3293 753 3307 767
rect 4213 753 4227 767
rect 4913 753 4927 767
rect 813 733 827 747
rect 473 693 487 707
rect 813 613 827 627
rect 473 593 487 607
rect 2753 733 2767 747
rect 3273 733 3287 747
rect 1973 693 1987 707
rect 2133 693 2147 707
rect 953 573 967 587
rect 2933 693 2947 707
rect 3433 733 3447 747
rect 3292 653 3306 667
rect 3314 653 3328 667
rect 3273 613 3287 627
rect 2933 573 2947 587
rect 3634 693 3648 707
rect 3433 613 3447 627
rect 5773 733 5787 747
rect 4393 693 4407 707
rect 4573 693 4587 707
rect 4913 693 4927 707
rect 5053 693 5067 707
rect 5213 693 5227 707
rect 5773 693 5787 707
rect 4393 573 4407 587
rect 4573 573 4587 587
rect 5413 633 5427 647
rect 5213 593 5227 607
rect 5593 573 5607 587
rect 1973 553 1987 567
rect 2133 553 2147 567
rect 2753 553 2767 567
rect 3313 553 3327 567
rect 3613 553 3627 567
rect 4213 553 4227 567
rect 5053 553 5067 567
rect 5413 553 5427 567
rect 5573 553 5587 567
rect 813 493 827 507
rect 1773 493 1787 507
rect 3314 493 3328 507
rect 3513 493 3527 507
rect 3832 493 3846 507
rect 3854 493 3868 507
rect 4034 493 4048 507
rect 974 453 988 467
rect 833 433 847 447
rect 833 373 847 387
rect 993 333 1007 347
rect 3093 473 3107 487
rect 3313 453 3327 467
rect 3093 393 3107 407
rect 3513 353 3527 367
rect 813 313 827 327
rect 1773 313 1787 327
rect 4214 473 4228 487
rect 5613 473 5627 487
rect 3873 333 3887 347
rect 4033 333 4047 347
rect 5493 453 5507 467
rect 5493 313 5507 327
rect 5993 453 6007 467
rect 5993 313 6007 327
rect 3833 293 3847 307
rect 4213 293 4227 307
rect 5613 293 5627 307
rect 714 233 728 247
rect 1333 233 1347 247
rect 2293 233 2307 247
rect 3873 233 3887 247
rect 6193 233 6207 247
rect 353 213 367 227
rect 692 213 706 227
rect 212 173 226 187
rect 213 73 227 87
rect 373 173 387 187
rect 373 133 387 147
rect 673 133 687 147
rect 673 73 687 87
rect 353 53 367 67
rect 854 213 868 227
rect 1153 213 1167 227
rect 1033 173 1047 187
rect 713 73 727 87
rect 853 73 867 87
rect 1033 73 1047 87
rect 1193 173 1207 187
rect 2153 213 2167 227
rect 1333 73 1347 87
rect 1193 53 1207 67
rect 3533 213 3547 227
rect 3213 173 3227 187
rect 3033 153 3047 167
rect 2293 73 2307 87
rect 3713 193 3727 207
rect 3693 173 3707 187
rect 3533 113 3547 127
rect 3213 73 3227 87
rect 3713 133 3727 147
rect 4933 213 4947 227
rect 3893 153 3907 167
rect 3873 113 3887 127
rect 3893 73 3907 87
rect 6033 173 6047 187
rect 6213 173 6227 187
rect 6193 113 6207 127
rect 6213 73 6227 87
rect 3693 53 3707 67
rect 4933 53 4947 67
rect 6033 53 6047 67
rect 693 33 707 47
rect 1153 33 1167 47
rect 2153 33 2167 47
rect 3032 33 3046 47
<< metal2 >>
rect 1067 6516 2293 6523
rect 2596 6516 3933 6523
rect 1507 6496 1693 6503
rect 2596 6503 2603 6516
rect 3987 6516 4013 6523
rect 6247 6516 6273 6523
rect 1867 6496 2603 6503
rect 2767 6496 2933 6503
rect 3267 6496 3413 6503
rect 5267 6496 5693 6503
rect 367 6476 553 6483
rect 567 6476 693 6483
rect 947 6476 1093 6483
rect 1296 6476 2093 6483
rect 436 6456 593 6463
rect 436 6427 443 6456
rect 607 6456 733 6463
rect 1296 6463 1303 6476
rect 2267 6476 2293 6483
rect 2307 6476 2613 6483
rect 2827 6476 2853 6483
rect 3187 6476 3573 6483
rect 4647 6476 4753 6483
rect 5867 6476 5933 6483
rect 5947 6476 5983 6483
rect 987 6456 1303 6463
rect 1176 6427 1183 6456
rect 1327 6456 1533 6463
rect 1547 6456 2213 6463
rect 2407 6456 2723 6463
rect 1493 6427 1507 6433
rect 2147 6436 2253 6443
rect 1853 6427 1867 6433
rect 2716 6427 2723 6456
rect 3547 6456 3653 6463
rect 3667 6456 3753 6463
rect 4687 6456 4713 6463
rect 5976 6447 5983 6476
rect 6027 6456 6073 6463
rect 6387 6456 6473 6463
rect 3327 6433 3333 6447
rect 5007 6436 5103 6443
rect 267 6416 353 6423
rect 607 6416 673 6423
rect 786 6413 792 6427
rect 828 6416 893 6423
rect 1047 6413 1053 6427
rect 1287 6416 1333 6423
rect 1587 6416 1653 6423
rect 1747 6416 1853 6423
rect 1907 6416 1973 6423
rect 2347 6416 2413 6423
rect 2567 6416 2673 6423
rect 3427 6416 3493 6423
rect 3587 6416 3673 6423
rect 3987 6413 3993 6427
rect 4807 6416 4913 6423
rect 5096 6407 5103 6436
rect 5567 6413 5573 6427
rect 6107 6416 6153 6423
rect 6440 6423 6453 6427
rect 6427 6416 6453 6423
rect 6440 6413 6453 6416
rect 5096 6396 5113 6407
rect 5100 6393 5113 6396
rect 5387 6393 5393 6407
rect 2287 6376 2353 6383
rect 2787 6376 2873 6383
rect 4247 6373 4253 6387
rect 4267 6376 4313 6383
rect 4400 6383 4413 6387
rect 4387 6376 4413 6383
rect 4400 6373 4413 6376
rect 5967 6376 6013 6383
rect 6207 6383 6220 6387
rect 6207 6376 6233 6383
rect 6207 6373 6220 6376
rect 3193 6367 3207 6373
rect 127 6356 193 6363
rect 1007 6356 1053 6363
rect 3060 6363 3073 6367
rect 2947 6356 3033 6363
rect 3047 6356 3073 6363
rect 3060 6353 3073 6356
rect 2507 6333 2513 6347
rect 2847 6336 2893 6343
rect 3087 6336 3213 6343
rect 3356 6343 3363 6373
rect 3767 6356 3833 6363
rect 5440 6363 5453 6367
rect 5427 6356 5453 6363
rect 5440 6353 5453 6356
rect 5827 6353 5833 6367
rect 6127 6356 6173 6363
rect 6033 6347 6047 6353
rect 6113 6347 6127 6353
rect 3227 6336 3363 6343
rect 3387 6336 3413 6343
rect 6033 6340 6053 6347
rect 6036 6336 6053 6340
rect 6040 6333 6053 6336
rect 147 6316 373 6323
rect 387 6316 513 6323
rect 527 6316 1273 6323
rect 1287 6316 1473 6323
rect 1687 6316 1833 6323
rect 1847 6316 2333 6323
rect 2507 6316 2533 6323
rect 2627 6316 2712 6323
rect 2748 6316 2773 6323
rect 3707 6316 3993 6323
rect 4907 6316 4953 6323
rect 5407 6316 5553 6323
rect 5687 6316 6153 6323
rect 3073 6307 3087 6313
rect 927 6296 993 6303
rect 1107 6296 1213 6303
rect 1387 6296 1753 6303
rect 2507 6296 2813 6303
rect 4027 6296 4353 6303
rect 4747 6296 4933 6303
rect 4947 6296 5093 6303
rect 5827 6296 5933 6303
rect 747 6276 813 6283
rect 1207 6276 1573 6283
rect 1756 6283 1763 6293
rect 1756 6276 2493 6283
rect 2516 6276 3193 6283
rect 687 6256 1033 6263
rect 1347 6256 1593 6263
rect 1887 6256 1953 6263
rect 2516 6263 2523 6276
rect 4127 6276 4473 6283
rect 4487 6276 4672 6283
rect 4696 6276 4993 6283
rect 4696 6267 4703 6276
rect 5227 6276 5473 6283
rect 1967 6256 2523 6263
rect 2827 6256 3813 6263
rect 4247 6256 4693 6263
rect 4887 6256 5053 6263
rect 5067 6256 5653 6263
rect 5847 6256 6253 6263
rect 6267 6256 6333 6263
rect 427 6236 473 6243
rect 487 6236 1153 6243
rect 1167 6236 1473 6243
rect 1567 6236 1733 6243
rect 1756 6240 2543 6243
rect 1756 6236 2547 6240
rect 247 6216 1253 6223
rect 1367 6216 1513 6223
rect 1756 6223 1763 6236
rect 2533 6227 2547 6236
rect 2707 6236 2753 6243
rect 2887 6236 3173 6243
rect 3187 6236 4433 6243
rect 4447 6236 4953 6243
rect 5007 6236 5113 6243
rect 5187 6236 5913 6243
rect 5927 6236 6313 6243
rect 1527 6216 1763 6223
rect 1787 6216 2512 6223
rect 2533 6220 2534 6227
rect 2587 6216 2833 6223
rect 2847 6216 3153 6223
rect 3167 6216 3633 6223
rect 3787 6216 4093 6223
rect 4427 6216 4593 6223
rect 4607 6216 4873 6223
rect 5047 6216 5148 6223
rect 5184 6213 5193 6227
rect 5247 6216 5293 6223
rect 5307 6216 5393 6223
rect 287 6196 613 6203
rect 1227 6196 1553 6203
rect 1967 6196 2013 6203
rect 2367 6196 2993 6203
rect 3056 6196 3373 6203
rect 3056 6187 3063 6196
rect 3427 6196 3473 6203
rect 3867 6196 3913 6203
rect 5331 6193 5333 6207
rect 5887 6196 6193 6203
rect 367 6176 393 6183
rect 407 6176 1013 6183
rect 1267 6176 1293 6183
rect 1407 6176 1513 6183
rect 1727 6176 1833 6183
rect 1847 6176 1993 6183
rect 2007 6176 2553 6183
rect 2576 6176 2613 6183
rect 687 6156 853 6163
rect 2576 6163 2583 6176
rect 2747 6176 3053 6183
rect 3327 6176 3453 6183
rect 3587 6176 3692 6183
rect 3728 6176 3873 6183
rect 3887 6176 4033 6183
rect 4047 6176 4073 6183
rect 4587 6176 4763 6183
rect 2376 6156 2583 6163
rect 107 6136 153 6143
rect 273 6143 287 6153
rect 2376 6147 2383 6156
rect 4107 6156 4233 6163
rect 4756 6147 4763 6176
rect 6107 6176 6183 6183
rect 6116 6156 6153 6163
rect 227 6136 263 6143
rect 273 6140 353 6143
rect 276 6136 353 6140
rect 256 6123 263 6136
rect 2087 6133 2093 6147
rect 2327 6136 2373 6143
rect 3487 6133 3493 6147
rect 3507 6143 3520 6147
rect 3507 6136 3533 6143
rect 3507 6133 3520 6136
rect 3627 6136 3693 6143
rect 6047 6133 6053 6147
rect 6116 6143 6123 6156
rect 6176 6163 6183 6176
rect 6176 6156 6203 6163
rect 6067 6136 6123 6143
rect 6196 6127 6203 6156
rect 6247 6156 6283 6163
rect 6276 6143 6283 6156
rect 6276 6136 6333 6143
rect 256 6116 293 6123
rect 807 6116 853 6123
rect 1307 6116 1373 6123
rect 1607 6116 1693 6123
rect 2107 6116 2153 6123
rect 2467 6113 2473 6127
rect 3127 6116 3193 6123
rect 4087 6116 4173 6123
rect 1587 6096 1653 6103
rect 1747 6103 1760 6107
rect 1747 6093 1763 6103
rect 5187 6093 5193 6107
rect 507 6076 573 6083
rect 667 6073 673 6087
rect 1027 6076 1073 6083
rect 1127 6076 1213 6083
rect 1227 6073 1233 6087
rect 1473 6083 1487 6093
rect 1756 6083 1763 6093
rect 1473 6080 1533 6083
rect 1476 6076 1533 6080
rect 1756 6076 1853 6083
rect 1967 6076 2013 6083
rect 2587 6076 2633 6083
rect 2747 6076 2793 6083
rect 3307 6076 3393 6083
rect 3487 6076 3553 6083
rect 3827 6073 3833 6087
rect 3927 6076 4013 6083
rect 4207 6073 4213 6087
rect 4487 6076 4553 6083
rect 4647 6076 4733 6083
rect 1447 6056 1493 6063
rect 1576 6056 1673 6063
rect 127 6036 353 6043
rect 867 6036 943 6043
rect 787 6016 913 6023
rect 936 6023 943 6036
rect 987 6036 1033 6043
rect 1576 6043 1583 6056
rect 2107 6063 2120 6067
rect 2107 6056 2133 6063
rect 2107 6053 2120 6056
rect 2187 6056 2263 6063
rect 1407 6036 1583 6043
rect 1907 6036 2093 6043
rect 2256 6043 2263 6056
rect 2256 6036 2393 6043
rect 2547 6036 2753 6043
rect 3256 6043 3263 6073
rect 4447 6063 4460 6067
rect 4447 6053 4463 6063
rect 2967 6036 3263 6043
rect 3787 6036 3853 6043
rect 3907 6036 4053 6043
rect 4067 6036 4233 6043
rect 4456 6043 4463 6053
rect 4596 6043 4603 6073
rect 5187 6056 5333 6063
rect 5716 6063 5723 6093
rect 6527 6076 6563 6083
rect 5607 6056 5723 6063
rect 4456 6036 4603 6043
rect 5896 6043 5903 6073
rect 5647 6036 5903 6043
rect 936 6016 963 6023
rect 687 5996 873 6003
rect 887 5996 933 6003
rect 956 6003 963 6016
rect 1327 6016 3213 6023
rect 3407 6016 3473 6023
rect 3947 6016 4013 6023
rect 5207 6016 5293 6023
rect 5947 6016 6213 6023
rect 956 5996 993 6003
rect 1013 6003 1027 6013
rect 1013 6000 1293 6003
rect 1016 5996 1293 6000
rect 1687 5996 1793 6003
rect 2067 5996 2153 6003
rect 2227 5996 2313 6003
rect 2387 5996 2433 6003
rect 2527 5996 3273 6003
rect 3496 5996 4473 6003
rect 867 5976 1093 5983
rect 1227 5976 2013 5983
rect 2147 5976 2293 5983
rect 2307 5976 2423 5983
rect 187 5956 233 5963
rect 247 5956 1772 5963
rect 1808 5956 2113 5963
rect 2207 5956 2393 5963
rect 2416 5963 2423 5976
rect 2507 5976 2573 5983
rect 2596 5976 2783 5983
rect 2416 5956 2452 5963
rect 2596 5963 2603 5976
rect 2488 5956 2603 5963
rect 2727 5956 2753 5963
rect 2776 5963 2783 5976
rect 3496 5983 3503 5996
rect 4767 5996 5173 6003
rect 5187 5996 5853 6003
rect 5867 5996 6013 6003
rect 3267 5976 3503 5983
rect 3976 5976 4193 5983
rect 2776 5956 3133 5963
rect 3976 5963 3983 5976
rect 4207 5976 4853 5983
rect 4936 5976 4993 5983
rect 3147 5956 3983 5963
rect 4147 5956 4253 5963
rect 4936 5963 4943 5976
rect 5047 5976 5073 5983
rect 5127 5976 5153 5983
rect 5467 5976 5893 5983
rect 6187 5976 6313 5983
rect 4487 5956 4943 5963
rect 5293 5967 5307 5973
rect 4967 5956 5193 5963
rect 5293 5960 5313 5967
rect 5296 5956 5313 5960
rect 5300 5953 5313 5956
rect 5447 5956 5553 5963
rect 5567 5956 5593 5963
rect 5787 5956 6053 5963
rect 116 5936 473 5943
rect 116 5907 123 5936
rect 687 5936 813 5943
rect 987 5936 1053 5943
rect 1267 5936 1353 5943
rect 1367 5936 1543 5943
rect 1536 5907 1543 5936
rect 1576 5936 1753 5943
rect 1576 5907 1583 5936
rect 2327 5936 2353 5943
rect 2827 5936 3023 5943
rect 2393 5907 2407 5913
rect 2553 5907 2567 5913
rect 3016 5907 3023 5936
rect 3047 5936 3173 5943
rect 3447 5936 3473 5943
rect 3527 5936 3963 5943
rect 3847 5916 3893 5923
rect 3633 5907 3647 5913
rect 3956 5907 3963 5936
rect 4247 5936 4273 5943
rect 4287 5936 4513 5943
rect 4587 5936 4953 5943
rect 4996 5936 5133 5943
rect 4253 5907 4267 5913
rect 4996 5907 5003 5936
rect 5147 5936 5253 5943
rect 5587 5936 5633 5943
rect 6027 5936 6113 5943
rect 6227 5936 6253 5943
rect 267 5896 313 5903
rect 607 5903 620 5907
rect 607 5896 633 5903
rect 607 5893 620 5896
rect 987 5896 1033 5903
rect 1307 5896 1373 5903
rect 1627 5896 1673 5903
rect 1887 5896 1933 5903
rect 2767 5896 2813 5903
rect 3507 5896 3553 5903
rect 3727 5896 3773 5903
rect 4007 5896 4093 5903
rect 4647 5903 4660 5907
rect 4647 5896 4673 5903
rect 4647 5893 4660 5896
rect 4767 5903 4780 5907
rect 4767 5896 4793 5903
rect 4767 5893 4780 5896
rect 5627 5896 5733 5903
rect 5827 5903 5840 5907
rect 5827 5896 5853 5903
rect 5827 5893 5840 5896
rect 6067 5896 6173 5903
rect 1036 5883 1043 5893
rect 1036 5876 1073 5883
rect 3567 5873 3573 5887
rect 2067 5853 2073 5867
rect 2127 5856 2213 5863
rect 2300 5863 2313 5867
rect 2287 5856 2313 5863
rect 2300 5853 2313 5856
rect 3167 5853 3173 5867
rect 3287 5856 3333 5863
rect 4847 5856 4912 5863
rect 4948 5853 4953 5867
rect 5160 5863 5173 5867
rect 5147 5856 5173 5863
rect 5160 5853 5173 5856
rect 5327 5856 5413 5863
rect 5427 5856 5493 5863
rect 6267 5856 6313 5863
rect 493 5847 507 5853
rect 707 5836 773 5843
rect 1156 5836 1233 5843
rect 1156 5823 1163 5836
rect 1447 5836 1513 5843
rect 2627 5836 2693 5843
rect 3820 5843 3833 5847
rect 3807 5836 3833 5843
rect 3820 5833 3833 5836
rect 4467 5836 4533 5843
rect 6060 5843 6073 5847
rect 6047 5836 6073 5843
rect 6060 5833 6073 5836
rect 1007 5816 1163 5823
rect 2067 5816 2093 5823
rect 2287 5813 2293 5827
rect 2467 5816 2493 5823
rect 4867 5816 5193 5823
rect 5416 5816 5533 5823
rect 267 5796 433 5803
rect 747 5796 913 5803
rect 967 5796 1353 5803
rect 1427 5796 1553 5803
rect 1567 5796 1613 5803
rect 1907 5796 2373 5803
rect 2387 5796 2653 5803
rect 2667 5796 2993 5803
rect 3007 5796 3553 5803
rect 3667 5796 3713 5803
rect 3947 5796 4193 5803
rect 4447 5796 4572 5803
rect 4608 5796 4993 5803
rect 5416 5803 5423 5816
rect 5753 5823 5767 5833
rect 5753 5816 5813 5823
rect 5827 5816 5853 5823
rect 6267 5816 6473 5823
rect 5047 5796 5423 5803
rect 5447 5796 5472 5803
rect 5508 5796 5573 5803
rect 5827 5793 5833 5807
rect 6027 5796 6193 5803
rect 1127 5776 1233 5783
rect 1767 5776 1853 5783
rect 1867 5776 2143 5783
rect 2136 5767 2143 5776
rect 2247 5776 2292 5783
rect 2328 5776 2353 5783
rect 2467 5776 2532 5783
rect 2568 5776 2673 5783
rect 2687 5776 2733 5783
rect 2747 5776 2873 5783
rect 2887 5776 3093 5783
rect 3107 5776 3153 5783
rect 3227 5776 3463 5783
rect 107 5756 133 5763
rect 847 5756 953 5763
rect 976 5756 1313 5763
rect 976 5743 983 5756
rect 1707 5756 1933 5763
rect 2136 5756 2153 5767
rect 2140 5753 2153 5756
rect 2347 5756 2472 5763
rect 2508 5756 2613 5763
rect 2766 5753 2767 5760
rect 2788 5756 3233 5763
rect 3247 5756 3433 5763
rect 3456 5763 3463 5776
rect 3527 5776 4153 5783
rect 4847 5776 5183 5783
rect 3456 5756 3583 5763
rect 2293 5747 2307 5753
rect 27 5736 983 5743
rect 1027 5736 2233 5743
rect 2507 5736 2533 5743
rect 2753 5743 2767 5753
rect 2753 5740 2893 5743
rect 2755 5736 2893 5740
rect 2987 5736 3253 5743
rect 3367 5736 3553 5743
rect 3576 5743 3583 5756
rect 3807 5756 3873 5763
rect 3927 5756 4213 5763
rect 4606 5753 4607 5760
rect 4628 5756 4653 5763
rect 4787 5756 5113 5763
rect 5176 5763 5183 5776
rect 5207 5776 6513 5783
rect 5176 5756 5233 5763
rect 5247 5756 5292 5763
rect 5313 5753 5314 5760
rect 5367 5756 5713 5763
rect 5727 5756 5873 5763
rect 5887 5756 6053 5763
rect 6107 5756 6173 5763
rect 4593 5747 4607 5753
rect 3576 5736 3963 5743
rect 707 5716 1883 5723
rect 867 5696 973 5703
rect 1367 5693 1373 5707
rect 1527 5696 1853 5703
rect 1876 5703 1883 5716
rect 2187 5716 2573 5723
rect 3207 5716 3513 5723
rect 3556 5723 3563 5733
rect 3556 5716 3933 5723
rect 1876 5696 2593 5703
rect 2616 5696 2913 5703
rect 367 5676 1213 5683
rect 1587 5676 1673 5683
rect 1747 5676 1813 5683
rect 1827 5676 1993 5683
rect 2007 5676 2053 5683
rect 2067 5676 2353 5683
rect 2616 5683 2623 5696
rect 3187 5696 3433 5703
rect 3627 5696 3673 5703
rect 3736 5696 3853 5703
rect 2536 5676 2623 5683
rect 367 5656 413 5663
rect 667 5656 1053 5663
rect 1067 5656 1303 5663
rect 1013 5636 1113 5643
rect 1013 5627 1027 5636
rect 1296 5627 1303 5656
rect 1487 5656 1613 5663
rect 1627 5656 1693 5663
rect 2536 5663 2543 5676
rect 2847 5676 2903 5683
rect 2107 5656 2543 5663
rect 2587 5656 2873 5663
rect 2896 5663 2903 5676
rect 3167 5676 3313 5683
rect 3736 5687 3743 5696
rect 3907 5693 3913 5707
rect 3956 5703 3963 5736
rect 3987 5736 4133 5743
rect 4147 5736 4453 5743
rect 4606 5740 4607 5747
rect 4667 5736 4813 5743
rect 4887 5736 5123 5743
rect 4267 5716 4833 5723
rect 4896 5716 5093 5723
rect 3956 5696 4273 5703
rect 4627 5696 4753 5703
rect 4896 5703 4903 5716
rect 5116 5723 5123 5736
rect 5313 5743 5327 5753
rect 5227 5740 5327 5743
rect 5227 5736 5323 5740
rect 5927 5736 6093 5743
rect 5116 5716 5233 5723
rect 5367 5716 6513 5723
rect 4767 5696 4903 5703
rect 4947 5696 5333 5703
rect 5747 5693 5753 5707
rect 6427 5696 6493 5703
rect 6373 5687 6387 5693
rect 3327 5676 3343 5683
rect 2896 5656 3313 5663
rect 3336 5663 3343 5676
rect 3367 5676 3733 5683
rect 4567 5676 4673 5683
rect 4687 5676 4853 5683
rect 4867 5676 4913 5683
rect 3336 5656 3753 5663
rect 3767 5656 3893 5663
rect 4507 5656 4613 5663
rect 4727 5656 4873 5663
rect 4967 5656 5033 5663
rect 5356 5656 5413 5663
rect 2087 5636 2173 5643
rect 3347 5633 3353 5647
rect 3747 5636 3793 5643
rect 4067 5636 4173 5643
rect 4407 5636 4473 5643
rect 3553 5627 3567 5633
rect 5356 5627 5363 5656
rect 5427 5656 5453 5663
rect 5667 5656 5703 5663
rect 5696 5643 5703 5656
rect 5727 5656 6093 5663
rect 6227 5656 6343 5663
rect 6336 5643 6343 5656
rect 6367 5656 6453 5663
rect 5696 5636 5807 5643
rect 6336 5636 6393 5643
rect 5793 5627 5807 5636
rect 347 5616 373 5623
rect 607 5616 673 5623
rect 807 5616 853 5623
rect 867 5616 933 5623
rect 1867 5616 1913 5623
rect 3307 5616 3352 5623
rect 3388 5613 3393 5627
rect 3747 5616 3833 5623
rect 3847 5616 3893 5623
rect 5007 5613 5013 5627
rect 6320 5623 6333 5627
rect 6307 5616 6333 5623
rect 6320 5613 6333 5616
rect 3433 5607 3447 5613
rect 6373 5607 6387 5613
rect 1067 5596 1093 5603
rect 1867 5593 1873 5607
rect 2027 5596 2073 5603
rect 2367 5593 2373 5607
rect 4107 5593 4113 5607
rect 4420 5603 4433 5607
rect 4407 5596 4433 5603
rect 4420 5593 4433 5596
rect 6107 5603 6120 5607
rect 6107 5596 6133 5603
rect 6107 5593 6120 5596
rect 6527 5596 6563 5603
rect 2856 5576 2933 5583
rect 287 5556 352 5563
rect 388 5553 393 5567
rect 447 5556 533 5563
rect 747 5553 753 5567
rect 1367 5556 1433 5563
rect 1487 5556 1553 5563
rect 1660 5563 1672 5567
rect 1647 5556 1672 5563
rect 1660 5553 1672 5556
rect 1708 5556 1753 5563
rect 2260 5563 2273 5567
rect 2247 5556 2273 5563
rect 2260 5553 2273 5556
rect 2856 5563 2863 5576
rect 3367 5576 3393 5583
rect 3887 5576 3923 5583
rect 2827 5556 2863 5563
rect 2887 5556 2973 5563
rect 3067 5556 3153 5563
rect 3587 5556 3633 5563
rect 3727 5556 3813 5563
rect 3827 5556 3893 5563
rect 3916 5563 3923 5576
rect 5916 5576 5953 5583
rect 3916 5556 3953 5563
rect 4007 5556 4053 5563
rect 4427 5556 4533 5563
rect 4587 5553 4593 5567
rect 4667 5563 4680 5567
rect 4667 5556 4693 5563
rect 4667 5553 4680 5556
rect 4787 5556 4833 5563
rect 4887 5556 4893 5563
rect 4907 5556 4933 5563
rect 5687 5556 5733 5563
rect 5916 5563 5923 5576
rect 5827 5556 5923 5563
rect 5947 5556 5993 5563
rect 6327 5556 6393 5563
rect 6447 5556 6493 5563
rect 573 5547 587 5553
rect 147 5516 293 5523
rect 487 5516 713 5523
rect 996 5523 1003 5553
rect 1153 5547 1167 5553
rect 727 5516 1003 5523
rect 1327 5516 1413 5523
rect 1596 5523 1603 5553
rect 1427 5516 1603 5523
rect 1936 5523 1943 5553
rect 1787 5516 1943 5523
rect 2007 5513 2013 5527
rect 2247 5516 2433 5523
rect 2676 5523 2683 5553
rect 3673 5547 3687 5553
rect 2527 5516 2683 5523
rect 2707 5516 3073 5523
rect 167 5496 253 5503
rect 267 5496 333 5503
rect 627 5496 833 5503
rect 847 5496 1173 5503
rect 1187 5496 1333 5503
rect 1867 5496 2093 5503
rect 2696 5503 2703 5513
rect 3373 5507 3387 5513
rect 2547 5496 2703 5503
rect 3047 5496 3333 5503
rect 3707 5516 4053 5523
rect 4527 5516 4633 5523
rect 4736 5516 4853 5523
rect 3613 5507 3627 5513
rect 3907 5496 4093 5503
rect 4107 5496 4193 5503
rect 4627 5493 4632 5507
rect 4668 5496 4713 5503
rect 127 5476 573 5483
rect 587 5476 993 5483
rect 1447 5476 1473 5483
rect 1547 5476 1633 5483
rect 1647 5476 1993 5483
rect 2347 5476 2393 5483
rect 2447 5476 2733 5483
rect 3127 5476 3393 5483
rect 3467 5476 3493 5483
rect 3587 5476 3693 5483
rect 3887 5476 4093 5483
rect 4347 5476 4413 5483
rect 4736 5483 4743 5516
rect 5387 5516 5433 5523
rect 5587 5516 5633 5523
rect 5647 5516 5773 5523
rect 6047 5516 6073 5523
rect 6087 5516 6133 5523
rect 6436 5523 6443 5553
rect 6407 5516 6443 5523
rect 4767 5496 4893 5503
rect 5127 5496 5183 5503
rect 4467 5476 4743 5483
rect 5176 5483 5183 5496
rect 5276 5496 5473 5503
rect 5276 5483 5283 5496
rect 5527 5496 5613 5503
rect 5807 5496 6033 5503
rect 6107 5496 6513 5503
rect 4807 5476 5143 5483
rect 5176 5476 5283 5483
rect 5136 5467 5143 5476
rect 5307 5476 5773 5483
rect 5987 5476 6093 5483
rect 6107 5476 6333 5483
rect 507 5456 553 5463
rect 1807 5456 1953 5463
rect 2147 5456 2533 5463
rect 2607 5456 2793 5463
rect 2867 5456 3273 5463
rect 3647 5456 3833 5463
rect 4007 5463 4020 5467
rect 4007 5453 4023 5463
rect 4047 5456 4253 5463
rect 4487 5456 4613 5463
rect 4687 5456 4833 5463
rect 4967 5456 5053 5463
rect 5147 5456 5273 5463
rect 5347 5456 5372 5463
rect 5408 5456 5713 5463
rect 5907 5456 6073 5463
rect 6267 5456 6453 5463
rect 347 5436 673 5443
rect 827 5436 853 5443
rect 907 5436 1153 5443
rect 1687 5436 1733 5443
rect 2047 5436 2633 5443
rect 2687 5436 3113 5443
rect 3187 5436 3312 5443
rect 3348 5436 3413 5443
rect 3427 5436 3473 5443
rect 3607 5436 3713 5443
rect 3727 5436 3913 5443
rect 4016 5443 4023 5453
rect 4016 5436 4053 5443
rect 4107 5436 4753 5443
rect 5007 5436 5353 5443
rect 5507 5436 5552 5443
rect 5588 5433 5593 5447
rect 5887 5436 5933 5443
rect 6287 5436 6313 5443
rect 447 5416 493 5423
rect 507 5416 653 5423
rect 667 5416 1293 5423
rect 1307 5416 1503 5423
rect 1247 5393 1253 5407
rect 1333 5387 1347 5393
rect 1496 5387 1503 5416
rect 1727 5416 1752 5423
rect 1788 5416 1843 5423
rect 1836 5387 1843 5416
rect 2287 5416 2413 5423
rect 2876 5416 2912 5423
rect 2633 5387 2647 5393
rect 2876 5387 2883 5416
rect 2948 5416 2973 5423
rect 3327 5416 3353 5423
rect 3367 5416 3433 5423
rect 3447 5416 3613 5423
rect 3807 5413 3812 5427
rect 3848 5416 3893 5423
rect 4187 5416 4213 5423
rect 4227 5416 4493 5423
rect 4507 5416 4573 5423
rect 4647 5416 4713 5423
rect 5027 5416 5053 5423
rect 5227 5416 5313 5423
rect 5356 5416 5393 5423
rect 3273 5407 3287 5413
rect 5356 5407 5363 5416
rect 5607 5413 5613 5427
rect 5707 5416 5853 5423
rect 6167 5416 6313 5423
rect 6387 5416 6433 5423
rect 4256 5396 4473 5403
rect 87 5376 133 5383
rect 547 5373 553 5387
rect 727 5373 733 5387
rect 987 5376 1033 5383
rect 1200 5383 1213 5387
rect 1187 5376 1213 5383
rect 1200 5373 1213 5376
rect 1587 5376 1653 5383
rect 1887 5376 1993 5383
rect 2940 5383 2953 5387
rect 2927 5376 2953 5383
rect 2940 5373 2953 5376
rect 3007 5376 3033 5383
rect 3327 5376 3393 5383
rect 3487 5376 3553 5383
rect 3567 5376 3633 5383
rect 3767 5376 3873 5383
rect 4256 5383 4263 5396
rect 5347 5396 5363 5407
rect 5347 5393 5360 5396
rect 5560 5403 5573 5407
rect 5547 5396 5573 5403
rect 5560 5393 5573 5396
rect 6527 5396 6563 5403
rect 6173 5387 6187 5393
rect 4187 5376 4263 5383
rect 4547 5376 4633 5383
rect 4687 5373 4693 5387
rect 5727 5383 5740 5387
rect 5727 5376 5753 5383
rect 5727 5373 5740 5376
rect 5807 5376 5893 5383
rect 6556 5376 6563 5396
rect 4453 5367 4467 5373
rect 807 5356 833 5363
rect 1427 5356 1453 5363
rect 3267 5336 3333 5343
rect 4087 5336 4133 5343
rect 4367 5336 4393 5343
rect 4407 5333 4413 5347
rect 4847 5336 4893 5343
rect 5227 5333 5233 5347
rect 5307 5336 5333 5343
rect 5527 5336 5593 5343
rect 280 5323 293 5327
rect 267 5316 293 5323
rect 280 5313 293 5316
rect 347 5323 360 5327
rect 347 5316 373 5323
rect 347 5313 360 5316
rect 767 5316 813 5323
rect 1407 5316 1473 5323
rect 1767 5316 1813 5323
rect 1387 5296 1413 5303
rect 1547 5296 1573 5303
rect 2156 5303 2163 5333
rect 2333 5327 2347 5333
rect 2473 5327 2487 5333
rect 2047 5296 2163 5303
rect 2307 5296 2523 5303
rect 407 5276 513 5283
rect 527 5276 1053 5283
rect 1067 5276 1093 5283
rect 1247 5276 2493 5283
rect 2516 5283 2523 5296
rect 3096 5303 3103 5333
rect 3507 5323 3520 5327
rect 3507 5316 3533 5323
rect 3507 5313 3520 5316
rect 3776 5316 3853 5323
rect 3213 5307 3227 5313
rect 3027 5296 3103 5303
rect 3147 5296 3173 5303
rect 3776 5303 3783 5316
rect 3667 5296 3783 5303
rect 4136 5303 4143 5333
rect 5953 5327 5967 5333
rect 4136 5296 4473 5303
rect 4967 5296 5053 5303
rect 5887 5296 5993 5303
rect 2516 5276 2833 5283
rect 2927 5276 2953 5283
rect 3067 5276 3093 5283
rect 3207 5276 3383 5283
rect 487 5256 693 5263
rect 1327 5256 1473 5263
rect 1727 5256 1803 5263
rect 813 5247 827 5253
rect 1796 5247 1803 5256
rect 3096 5263 3103 5273
rect 2127 5256 3103 5263
rect 3167 5256 3193 5263
rect 3376 5263 3383 5276
rect 3407 5276 3573 5283
rect 3627 5276 3973 5283
rect 4027 5276 4293 5283
rect 4316 5276 4653 5283
rect 3376 5256 3433 5263
rect 3707 5256 3733 5263
rect 4316 5263 4323 5276
rect 5087 5276 5213 5283
rect 5287 5276 5313 5283
rect 5667 5276 5813 5283
rect 5867 5276 5953 5283
rect 6407 5276 6453 5283
rect 4067 5256 4323 5263
rect 4487 5256 4763 5263
rect 4756 5247 4763 5256
rect 4987 5256 5293 5263
rect 5727 5256 5953 5263
rect 6087 5256 6313 5263
rect 1247 5236 1413 5243
rect 1427 5236 1533 5243
rect 1807 5236 1913 5243
rect 2087 5236 2393 5243
rect 2507 5236 2933 5243
rect 3227 5233 3233 5247
rect 3387 5236 3453 5243
rect 3546 5233 3547 5240
rect 3568 5236 3593 5243
rect 3807 5236 3873 5243
rect 4067 5243 4080 5247
rect 4067 5236 4453 5243
rect 4067 5233 4083 5236
rect 4567 5236 4723 5243
rect 4756 5236 4773 5247
rect 1207 5216 1393 5223
rect 1867 5216 1973 5223
rect 2136 5220 2153 5223
rect 2133 5216 2153 5220
rect 2133 5207 2147 5216
rect 2167 5216 2693 5223
rect 3087 5216 3353 5223
rect 3533 5223 3547 5233
rect 4076 5227 4083 5233
rect 4716 5227 4723 5236
rect 4760 5233 4773 5236
rect 4827 5236 5183 5243
rect 3533 5220 4073 5223
rect 3535 5216 4073 5220
rect 4207 5216 4703 5223
rect 307 5196 413 5203
rect 1307 5196 1813 5203
rect 2427 5196 2653 5203
rect 2667 5196 3193 5203
rect 3276 5196 4563 5203
rect 3276 5187 3283 5196
rect 127 5176 313 5183
rect 547 5176 593 5183
rect 747 5176 933 5183
rect 987 5176 1053 5183
rect 1107 5173 1113 5187
rect 1447 5173 1453 5187
rect 1547 5176 1793 5183
rect 1927 5176 2013 5183
rect 2027 5176 2253 5183
rect 2267 5176 2333 5183
rect 2587 5176 2633 5183
rect 2767 5176 2993 5183
rect 3267 5176 3283 5187
rect 3267 5173 3280 5176
rect 3307 5176 3393 5183
rect 3467 5176 3713 5183
rect 3787 5176 3933 5183
rect 3987 5176 4453 5183
rect 4556 5183 4563 5196
rect 4587 5196 4633 5203
rect 4696 5203 4703 5216
rect 4727 5216 5073 5223
rect 5176 5223 5183 5236
rect 5207 5236 5553 5243
rect 5176 5216 5533 5223
rect 5707 5216 5773 5223
rect 5887 5216 5913 5223
rect 6307 5216 6473 5223
rect 4696 5196 4993 5203
rect 6247 5196 6413 5203
rect 6427 5196 6453 5203
rect 4556 5176 5813 5183
rect 5827 5176 6153 5183
rect 6387 5176 6473 5183
rect 207 5156 273 5163
rect 287 5156 633 5163
rect 647 5156 1153 5163
rect 1167 5156 1473 5163
rect 2247 5156 2293 5163
rect 2787 5156 3053 5163
rect 3107 5156 3552 5163
rect 3588 5156 3633 5163
rect 3647 5156 3693 5163
rect 3827 5156 3973 5163
rect 4156 5156 4252 5163
rect 87 5136 113 5143
rect 167 5136 233 5143
rect 247 5136 533 5143
rect 547 5136 1113 5143
rect 1127 5136 1193 5143
rect 1207 5136 1372 5143
rect 1408 5136 1513 5143
rect 1527 5136 1613 5143
rect 1887 5136 2093 5143
rect 2207 5136 2433 5143
rect 2547 5136 2612 5143
rect 2648 5136 3293 5143
rect 3347 5136 3373 5143
rect 3527 5136 3643 5143
rect 507 5116 607 5123
rect 593 5107 607 5116
rect 2687 5116 2733 5123
rect 2747 5113 2752 5127
rect 2788 5116 3023 5123
rect 327 5096 433 5103
rect 767 5096 873 5103
rect 980 5103 993 5107
rect 967 5096 993 5103
rect 980 5093 993 5096
rect 2927 5096 2953 5103
rect 3016 5087 3023 5116
rect 3636 5123 3643 5136
rect 3667 5136 3892 5143
rect 4156 5143 4163 5156
rect 4288 5156 4433 5163
rect 4607 5156 4773 5163
rect 4787 5156 4853 5163
rect 5707 5156 5913 5163
rect 6167 5156 6253 5163
rect 3928 5136 4163 5143
rect 4187 5136 4373 5143
rect 4427 5136 4813 5143
rect 5436 5136 5633 5143
rect 3507 5116 3623 5123
rect 3636 5116 3673 5123
rect 3067 5096 3113 5103
rect 3616 5087 3623 5116
rect 4087 5116 4143 5123
rect 3887 5096 3933 5103
rect 4136 5103 4143 5116
rect 4467 5116 4683 5123
rect 4136 5096 4213 5103
rect 4307 5096 4353 5103
rect 4676 5087 4683 5116
rect 4707 5116 4793 5123
rect 5436 5123 5443 5136
rect 6247 5136 6343 5143
rect 5373 5116 5443 5123
rect 5373 5107 5387 5116
rect 5627 5116 5653 5123
rect 5667 5116 5692 5123
rect 5728 5116 5753 5123
rect 5807 5113 5813 5127
rect 6336 5107 6343 5136
rect 5267 5096 5333 5103
rect 6047 5103 6060 5107
rect 6047 5096 6073 5103
rect 6047 5093 6060 5096
rect 5013 5087 5027 5093
rect -24 5076 13 5083
rect 2627 5076 2673 5083
rect 2867 5076 2913 5083
rect 4027 5076 4093 5083
rect 4447 5076 4513 5083
rect 4767 5076 4813 5083
rect 2607 5056 2633 5063
rect 3356 5056 3413 5063
rect 87 5033 93 5047
rect 407 5036 453 5043
rect 747 5036 793 5043
rect 1127 5036 1213 5043
rect 1267 5036 1333 5043
rect 1487 5036 1533 5043
rect 1627 5036 1713 5043
rect 1807 5036 1853 5043
rect 2080 5043 2093 5047
rect 2067 5036 2093 5043
rect 2080 5033 2093 5036
rect 2187 5033 2193 5047
rect 2447 5036 2553 5043
rect 3147 5036 3213 5043
rect 3356 5043 3363 5056
rect 3327 5036 3363 5043
rect 3387 5036 3453 5043
rect 3687 5036 3793 5043
rect 3847 5036 3912 5043
rect 3948 5033 3954 5047
rect 4227 5033 4233 5047
rect 4387 5033 4393 5047
rect 5127 5036 5193 5043
rect 5307 5036 5353 5043
rect 5407 5036 5433 5043
rect 5447 5033 5453 5047
rect 5520 5043 5533 5047
rect 5507 5036 5533 5043
rect 5520 5033 5533 5036
rect 5947 5036 6013 5043
rect 6127 5036 6213 5043
rect 293 5027 307 5033
rect 613 5027 627 5033
rect 893 5027 907 5033
rect 1467 5016 1493 5023
rect 147 4996 193 5003
rect 267 4996 313 5003
rect 507 4996 573 5003
rect 1227 4996 1253 5003
rect 1307 4996 1333 5003
rect 1567 4996 1713 5003
rect 1856 4996 1893 5003
rect 547 4973 553 4987
rect 1467 4976 1633 4983
rect 1647 4976 1753 4983
rect 1856 4983 1863 4996
rect 1907 4996 2033 5003
rect 2087 4996 2133 5003
rect 2376 5003 2383 5033
rect 2807 5023 2820 5027
rect 2807 5016 2833 5023
rect 2807 5013 2820 5016
rect 2887 5013 2892 5027
rect 2913 5013 2914 5020
rect 2987 5013 2993 5027
rect 5247 5016 5313 5023
rect 5807 5016 5873 5023
rect 6367 5016 6513 5023
rect 2873 5007 2887 5013
rect 2913 5007 2927 5013
rect 2307 4996 2383 5003
rect 2527 4996 2553 5003
rect 2567 4996 2693 5003
rect 2926 5000 2927 5007
rect 2948 4993 2953 5007
rect 1807 4976 1863 4983
rect 1887 4976 2313 4983
rect 2996 4983 3003 5013
rect 3087 4996 3233 5003
rect 3247 4996 3333 5003
rect 3687 4996 3853 5003
rect 3927 4996 4033 5003
rect 4207 4996 4693 5003
rect 5167 4996 5253 5003
rect 5267 4996 5473 5003
rect 5987 4996 6073 5003
rect 2647 4976 3153 4983
rect 3167 4976 3253 4983
rect 3347 4976 3372 4983
rect 3408 4976 3933 4983
rect 4087 4976 4113 4983
rect 4527 4976 4593 4983
rect 4647 4976 4733 4983
rect 5107 4976 5253 4983
rect 5347 4976 5413 4983
rect 5467 4976 5673 4983
rect 5727 4976 5893 4983
rect 5907 4976 6113 4983
rect 907 4956 1673 4963
rect 2047 4956 2413 4963
rect 2847 4956 2953 4963
rect 3047 4956 3573 4963
rect 3627 4956 4033 4963
rect 4247 4956 4413 4963
rect 4456 4956 4613 4963
rect 187 4936 393 4943
rect 987 4936 1233 4943
rect 1467 4936 1533 4943
rect 1587 4936 1693 4943
rect 1707 4936 2193 4943
rect 2247 4936 2373 4943
rect 2927 4936 3053 4943
rect 3247 4936 3293 4943
rect 3647 4936 3953 4943
rect 4127 4936 4313 4943
rect 2233 4927 2247 4933
rect 307 4916 473 4923
rect 487 4916 653 4923
rect 867 4916 1013 4923
rect 1747 4916 2153 4923
rect 2327 4916 2903 4923
rect 107 4896 153 4903
rect 427 4896 613 4903
rect 627 4896 713 4903
rect 1187 4896 1293 4903
rect 1307 4896 1492 4903
rect 1528 4896 1613 4903
rect 2127 4896 2232 4903
rect 2268 4896 2613 4903
rect 2747 4896 2873 4903
rect 2896 4903 2903 4916
rect 2987 4916 3013 4923
rect 3087 4916 3133 4923
rect 3207 4916 3363 4923
rect 2896 4896 2993 4903
rect 3007 4896 3073 4903
rect 3356 4903 3363 4916
rect 3547 4916 4233 4923
rect 4456 4923 4463 4956
rect 4827 4956 5053 4963
rect 5067 4956 5313 4963
rect 5447 4956 5613 4963
rect 6107 4956 6253 4963
rect 4487 4936 4563 4943
rect 4556 4927 4563 4936
rect 4707 4936 5293 4943
rect 6313 4943 6327 4953
rect 6067 4940 6327 4943
rect 6067 4936 6323 4940
rect 4456 4916 4493 4923
rect 4567 4916 4673 4923
rect 4747 4916 4833 4923
rect 4887 4916 4933 4923
rect 4947 4916 5193 4923
rect 5216 4916 5433 4923
rect 3356 4896 3692 4903
rect 3728 4896 3783 4903
rect 467 4876 493 4883
rect 2247 4876 2273 4883
rect 2407 4876 2453 4883
rect 2547 4876 2653 4883
rect 2856 4876 2913 4883
rect 1853 4867 1867 4873
rect 147 4856 253 4863
rect 387 4853 393 4867
rect 1027 4856 1093 4863
rect 1247 4863 1260 4867
rect 1247 4856 1273 4863
rect 1247 4853 1260 4856
rect 1507 4856 1553 4863
rect 2027 4856 2093 4863
rect 2187 4853 2192 4867
rect 2228 4856 2333 4863
rect 2747 4863 2760 4867
rect 2856 4863 2863 4876
rect 3776 4883 3783 4896
rect 3907 4896 4133 4903
rect 4547 4896 4593 4903
rect 4647 4896 4713 4903
rect 4727 4896 4893 4903
rect 5027 4896 5093 4903
rect 5216 4903 5223 4916
rect 5487 4916 5652 4923
rect 5688 4916 5713 4923
rect 5787 4916 5883 4923
rect 5876 4907 5883 4916
rect 6287 4916 6493 4923
rect 5147 4896 5223 4903
rect 5747 4896 5852 4903
rect 5888 4896 6083 4903
rect 3776 4876 3833 4883
rect 3573 4867 3587 4873
rect 6076 4867 6083 4896
rect 2747 4856 2773 4863
rect 2827 4856 2863 4863
rect 2747 4853 2760 4856
rect 2927 4856 2993 4863
rect 3467 4856 3533 4863
rect 3967 4856 4033 4863
rect 4187 4856 4233 4863
rect 4487 4856 4593 4863
rect 4647 4856 4753 4863
rect 5007 4856 5073 4863
rect 5187 4856 5213 4863
rect 5347 4856 5433 4863
rect 5667 4856 5713 4863
rect 1187 4833 1193 4847
rect 1747 4836 1793 4843
rect 2867 4833 2873 4847
rect 747 4816 833 4823
rect 887 4816 953 4823
rect 1707 4816 1793 4823
rect 2687 4816 2753 4823
rect 3147 4816 3233 4823
rect 4907 4813 4913 4827
rect 5207 4823 5220 4827
rect 5207 4816 5233 4823
rect 5207 4813 5220 4816
rect 5607 4816 5693 4823
rect 6187 4816 6233 4823
rect 6287 4816 6393 4823
rect 3313 4807 3327 4813
rect 5273 4807 5287 4813
rect 167 4796 273 4803
rect 567 4793 573 4807
rect 1207 4796 1253 4803
rect 2927 4796 2973 4803
rect 4027 4796 4073 4803
rect 4467 4796 4533 4803
rect 4787 4796 4873 4803
rect 5107 4796 5203 4803
rect 987 4776 1053 4783
rect 127 4756 173 4763
rect 307 4756 493 4763
rect 507 4756 733 4763
rect 1167 4756 1213 4763
rect 1436 4763 1443 4793
rect 2447 4776 2633 4783
rect 3067 4776 3373 4783
rect 3787 4776 3873 4783
rect 4156 4767 4163 4793
rect 4807 4776 5013 4783
rect 5196 4783 5203 4796
rect 5196 4776 5253 4783
rect 5267 4776 5313 4783
rect 5507 4776 5553 4783
rect 5687 4773 5693 4787
rect 6147 4776 6213 4783
rect 1267 4756 1443 4763
rect 1507 4756 1612 4763
rect 1648 4756 2073 4763
rect 2087 4756 2193 4763
rect 2367 4756 2453 4763
rect 2767 4756 3112 4763
rect 3148 4756 3193 4763
rect 3367 4756 3813 4763
rect 3867 4756 3893 4763
rect 3947 4756 4073 4763
rect 4156 4756 4173 4767
rect 4160 4753 4173 4756
rect 4467 4756 4493 4763
rect 4547 4756 5333 4763
rect 5407 4756 5453 4763
rect 5676 4756 6373 4763
rect 1527 4736 1673 4743
rect 1687 4736 1713 4743
rect 1807 4736 2373 4743
rect 2396 4736 2553 4743
rect 747 4716 853 4723
rect 927 4716 1493 4723
rect 1547 4716 2292 4723
rect 2396 4723 2403 4736
rect 2576 4736 2733 4743
rect 2328 4716 2403 4723
rect 2576 4723 2583 4736
rect 2747 4736 2923 4743
rect 2427 4716 2583 4723
rect 2627 4716 2793 4723
rect 2887 4713 2893 4727
rect 2916 4723 2923 4736
rect 2967 4736 3103 4743
rect 2916 4716 3033 4723
rect 3047 4716 3073 4723
rect 3096 4723 3103 4736
rect 3187 4736 3452 4743
rect 3488 4736 3583 4743
rect 3096 4716 3352 4723
rect 3388 4716 3553 4723
rect 3576 4723 3583 4736
rect 3647 4733 3652 4747
rect 3688 4736 4213 4743
rect 4687 4736 4793 4743
rect 5676 4747 5683 4756
rect 4847 4736 4973 4743
rect 4987 4736 5613 4743
rect 5627 4736 5673 4743
rect 5727 4736 6133 4743
rect 3576 4716 3773 4723
rect 3796 4716 3833 4723
rect 1067 4696 1393 4703
rect 1847 4696 2033 4703
rect 2407 4696 2693 4703
rect 3796 4703 3803 4716
rect 3887 4716 4473 4723
rect 4547 4716 4693 4723
rect 4807 4716 5153 4723
rect 5207 4716 5573 4723
rect 2907 4696 3803 4703
rect 807 4676 833 4683
rect 1227 4676 1533 4683
rect 1987 4676 2053 4683
rect 2467 4676 3133 4683
rect 3367 4676 3432 4683
rect 3468 4676 3773 4683
rect 3796 4683 3803 4696
rect 3827 4696 4273 4703
rect 4327 4696 4493 4703
rect 4747 4696 4893 4703
rect 5007 4696 5373 4703
rect 5387 4696 5913 4703
rect 3796 4676 5133 4683
rect 5447 4676 6153 4683
rect 687 4656 733 4663
rect 747 4656 1173 4663
rect 1267 4656 1592 4663
rect 1628 4656 1953 4663
rect 2147 4656 2252 4663
rect 2288 4653 2293 4667
rect 2367 4656 2633 4663
rect 2887 4656 2972 4663
rect 3008 4656 3133 4663
rect 267 4636 433 4643
rect 527 4636 813 4643
rect 1007 4636 1693 4643
rect 1993 4640 2007 4653
rect 3327 4656 3453 4663
rect 3193 4647 3207 4653
rect 3496 4656 3703 4663
rect 1996 4627 2003 4640
rect 2727 4636 2853 4643
rect 2867 4636 2893 4643
rect 2967 4636 3053 4643
rect 3496 4643 3503 4656
rect 3447 4636 3503 4643
rect 3647 4633 3653 4647
rect 3696 4643 3703 4656
rect 3747 4656 3793 4663
rect 3867 4656 4013 4663
rect 4027 4656 4383 4663
rect 4376 4647 4383 4656
rect 4647 4656 4872 4663
rect 4908 4656 5193 4663
rect 5287 4656 5713 4663
rect 5847 4656 5973 4663
rect 3696 4636 3733 4643
rect 3787 4636 3913 4643
rect 3967 4636 4053 4643
rect 4387 4636 4593 4643
rect 4847 4636 5233 4643
rect 5467 4633 5473 4647
rect 5547 4636 5733 4643
rect 5747 4636 6053 4643
rect 6247 4636 6313 4643
rect 327 4616 373 4623
rect 507 4616 573 4623
rect 787 4616 833 4623
rect 947 4616 1213 4623
rect 1287 4616 1553 4623
rect 1567 4616 1953 4623
rect 2007 4616 2033 4623
rect 2767 4616 3173 4623
rect 3247 4616 3333 4623
rect 4287 4616 4533 4623
rect 5027 4616 5093 4623
rect 5307 4616 5393 4623
rect 6147 4616 6293 4623
rect -24 4596 13 4603
rect 1100 4603 1113 4607
rect 1093 4593 1113 4603
rect 1327 4596 1513 4603
rect 1707 4596 1873 4603
rect 2167 4596 2223 4603
rect 1093 4587 1107 4593
rect 487 4576 533 4583
rect 1393 4567 1407 4573
rect 2216 4567 2223 4596
rect 3567 4596 3633 4603
rect 3767 4596 3813 4603
rect 4267 4596 4333 4603
rect 2853 4587 2867 4593
rect 5396 4587 5403 4613
rect 6013 4596 6113 4603
rect 6013 4587 6027 4596
rect 2767 4573 2773 4587
rect 2947 4576 2993 4583
rect 3087 4576 3133 4583
rect 3787 4576 3853 4583
rect 5467 4576 5513 4583
rect 5880 4583 5893 4587
rect 5867 4576 5893 4583
rect 5880 4573 5893 4576
rect -24 4556 13 4563
rect 207 4556 253 4563
rect 827 4556 893 4563
rect 1636 4556 1713 4563
rect 1636 4547 1643 4556
rect 1927 4556 1993 4563
rect 3207 4556 3253 4563
rect 4607 4556 4673 4563
rect 6367 4556 6413 4563
rect 4596 4547 4603 4553
rect 27 4533 33 4547
rect 1627 4536 1643 4547
rect 1627 4533 1640 4536
rect 2107 4536 2133 4543
rect 4587 4536 4603 4547
rect 4587 4533 4600 4536
rect 107 4516 233 4523
rect 427 4516 493 4523
rect 647 4516 713 4523
rect 1227 4513 1233 4527
rect 1467 4516 1573 4523
rect 1947 4516 1993 4523
rect 2067 4516 2153 4523
rect 2307 4516 2413 4523
rect 2647 4516 2693 4523
rect 3180 4523 3192 4527
rect 2787 4516 2873 4523
rect 3167 4516 3192 4523
rect 3180 4513 3192 4516
rect 3228 4516 3273 4523
rect 3327 4513 3333 4527
rect 3780 4523 3793 4527
rect 3587 4516 3713 4523
rect 3767 4516 3793 4523
rect 3780 4513 3793 4516
rect 3847 4523 3860 4527
rect 3847 4516 3873 4523
rect 3847 4513 3860 4516
rect 4447 4516 4533 4523
rect 4787 4523 4800 4527
rect 4787 4516 4813 4523
rect 4787 4513 4800 4516
rect 4867 4516 4973 4523
rect 5167 4516 5233 4523
rect 5887 4516 5953 4523
rect 27 4476 473 4483
rect 596 4483 603 4513
rect 527 4476 603 4483
rect 767 4476 893 4483
rect 1076 4483 1083 4513
rect 2733 4507 2747 4513
rect 3013 4507 3027 4513
rect 1787 4496 1853 4503
rect 2096 4496 2193 4503
rect 1076 4476 1152 4483
rect 1188 4476 1313 4483
rect 1827 4476 1873 4483
rect 2096 4483 2103 4496
rect 2247 4496 2293 4503
rect 2927 4496 2953 4503
rect 3607 4496 3673 4503
rect 2047 4476 2103 4483
rect 2667 4476 3213 4483
rect 3287 4476 3353 4483
rect 3467 4476 3493 4483
rect 3647 4476 3723 4483
rect 1107 4456 1253 4463
rect 1427 4456 1473 4463
rect 1487 4456 1633 4463
rect 1896 4456 2173 4463
rect 1896 4447 1903 4456
rect 2247 4456 2313 4463
rect 2627 4456 2913 4463
rect 2967 4456 3193 4463
rect 3247 4456 3353 4463
rect 3447 4456 3493 4463
rect 3587 4456 3693 4463
rect 3716 4463 3723 4476
rect 3996 4483 4003 4513
rect 4353 4507 4367 4513
rect 3747 4476 4003 4483
rect 4396 4483 4403 4513
rect 4287 4476 4403 4483
rect 4416 4476 4693 4483
rect 3716 4456 3873 4463
rect 3987 4456 4033 4463
rect 4416 4463 4423 4476
rect 4787 4476 4833 4483
rect 5116 4483 5123 4513
rect 5693 4507 5707 4513
rect 5993 4507 6007 4513
rect 4967 4476 5123 4483
rect 5147 4476 5293 4483
rect 5547 4476 5953 4483
rect 5967 4476 6113 4483
rect 4307 4456 4423 4463
rect 4487 4456 4613 4463
rect 4727 4456 4853 4463
rect 4947 4456 5093 4463
rect 5107 4456 5253 4463
rect 5347 4456 5573 4463
rect 5767 4456 5993 4463
rect 1047 4436 1213 4443
rect 1367 4436 1493 4443
rect 1627 4436 1893 4443
rect 1967 4436 2523 4443
rect 147 4416 2273 4423
rect 2347 4416 2433 4423
rect 2516 4423 2523 4436
rect 2547 4436 2733 4443
rect 2867 4436 3113 4443
rect 3267 4436 3333 4443
rect 3407 4436 4653 4443
rect 4847 4436 5013 4443
rect 5036 4436 5183 4443
rect 2516 4416 2733 4423
rect 2747 4416 3153 4423
rect 3307 4416 3413 4423
rect 3436 4416 3472 4423
rect 707 4396 773 4403
rect 787 4396 1033 4403
rect 1127 4396 1173 4403
rect 1347 4396 1373 4403
rect 1387 4396 1733 4403
rect 1867 4393 1873 4407
rect 1967 4396 1993 4403
rect 2007 4396 2053 4403
rect 2187 4396 2253 4403
rect 2527 4396 2673 4403
rect 3007 4396 3313 4403
rect 3436 4403 3443 4416
rect 3508 4416 3552 4423
rect 3588 4416 3773 4423
rect 5036 4423 5043 4436
rect 4147 4416 5043 4423
rect 5067 4416 5153 4423
rect 5176 4423 5183 4436
rect 5176 4416 5793 4423
rect 3367 4396 3443 4403
rect 3707 4396 4173 4403
rect 4247 4396 4293 4403
rect 4367 4396 4553 4403
rect 4567 4396 5653 4403
rect 5667 4396 6293 4403
rect 247 4376 333 4383
rect 747 4376 853 4383
rect 816 4347 823 4376
rect 947 4376 1193 4383
rect 1256 4376 1312 4383
rect 1256 4347 1263 4376
rect 1348 4376 1427 4383
rect 1413 4367 1427 4376
rect 1687 4376 1752 4383
rect 1788 4376 1833 4383
rect 2047 4376 2213 4383
rect 3227 4376 3353 4383
rect 3707 4376 3893 4383
rect 4087 4376 4513 4383
rect 4527 4376 4753 4383
rect 4827 4376 5213 4383
rect 5487 4376 5513 4383
rect 5567 4376 5753 4383
rect 5807 4376 6063 4383
rect 2507 4356 2533 4363
rect 3967 4356 4193 4363
rect 3773 4347 3787 4353
rect 4933 4347 4947 4353
rect 6056 4347 6063 4376
rect 6156 4367 6163 4396
rect 6307 4396 6353 4403
rect 6276 4376 6313 4383
rect 6276 4363 6283 4376
rect 6387 4376 6433 4383
rect 6207 4356 6283 4363
rect 267 4336 313 4343
rect 587 4336 693 4343
rect 1127 4336 1213 4343
rect 1527 4336 1613 4343
rect 1707 4336 1793 4343
rect 2260 4343 2273 4347
rect 2247 4336 2273 4343
rect 2260 4333 2273 4336
rect 3100 4343 3112 4347
rect 2967 4336 3033 4343
rect 3087 4336 3112 4343
rect 3100 4333 3112 4336
rect 3148 4336 3213 4343
rect 3327 4336 3373 4343
rect 3687 4336 3733 4343
rect 4507 4336 4573 4343
rect 4667 4333 4673 4347
rect 5280 4343 5292 4347
rect 5267 4336 5292 4343
rect 5280 4333 5292 4336
rect 5328 4336 5413 4343
rect 5507 4333 5513 4347
rect 5647 4336 5693 4343
rect 5787 4336 5853 4343
rect 5920 4343 5932 4347
rect 5907 4336 5932 4343
rect 5920 4333 5932 4336
rect 5968 4333 5973 4347
rect 6407 4336 6473 4343
rect 447 4316 473 4323
rect 47 4296 93 4303
rect 1687 4293 1693 4307
rect 2927 4293 2933 4307
rect 3847 4296 3933 4303
rect 4167 4303 4180 4307
rect 4167 4296 4193 4303
rect 4167 4293 4180 4296
rect 6087 4296 6173 4303
rect 1433 4287 1447 4293
rect 1953 4287 1967 4293
rect 2633 4287 2647 4293
rect 847 4276 913 4283
rect 967 4276 1053 4283
rect 2280 4283 2293 4287
rect 2267 4276 2293 4283
rect 2280 4273 2293 4276
rect 4807 4276 4953 4283
rect 5407 4276 5473 4283
rect 5940 4283 5953 4287
rect 5927 4276 5953 4283
rect 5940 4273 5953 4276
rect 1007 4256 1053 4263
rect 1407 4256 1453 4263
rect 1467 4256 1493 4263
rect 1836 4256 2093 4263
rect 207 4236 233 4243
rect 387 4236 573 4243
rect 727 4236 933 4243
rect 947 4236 973 4243
rect 1836 4243 1843 4256
rect 2507 4256 2573 4263
rect 2587 4256 2713 4263
rect 2927 4256 2993 4263
rect 4087 4256 4113 4263
rect 4427 4256 4453 4263
rect 1047 4236 1843 4243
rect 1856 4236 1973 4243
rect 327 4216 553 4223
rect 1067 4216 1133 4223
rect 1247 4216 1353 4223
rect 1367 4216 1773 4223
rect 1856 4223 1863 4236
rect 2067 4236 2133 4243
rect 2547 4236 2633 4243
rect 3187 4236 3233 4243
rect 3413 4243 3427 4253
rect 3387 4240 3427 4243
rect 3387 4236 3423 4240
rect 3667 4236 3833 4243
rect 3907 4236 4163 4243
rect 1827 4216 1863 4223
rect 1927 4216 2033 4223
rect 2087 4216 2153 4223
rect 2516 4216 2593 4223
rect 1207 4196 1253 4203
rect 1327 4193 1333 4207
rect 1887 4196 2173 4203
rect 2516 4203 2523 4216
rect 2940 4223 2953 4227
rect 2807 4216 2863 4223
rect 2307 4196 2523 4203
rect 2547 4196 2833 4203
rect 2856 4203 2863 4216
rect 2936 4214 2953 4223
rect 3067 4216 3153 4223
rect 2936 4213 2960 4214
rect 3207 4216 3253 4223
rect 3327 4216 3413 4223
rect 4156 4223 4163 4236
rect 4387 4236 4433 4243
rect 4527 4236 4553 4243
rect 4667 4236 4713 4243
rect 4787 4236 4813 4243
rect 5096 4243 5103 4273
rect 5187 4256 5213 4263
rect 5096 4236 5233 4243
rect 5396 4243 5403 4273
rect 5873 4267 5887 4273
rect 5287 4236 5403 4243
rect 5447 4236 6313 4243
rect 4156 4216 4353 4223
rect 4367 4216 4413 4223
rect 4987 4216 5113 4223
rect 5127 4216 5503 4223
rect 2936 4203 2943 4213
rect 5496 4207 5503 4216
rect 5567 4216 5753 4223
rect 5887 4216 6173 4223
rect 6187 4216 6353 4223
rect 2960 4206 2973 4207
rect 2856 4196 2943 4203
rect 287 4176 393 4183
rect 407 4176 1813 4183
rect 2967 4193 2973 4206
rect 3067 4196 3292 4203
rect 3328 4196 3432 4203
rect 3468 4196 3573 4203
rect 3587 4196 3692 4203
rect 3728 4196 4183 4203
rect 2956 4183 2963 4192
rect 2127 4176 2963 4183
rect 3167 4176 3193 4183
rect 3247 4176 3493 4183
rect 3507 4176 3753 4183
rect 3767 4176 4153 4183
rect 4176 4183 4183 4196
rect 4207 4196 4553 4203
rect 4567 4196 4913 4203
rect 5027 4196 5313 4203
rect 5356 4196 5432 4203
rect 4176 4176 4273 4183
rect 4287 4176 4633 4183
rect 4707 4176 5053 4183
rect 5356 4183 5363 4196
rect 5468 4193 5472 4207
rect 5508 4196 5533 4203
rect 5587 4196 5693 4203
rect 5747 4196 5913 4203
rect 5067 4176 5363 4183
rect 5387 4176 5553 4183
rect 867 4156 1313 4163
rect 1467 4156 1913 4163
rect 2067 4156 2183 4163
rect 547 4136 1173 4143
rect 1307 4136 1433 4143
rect 1487 4136 1573 4143
rect 1647 4136 1953 4143
rect 2007 4136 2053 4143
rect 2127 4136 2153 4143
rect 2176 4143 2183 4156
rect 2267 4156 2452 4163
rect 2488 4156 2933 4163
rect 3047 4156 3112 4163
rect 3148 4156 3283 4163
rect 3276 4147 3283 4156
rect 3327 4156 3373 4163
rect 3396 4156 4053 4163
rect 2176 4136 2533 4143
rect 2627 4136 2652 4143
rect 2688 4136 2792 4143
rect 2828 4136 2973 4143
rect 3027 4136 3053 4143
rect 3107 4136 3193 4143
rect 3396 4143 3403 4156
rect 4127 4156 4373 4163
rect 4427 4156 4873 4163
rect 5027 4156 6193 4163
rect 3287 4136 3403 4143
rect 3687 4136 3713 4143
rect 3727 4136 4043 4143
rect 947 4116 1273 4123
rect 1667 4116 1693 4123
rect 1787 4116 1933 4123
rect 1987 4116 2073 4123
rect 2096 4116 2543 4123
rect 367 4096 453 4103
rect 567 4096 733 4103
rect 827 4096 893 4103
rect 1407 4096 1533 4103
rect 1547 4096 1733 4103
rect 1867 4096 1913 4103
rect 1927 4096 2013 4103
rect 2096 4103 2103 4116
rect 2027 4096 2103 4103
rect 2187 4096 2513 4103
rect 2536 4103 2543 4116
rect 2687 4116 2873 4123
rect 2896 4116 3132 4123
rect 2896 4103 2903 4116
rect 3168 4116 3323 4123
rect 2536 4096 2903 4103
rect 3027 4096 3052 4103
rect 3088 4096 3123 4103
rect 927 4076 1033 4083
rect 1107 4076 1173 4083
rect 2227 4076 2333 4083
rect 3007 4073 3013 4087
rect 3116 4083 3123 4096
rect 3147 4096 3293 4103
rect 3316 4103 3323 4116
rect 3347 4116 3493 4123
rect 4036 4123 4043 4136
rect 4547 4136 4593 4143
rect 4687 4136 4793 4143
rect 5187 4136 5503 4143
rect 5496 4127 5503 4136
rect 5607 4136 5833 4143
rect 6127 4136 6373 4143
rect 4036 4116 4173 4123
rect 4767 4116 4833 4123
rect 4927 4116 5053 4123
rect 5067 4116 5453 4123
rect 5507 4116 5633 4123
rect 5867 4116 6053 4123
rect 6067 4116 6153 4123
rect 3316 4096 4233 4103
rect 4567 4096 4793 4103
rect 4887 4096 4973 4103
rect 5147 4096 5193 4103
rect 5267 4096 5913 4103
rect 5927 4096 5953 4103
rect 6167 4096 6463 4103
rect 3116 4076 3153 4083
rect 3427 4076 3453 4083
rect 3636 4076 3773 4083
rect 107 4056 153 4063
rect 287 4056 313 4063
rect 687 4056 733 4063
rect 807 4053 813 4067
rect 1247 4056 1293 4063
rect 1447 4056 1493 4063
rect 2367 4063 2380 4067
rect 2367 4056 2393 4063
rect 2367 4053 2380 4056
rect 2447 4056 2513 4063
rect 3636 4047 3643 4076
rect 4227 4076 4313 4083
rect 4647 4076 4893 4083
rect 5373 4067 5387 4073
rect 6456 4067 6463 4096
rect 3687 4056 3713 4063
rect 4607 4053 4613 4067
rect 4887 4056 4933 4063
rect 4987 4056 5053 4063
rect 5247 4053 5253 4067
rect 5787 4053 5793 4067
rect 5900 4063 5913 4067
rect 5887 4056 5913 4063
rect 5900 4053 5913 4056
rect 907 4036 953 4043
rect 1007 4036 1113 4043
rect 1747 4036 1813 4043
rect 2087 4043 2100 4047
rect 2087 4036 2113 4043
rect 2087 4033 2100 4036
rect 2247 4043 2260 4047
rect 2247 4036 2273 4043
rect 2247 4033 2260 4036
rect 3587 4036 3633 4043
rect 4307 4033 4313 4047
rect 4447 4033 4453 4047
rect 4467 4036 4553 4043
rect 327 3996 373 4003
rect 427 3996 533 4003
rect 747 3996 793 4003
rect 1187 4003 1200 4007
rect 1187 3996 1213 4003
rect 1187 3993 1200 3996
rect 1347 4003 1360 4007
rect 1347 3996 1373 4003
rect 1347 3993 1360 3996
rect 1527 3996 1572 4003
rect 1608 3996 1673 4003
rect 2007 3996 2053 4003
rect 2227 3993 2233 4007
rect 2440 4003 2452 4007
rect 2427 3996 2452 4003
rect 2440 3993 2452 3996
rect 2488 3996 2533 4003
rect 2853 4003 2867 4013
rect 2747 4000 2867 4003
rect 2747 3996 2863 4000
rect 3247 3996 3293 4003
rect 3307 3993 3313 4007
rect 3367 3996 3403 4003
rect 256 3963 263 3993
rect 2613 3987 2627 3993
rect 3073 3987 3087 3993
rect 2787 3976 2853 3983
rect 3396 3983 3403 3996
rect 3427 3996 3513 4003
rect 3567 3996 3613 4003
rect 4093 4003 4107 4013
rect 3987 4000 4107 4003
rect 3987 3996 4103 4000
rect 5067 3996 5113 4003
rect 5527 3996 5613 4003
rect 5707 3996 5773 4003
rect 6067 3996 6133 4003
rect 6327 3996 6373 4003
rect 3396 3976 3473 3983
rect 4027 3976 4093 3983
rect 4787 3976 4833 3983
rect 207 3956 263 3963
rect 707 3956 833 3963
rect 847 3956 893 3963
rect 1187 3953 1193 3967
rect 1487 3956 1693 3963
rect 1747 3956 2333 3963
rect 2507 3956 3313 3963
rect 3467 3956 3513 3963
rect 3587 3956 3733 3963
rect 3927 3956 3953 3963
rect 4007 3956 4413 3963
rect 4427 3956 4533 3963
rect 127 3936 153 3943
rect 167 3936 1093 3943
rect 1107 3936 1252 3943
rect 1288 3936 2353 3943
rect 2467 3936 2673 3943
rect 2767 3936 2913 3943
rect 2927 3936 3333 3943
rect 3347 3936 3573 3943
rect 3667 3936 3713 3943
rect 3867 3936 3953 3943
rect 4047 3936 4072 3943
rect 4108 3936 4153 3943
rect 4167 3936 4293 3943
rect 4307 3936 4433 3943
rect 4686 3933 4687 3940
rect 4776 3943 4783 3973
rect 4956 3963 4963 3993
rect 5567 3976 5613 3983
rect 4956 3956 5073 3963
rect 5087 3956 5353 3963
rect 5367 3956 5573 3963
rect 5627 3956 5703 3963
rect 4708 3936 4783 3943
rect 4807 3936 5093 3943
rect 5107 3936 5153 3943
rect 5167 3936 5273 3943
rect 5287 3936 5413 3943
rect 5567 3936 5592 3943
rect 5628 3936 5653 3943
rect 5696 3943 5703 3956
rect 5816 3963 5823 3993
rect 5727 3956 5823 3963
rect 5867 3956 5913 3963
rect 5976 3963 5983 3993
rect 6013 3987 6027 3993
rect 5976 3956 6053 3963
rect 6147 3956 6213 3963
rect 6387 3956 6453 3963
rect 5696 3936 5752 3943
rect 5788 3933 5793 3947
rect 5807 3936 5933 3943
rect 527 3916 613 3923
rect 627 3916 1113 3923
rect 1136 3916 2292 3923
rect 247 3896 453 3903
rect 467 3896 913 3903
rect 967 3896 993 3903
rect 1136 3903 1143 3916
rect 2328 3916 2453 3923
rect 2507 3916 2612 3923
rect 2648 3916 2713 3923
rect 2767 3916 2993 3923
rect 3327 3916 3423 3923
rect 1047 3896 1143 3903
rect 1307 3896 2372 3903
rect 2408 3896 2553 3903
rect 2607 3896 2653 3903
rect 2667 3896 2723 3903
rect 807 3876 873 3883
rect 1407 3876 1833 3883
rect 1847 3876 2053 3883
rect 2307 3873 2312 3887
rect 2348 3876 2633 3883
rect 2716 3883 2723 3896
rect 2747 3896 2812 3903
rect 2848 3896 2893 3903
rect 2907 3896 3213 3903
rect 3347 3896 3373 3903
rect 3416 3903 3423 3916
rect 3447 3916 3553 3923
rect 3776 3916 3913 3923
rect 3776 3903 3783 3916
rect 3987 3916 4473 3923
rect 4673 3923 4687 3933
rect 4673 3920 4753 3923
rect 4675 3916 4753 3920
rect 4807 3916 5013 3923
rect 5067 3916 5253 3923
rect 5327 3916 5393 3923
rect 3416 3896 3783 3903
rect 3807 3896 4223 3903
rect 2716 3876 2753 3883
rect 3267 3876 3293 3883
rect 4216 3883 4223 3896
rect 4247 3896 4593 3903
rect 4987 3900 5043 3903
rect 4987 3896 5047 3900
rect 5033 3887 5047 3896
rect 5247 3896 5313 3903
rect 5327 3896 5613 3903
rect 5767 3896 6113 3903
rect 4216 3876 4513 3883
rect 4667 3876 4693 3883
rect 4847 3876 4892 3883
rect 4928 3876 4953 3883
rect 5267 3876 5633 3883
rect 5827 3876 6053 3883
rect 6393 3867 6407 3873
rect 567 3856 653 3863
rect 1947 3856 2332 3863
rect 687 3836 733 3843
rect 913 3827 927 3833
rect 2096 3827 2103 3856
rect 2368 3856 2473 3863
rect 2527 3856 2623 3863
rect 2616 3827 2623 3856
rect 3147 3856 3192 3863
rect 3228 3856 3333 3863
rect 4687 3856 4733 3863
rect 4747 3856 4793 3863
rect 5047 3856 5193 3863
rect 5207 3856 5273 3863
rect 5487 3856 5652 3863
rect 5688 3856 5713 3863
rect 6013 3847 6027 3853
rect 3087 3836 3133 3843
rect 6136 3856 6252 3863
rect 6136 3827 6143 3856
rect 6288 3856 6313 3863
rect 67 3816 113 3823
rect 267 3816 333 3823
rect 427 3816 492 3823
rect 528 3816 573 3823
rect 1147 3816 1213 3823
rect 1267 3816 1373 3823
rect 1567 3816 1653 3823
rect 1827 3813 1833 3827
rect 2007 3813 2013 3827
rect 2267 3816 2313 3823
rect 2487 3816 2573 3823
rect 3307 3816 3353 3823
rect 5127 3816 5193 3823
rect 5216 3816 5273 3823
rect 653 3807 667 3813
rect 4567 3796 4593 3803
rect 5216 3803 5223 3816
rect 5467 3816 5553 3823
rect 5666 3813 5673 3827
rect 5840 3823 5853 3827
rect 5827 3816 5853 3823
rect 5840 3813 5853 3816
rect 5987 3813 5993 3827
rect 6307 3814 6313 3827
rect 6307 3813 6320 3814
rect 5187 3796 5223 3803
rect 5693 3787 5707 3793
rect 767 3776 853 3783
rect 1100 3783 1113 3787
rect 1087 3776 1113 3783
rect 1100 3773 1113 3776
rect 1720 3783 1733 3787
rect 1707 3776 1733 3783
rect 1720 3773 1733 3776
rect 1807 3773 1813 3787
rect 1967 3773 1973 3787
rect 2487 3776 2513 3783
rect 4307 3776 4353 3783
rect 4847 3776 4933 3783
rect 4987 3776 5033 3783
rect 6367 3773 6373 3787
rect 6387 3776 6433 3783
rect 3013 3767 3027 3773
rect 1187 3753 1193 3767
rect 1287 3756 1353 3763
rect 1527 3753 1533 3767
rect 2127 3756 2193 3763
rect 2547 3753 2553 3767
rect 747 3736 773 3743
rect 987 3736 1053 3743
rect 2593 3743 2607 3753
rect 2593 3736 2633 3743
rect 3087 3736 3133 3743
rect 4216 3743 4223 3773
rect 4587 3756 4653 3763
rect 4748 3763 4760 3767
rect 4748 3756 4773 3763
rect 4748 3753 4760 3756
rect 5147 3756 5253 3763
rect 5660 3763 5673 3767
rect 5647 3756 5673 3763
rect 5660 3753 5673 3756
rect 4107 3736 4223 3743
rect 6393 3747 6407 3753
rect 147 3716 313 3723
rect 327 3716 453 3723
rect 607 3716 853 3723
rect 867 3716 893 3723
rect 947 3716 1093 3723
rect 1147 3716 1193 3723
rect 1247 3716 1453 3723
rect 1747 3716 1913 3723
rect 1987 3716 2133 3723
rect 2247 3716 2393 3723
rect 2447 3716 2473 3723
rect 3207 3716 3293 3723
rect 4447 3716 4493 3723
rect 4567 3716 4592 3723
rect 4628 3716 4693 3723
rect 4767 3716 4833 3723
rect 4947 3716 5133 3723
rect 5307 3716 5433 3723
rect 5567 3716 5733 3723
rect 5747 3716 5913 3723
rect 67 3696 233 3703
rect 507 3696 1493 3703
rect 2287 3696 2313 3703
rect 2436 3703 2443 3713
rect 6013 3707 6027 3713
rect 2327 3696 2443 3703
rect 3247 3696 3373 3703
rect 4807 3696 4913 3703
rect 5347 3696 5473 3703
rect 5727 3696 5753 3703
rect 5767 3696 5953 3703
rect 287 3676 333 3683
rect 347 3676 393 3683
rect 1067 3676 1153 3683
rect 2267 3676 2312 3683
rect 2348 3676 2413 3683
rect 2567 3676 2733 3683
rect 2847 3676 3113 3683
rect 3127 3676 3433 3683
rect 3447 3676 3853 3683
rect 3867 3676 4093 3683
rect 4167 3676 4572 3683
rect 4608 3676 4683 3683
rect 107 3656 553 3663
rect 1487 3656 1513 3663
rect 1867 3656 2143 3663
rect 267 3636 473 3643
rect 787 3636 933 3643
rect 2136 3643 2143 3656
rect 2336 3656 2533 3663
rect 2136 3636 2273 3643
rect 2336 3643 2343 3656
rect 2867 3656 3153 3663
rect 3587 3656 3673 3663
rect 3927 3656 3993 3663
rect 4096 3656 4653 3663
rect 2287 3636 2343 3643
rect 2367 3636 2473 3643
rect 2496 3636 2713 3643
rect 747 3616 853 3623
rect 867 3616 1253 3623
rect 2496 3623 2503 3636
rect 2907 3636 3033 3643
rect 3576 3643 3583 3653
rect 3056 3636 3583 3643
rect 2127 3616 2503 3623
rect 3056 3623 3063 3636
rect 3627 3636 3933 3643
rect 4096 3643 4103 3656
rect 4676 3663 4683 3676
rect 5287 3676 5553 3683
rect 5667 3676 5693 3683
rect 5736 3676 5813 3683
rect 5736 3663 5743 3676
rect 5907 3676 6473 3683
rect 4676 3656 5743 3663
rect 5847 3656 6073 3663
rect 6467 3656 6493 3663
rect 4027 3636 4103 3643
rect 4127 3636 4693 3643
rect 4907 3636 4933 3643
rect 4947 3636 5093 3643
rect 2527 3616 3063 3623
rect 3147 3616 3233 3623
rect 3667 3616 4353 3623
rect 4507 3616 4613 3623
rect 4667 3616 4993 3623
rect 5767 3616 5933 3623
rect 5947 3616 6013 3623
rect 6227 3616 6273 3623
rect 876 3596 1373 3603
rect 87 3576 193 3583
rect 327 3576 413 3583
rect 427 3576 513 3583
rect 607 3576 833 3583
rect 876 3583 883 3596
rect 1427 3596 1533 3603
rect 1547 3596 1653 3603
rect 1827 3596 2513 3603
rect 3427 3596 3513 3603
rect 4067 3596 4253 3603
rect 4267 3596 4463 3603
rect 847 3576 883 3583
rect 907 3576 973 3583
rect 1267 3576 1553 3583
rect 1627 3576 1833 3583
rect 2347 3576 2393 3583
rect 2767 3576 2853 3583
rect 3187 3576 3253 3583
rect 3267 3576 3453 3583
rect 3567 3576 3593 3583
rect 4047 3576 4433 3583
rect 4456 3583 4463 3596
rect 4587 3596 5712 3603
rect 5748 3596 5893 3603
rect 4456 3576 4743 3583
rect 2493 3567 2507 3573
rect 4736 3567 4743 3576
rect 4787 3576 5033 3583
rect 5347 3576 5493 3583
rect 5607 3576 5833 3583
rect 5967 3576 5993 3583
rect 6087 3576 6212 3583
rect 6248 3576 6513 3583
rect 2827 3556 2863 3563
rect 1927 3536 1953 3543
rect 2187 3533 2193 3547
rect 2327 3536 2373 3543
rect 2480 3543 2493 3547
rect 2467 3536 2493 3543
rect 2480 3533 2493 3536
rect 2856 3543 2863 3556
rect 3047 3556 3093 3563
rect 4847 3556 4893 3563
rect 5567 3556 5667 3563
rect 4733 3547 4747 3553
rect 2856 3536 2913 3543
rect 3247 3533 3253 3547
rect 5047 3536 5093 3543
rect 5653 3547 5667 3556
rect 5767 3536 5853 3543
rect 6307 3533 6313 3547
rect 6327 3543 6340 3547
rect 6327 3536 6353 3543
rect 6327 3533 6340 3536
rect 147 3516 233 3523
rect 447 3513 453 3527
rect 976 3516 1053 3523
rect 1067 3516 1173 3523
rect 976 3507 983 3516
rect 1727 3516 1793 3523
rect 3827 3513 3833 3527
rect 4087 3516 4153 3523
rect 4867 3516 4953 3523
rect 5107 3516 5173 3523
rect 5587 3516 5613 3523
rect 967 3496 983 3507
rect 967 3493 980 3496
rect 2487 3496 2533 3503
rect 4907 3496 4973 3503
rect 5727 3496 5753 3503
rect 307 3476 373 3483
rect 567 3476 613 3483
rect 847 3476 913 3483
rect 1387 3473 1393 3487
rect 1567 3476 1613 3483
rect 1867 3473 1873 3487
rect 2027 3476 2113 3483
rect 2447 3473 2453 3487
rect 2627 3476 2713 3483
rect 2867 3483 2880 3487
rect 2920 3483 2933 3487
rect 2867 3476 2893 3483
rect 2907 3476 2933 3483
rect 2867 3473 2880 3476
rect 2920 3473 2933 3476
rect 3187 3476 3233 3483
rect 3367 3476 3453 3483
rect 3547 3476 3633 3483
rect 3967 3476 4013 3483
rect 4427 3476 4533 3483
rect 4607 3473 4613 3487
rect 4727 3476 4793 3483
rect 4927 3476 5013 3483
rect 5027 3476 5153 3483
rect 5227 3476 5273 3483
rect 5367 3476 5473 3483
rect 5700 3486 5720 3487
rect 5700 3483 5713 3486
rect 5687 3476 5713 3483
rect 5700 3473 5713 3476
rect 756 3443 763 3473
rect 647 3436 763 3443
rect 827 3436 873 3443
rect 1236 3443 1243 3473
rect 2507 3456 2533 3463
rect 887 3436 943 3443
rect 1236 3436 1413 3443
rect 867 3416 913 3423
rect 936 3423 943 3436
rect 1427 3436 1573 3443
rect 1587 3436 1673 3443
rect 1827 3436 2233 3443
rect 2527 3436 2573 3443
rect 2907 3436 2953 3443
rect 3047 3436 3093 3443
rect 3316 3443 3323 3473
rect 5513 3467 5527 3473
rect 5827 3473 5833 3487
rect 6067 3476 6093 3483
rect 6107 3476 6153 3483
rect 6247 3476 6293 3483
rect 3287 3436 3323 3443
rect 3347 3436 3593 3443
rect 4047 3436 4393 3443
rect 4527 3436 4633 3443
rect 4687 3436 4773 3443
rect 5167 3436 5313 3443
rect 5567 3436 5753 3443
rect 5887 3436 5953 3443
rect 5967 3436 6013 3443
rect 6127 3436 6193 3443
rect 936 3416 1093 3423
rect 1687 3416 2033 3423
rect 2047 3416 2373 3423
rect 2647 3416 2703 3423
rect 607 3396 1313 3403
rect 1927 3396 2033 3403
rect 2287 3396 2513 3403
rect 2567 3396 2673 3403
rect 2696 3403 2703 3416
rect 2787 3416 2963 3423
rect 2696 3396 2793 3403
rect 2956 3403 2963 3416
rect 3176 3416 3353 3423
rect 2956 3396 2992 3403
rect 3176 3403 3183 3416
rect 3467 3416 3493 3423
rect 3947 3416 4173 3423
rect 4187 3416 4293 3423
rect 4467 3416 4613 3423
rect 4627 3416 4873 3423
rect 5047 3416 5173 3423
rect 5527 3416 5593 3423
rect 5687 3416 5733 3423
rect 6227 3416 6272 3423
rect 6308 3416 6333 3423
rect 3028 3396 3183 3403
rect 3307 3396 3393 3403
rect 4647 3396 4813 3403
rect 5007 3396 5053 3403
rect 5627 3396 5893 3403
rect 5907 3396 5993 3403
rect 727 3376 773 3383
rect 787 3376 1033 3383
rect 1107 3376 1253 3383
rect 1347 3376 1813 3383
rect 1887 3376 2013 3383
rect 2027 3376 2153 3383
rect 2193 3373 2194 3380
rect 2727 3376 3313 3383
rect 3847 3376 4203 3383
rect 2193 3367 2207 3373
rect 2333 3367 2347 3373
rect 467 3356 733 3363
rect 1167 3356 1273 3363
rect 1387 3356 1973 3363
rect 2127 3356 2172 3363
rect 2193 3360 2194 3367
rect 2467 3356 2572 3363
rect 2608 3356 2713 3363
rect 2927 3356 3013 3363
rect 3287 3356 3353 3363
rect 3407 3356 3473 3363
rect 3487 3356 3533 3363
rect 3727 3356 3752 3363
rect 3788 3356 3903 3363
rect 3896 3347 3903 3356
rect 4067 3356 4113 3363
rect 4167 3353 4173 3367
rect 4196 3363 4203 3376
rect 4227 3376 4413 3383
rect 4807 3376 4953 3383
rect 5080 3383 5093 3387
rect 5075 3380 5093 3383
rect 5073 3374 5093 3380
rect 5073 3373 5100 3374
rect 5167 3376 5193 3383
rect 5427 3376 5893 3383
rect 5073 3367 5087 3373
rect 4196 3356 4513 3363
rect 4536 3356 4573 3363
rect 107 3336 193 3343
rect 207 3336 253 3343
rect 447 3336 533 3343
rect 987 3336 1013 3343
rect 1027 3336 1353 3343
rect 1887 3336 1933 3343
rect 1947 3336 2093 3343
rect 2267 3336 2333 3343
rect 2507 3336 2633 3343
rect 2767 3336 2803 3343
rect 940 3323 953 3327
rect 927 3316 953 3323
rect 940 3313 953 3316
rect 1547 3316 1613 3323
rect 2327 3316 2393 3323
rect 593 3307 607 3313
rect 1333 3307 1347 3313
rect 2593 3307 2607 3313
rect 2796 3307 2803 3336
rect 3647 3336 3833 3343
rect 3907 3336 4073 3343
rect 4536 3343 4543 3356
rect 4647 3356 4673 3363
rect 4847 3356 4933 3363
rect 4987 3356 5052 3363
rect 5086 3360 5087 3367
rect 5108 3356 5293 3363
rect 5387 3356 5633 3363
rect 5907 3356 5953 3363
rect 6187 3356 6273 3363
rect 6407 3353 6413 3367
rect 4147 3336 4183 3343
rect 3127 3316 3153 3323
rect 4176 3323 4183 3336
rect 4293 3336 4543 3343
rect 4293 3327 4307 3336
rect 4567 3336 4593 3343
rect 4707 3336 4753 3343
rect 4847 3336 5133 3343
rect 5147 3336 5233 3343
rect 5747 3336 5773 3343
rect 6027 3336 6093 3343
rect 6267 3336 6293 3343
rect 4176 3316 4253 3323
rect 67 3296 113 3303
rect 307 3293 313 3307
rect 427 3296 473 3303
rect 647 3296 753 3303
rect 1087 3296 1173 3303
rect 1387 3296 1473 3303
rect 1707 3296 1733 3303
rect 1987 3296 2033 3303
rect 2147 3296 2193 3303
rect 2287 3296 2353 3303
rect 2467 3296 2533 3303
rect 3247 3296 3273 3303
rect 3447 3296 3473 3303
rect 3880 3303 3893 3307
rect 3867 3296 3893 3303
rect 3880 3293 3893 3296
rect 4147 3296 4213 3303
rect 4747 3296 4833 3303
rect 5007 3296 5093 3303
rect 5187 3293 5193 3307
rect 5347 3296 5413 3303
rect 5507 3296 5573 3303
rect 5840 3303 5853 3307
rect 5827 3296 5853 3303
rect 5840 3293 5853 3296
rect 6160 3303 6172 3307
rect 6147 3296 6172 3303
rect 6160 3293 6172 3296
rect 6208 3296 6293 3303
rect 6427 3303 6440 3307
rect 6427 3296 6453 3303
rect 6427 3293 6440 3296
rect 2027 3276 2053 3283
rect 5047 3276 5073 3283
rect 907 3256 973 3263
rect 1527 3256 1573 3263
rect 1687 3256 1733 3263
rect 2187 3253 2193 3267
rect 3647 3253 3653 3267
rect 3727 3256 3813 3263
rect 3987 3256 4052 3263
rect 4088 3253 4093 3267
rect 4480 3263 4492 3267
rect 4467 3256 4492 3263
rect 4480 3253 4492 3256
rect 4528 3253 4533 3267
rect 6407 3256 6433 3263
rect 3373 3247 3387 3253
rect 4273 3247 4287 3253
rect 1227 3236 1313 3243
rect 1807 3236 1873 3243
rect 2007 3236 2073 3243
rect 2787 3236 2883 3243
rect 673 3227 687 3233
rect 987 3213 993 3227
rect 2827 3216 2853 3223
rect 2876 3223 2883 3236
rect 2876 3216 2973 3223
rect 3236 3220 3453 3223
rect 3233 3216 3453 3220
rect 3233 3207 3247 3216
rect 3907 3216 3973 3223
rect 4067 3216 4233 3223
rect 4456 3223 4463 3253
rect 4567 3233 4573 3247
rect 4587 3236 4633 3243
rect 4767 3236 4853 3243
rect 5167 3236 5233 3243
rect 4327 3216 4463 3223
rect 4627 3226 4640 3227
rect 4627 3213 4633 3226
rect 5976 3223 5983 3253
rect 6473 3227 6487 3233
rect 5976 3216 6073 3223
rect 6400 3223 6413 3227
rect 6236 3216 6283 3223
rect 227 3196 273 3203
rect 407 3196 533 3203
rect 1167 3196 1533 3203
rect 1927 3196 2113 3203
rect 2207 3196 2293 3203
rect 2367 3193 2373 3207
rect 2427 3196 2473 3203
rect 2547 3196 2913 3203
rect 3287 3196 3773 3203
rect 4307 3196 4533 3203
rect 4547 3196 4693 3203
rect 4827 3196 5113 3203
rect 5247 3196 5273 3203
rect 5667 3196 5733 3203
rect 5747 3196 5933 3203
rect 6236 3203 6243 3216
rect 6167 3196 6243 3203
rect 6276 3203 6283 3216
rect 6396 3213 6413 3223
rect 6396 3203 6403 3213
rect 6276 3196 6403 3203
rect 147 3176 233 3183
rect 247 3176 633 3183
rect 787 3176 833 3183
rect 1347 3176 1453 3183
rect 2347 3176 2493 3183
rect 2596 3176 2953 3183
rect 673 3167 687 3173
rect 927 3156 953 3163
rect 1167 3156 1473 3163
rect 2596 3163 2603 3176
rect 3307 3176 3373 3183
rect 3467 3176 3653 3183
rect 3936 3176 4333 3183
rect 2027 3156 2603 3163
rect 3207 3156 3513 3163
rect 3936 3163 3943 3176
rect 4387 3176 4453 3183
rect 4587 3176 4793 3183
rect 4807 3176 4973 3183
rect 5047 3173 5053 3187
rect 5267 3176 5413 3183
rect 5427 3176 5563 3183
rect 3607 3156 3943 3163
rect 4127 3156 4173 3163
rect 4887 3156 5013 3163
rect 5087 3156 5153 3163
rect 5407 3156 5453 3163
rect 5556 3163 5563 3176
rect 5587 3176 5753 3183
rect 5767 3176 5893 3183
rect 5556 3156 5673 3163
rect 5827 3156 5853 3163
rect 6007 3156 6193 3163
rect 6367 3156 6513 3163
rect 2387 3136 2453 3143
rect 2527 3136 2893 3143
rect 2967 3136 3753 3143
rect 3927 3136 4163 3143
rect 4156 3127 4163 3136
rect 4367 3136 4683 3143
rect 1147 3116 1353 3123
rect 2627 3116 3793 3123
rect 3847 3116 4053 3123
rect 4167 3116 4593 3123
rect 4640 3123 4653 3127
rect 4636 3113 4653 3123
rect 4676 3123 4683 3136
rect 4707 3136 4933 3143
rect 5067 3136 5393 3143
rect 4676 3116 5773 3123
rect 5887 3116 6033 3123
rect 6107 3116 6233 3123
rect 247 3096 573 3103
rect 827 3096 1253 3103
rect 2227 3096 2253 3103
rect 2507 3093 2512 3107
rect 2548 3096 2573 3103
rect 2827 3096 2913 3103
rect 2967 3096 4393 3103
rect 4636 3103 4643 3113
rect 4527 3096 4643 3103
rect 4707 3096 4913 3103
rect 5007 3096 5033 3103
rect 5827 3096 6353 3103
rect 6467 3093 6472 3107
rect 6508 3093 6513 3107
rect 767 3076 1073 3083
rect 1487 3076 1613 3083
rect 1667 3076 1973 3083
rect 2207 3076 2433 3083
rect 2616 3080 2773 3083
rect 2613 3076 2773 3080
rect 2613 3067 2627 3076
rect 2787 3076 2813 3083
rect 2907 3076 3213 3083
rect 3827 3076 4113 3083
rect 4267 3076 4433 3083
rect 4447 3076 4713 3083
rect 4947 3076 5073 3083
rect 5487 3076 5793 3083
rect 5807 3076 6013 3083
rect 6087 3076 6133 3083
rect 6227 3076 6293 3083
rect 67 3056 93 3063
rect 847 3056 873 3063
rect 947 3056 1393 3063
rect 1587 3056 1693 3063
rect 1787 3056 1913 3063
rect 2347 3056 2373 3063
rect 2427 3056 2452 3063
rect 2488 3056 2513 3063
rect 2667 3056 2953 3063
rect 4067 3056 4173 3063
rect 4227 3056 4293 3063
rect 4307 3056 4453 3063
rect 4467 3056 5013 3063
rect 5207 3056 5373 3063
rect 5387 3056 5533 3063
rect 5727 3056 5873 3063
rect 5987 3053 5993 3067
rect 6167 3056 6213 3063
rect 6327 3056 6373 3063
rect 2136 3036 2233 3043
rect 887 3016 953 3023
rect 1107 3016 1173 3023
rect 1547 3016 1613 3023
rect 2136 3007 2143 3036
rect 2727 3036 2803 3043
rect 2207 3016 2233 3023
rect 2487 3016 2533 3023
rect 2796 3007 2803 3036
rect 2847 3036 2883 3043
rect 2876 3023 2883 3036
rect 3976 3036 4033 3043
rect 2876 3016 2933 3023
rect 3027 3023 3040 3027
rect 3027 3016 3053 3023
rect 3027 3013 3040 3016
rect 3447 3016 3533 3023
rect 3976 3007 3983 3036
rect 4027 3016 4073 3023
rect 4833 3027 4847 3033
rect 4527 3023 4540 3027
rect 4527 3016 4553 3023
rect 4527 3013 4540 3016
rect 4667 3016 4733 3023
rect 6427 3016 6513 3023
rect 167 2996 233 3003
rect 587 3003 600 3007
rect 587 2996 613 3003
rect 587 2993 600 2996
rect 1907 2996 1953 3003
rect 3687 2993 3693 3007
rect 3867 2996 3913 3003
rect 3987 2996 4073 3003
rect 4967 2996 4993 3003
rect 2507 2976 2553 2983
rect 6447 2976 6493 2983
rect 4853 2967 4867 2973
rect 247 2956 293 2963
rect 707 2956 813 2963
rect 960 2963 973 2967
rect 947 2956 973 2963
rect 960 2953 973 2956
rect 1140 2963 1153 2967
rect 1127 2956 1153 2963
rect 1140 2953 1153 2956
rect 1247 2956 1333 2963
rect 1527 2956 1593 2963
rect 2227 2963 2240 2967
rect 2227 2956 2253 2963
rect 2227 2953 2240 2956
rect 2867 2956 2913 2963
rect 3007 2956 3053 2963
rect 3067 2953 3073 2967
rect 3127 2956 3173 2963
rect 3467 2956 3513 2963
rect 3847 2956 3893 2963
rect 4147 2956 4213 2963
rect 4627 2953 4633 2967
rect 5107 2956 5153 2963
rect 5407 2956 5473 2963
rect 5567 2956 5653 2963
rect 5747 2956 5813 2963
rect 5907 2953 5913 2967
rect 5927 2956 5973 2963
rect 6100 2963 6113 2967
rect 6087 2956 6113 2963
rect 6100 2953 6113 2956
rect 6287 2956 6353 2963
rect 347 2916 393 2923
rect 456 2923 463 2953
rect 456 2916 813 2923
rect 867 2916 1093 2923
rect 1376 2923 1383 2953
rect 1107 2916 1653 2923
rect 1676 2923 1683 2953
rect 1747 2936 1773 2943
rect 1676 2916 1813 2923
rect 1836 2923 1843 2953
rect 2593 2947 2607 2953
rect 1836 2916 2733 2923
rect 2813 2923 2827 2933
rect 2813 2916 3213 2923
rect 3516 2923 3523 2953
rect 4273 2947 4287 2953
rect 3516 2916 3653 2923
rect 4416 2923 4423 2953
rect 4847 2936 4873 2943
rect 4416 2916 4533 2923
rect 4587 2916 4653 2923
rect 4707 2916 4732 2923
rect 4768 2916 4833 2923
rect 4936 2923 4943 2953
rect 4993 2947 5007 2953
rect 5233 2947 5247 2953
rect 6193 2947 6207 2953
rect 5947 2936 6003 2943
rect 4936 2916 5413 2923
rect 5427 2916 5473 2923
rect 5487 2916 5693 2923
rect 5807 2916 5853 2923
rect 5996 2923 6003 2936
rect 5996 2916 6033 2923
rect 6247 2916 6273 2923
rect 6367 2916 6393 2923
rect 267 2896 553 2903
rect 807 2896 933 2903
rect 1067 2896 1113 2903
rect 2087 2896 2453 2903
rect 2526 2893 2527 2900
rect 2548 2893 2553 2907
rect 2727 2896 2973 2903
rect 3447 2896 3493 2903
rect 3587 2896 3613 2903
rect 3627 2896 3933 2903
rect 4267 2896 4353 2903
rect 4527 2896 4553 2903
rect 4607 2896 4813 2903
rect 4866 2893 4867 2900
rect 4888 2896 5073 2903
rect 5167 2896 5353 2903
rect 5367 2896 5513 2903
rect 5887 2896 5973 2903
rect 6127 2893 6132 2907
rect 6168 2893 6173 2907
rect 6267 2896 6293 2903
rect 2513 2887 2527 2893
rect 467 2876 1013 2883
rect 1027 2876 1073 2883
rect 1347 2876 1633 2883
rect 1647 2876 1733 2883
rect 1747 2876 2093 2883
rect 2267 2876 2393 2883
rect 2607 2876 2773 2883
rect 2907 2876 3153 2883
rect 3207 2876 3263 2883
rect 507 2856 1113 2863
rect 2367 2856 2413 2863
rect 3047 2856 3233 2863
rect 3256 2863 3263 2876
rect 3287 2876 3773 2883
rect 4087 2876 4493 2883
rect 4853 2883 4867 2893
rect 6367 2896 6453 2903
rect 4547 2876 5053 2883
rect 5127 2876 5193 2883
rect 5267 2876 5433 2883
rect 5487 2876 5573 2883
rect 5587 2876 5733 2883
rect 5987 2876 6293 2883
rect 6307 2876 6413 2883
rect 3256 2856 3533 2863
rect 3587 2856 3853 2863
rect 3907 2856 4283 2863
rect 187 2836 573 2843
rect 907 2836 953 2843
rect 967 2836 1553 2843
rect 1607 2836 1693 2843
rect 1707 2836 2073 2843
rect 2267 2836 2313 2843
rect 2387 2836 2593 2843
rect 2707 2836 2733 2843
rect 3127 2836 3273 2843
rect 4276 2843 4283 2856
rect 4407 2856 4593 2863
rect 4707 2856 4792 2863
rect 4828 2856 4873 2863
rect 5087 2856 5593 2863
rect 6007 2856 6313 2863
rect 3507 2836 3903 2843
rect 4276 2836 4452 2843
rect 267 2816 313 2823
rect 407 2816 613 2823
rect 1787 2816 1833 2823
rect 1987 2816 2013 2823
rect 2027 2816 2133 2823
rect 2287 2816 2312 2823
rect 753 2807 767 2813
rect 2348 2816 2453 2823
rect 2616 2816 2713 2823
rect 1553 2787 1567 2793
rect 1993 2787 2007 2793
rect 2616 2787 2623 2816
rect 3527 2816 3713 2823
rect 3767 2816 3853 2823
rect 3896 2823 3903 2836
rect 4488 2840 4683 2843
rect 4488 2836 4687 2840
rect 4673 2827 4687 2836
rect 4927 2836 4993 2843
rect 5007 2833 5013 2847
rect 5167 2836 5213 2843
rect 5587 2836 5633 2843
rect 5847 2836 5973 2843
rect 5987 2836 6193 2843
rect 6347 2836 6393 2843
rect 3896 2816 4293 2823
rect 4587 2816 4633 2823
rect 4747 2816 4793 2823
rect 4907 2816 4953 2823
rect 4996 2816 5133 2823
rect 4147 2796 4173 2803
rect 4053 2787 4067 2793
rect 4996 2787 5003 2816
rect 5407 2816 5432 2823
rect 5468 2816 5573 2823
rect 6207 2816 6313 2823
rect 6327 2816 6353 2823
rect 6173 2787 6187 2793
rect 387 2776 453 2783
rect 507 2773 513 2787
rect 607 2776 693 2783
rect 747 2776 833 2783
rect 1107 2776 1172 2783
rect 1387 2776 1493 2783
rect 1900 2783 1913 2787
rect 1887 2776 1913 2783
rect 1900 2773 1913 2776
rect 2207 2776 2253 2783
rect 2380 2783 2393 2787
rect 2367 2776 2393 2783
rect 2380 2773 2393 2776
rect 2800 2783 2813 2787
rect 2787 2776 2813 2783
rect 2800 2773 2813 2776
rect 3527 2776 3573 2783
rect 3587 2776 3633 2783
rect 4247 2776 4353 2783
rect 4407 2776 4473 2783
rect 4860 2783 4873 2787
rect 4847 2776 4873 2783
rect 4860 2773 4873 2776
rect 5147 2776 5253 2783
rect 5507 2776 5553 2783
rect 5607 2783 5620 2787
rect 5607 2776 5633 2783
rect 5607 2773 5620 2776
rect 5727 2776 5793 2783
rect 6027 2773 6033 2787
rect 6387 2776 6433 2783
rect 4707 2756 4753 2763
rect 4900 2763 4913 2767
rect 4896 2753 4913 2763
rect 5887 2756 5933 2763
rect 127 2736 193 2743
rect 747 2733 753 2747
rect 1727 2736 1773 2743
rect 3667 2736 3713 2743
rect 3907 2736 3973 2743
rect 4087 2736 4133 2743
rect 4567 2736 4633 2743
rect 4896 2743 4903 2753
rect 4867 2736 4903 2743
rect 5347 2736 5393 2743
rect 247 2716 313 2723
rect 627 2716 673 2723
rect 907 2716 973 2723
rect 2267 2723 2280 2727
rect 2267 2716 2293 2723
rect 2267 2713 2280 2716
rect 2387 2716 2473 2723
rect 107 2696 133 2703
rect 296 2696 333 2703
rect 296 2683 303 2696
rect 207 2676 303 2683
rect 327 2676 533 2683
rect 647 2676 813 2683
rect 1087 2676 1213 2683
rect 1236 2683 1243 2713
rect 2687 2696 2733 2703
rect 3216 2703 3223 2733
rect 3547 2716 3593 2723
rect 4347 2723 4360 2727
rect 4347 2716 4373 2723
rect 4347 2713 4360 2716
rect 4427 2713 4433 2727
rect 4687 2716 4733 2723
rect 3147 2696 3203 2703
rect 3216 2696 3293 2703
rect 1236 2676 1393 2683
rect 1827 2676 1973 2683
rect 2027 2676 2113 2683
rect 2167 2676 2293 2683
rect 2316 2676 2393 2683
rect 1187 2656 1353 2663
rect 1376 2656 1933 2663
rect 547 2636 1073 2643
rect 1207 2636 1293 2643
rect 1376 2643 1383 2656
rect 2067 2656 2193 2663
rect 2316 2663 2323 2676
rect 2527 2676 2793 2683
rect 3196 2683 3203 2696
rect 4516 2696 4643 2703
rect 3196 2676 3253 2683
rect 3507 2673 3513 2687
rect 3727 2676 3813 2683
rect 3867 2676 4113 2683
rect 4187 2676 4233 2683
rect 4247 2676 4263 2683
rect 2247 2656 2323 2663
rect 2347 2656 2693 2663
rect 3056 2656 3173 2663
rect 1307 2636 1383 2643
rect 1427 2636 1553 2643
rect 1867 2636 1993 2643
rect 2127 2636 2753 2643
rect 3056 2643 3063 2656
rect 3496 2656 4053 2663
rect 2847 2636 3063 2643
rect 3107 2636 3433 2643
rect 3496 2643 3503 2656
rect 4256 2667 4263 2676
rect 4287 2676 4432 2683
rect 4516 2683 4523 2696
rect 4468 2676 4523 2683
rect 4547 2683 4560 2687
rect 4636 2683 4643 2696
rect 4547 2680 4563 2683
rect 4547 2673 4567 2680
rect 4636 2676 4853 2683
rect 4907 2676 5093 2683
rect 5167 2676 5273 2683
rect 5827 2676 5993 2683
rect 6307 2676 6353 2683
rect 4553 2667 4567 2673
rect 4147 2656 4173 2663
rect 4187 2656 4213 2663
rect 4256 2666 4280 2667
rect 4256 2656 4273 2666
rect 4260 2653 4273 2656
rect 4687 2656 4933 2663
rect 5047 2656 5253 2663
rect 5667 2656 5853 2663
rect 3456 2636 3503 2643
rect 1067 2616 1433 2623
rect 1447 2616 1873 2623
rect 1947 2616 2393 2623
rect 2547 2616 2573 2623
rect 2647 2616 2692 2623
rect 2728 2616 2893 2623
rect 3267 2616 3313 2623
rect 3456 2623 3463 2636
rect 3947 2636 4013 2643
rect 4067 2636 4132 2643
rect 4168 2636 4233 2643
rect 4527 2636 4613 2643
rect 4887 2636 5113 2643
rect 5127 2636 5313 2643
rect 5587 2636 5633 2643
rect 5727 2636 6513 2643
rect 3327 2616 3463 2623
rect 3687 2616 3744 2623
rect 1287 2596 1533 2603
rect 1707 2596 3093 2603
rect 3527 2596 3653 2603
rect 3737 2587 3744 2616
rect 4127 2616 4193 2623
rect 4407 2616 4473 2623
rect 4487 2616 4693 2623
rect 4747 2616 4873 2623
rect 5407 2616 5433 2623
rect 5967 2616 6413 2623
rect 3807 2596 4153 2603
rect 4307 2596 4593 2603
rect 4787 2596 4933 2603
rect 5327 2596 5413 2603
rect 5787 2596 5973 2603
rect 6107 2596 6133 2603
rect 507 2576 893 2583
rect 947 2576 973 2583
rect 1267 2576 1333 2583
rect 1347 2576 1373 2583
rect 1387 2576 2243 2583
rect 2236 2567 2243 2576
rect 2407 2573 2412 2587
rect 2448 2576 2493 2583
rect 2567 2576 2793 2583
rect 2816 2576 3063 2583
rect 147 2556 333 2563
rect 347 2556 793 2563
rect 996 2556 1193 2563
rect 187 2536 293 2543
rect 687 2536 773 2543
rect 787 2536 853 2543
rect 996 2543 1003 2556
rect 1407 2556 1433 2563
rect 2147 2556 2212 2563
rect 2248 2556 2353 2563
rect 2407 2556 2553 2563
rect 2816 2563 2823 2576
rect 3056 2567 3063 2576
rect 3167 2576 3712 2583
rect 3787 2576 3913 2583
rect 4047 2576 4113 2583
rect 4207 2573 4213 2587
rect 4467 2576 4553 2583
rect 4647 2576 4733 2583
rect 4827 2576 5093 2583
rect 5147 2576 5212 2583
rect 5248 2576 5373 2583
rect 5427 2576 5573 2583
rect 6087 2576 6293 2583
rect 2567 2556 2823 2563
rect 2867 2560 2963 2563
rect 2867 2556 2967 2560
rect 947 2536 1003 2543
rect 1027 2536 1153 2543
rect 1396 2543 1403 2553
rect 2953 2547 2967 2556
rect 3067 2556 3113 2563
rect 3207 2556 3753 2563
rect 3767 2556 3973 2563
rect 4087 2556 4153 2563
rect 4216 2563 4223 2573
rect 4216 2556 4613 2563
rect 4627 2556 4973 2563
rect 5207 2556 5613 2563
rect 6167 2556 6213 2563
rect 1227 2536 1403 2543
rect 1767 2536 1973 2543
rect 1987 2536 2013 2543
rect 2067 2536 2373 2543
rect 2427 2536 2613 2543
rect 2667 2536 2713 2543
rect 2827 2536 2913 2543
rect 3367 2536 3532 2543
rect 3568 2533 3572 2547
rect 3608 2536 3853 2543
rect 3927 2536 4073 2543
rect 4327 2536 4373 2543
rect 4427 2536 4493 2543
rect 4647 2536 4712 2543
rect 4748 2536 4913 2543
rect 4927 2536 5173 2543
rect 5216 2536 5513 2543
rect 1147 2516 1203 2523
rect 1196 2487 1203 2516
rect 1327 2516 1403 2523
rect 1396 2487 1403 2516
rect 2176 2516 2433 2523
rect 2176 2487 2183 2516
rect 2547 2513 2553 2527
rect 3647 2516 3753 2523
rect 4927 2516 4993 2523
rect 5107 2514 5113 2527
rect 5100 2513 5113 2514
rect 5216 2507 5223 2536
rect 5647 2536 5793 2543
rect 5927 2536 6033 2543
rect 6047 2536 6233 2543
rect 5516 2523 5523 2533
rect 5516 2516 5733 2523
rect 2387 2493 2393 2507
rect 3420 2503 3432 2507
rect 3407 2496 3432 2503
rect 3420 2493 3432 2496
rect 3468 2496 3533 2503
rect 3547 2496 3633 2503
rect 3747 2496 3793 2503
rect 3927 2493 3933 2507
rect 4207 2496 4253 2503
rect 4727 2496 4793 2503
rect 5107 2496 5133 2503
rect 5867 2496 5933 2503
rect 6327 2496 6393 2503
rect 827 2476 913 2483
rect 1447 2476 1513 2483
rect 1927 2476 1973 2483
rect 2107 2476 2173 2483
rect 2287 2476 2333 2483
rect 3167 2476 3233 2483
rect 3667 2473 3673 2487
rect 4567 2476 4633 2483
rect 2447 2453 2453 2467
rect 5076 2456 5113 2463
rect 107 2433 113 2447
rect 207 2436 273 2443
rect 367 2436 433 2443
rect 627 2436 673 2443
rect 780 2443 793 2447
rect 767 2436 793 2443
rect 780 2433 793 2436
rect 987 2436 1013 2443
rect 1027 2433 1033 2447
rect 1587 2433 1593 2447
rect 2027 2433 2033 2447
rect 2107 2436 2153 2443
rect 2427 2436 2493 2443
rect 2627 2433 2633 2447
rect 3487 2443 3500 2447
rect 3487 2436 3513 2443
rect 3527 2436 3592 2443
rect 3487 2433 3500 2436
rect 3628 2433 3633 2447
rect 3827 2436 3873 2443
rect 3947 2433 3953 2447
rect 3967 2436 4033 2443
rect 4127 2433 4133 2447
rect 4407 2433 4413 2447
rect 4707 2436 4773 2443
rect 4867 2436 4933 2443
rect 5076 2443 5083 2456
rect 5047 2436 5083 2443
rect 5107 2436 5193 2443
rect 5347 2436 5413 2443
rect 5907 2433 5913 2447
rect 5987 2436 6053 2443
rect 113 2427 127 2433
rect 1733 2427 1747 2433
rect 2953 2427 2967 2433
rect 3093 2427 3107 2433
rect 4813 2427 4827 2433
rect 5293 2427 5307 2433
rect 6247 2436 6293 2443
rect 3747 2416 3773 2423
rect 4906 2413 4907 2420
rect 2133 2407 2147 2413
rect 167 2396 313 2403
rect 327 2396 352 2403
rect 388 2396 453 2403
rect 467 2396 573 2403
rect 1467 2396 1853 2403
rect 1927 2396 1993 2403
rect 2207 2396 2273 2403
rect 2327 2396 2413 2403
rect 2487 2396 3193 2403
rect 3307 2396 3433 2403
rect 3447 2393 3453 2407
rect 3527 2396 3572 2403
rect 3608 2396 4053 2403
rect 4067 2396 4333 2403
rect 4487 2396 4613 2403
rect 4727 2396 4753 2403
rect 4767 2396 4833 2403
rect 4893 2403 4907 2413
rect 4847 2400 4907 2403
rect 4913 2413 4914 2420
rect 5107 2416 5133 2423
rect 4913 2407 4927 2413
rect 4847 2396 4902 2400
rect 4967 2396 5033 2403
rect 5127 2396 5353 2403
rect 5507 2396 5533 2403
rect 5727 2396 5773 2403
rect 6127 2393 6193 2400
rect 487 2376 533 2383
rect 696 2376 813 2383
rect 427 2356 593 2363
rect 696 2363 703 2376
rect 1767 2376 1813 2383
rect 2236 2376 2413 2383
rect 607 2356 703 2363
rect 1107 2356 1273 2363
rect 2236 2363 2243 2376
rect 2547 2376 2573 2383
rect 2667 2376 2833 2383
rect 2880 2383 2892 2387
rect 2876 2373 2892 2383
rect 2928 2376 3093 2383
rect 3167 2376 3473 2383
rect 3567 2376 3713 2383
rect 3767 2376 4113 2383
rect 4227 2376 4253 2383
rect 4307 2373 4313 2387
rect 4467 2376 4653 2383
rect 4707 2376 5433 2383
rect 5807 2376 5853 2383
rect 6167 2376 6213 2383
rect 1567 2356 2243 2363
rect 2267 2356 2433 2363
rect 2447 2356 2613 2363
rect 2876 2363 2883 2373
rect 2627 2356 2883 2363
rect 2896 2356 3093 2363
rect 807 2336 893 2343
rect 907 2336 1013 2343
rect 1036 2336 1193 2343
rect 1036 2327 1043 2336
rect 1207 2336 1373 2343
rect 1387 2336 1833 2343
rect 1847 2336 2193 2343
rect 2427 2336 2553 2343
rect 2896 2343 2903 2356
rect 3196 2360 3653 2363
rect 3193 2356 3653 2360
rect 2567 2336 2903 2343
rect 2916 2336 3153 2343
rect 787 2316 853 2323
rect 867 2316 933 2323
rect 1020 2326 1043 2327
rect 1027 2316 1043 2326
rect 1027 2313 1040 2316
rect 1067 2316 1233 2323
rect 1507 2316 1692 2323
rect 1728 2316 1793 2323
rect 1907 2316 2332 2323
rect 2368 2316 2473 2323
rect 2607 2316 2733 2323
rect 2916 2323 2923 2336
rect 3193 2347 3207 2356
rect 3667 2356 4013 2363
rect 4087 2356 4193 2363
rect 4296 2356 4533 2363
rect 3207 2336 3313 2343
rect 4296 2343 4303 2356
rect 4987 2356 5153 2363
rect 5307 2356 5453 2363
rect 5467 2356 5613 2363
rect 5847 2356 6033 2363
rect 3727 2336 4303 2343
rect 4347 2336 4373 2343
rect 4427 2336 5113 2343
rect 5156 2343 5163 2353
rect 5156 2336 5313 2343
rect 5607 2336 5653 2343
rect 5716 2340 6213 2343
rect 5713 2336 6213 2340
rect 2827 2316 2923 2323
rect 5713 2327 5727 2336
rect 3007 2316 3153 2323
rect 3267 2316 3373 2323
rect 3387 2316 3413 2323
rect 3427 2316 3593 2323
rect 3927 2316 3973 2323
rect 4247 2316 4433 2323
rect 4607 2316 4813 2323
rect 4827 2316 4853 2323
rect 4867 2316 4993 2323
rect 5107 2316 5173 2323
rect 5227 2316 5253 2323
rect 5347 2316 5433 2323
rect 5767 2316 5893 2323
rect 6047 2316 6233 2323
rect 6247 2316 6313 2323
rect 567 2296 743 2303
rect 736 2267 743 2296
rect 1227 2296 1353 2303
rect 1367 2296 1473 2303
rect 1487 2296 1593 2303
rect 1647 2296 1733 2303
rect 2216 2296 2293 2303
rect 2216 2283 2223 2296
rect 2647 2296 2713 2303
rect 2807 2296 2833 2303
rect 2887 2296 2993 2303
rect 3067 2296 3113 2303
rect 3667 2296 3773 2303
rect 4347 2296 4513 2303
rect 4947 2296 5193 2303
rect 5247 2296 5373 2303
rect 5687 2296 5873 2303
rect 5887 2296 6003 2303
rect 2187 2276 2223 2283
rect 3447 2276 3553 2283
rect 3647 2276 3693 2283
rect 2853 2267 2867 2273
rect 5833 2267 5847 2273
rect 5996 2267 6003 2296
rect 6187 2296 6273 2303
rect 6387 2296 6433 2303
rect 6213 2267 6227 2273
rect 147 2253 153 2267
rect 507 2256 573 2263
rect 587 2256 633 2263
rect 947 2256 1033 2263
rect 1407 2256 1453 2263
rect 1547 2256 1633 2263
rect 1700 2263 1713 2267
rect 1687 2256 1713 2263
rect 1700 2253 1713 2256
rect 2107 2253 2113 2267
rect 2307 2256 2393 2263
rect 2667 2253 2673 2267
rect 2927 2256 3033 2263
rect 3267 2256 3293 2263
rect 3467 2256 3513 2263
rect 4127 2256 4213 2263
rect 4367 2256 4413 2263
rect 4507 2256 4573 2263
rect 4907 2256 4953 2263
rect 5047 2256 5113 2263
rect 5207 2256 5273 2263
rect 5287 2256 5333 2263
rect 5427 2256 5493 2263
rect 5627 2256 5693 2263
rect 6267 2256 6333 2263
rect 4747 2236 4773 2243
rect 827 2216 873 2223
rect 3107 2216 3173 2223
rect 3847 2216 3913 2223
rect 4087 2216 4133 2223
rect 127 2196 213 2203
rect 1307 2203 1320 2207
rect 1307 2196 1333 2203
rect 1307 2193 1320 2196
rect 1680 2203 1693 2207
rect 1667 2196 1693 2203
rect 1680 2193 1693 2196
rect 1947 2196 2033 2203
rect 2247 2196 2333 2203
rect 2547 2196 2633 2203
rect 253 2187 267 2193
rect 3356 2183 3363 2213
rect 3107 2176 3363 2183
rect 3407 2176 3433 2183
rect 3447 2176 3533 2183
rect 3576 2183 3583 2213
rect 3753 2207 3767 2213
rect 4633 2207 4647 2213
rect 4467 2193 4473 2207
rect 5487 2196 5553 2203
rect 3576 2176 3673 2183
rect 3807 2176 4113 2183
rect 5347 2176 5373 2183
rect 447 2156 553 2163
rect 627 2156 713 2163
rect 727 2156 1133 2163
rect 1207 2156 1313 2163
rect 1407 2156 1693 2163
rect 1827 2156 1953 2163
rect 2147 2156 2433 2163
rect 2456 2156 2693 2163
rect 1196 2143 1203 2153
rect 1047 2136 1203 2143
rect 1487 2136 1713 2143
rect 2127 2136 2352 2143
rect 2456 2143 2463 2156
rect 2707 2156 2913 2163
rect 3007 2156 3353 2163
rect 3947 2156 4353 2163
rect 4507 2156 4973 2163
rect 5207 2156 5533 2163
rect 6167 2156 6253 2163
rect 6307 2156 6393 2163
rect 6407 2156 6513 2163
rect 2388 2136 2463 2143
rect 2667 2136 2853 2143
rect 2907 2136 3013 2143
rect 3027 2136 3093 2143
rect 3207 2136 3263 2143
rect 727 2116 913 2123
rect 927 2116 1393 2123
rect 1447 2116 2053 2123
rect 2316 2116 2393 2123
rect 287 2096 573 2103
rect 587 2096 813 2103
rect 1436 2103 1443 2113
rect 907 2096 1443 2103
rect 2316 2103 2323 2116
rect 2627 2116 2673 2123
rect 2847 2116 3103 2123
rect 1707 2096 2323 2103
rect 2347 2096 2733 2103
rect 2807 2096 2923 2103
rect 887 2076 972 2083
rect 1008 2076 1563 2083
rect 987 2056 1093 2063
rect 1556 2063 1563 2076
rect 1667 2076 2313 2083
rect 2367 2076 2533 2083
rect 2547 2076 2633 2083
rect 2707 2076 2773 2083
rect 2916 2083 2923 2096
rect 2987 2096 3053 2103
rect 3096 2103 3103 2116
rect 3167 2116 3233 2123
rect 3256 2123 3263 2136
rect 3287 2136 3433 2143
rect 3527 2136 3653 2143
rect 4007 2136 4053 2143
rect 4147 2136 4193 2143
rect 4327 2136 4453 2143
rect 4567 2136 4633 2143
rect 4647 2136 4833 2143
rect 4927 2136 5093 2143
rect 5116 2136 5433 2143
rect 3256 2116 3452 2123
rect 3488 2116 3553 2123
rect 3667 2116 3753 2123
rect 3767 2116 3893 2123
rect 4136 2123 4143 2133
rect 4047 2116 4143 2123
rect 4247 2116 4492 2123
rect 4528 2116 4613 2123
rect 4687 2116 4733 2123
rect 4907 2116 4973 2123
rect 5116 2123 5123 2136
rect 5507 2136 5533 2143
rect 5907 2136 5953 2143
rect 6156 2143 6163 2153
rect 6027 2136 6163 2143
rect 5027 2116 5123 2123
rect 5147 2116 5473 2123
rect 5487 2116 5693 2123
rect 6067 2116 6173 2123
rect 6187 2116 6233 2123
rect 3096 2096 3463 2103
rect 3456 2087 3463 2096
rect 4236 2103 4243 2113
rect 3547 2096 4243 2103
rect 4607 2096 4713 2103
rect 4947 2096 5253 2103
rect 5387 2096 5593 2103
rect 2916 2076 3413 2083
rect 3467 2076 3613 2083
rect 3727 2076 3833 2083
rect 4367 2076 5013 2083
rect 5447 2076 5513 2083
rect 5627 2076 5733 2083
rect 4173 2067 4187 2073
rect 1556 2056 2593 2063
rect 2687 2056 2732 2063
rect 2768 2056 2813 2063
rect 3027 2056 3213 2063
rect 3227 2056 3493 2063
rect 3647 2056 3773 2063
rect 4427 2053 4432 2067
rect 4468 2056 4733 2063
rect 4827 2056 5072 2063
rect 5108 2056 5193 2063
rect 5247 2053 5253 2067
rect 5427 2056 5493 2063
rect 5567 2056 5713 2063
rect 5807 2056 5853 2063
rect 127 2036 613 2043
rect 1147 2036 1253 2043
rect 1267 2036 2013 2043
rect 2067 2036 2723 2043
rect 447 2016 533 2023
rect 547 2016 673 2023
rect 687 2016 793 2023
rect 947 2016 1172 2023
rect 1208 2016 1293 2023
rect 1687 2016 1813 2023
rect 1967 2016 2033 2023
rect 2227 2016 2293 2023
rect 2587 2016 2693 2023
rect 2716 2023 2723 2036
rect 2847 2033 2853 2047
rect 2927 2036 3933 2043
rect 4047 2036 4113 2043
rect 4207 2036 4513 2043
rect 4587 2036 4653 2043
rect 4667 2036 4752 2043
rect 4788 2036 4853 2043
rect 4967 2036 5813 2043
rect 6367 2036 6433 2043
rect 2716 2016 3313 2023
rect 3367 2016 3393 2023
rect 3447 2016 3513 2023
rect 4147 2016 4253 2023
rect 4387 2016 4413 2023
rect 4467 2016 4493 2023
rect 4627 2016 5003 2023
rect 2187 1996 2233 2003
rect 2487 1996 2573 2003
rect 2867 1996 3133 2003
rect 3156 1996 3253 2003
rect 107 1976 193 1983
rect 347 1976 413 1983
rect 1007 1976 1093 1983
rect 3156 1967 3163 1996
rect 4867 1996 4933 2003
rect 4996 2003 5003 2016
rect 5067 2016 5113 2023
rect 5187 2016 5233 2023
rect 5307 2016 5453 2023
rect 5508 2016 5653 2023
rect 5907 2013 6113 2020
rect 6207 2016 6273 2023
rect 6327 2016 6413 2023
rect 4996 1996 5073 2003
rect 4007 1976 4033 1983
rect 4367 1976 4433 1983
rect 4827 1976 4873 1983
rect 4953 1967 4967 1973
rect 5213 1967 5227 1973
rect 667 1956 733 1963
rect 1567 1956 1613 1963
rect 1887 1953 1893 1967
rect 2187 1956 2273 1963
rect 2447 1963 2460 1967
rect 2447 1956 2473 1963
rect 2447 1953 2460 1956
rect 3107 1953 3113 1967
rect 4247 1956 4313 1963
rect 5007 1956 5053 1963
rect 5240 1963 5253 1967
rect 5236 1953 5253 1963
rect 1667 1936 1733 1943
rect 2747 1933 2753 1947
rect 3267 1934 3273 1947
rect 3267 1933 3280 1934
rect 3707 1936 3733 1943
rect 5236 1947 5243 1953
rect 6127 1953 6213 1960
rect 4147 1936 4173 1943
rect 4767 1936 4793 1943
rect 5227 1936 5243 1947
rect 5227 1933 5240 1936
rect 807 1916 873 1923
rect 1167 1916 1233 1923
rect 1327 1916 1413 1923
rect 233 1907 247 1913
rect 207 1876 273 1883
rect 556 1883 563 1913
rect 447 1876 563 1883
rect 1116 1883 1123 1913
rect 1453 1907 1467 1913
rect 2067 1913 2073 1927
rect 2347 1916 2453 1923
rect 2627 1923 2640 1927
rect 2627 1916 2653 1923
rect 2627 1913 2640 1916
rect 2807 1913 2813 1927
rect 2987 1913 2993 1927
rect 3287 1916 3333 1923
rect 3647 1916 3733 1923
rect 3227 1896 3293 1903
rect 1116 1876 1493 1883
rect 1747 1876 2013 1883
rect 2587 1876 3003 1883
rect 327 1856 473 1863
rect 767 1856 1073 1863
rect 1607 1856 1833 1863
rect 1847 1856 2293 1863
rect 2607 1856 2773 1863
rect 2996 1867 3003 1876
rect 3247 1876 3373 1883
rect 3476 1883 3483 1913
rect 3827 1916 3893 1923
rect 3947 1916 4013 1923
rect 4107 1916 4173 1923
rect 4507 1916 4553 1923
rect 4687 1913 4693 1927
rect 5187 1913 5193 1927
rect 5427 1913 5433 1927
rect 5527 1923 5540 1927
rect 5527 1916 5553 1923
rect 5527 1913 5540 1916
rect 5667 1916 5713 1923
rect 5967 1916 6053 1923
rect 5913 1907 5927 1913
rect 6387 1916 6433 1923
rect 4280 1903 4293 1907
rect 4267 1896 4293 1903
rect 4280 1893 4293 1896
rect 4573 1887 4587 1893
rect 3476 1876 3593 1883
rect 3607 1876 3693 1883
rect 3847 1876 3913 1883
rect 4027 1876 4073 1883
rect 4427 1876 4513 1883
rect 4627 1876 4833 1883
rect 5087 1876 5153 1883
rect 5227 1873 5233 1887
rect 5247 1876 5273 1883
rect 5467 1876 5733 1883
rect 6147 1876 6253 1883
rect 6427 1876 6493 1883
rect 2787 1856 2853 1863
rect 3007 1856 3133 1863
rect 3207 1856 3253 1863
rect 3427 1856 3493 1863
rect 3647 1856 3773 1863
rect 3827 1856 3993 1863
rect 4187 1856 4292 1863
rect 4313 1853 4314 1860
rect 4567 1856 4633 1863
rect 4676 1856 4933 1863
rect 1287 1836 1733 1843
rect 1787 1836 1953 1843
rect 2027 1836 2153 1843
rect 2547 1836 2713 1843
rect 2787 1836 2913 1843
rect 3107 1836 3333 1843
rect 3527 1836 3843 1843
rect 247 1816 332 1823
rect 368 1816 493 1823
rect 507 1816 613 1823
rect 627 1816 793 1823
rect 807 1816 933 1823
rect 1227 1816 1653 1823
rect 1696 1820 2173 1823
rect 1693 1816 2173 1820
rect 1693 1807 1707 1816
rect 2407 1816 3033 1823
rect 3127 1816 3813 1823
rect 207 1793 213 1807
rect 407 1796 543 1803
rect 536 1787 543 1796
rect 1347 1796 1533 1803
rect 1747 1796 1913 1803
rect 2067 1796 2093 1803
rect 2187 1796 2953 1803
rect 3027 1796 3053 1803
rect 3107 1793 3112 1807
rect 3148 1796 3193 1803
rect 3247 1796 3373 1803
rect 3396 1796 3533 1803
rect 127 1776 193 1783
rect 547 1776 653 1783
rect 667 1776 813 1783
rect 1387 1773 1393 1787
rect 1456 1776 1553 1783
rect 1273 1747 1287 1753
rect 1456 1747 1463 1776
rect 1647 1776 1692 1783
rect 1728 1776 1773 1783
rect 1827 1776 1853 1783
rect 1956 1776 2033 1783
rect 1593 1747 1607 1753
rect 1956 1747 1963 1776
rect 2047 1776 2192 1783
rect 2228 1773 2233 1787
rect 2387 1776 2573 1783
rect 2647 1776 2692 1783
rect 2728 1776 2923 1783
rect 2593 1747 2607 1753
rect 2753 1747 2767 1753
rect 2916 1747 2923 1776
rect 3147 1776 3253 1783
rect 3396 1783 3403 1796
rect 3687 1796 3753 1803
rect 3836 1803 3843 1836
rect 4033 1843 4047 1853
rect 3947 1840 4047 1843
rect 3947 1836 4043 1840
rect 4313 1843 4327 1853
rect 4287 1840 4327 1843
rect 4287 1836 4323 1840
rect 4676 1843 4683 1856
rect 4976 1856 5093 1863
rect 4976 1847 4983 1856
rect 5247 1853 5253 1867
rect 5607 1856 5793 1863
rect 6047 1856 6313 1863
rect 4347 1836 4683 1843
rect 4707 1836 4833 1843
rect 4887 1836 4973 1843
rect 5027 1836 5313 1843
rect 5327 1836 5453 1843
rect 6107 1836 6193 1843
rect 6307 1836 6453 1843
rect 3907 1816 4033 1823
rect 4087 1816 4213 1823
rect 4487 1816 4773 1823
rect 4787 1816 5373 1823
rect 5587 1816 5753 1823
rect 5767 1816 6153 1823
rect 6167 1816 6453 1823
rect 3836 1796 3863 1803
rect 3856 1787 3863 1796
rect 3887 1796 4333 1803
rect 4376 1796 4693 1803
rect 4376 1787 4383 1796
rect 4707 1796 4793 1803
rect 4847 1796 5013 1803
rect 5087 1796 5133 1803
rect 5207 1796 5353 1803
rect 5367 1796 5493 1803
rect 5807 1796 6193 1803
rect 6316 1796 6473 1803
rect 6316 1787 6323 1796
rect 3307 1776 3403 1783
rect 3487 1776 3573 1783
rect 3707 1776 3843 1783
rect 3856 1776 3873 1787
rect 3407 1756 3433 1763
rect 3836 1763 3843 1776
rect 3860 1773 3873 1776
rect 3927 1773 3933 1787
rect 4267 1776 4373 1783
rect 4447 1776 4593 1783
rect 4616 1776 4753 1783
rect 3833 1756 3913 1763
rect 3833 1747 3847 1756
rect 4427 1756 4453 1763
rect 4616 1763 4623 1776
rect 4836 1776 4973 1783
rect 4567 1756 4623 1763
rect 247 1736 313 1743
rect 527 1736 573 1743
rect 927 1736 993 1743
rect 1747 1743 1760 1747
rect 1747 1736 1773 1743
rect 1747 1733 1760 1736
rect 2047 1736 2113 1743
rect 2187 1736 2253 1743
rect 2447 1736 2493 1743
rect 2820 1743 2833 1747
rect 2807 1736 2833 1743
rect 2820 1733 2833 1736
rect 3387 1736 3473 1743
rect 3747 1736 3793 1743
rect 3887 1736 3973 1743
rect 3987 1736 4073 1743
rect 4287 1736 4333 1743
rect 4836 1747 4843 1776
rect 4987 1776 5053 1783
rect 5107 1776 5343 1783
rect 5336 1747 5343 1776
rect 5487 1776 5573 1783
rect 5747 1776 6123 1783
rect 6116 1747 6123 1776
rect 6247 1776 6313 1783
rect 6427 1776 6493 1783
rect 6453 1747 6467 1753
rect 4527 1733 4532 1747
rect 4568 1736 4653 1743
rect 5547 1733 5553 1747
rect 5847 1736 5933 1743
rect 6207 1736 6253 1743
rect 6307 1736 6413 1743
rect 193 1727 207 1733
rect 2667 1716 2713 1723
rect 3367 1716 3393 1723
rect 387 1696 453 1703
rect 687 1696 733 1703
rect 880 1703 893 1707
rect 867 1696 893 1703
rect 880 1693 893 1696
rect 1547 1696 1573 1703
rect 2027 1696 2053 1703
rect 2187 1696 2233 1703
rect 2853 1707 2867 1713
rect 3067 1693 3073 1707
rect 3207 1693 3213 1707
rect 5587 1696 5633 1703
rect 3653 1687 3667 1693
rect 4033 1687 4047 1693
rect 87 1673 93 1687
rect 1127 1676 1213 1683
rect 1487 1676 1553 1683
rect 1680 1683 1693 1687
rect 1667 1676 1693 1683
rect 1680 1673 1693 1676
rect 1847 1676 1893 1683
rect 2227 1686 2240 1687
rect 2227 1673 2233 1686
rect 2847 1676 2893 1683
rect 3347 1676 3413 1683
rect 1327 1653 1333 1667
rect 1507 1656 1573 1663
rect 2627 1656 2693 1663
rect 3087 1656 3173 1663
rect 3547 1656 3733 1663
rect 4036 1656 4053 1663
rect 267 1636 353 1643
rect 1147 1636 1273 1643
rect 1287 1636 1333 1643
rect 1387 1636 1433 1643
rect 1487 1636 1713 1643
rect 1807 1636 2172 1643
rect 2208 1636 2813 1643
rect 2887 1633 2893 1647
rect 2967 1636 3113 1643
rect 3267 1636 3312 1643
rect 3348 1636 3493 1643
rect 3587 1636 3643 1643
rect 1507 1616 1713 1623
rect 1867 1616 2053 1623
rect 2187 1616 2653 1623
rect 2707 1616 2733 1623
rect 2867 1613 2873 1627
rect 2927 1616 3193 1623
rect 3527 1616 3573 1623
rect 3587 1616 3613 1623
rect 3636 1623 3643 1636
rect 3707 1636 3853 1643
rect 3867 1636 3893 1643
rect 4036 1643 4043 1656
rect 4067 1656 4093 1663
rect 4136 1663 4143 1693
rect 5513 1687 5527 1693
rect 5787 1676 5873 1683
rect 5967 1676 6053 1683
rect 4136 1656 4253 1663
rect 4387 1656 4413 1663
rect 5036 1656 5073 1663
rect 3947 1636 4043 1643
rect 4287 1636 4333 1643
rect 4416 1643 4423 1653
rect 4416 1636 4633 1643
rect 4767 1636 4953 1643
rect 5036 1643 5043 1656
rect 4967 1636 5043 1643
rect 5067 1636 5112 1643
rect 5148 1636 5173 1643
rect 6007 1636 6093 1643
rect 6107 1636 6133 1643
rect 6367 1636 6413 1643
rect 6467 1636 6493 1643
rect 3636 1616 3753 1623
rect 3767 1616 3873 1623
rect 3927 1626 3940 1627
rect 3927 1613 3933 1626
rect 3987 1616 4012 1623
rect 4048 1613 4053 1627
rect 4267 1616 4453 1623
rect 4527 1616 4633 1623
rect 1307 1596 1333 1603
rect 1547 1593 1553 1607
rect 1607 1596 1633 1603
rect 1707 1596 1933 1603
rect 2067 1593 2073 1607
rect 2147 1596 2313 1603
rect 2327 1596 2453 1603
rect 2467 1596 2493 1603
rect 2646 1593 2647 1600
rect 987 1576 1573 1583
rect 1727 1576 2193 1583
rect 2247 1576 2332 1583
rect 2368 1576 2553 1583
rect 2633 1583 2647 1593
rect 2668 1596 2873 1603
rect 3056 1596 3333 1603
rect 2633 1580 2713 1583
rect 2635 1576 2713 1580
rect 3056 1583 3063 1596
rect 3407 1593 3413 1607
rect 3567 1596 3612 1603
rect 3648 1596 3733 1603
rect 3787 1596 3953 1603
rect 4133 1603 4147 1613
rect 4727 1616 4993 1623
rect 5007 1616 5153 1623
rect 5207 1616 5393 1623
rect 5516 1616 5653 1623
rect 3967 1600 4147 1603
rect 3967 1596 4143 1600
rect 4167 1596 4593 1603
rect 4607 1596 4853 1603
rect 5516 1603 5523 1616
rect 4967 1596 5523 1603
rect 5547 1593 5553 1607
rect 6207 1596 6353 1603
rect 6367 1596 6473 1603
rect 2827 1576 3063 1583
rect 3087 1576 3133 1583
rect 3187 1576 3453 1583
rect 3527 1576 3733 1583
rect 3756 1576 5833 1583
rect 87 1556 273 1563
rect 1027 1563 1040 1567
rect 1027 1553 1043 1563
rect 1547 1556 1673 1563
rect 1696 1556 1793 1563
rect 1036 1543 1043 1553
rect 206 1533 207 1540
rect 1036 1536 1273 1543
rect 1607 1536 1633 1543
rect 1696 1543 1703 1556
rect 2067 1556 2203 1563
rect 1647 1536 1703 1543
rect 1727 1536 2173 1543
rect 2196 1543 2203 1556
rect 2287 1556 2413 1563
rect 3756 1563 3763 1576
rect 6227 1576 6293 1583
rect 2427 1556 3763 1563
rect 3787 1556 3993 1563
rect 4007 1556 4173 1563
rect 4287 1556 4353 1563
rect 4367 1556 4673 1563
rect 4687 1556 4813 1563
rect 5047 1556 5133 1563
rect 5156 1556 5193 1563
rect 2196 1536 2773 1543
rect 3047 1536 3353 1543
rect 3507 1536 3593 1543
rect 3607 1536 3653 1543
rect 3747 1536 3913 1543
rect 4327 1536 4413 1543
rect 4467 1536 4552 1543
rect 4588 1536 4612 1543
rect 5156 1543 5163 1556
rect 5247 1556 5313 1563
rect 4648 1536 5163 1543
rect 5227 1536 5413 1543
rect 5627 1536 5713 1543
rect 6247 1536 6273 1543
rect 6287 1536 6393 1543
rect 193 1527 207 1533
rect 4153 1527 4167 1533
rect 206 1520 207 1527
rect 228 1516 373 1523
rect 587 1516 953 1523
rect 1647 1516 1883 1523
rect 467 1496 612 1503
rect 648 1496 793 1503
rect 807 1496 913 1503
rect 927 1496 1033 1503
rect 1087 1496 1713 1503
rect 1787 1496 1853 1503
rect 1876 1503 1883 1516
rect 2227 1516 2393 1523
rect 2487 1516 2893 1523
rect 2947 1516 3093 1523
rect 3147 1516 3253 1523
rect 3567 1516 3652 1523
rect 3688 1516 3793 1523
rect 4207 1516 4253 1523
rect 4407 1516 4513 1523
rect 4527 1516 4733 1523
rect 5007 1516 5173 1523
rect 5187 1516 5353 1523
rect 5547 1516 5633 1523
rect 6307 1516 6493 1523
rect 1876 1496 2863 1503
rect 173 1487 187 1493
rect 2487 1476 2703 1483
rect 1493 1467 1507 1473
rect 167 1456 193 1463
rect 627 1456 713 1463
rect 1027 1456 1073 1463
rect 1927 1453 1933 1467
rect 2073 1447 2087 1453
rect 2696 1447 2703 1476
rect 2856 1467 2863 1496
rect 2887 1496 3293 1503
rect 3307 1496 3692 1503
rect 3728 1496 3773 1503
rect 3927 1496 3973 1503
rect 4087 1496 4293 1503
rect 4767 1496 4793 1503
rect 5167 1496 5193 1503
rect 5267 1496 5313 1503
rect 5627 1496 5693 1503
rect 6267 1496 6393 1503
rect 5736 1476 5833 1483
rect 2867 1456 2933 1463
rect 3247 1456 3293 1463
rect 3487 1456 3553 1463
rect 3620 1463 3633 1467
rect 3607 1456 3633 1463
rect 3620 1453 3633 1456
rect 4167 1463 4180 1467
rect 4167 1456 4193 1463
rect 4167 1453 4180 1456
rect 4287 1456 4353 1463
rect 5587 1456 5633 1463
rect 5736 1447 5743 1476
rect 5847 1476 5973 1483
rect 6327 1476 6513 1483
rect 6353 1447 6367 1453
rect 2507 1443 2520 1447
rect 2507 1436 2533 1443
rect 2507 1433 2520 1436
rect 2907 1436 2973 1443
rect 3787 1436 3833 1443
rect 4607 1436 4673 1443
rect 4987 1436 5013 1443
rect 5920 1443 5933 1447
rect 5907 1436 5933 1443
rect 5920 1433 5933 1436
rect 3367 1416 3393 1423
rect 3667 1413 3673 1427
rect 5327 1413 5333 1427
rect 5647 1413 5653 1427
rect 307 1396 352 1403
rect 388 1403 400 1407
rect 388 1396 413 1403
rect 388 1393 400 1396
rect 507 1396 593 1403
rect 827 1396 913 1403
rect 1240 1403 1253 1407
rect 1227 1396 1253 1403
rect 1240 1393 1253 1396
rect 1307 1396 1353 1403
rect 1367 1396 1433 1403
rect 1527 1396 1613 1403
rect 1747 1393 1753 1407
rect 1867 1403 1880 1407
rect 1867 1396 1893 1403
rect 1867 1393 1880 1396
rect 2147 1396 2233 1403
rect 2287 1396 2333 1403
rect 2427 1396 2513 1403
rect 3767 1396 3813 1403
rect 4267 1393 4273 1407
rect 4587 1396 4693 1403
rect 4800 1403 4813 1407
rect 4787 1396 4813 1403
rect 4800 1393 4813 1396
rect 4947 1396 4993 1403
rect 5087 1396 5153 1403
rect 5280 1403 5293 1407
rect 5267 1396 5293 1403
rect 5280 1393 5293 1396
rect 5427 1396 5493 1403
rect 5567 1396 5653 1403
rect 5987 1396 6033 1403
rect 6207 1396 6293 1403
rect 6427 1396 6493 1403
rect 133 1387 147 1393
rect 186 1353 187 1360
rect 267 1356 313 1363
rect 416 1363 423 1393
rect 593 1387 607 1393
rect 773 1387 787 1393
rect 3153 1387 3167 1393
rect 2607 1373 2613 1387
rect 2667 1373 2673 1387
rect 3313 1387 3327 1393
rect 3373 1387 3387 1393
rect 3627 1376 3693 1383
rect 416 1356 913 1363
rect 927 1356 1013 1363
rect 1247 1356 1333 1363
rect 1347 1356 1813 1363
rect 1827 1356 2013 1363
rect 2267 1356 2473 1363
rect 2567 1356 2613 1363
rect 2827 1356 2873 1363
rect 3247 1356 3373 1363
rect 3387 1356 3493 1363
rect 3647 1356 3713 1363
rect 3896 1363 3903 1393
rect 4053 1387 4067 1393
rect 4373 1387 4387 1393
rect 4127 1376 4153 1383
rect 4167 1373 4173 1387
rect 4733 1387 4747 1393
rect 5307 1373 5312 1387
rect 5348 1373 5353 1387
rect 3896 1356 4593 1363
rect 4727 1356 4773 1363
rect 4907 1356 4973 1363
rect 5167 1356 5373 1363
rect 5396 1356 5513 1363
rect 173 1347 187 1353
rect 186 1340 187 1347
rect 208 1333 213 1347
rect 367 1336 453 1343
rect 1287 1336 1373 1343
rect 1587 1336 1693 1343
rect 1907 1336 2093 1343
rect 2627 1336 2653 1343
rect 2707 1336 2733 1343
rect 2787 1336 2913 1343
rect 2967 1336 3153 1343
rect 3176 1336 3312 1343
rect 127 1316 413 1323
rect 1187 1316 1293 1323
rect 1447 1316 1533 1323
rect 2027 1316 2193 1323
rect 2207 1316 2293 1323
rect 2307 1316 2433 1323
rect 2447 1316 3053 1323
rect 3176 1323 3183 1336
rect 3348 1336 3372 1343
rect 3408 1333 3413 1347
rect 3427 1336 3633 1343
rect 3767 1336 3793 1343
rect 4067 1336 4413 1343
rect 4427 1336 4473 1343
rect 4487 1336 4513 1343
rect 4587 1336 4613 1343
rect 4707 1336 4873 1343
rect 4927 1336 5013 1343
rect 5027 1336 5233 1343
rect 5396 1343 5403 1356
rect 5667 1356 5873 1363
rect 5887 1356 6053 1363
rect 5247 1336 5403 1343
rect 5547 1336 5613 1343
rect 5667 1336 5793 1343
rect 6187 1336 6373 1343
rect 3076 1316 3183 1323
rect 147 1296 453 1303
rect 1296 1303 1303 1313
rect 1296 1296 1793 1303
rect 1807 1296 2053 1303
rect 2147 1296 2283 1303
rect 2276 1287 2283 1296
rect 2907 1296 2953 1303
rect 3007 1296 3053 1303
rect 3076 1303 3083 1316
rect 3227 1316 3273 1323
rect 3327 1316 4213 1323
rect 4227 1316 4433 1323
rect 4827 1316 4853 1323
rect 4867 1316 5093 1323
rect 5307 1316 5893 1323
rect 6007 1316 6133 1323
rect 6347 1316 6493 1323
rect 3067 1296 3083 1303
rect 4027 1296 4073 1303
rect 4187 1296 4333 1303
rect 4387 1296 4793 1303
rect 4807 1296 5033 1303
rect 5047 1296 5173 1303
rect 5747 1296 5933 1303
rect 5947 1296 6173 1303
rect 6247 1296 6413 1303
rect 407 1276 473 1283
rect 1147 1276 1313 1283
rect 1327 1276 1353 1283
rect 1407 1276 1493 1283
rect 1567 1276 1613 1283
rect 1956 1276 2233 1283
rect 213 1267 227 1273
rect 436 1256 533 1263
rect 436 1227 443 1256
rect 747 1256 773 1263
rect 1176 1256 1233 1263
rect 1176 1227 1183 1256
rect 1956 1263 1963 1276
rect 2287 1276 2393 1283
rect 2747 1276 2833 1283
rect 3227 1276 3673 1283
rect 3687 1276 3753 1283
rect 3907 1276 3933 1283
rect 4207 1276 4233 1283
rect 4287 1276 4373 1283
rect 4747 1276 4913 1283
rect 4967 1273 4972 1287
rect 5008 1276 5373 1283
rect 5387 1276 5472 1283
rect 5508 1276 5833 1283
rect 5847 1276 6153 1283
rect 6236 1276 6433 1283
rect 1607 1256 1963 1263
rect 2387 1256 2553 1263
rect 2727 1256 2773 1263
rect 2887 1256 3073 1263
rect 3127 1256 3293 1263
rect 3307 1256 3333 1263
rect 3407 1256 3553 1263
rect 3636 1256 3713 1263
rect 2087 1236 2153 1243
rect 3636 1227 3643 1256
rect 3827 1256 3993 1263
rect 4007 1256 4113 1263
rect 4207 1256 4253 1263
rect 4307 1256 4353 1263
rect 4856 1256 4953 1263
rect 4167 1236 4233 1243
rect 4856 1243 4863 1256
rect 5087 1256 5133 1263
rect 5327 1256 5353 1263
rect 5416 1256 5473 1263
rect 4767 1236 4863 1243
rect 5416 1227 5423 1256
rect 5576 1256 5753 1263
rect 5576 1227 5583 1256
rect 5767 1256 5993 1263
rect 6236 1263 6243 1276
rect 6056 1256 6243 1263
rect 6056 1227 6063 1256
rect 6267 1256 6363 1263
rect 6193 1227 6207 1233
rect 6356 1227 6363 1256
rect 127 1213 133 1227
rect 200 1223 213 1227
rect 187 1216 213 1223
rect 200 1213 213 1216
rect 307 1216 393 1223
rect 907 1216 953 1223
rect 1067 1216 1133 1223
rect 1307 1223 1320 1227
rect 1307 1216 1333 1223
rect 1307 1213 1320 1216
rect 1720 1223 1733 1227
rect 1707 1216 1733 1223
rect 1720 1213 1733 1216
rect 1880 1223 1893 1227
rect 1867 1216 1893 1223
rect 1880 1213 1893 1216
rect 2520 1223 2533 1227
rect 2507 1216 2533 1223
rect 2520 1213 2533 1216
rect 2647 1216 2712 1223
rect 2733 1213 2734 1220
rect 2800 1223 2812 1227
rect 2787 1216 2812 1223
rect 2800 1213 2812 1216
rect 2848 1216 2913 1223
rect 3087 1216 3133 1223
rect 3327 1213 3333 1227
rect 3527 1216 3593 1223
rect 3807 1216 3913 1223
rect 4307 1213 4312 1227
rect 4348 1216 4393 1223
rect 4527 1216 4593 1223
rect 4927 1216 4993 1223
rect 5087 1213 5093 1227
rect 5227 1216 5333 1223
rect 5467 1216 5533 1223
rect 5687 1213 5693 1227
rect 5827 1216 5873 1223
rect 2733 1207 2747 1213
rect 647 1176 713 1183
rect 1527 1176 1593 1183
rect 2200 1183 2213 1187
rect 2187 1176 2213 1183
rect 2200 1173 2213 1176
rect 2347 1176 2393 1183
rect 4327 1176 4373 1183
rect 4747 1176 4813 1183
rect 1993 1167 2007 1173
rect 4133 1167 4147 1173
rect 4453 1167 4467 1173
rect 547 1156 593 1163
rect 1367 1156 1473 1163
rect 3207 1156 3273 1163
rect 3507 1156 3573 1163
rect 4627 1156 4693 1163
rect 5067 1156 5153 1163
rect 5947 1156 5993 1163
rect 187 1136 213 1143
rect 227 1136 253 1143
rect 787 1136 813 1143
rect 3653 1143 3667 1153
rect 3653 1136 3753 1143
rect 4027 1136 4153 1143
rect 4367 1136 4493 1143
rect 507 1113 512 1127
rect 548 1116 873 1123
rect 887 1116 993 1123
rect 1147 1116 1353 1123
rect 1647 1116 1793 1123
rect 1847 1116 2532 1123
rect 2568 1116 2653 1123
rect 2727 1113 2733 1127
rect 2807 1116 2843 1123
rect 247 1096 313 1103
rect 967 1096 1193 1103
rect 1287 1096 1313 1103
rect 1327 1096 1493 1103
rect 1547 1096 1653 1103
rect 1667 1096 1813 1103
rect 2487 1096 2813 1103
rect 2836 1103 2843 1116
rect 2947 1116 3053 1123
rect 3096 1120 3473 1123
rect 3093 1116 3473 1120
rect 3093 1107 3107 1116
rect 3547 1116 3653 1123
rect 3707 1116 3853 1123
rect 3927 1116 4193 1123
rect 4207 1116 4312 1123
rect 4348 1116 4373 1123
rect 4907 1116 4973 1123
rect 4987 1116 5013 1123
rect 5207 1116 5313 1123
rect 5367 1116 5553 1123
rect 5867 1116 6033 1123
rect 2836 1096 2913 1103
rect 2927 1096 3013 1103
rect 3147 1096 3173 1103
rect 3347 1096 3413 1103
rect 3427 1096 3833 1103
rect 3947 1096 4073 1103
rect 4207 1096 4233 1103
rect 4287 1096 4373 1103
rect 4476 1096 4753 1103
rect 987 1076 1033 1083
rect 1187 1076 1333 1083
rect 1687 1076 1833 1083
rect 2007 1076 2253 1083
rect 2527 1076 2833 1083
rect 2847 1076 3432 1083
rect 3468 1076 3692 1083
rect 3728 1076 4053 1083
rect 4476 1083 4483 1096
rect 5487 1096 5513 1103
rect 5596 1096 5713 1103
rect 4107 1076 4483 1083
rect 5313 1087 5327 1093
rect 5407 1076 5452 1083
rect 5596 1083 5603 1096
rect 5907 1096 6213 1103
rect 6227 1096 6333 1103
rect 5488 1076 5603 1083
rect 5716 1083 5723 1093
rect 5716 1076 6253 1083
rect 6267 1076 6293 1083
rect 5633 1067 5647 1073
rect 1356 1056 1393 1063
rect 627 1036 793 1043
rect 807 1036 1033 1043
rect 1356 1043 1363 1056
rect 1507 1056 1633 1063
rect 1707 1056 2853 1063
rect 2867 1056 3843 1063
rect 1047 1036 1363 1043
rect 1387 1036 2873 1043
rect 3287 1036 3393 1043
rect 3836 1043 3843 1056
rect 3967 1056 4393 1063
rect 4416 1056 5133 1063
rect 3527 1036 3623 1043
rect 3836 1036 4333 1043
rect 2227 1016 2373 1023
rect 2467 1016 2493 1023
rect 2967 1016 3033 1023
rect 3167 1016 3293 1023
rect 3427 1013 3433 1027
rect 3567 1016 3593 1023
rect 3616 1023 3623 1036
rect 4416 1043 4423 1056
rect 5647 1056 5673 1063
rect 6007 1056 6153 1063
rect 4347 1036 4423 1043
rect 4467 1036 4553 1043
rect 4787 1036 5473 1043
rect 6107 1036 6253 1043
rect 3616 1016 3733 1023
rect 3747 1016 4013 1023
rect 4187 1016 4293 1023
rect 5027 1016 5093 1023
rect 1733 1007 1747 1013
rect 607 996 773 1003
rect 787 996 1073 1003
rect 1087 996 1433 1003
rect 1447 996 1533 1003
rect 2127 996 2333 1003
rect 2407 996 2593 1003
rect 2667 996 2713 1003
rect 2907 996 3093 1003
rect 3287 993 3293 1007
rect 3307 996 3383 1003
rect 167 976 633 983
rect 647 973 653 987
rect 747 976 873 983
rect 1127 976 1193 983
rect 1667 976 1813 983
rect 2027 976 2133 983
rect 2147 976 2493 983
rect 2647 976 2743 983
rect 2736 947 2743 976
rect 2827 976 3013 983
rect 3087 976 3193 983
rect 3207 976 3253 983
rect 3307 973 3313 987
rect 3376 983 3383 996
rect 3407 996 3693 1003
rect 3907 996 3933 1003
rect 4147 996 4212 1003
rect 4248 996 4473 1003
rect 4687 996 4733 1003
rect 4787 996 4833 1003
rect 4947 996 5073 1003
rect 6027 996 6053 1003
rect 6067 996 6293 1003
rect 3376 976 3453 983
rect 4067 976 4133 983
rect 4147 976 4253 983
rect 4367 976 4393 983
rect 4407 976 4633 983
rect 4727 976 4893 983
rect 4907 976 5093 983
rect 5547 976 5593 983
rect 5607 973 5613 987
rect 5827 976 5893 983
rect 6227 976 6473 983
rect 3867 956 4093 963
rect 327 936 373 943
rect 1287 936 1373 943
rect 2467 936 2533 943
rect 3107 936 3153 943
rect 3720 943 3733 947
rect 3707 936 3733 943
rect 3720 933 3733 936
rect 4347 936 4393 943
rect 5147 936 5253 943
rect 5587 936 5633 943
rect 5787 936 5813 943
rect 1887 916 1953 923
rect 4687 913 4693 927
rect 4387 896 4413 903
rect 207 876 253 883
rect 387 876 433 883
rect 447 876 512 883
rect 548 873 553 887
rect 727 873 733 887
rect 847 876 893 883
rect 1027 883 1040 887
rect 1027 876 1053 883
rect 1027 873 1040 876
rect 1527 876 1593 883
rect 1847 876 1933 883
rect 2047 876 2113 883
rect 2327 876 2393 883
rect 2507 876 2573 883
rect 2987 873 2993 887
rect 3227 873 3232 887
rect 3268 876 3333 883
rect 3427 876 3453 883
rect 3547 876 3633 883
rect 4327 873 4333 887
rect 4407 876 4453 883
rect 4627 876 4713 883
rect 4807 876 4853 883
rect 4967 873 4973 887
rect 5127 876 5173 883
rect 5647 876 5713 883
rect 5767 873 5773 887
rect 5927 876 5973 883
rect 6067 876 6153 883
rect 6247 873 6253 887
rect 6407 876 6453 883
rect 1213 867 1227 873
rect 327 863 340 867
rect 327 854 343 863
rect 320 853 343 854
rect 1633 867 1647 873
rect 2113 867 2127 873
rect 287 836 313 843
rect 336 843 343 853
rect 1733 847 1747 853
rect 336 836 453 843
rect 527 836 572 843
rect 608 836 653 843
rect 827 836 893 843
rect 1187 836 1273 843
rect 1987 836 2093 843
rect 2276 843 2283 873
rect 2433 867 2447 873
rect 2107 836 2283 843
rect 2296 836 2363 843
rect 127 816 353 823
rect 367 816 533 823
rect 576 823 583 833
rect 576 816 753 823
rect 987 816 1213 823
rect 1407 816 1453 823
rect 2296 823 2303 836
rect 1467 816 2303 823
rect 2327 813 2333 827
rect 2356 823 2363 836
rect 2407 836 2753 843
rect 2876 843 2883 873
rect 3493 867 3507 873
rect 2767 836 2883 843
rect 3027 836 3173 843
rect 3227 836 3363 843
rect 2356 816 2433 823
rect 2547 816 2633 823
rect 3047 816 3093 823
rect 3287 816 3333 823
rect 3356 823 3363 836
rect 3387 836 3533 843
rect 3587 836 3673 843
rect 3687 836 3793 843
rect 3836 843 3843 873
rect 4113 867 4127 873
rect 4667 856 4733 863
rect 3836 836 4153 843
rect 4167 836 4273 843
rect 4367 833 4373 847
rect 4867 836 4913 843
rect 4927 836 5053 843
rect 5276 843 5283 873
rect 5413 867 5427 873
rect 5276 836 5573 843
rect 5596 843 5603 873
rect 5827 853 5833 867
rect 5596 836 6053 843
rect 6067 836 6353 843
rect 4673 827 4687 833
rect 3356 816 3412 823
rect 3448 813 3453 827
rect 4227 816 4553 823
rect 4686 820 4687 827
rect 4708 813 4713 827
rect 5367 816 5873 823
rect 5987 816 6033 823
rect 207 796 473 803
rect 487 796 673 803
rect 767 796 853 803
rect 1847 796 2233 803
rect 2247 796 2793 803
rect 2847 796 2993 803
rect 3007 796 3052 803
rect 3088 796 3553 803
rect 4367 796 4773 803
rect 5267 796 5373 803
rect 5427 796 5533 803
rect 5547 796 5693 803
rect 5766 793 5767 800
rect 5788 796 6013 803
rect 6027 796 6113 803
rect 307 776 413 783
rect 427 776 833 783
rect 1827 776 1973 783
rect 1987 776 2032 783
rect 2068 776 2553 783
rect 2607 776 2693 783
rect 2867 776 3273 783
rect 3287 776 3493 783
rect 3787 776 3933 783
rect 4127 776 4273 783
rect 4287 776 4673 783
rect 4687 776 4793 783
rect 4927 776 5073 783
rect 5187 776 5293 783
rect 5447 776 5513 783
rect 5567 776 5593 783
rect 5753 783 5767 793
rect 5753 780 5813 783
rect 5755 776 5813 780
rect 127 756 553 763
rect 567 756 713 763
rect 967 756 1173 763
rect 1607 756 2193 763
rect 2207 756 2653 763
rect 2727 756 2773 763
rect 2927 756 3213 763
rect 3307 756 4213 763
rect 4427 756 4513 763
rect 4527 756 4653 763
rect 4827 756 4873 763
rect 4927 760 4963 763
rect 4927 756 4967 760
rect 4953 747 4967 756
rect 4987 756 5393 763
rect 5407 756 5453 763
rect 5467 756 5613 763
rect 5787 756 5873 763
rect 167 736 373 743
rect 827 736 873 743
rect 887 736 1033 743
rect 1047 736 1233 743
rect 1287 736 1413 743
rect 1707 736 1873 743
rect 1947 736 1993 743
rect 2407 736 2493 743
rect 2647 736 2673 743
rect 2767 736 3073 743
rect 3247 736 3273 743
rect 3447 736 3713 743
rect 3727 736 3773 743
rect 3816 736 3903 743
rect 233 707 247 713
rect 1276 707 1283 733
rect 2567 716 2623 723
rect 407 696 473 703
rect 587 696 653 703
rect 940 703 953 707
rect 927 696 953 703
rect 940 693 953 696
rect 1107 693 1113 707
rect 1347 696 1393 703
rect 1507 696 1553 703
rect 1847 703 1860 707
rect 1847 696 1873 703
rect 1847 693 1860 696
rect 1927 696 1973 703
rect 2120 703 2133 707
rect 2107 696 2133 703
rect 2120 693 2133 696
rect 2327 703 2340 707
rect 2327 696 2353 703
rect 2327 693 2340 696
rect 2527 696 2593 703
rect 2616 703 2623 716
rect 3067 716 3113 723
rect 3780 723 3793 727
rect 3776 713 3793 723
rect 2616 696 2673 703
rect 2807 693 2813 707
rect 2947 693 2953 707
rect 3247 696 3273 703
rect 3547 696 3612 703
rect 3648 693 3653 707
rect 3776 703 3783 713
rect 3816 707 3823 736
rect 3896 723 3903 736
rect 3927 736 3973 743
rect 4087 736 4163 743
rect 3896 716 3953 723
rect 4156 707 4163 736
rect 4347 736 4593 743
rect 4607 736 4633 743
rect 4656 736 4913 743
rect 4656 707 4663 736
rect 4967 736 5053 743
rect 5667 736 5733 743
rect 5787 736 5813 743
rect 6027 736 6053 743
rect 6156 736 6413 743
rect 6156 707 6163 736
rect 3707 696 3783 703
rect 3867 693 3873 707
rect 4027 693 4033 707
rect 4207 696 4313 703
rect 4407 696 4473 703
rect 4527 696 4573 703
rect 4847 696 4913 703
rect 5007 696 5053 703
rect 5167 696 5213 703
rect 5340 703 5353 707
rect 5327 696 5353 703
rect 5340 693 5353 696
rect 5507 696 5553 703
rect 5667 696 5773 703
rect 5867 693 5873 707
rect 5947 703 5960 707
rect 5947 696 5973 703
rect 5947 693 5960 696
rect 6207 696 6293 703
rect 2607 676 2633 683
rect 3267 676 3313 683
rect 2127 656 2213 663
rect 2927 656 2973 663
rect 3306 653 3307 660
rect 3328 663 3340 667
rect 3328 656 3353 663
rect 3328 653 3340 656
rect 733 647 747 653
rect 3173 647 3187 653
rect 2747 636 2833 643
rect 3293 647 3307 653
rect 3407 636 3473 643
rect 5427 633 5433 647
rect 5527 636 5633 643
rect 96 603 103 633
rect 253 623 267 633
rect 253 616 353 623
rect 667 616 813 623
rect 1807 616 1833 623
rect 2947 616 3033 623
rect 3047 616 3133 623
rect 3287 616 3433 623
rect 96 596 253 603
rect 487 596 853 603
rect 867 596 983 603
rect 647 576 953 583
rect 976 583 983 596
rect 1007 596 1413 603
rect 1587 596 1893 603
rect 1907 596 2113 603
rect 2247 596 2533 603
rect 2707 596 2973 603
rect 2987 596 3233 603
rect 3247 596 3753 603
rect 3767 596 4133 603
rect 4547 596 4673 603
rect 4687 596 4833 603
rect 4987 596 5013 603
rect 5027 596 5133 603
rect 5227 596 5273 603
rect 5287 596 5413 603
rect 5607 596 5633 603
rect 6047 596 6173 603
rect 6187 596 6353 603
rect 976 576 1053 583
rect 1067 576 1213 583
rect 1627 576 1693 583
rect 2427 576 2613 583
rect 2627 576 2733 583
rect 2947 576 3093 583
rect 3227 576 3793 583
rect 3807 576 3993 583
rect 4007 576 4393 583
rect 4587 576 4813 583
rect 5327 576 5373 583
rect 5387 576 5473 583
rect 5607 576 5673 583
rect 5887 576 6313 583
rect 6327 576 6393 583
rect 907 556 933 563
rect 947 556 1493 563
rect 1516 556 1973 563
rect 487 536 1333 543
rect 1516 543 1523 556
rect 2067 556 2133 563
rect 2707 556 2753 563
rect 2847 556 3313 563
rect 3627 553 3633 567
rect 3687 556 3833 563
rect 3847 556 4173 563
rect 4227 556 4673 563
rect 5067 556 5233 563
rect 5427 556 5493 563
rect 5507 556 5573 563
rect 5987 556 6133 563
rect 1447 536 1523 543
rect 1587 536 1733 543
rect 2007 536 2073 543
rect 2087 536 2553 543
rect 3887 536 4193 543
rect 4727 536 4933 543
rect 5236 543 5243 553
rect 5236 536 5593 543
rect 5667 536 6033 543
rect 127 516 233 523
rect 247 516 293 523
rect 307 516 1013 523
rect 1107 516 1253 523
rect 1267 516 1753 523
rect 2107 516 2493 523
rect 3067 516 3433 523
rect 3447 516 3543 523
rect 747 496 813 503
rect 1407 496 1773 503
rect 1787 496 2053 503
rect 2387 496 2513 503
rect 2567 496 3292 503
rect 3328 496 3513 503
rect 3536 503 3543 516
rect 3567 516 5933 523
rect 3536 496 3832 503
rect 3868 496 3913 503
rect 3967 496 4012 503
rect 4048 496 4073 503
rect 4147 496 5793 503
rect 787 476 1093 483
rect 1247 476 1353 483
rect 1367 476 2933 483
rect 3027 476 3093 483
rect 3187 476 3273 483
rect 3287 476 3713 483
rect 3727 476 4093 483
rect 4206 473 4207 480
rect 4228 476 4393 483
rect 4407 476 4753 483
rect 5627 476 5733 483
rect 5747 476 6193 483
rect 6207 476 6393 483
rect 167 456 273 463
rect 607 456 952 463
rect 988 456 1173 463
rect 1187 456 1433 463
rect 1527 456 1693 463
rect 1887 456 3313 463
rect 3467 456 3523 463
rect 687 436 713 443
rect 847 436 873 443
rect 1787 436 1813 443
rect 2367 436 2523 443
rect 1120 423 1133 427
rect 1107 416 1133 423
rect 1120 413 1133 416
rect 2373 407 2387 413
rect 2516 407 2523 436
rect 3516 423 3523 456
rect 3547 456 4133 463
rect 4193 463 4207 473
rect 4193 460 4253 463
rect 4196 456 4253 460
rect 4427 456 4613 463
rect 4807 456 5113 463
rect 5407 456 5433 463
rect 5507 456 5573 463
rect 5587 456 5753 463
rect 6007 456 6313 463
rect 4207 436 4303 443
rect 3516 416 3593 423
rect 4296 407 4303 436
rect 5947 436 5973 443
rect 5767 416 5833 423
rect 6347 413 6353 427
rect 5113 407 5127 413
rect 307 396 353 403
rect 1267 396 1313 403
rect 3107 396 3173 403
rect 4660 403 4673 407
rect 4647 396 4673 403
rect 4660 393 4673 396
rect 4847 396 4913 403
rect 6067 396 6113 403
rect 807 376 833 383
rect 3827 376 3873 383
rect 4007 376 4053 383
rect 467 356 533 363
rect 927 356 993 363
rect 1087 356 1153 363
rect 1247 356 1293 363
rect 1347 363 1360 367
rect 1347 356 1373 363
rect 1347 353 1360 356
rect 1467 356 1513 363
rect 1607 356 1633 363
rect 1727 356 1773 363
rect 2067 356 2143 363
rect 136 323 143 353
rect 573 347 587 353
rect 753 347 767 353
rect 987 333 993 347
rect 1587 336 1613 343
rect 136 316 413 323
rect 727 316 813 323
rect 827 316 853 323
rect 1716 323 1723 353
rect 1427 316 1723 323
rect 1787 316 1813 323
rect 1856 323 1863 353
rect 2136 347 2143 356
rect 2227 353 2233 367
rect 2747 356 2833 363
rect 2947 356 2993 363
rect 2136 336 2153 347
rect 2140 333 2153 336
rect 1856 316 2013 323
rect 2187 316 2313 323
rect 2676 323 2683 353
rect 3527 356 3613 363
rect 3887 363 3900 367
rect 3887 356 3913 363
rect 3887 353 3900 356
rect 5147 356 5233 363
rect 5327 356 5413 363
rect 5507 356 5553 363
rect 5607 356 5693 363
rect 5807 356 5893 363
rect 6127 356 6173 363
rect 3413 347 3427 353
rect 2607 316 2683 323
rect 2907 316 2993 323
rect 3047 316 3493 323
rect 3776 323 3783 353
rect 4133 347 4147 353
rect 4433 347 4447 353
rect 3867 333 3873 347
rect 3987 336 4033 343
rect 4047 333 4053 347
rect 3507 316 4233 323
rect 4347 316 4613 323
rect 4776 323 4783 353
rect 4947 336 5053 343
rect 4627 316 4783 323
rect 5407 316 5493 323
rect 5947 316 5993 323
rect 627 296 753 303
rect 807 296 1033 303
rect 1047 296 1193 303
rect 1207 296 1453 303
rect 1807 296 2093 303
rect 2147 296 2353 303
rect 2407 296 2873 303
rect 3147 296 3733 303
rect 4227 296 4273 303
rect 4296 296 4673 303
rect 107 276 373 283
rect 387 276 573 283
rect 727 276 893 283
rect 907 276 1873 283
rect 2007 276 2183 283
rect 147 256 433 263
rect 713 253 714 260
rect 847 256 1093 263
rect 1587 256 2013 263
rect 2176 263 2183 276
rect 2276 276 2513 283
rect 2276 263 2283 276
rect 2667 276 2793 283
rect 2847 276 3533 283
rect 3607 276 3813 283
rect 3833 283 3847 293
rect 4296 283 4303 296
rect 4847 296 4893 303
rect 4907 296 5093 303
rect 5527 296 5613 303
rect 5727 296 5973 303
rect 3833 280 4303 283
rect 3836 276 4303 280
rect 4387 276 4453 283
rect 4467 276 4573 283
rect 5167 276 5193 283
rect 5447 276 6073 283
rect 2176 256 2283 263
rect 2356 256 2393 263
rect 713 247 727 253
rect 567 236 692 243
rect 713 240 714 247
rect 887 236 1053 243
rect 1347 233 1353 247
rect 1547 236 2133 243
rect 2356 243 2363 256
rect 2867 256 2953 263
rect 2967 256 3053 263
rect 3107 256 3273 263
rect 3387 256 3693 263
rect 3747 256 3893 263
rect 3916 256 4153 263
rect 2307 236 2363 243
rect 2387 236 2413 243
rect 2427 236 2473 243
rect 2487 236 3173 243
rect 3187 236 3333 243
rect 3427 236 3473 243
rect 3487 236 3633 243
rect 3647 236 3813 243
rect 3916 243 3923 256
rect 4167 256 5313 263
rect 5487 256 5633 263
rect 3887 236 3923 243
rect 4007 236 4433 243
rect 4607 236 4833 243
rect 5027 236 5533 243
rect 5767 236 5953 243
rect 5967 236 6112 243
rect 6148 236 6193 243
rect 307 216 353 223
rect 447 216 473 223
rect 667 216 692 223
rect 728 216 832 223
rect 868 216 973 223
rect 1127 216 1153 223
rect 1307 216 1593 223
rect 1607 216 2033 223
rect 2167 216 2233 223
rect 2307 216 2693 223
rect 2767 216 3193 223
rect 3447 216 3533 223
rect 3996 223 4003 233
rect 3687 216 4003 223
rect 4107 216 4193 223
rect 4387 216 4653 223
rect 4667 216 4883 223
rect 373 187 387 193
rect 1033 187 1047 193
rect 1273 196 1373 203
rect 1273 187 1287 196
rect 1793 187 1807 193
rect 2193 187 2207 193
rect 2793 187 2807 193
rect 3707 193 3713 207
rect 2993 187 3007 193
rect 4876 187 4883 216
rect 4947 216 5133 223
rect 5227 216 5323 223
rect 5316 187 5323 216
rect 5367 216 5693 223
rect 5496 187 5503 216
rect 5987 216 6143 223
rect 6136 187 6143 216
rect 127 176 212 183
rect 248 173 253 187
rect 487 176 553 183
rect 576 176 613 183
rect 347 156 393 163
rect 576 163 583 176
rect 707 176 753 183
rect 847 176 933 183
rect 1207 183 1220 187
rect 1207 176 1233 183
rect 1207 173 1220 176
rect 1447 176 1533 183
rect 1627 176 1713 183
rect 1847 176 1873 183
rect 1980 183 1993 187
rect 1967 176 1993 183
rect 1980 173 1993 176
rect 2247 176 2313 183
rect 2407 173 2413 187
rect 2567 176 2633 183
rect 3167 176 3213 183
rect 3347 176 3433 183
rect 3547 176 3593 183
rect 3707 176 3773 183
rect 3907 176 3953 183
rect 4047 183 4060 187
rect 4047 176 4073 183
rect 4047 173 4060 176
rect 4127 176 4173 183
rect 4440 183 4453 187
rect 4427 176 4453 183
rect 4440 173 4453 176
rect 4707 173 4713 187
rect 4967 176 5033 183
rect 5207 176 5273 183
rect 5547 176 5653 183
rect 6020 183 6033 187
rect 6007 176 6033 183
rect 6020 173 6033 176
rect 6227 176 6273 183
rect 516 156 583 163
rect 516 147 523 156
rect 1027 156 1073 163
rect 1327 156 1353 163
rect 2887 156 2913 163
rect 3047 156 3073 163
rect 3687 156 3713 163
rect 3867 156 3893 163
rect 507 136 523 147
rect 507 133 520 136
rect 687 133 693 147
rect 1147 136 1193 143
rect 3027 136 3093 143
rect 3307 133 3313 147
rect 3727 133 3733 147
rect 4447 136 4533 143
rect 373 127 387 133
rect 527 116 593 123
rect 687 116 733 123
rect 1047 116 1093 123
rect 1107 116 1213 123
rect 2087 116 2173 123
rect 2687 116 2773 123
rect 3547 116 3613 123
rect 4267 116 4313 123
rect 5767 116 5813 123
rect 5827 116 5893 123
rect 6347 116 6433 123
rect 3873 107 3887 113
rect 3227 96 3373 103
rect 4093 103 4107 113
rect 6193 107 6207 113
rect 4007 96 4107 103
rect 4767 96 4813 103
rect 6047 96 6093 103
rect 227 76 273 83
rect 647 76 673 83
rect 727 76 773 83
rect 827 76 853 83
rect 907 76 953 83
rect 1007 76 1033 83
rect 1056 76 1203 83
rect 1056 63 1063 76
rect 1196 67 1203 76
rect 1267 76 1333 83
rect 1347 76 1413 83
rect 1467 76 1553 83
rect 1736 76 1893 83
rect 1736 67 1743 76
rect 2307 76 2413 83
rect 2436 76 3213 83
rect 367 56 1063 63
rect 1207 56 1733 63
rect 1787 56 1933 63
rect 2436 63 2443 76
rect 3507 76 3653 83
rect 3727 76 3833 83
rect 3907 76 3973 83
rect 4607 76 4893 83
rect 5067 76 5333 83
rect 5347 76 5673 83
rect 5687 76 6213 83
rect 1947 56 2443 63
rect 2867 56 2973 63
rect 2987 56 3693 63
rect 3807 56 3933 63
rect 3947 56 4933 63
rect 5187 56 6033 63
rect 707 36 1033 43
rect 1167 36 1293 43
rect 1307 36 2053 43
rect 2167 36 2513 43
rect 2527 36 3032 43
rect 3068 36 4173 43
rect 247 16 853 23
rect 2107 16 2373 23
rect 2547 16 2693 23
rect 2707 16 3112 23
rect 3148 16 3533 23
rect 3587 16 3673 23
rect 3747 16 4953 23
rect 5147 16 5173 23
<< m3contact >>
rect 1053 6513 1067 6527
rect 2293 6513 2307 6527
rect 1493 6493 1507 6507
rect 1693 6493 1707 6507
rect 1853 6493 1867 6507
rect 3933 6513 3947 6527
rect 3973 6513 3987 6527
rect 4013 6513 4027 6527
rect 6233 6513 6247 6527
rect 6273 6513 6287 6527
rect 2753 6493 2767 6507
rect 2933 6493 2947 6507
rect 3253 6493 3267 6507
rect 3413 6493 3427 6507
rect 5253 6493 5267 6507
rect 5693 6493 5707 6507
rect 553 6473 567 6487
rect 693 6473 707 6487
rect 933 6473 947 6487
rect 1093 6473 1107 6487
rect 593 6453 607 6467
rect 733 6453 747 6467
rect 973 6453 987 6467
rect 2093 6473 2107 6487
rect 2253 6473 2267 6487
rect 2293 6473 2307 6487
rect 2813 6473 2827 6487
rect 2853 6473 2867 6487
rect 3173 6473 3187 6487
rect 3573 6473 3587 6487
rect 4633 6473 4647 6487
rect 4753 6473 4767 6487
rect 5853 6473 5867 6487
rect 5933 6473 5947 6487
rect 1313 6453 1327 6467
rect 1533 6453 1547 6467
rect 2213 6453 2227 6467
rect 2393 6453 2407 6467
rect 1493 6433 1507 6447
rect 1853 6433 1867 6447
rect 2133 6433 2147 6447
rect 2293 6433 2307 6447
rect 3533 6453 3547 6467
rect 3653 6453 3667 6467
rect 3753 6453 3767 6467
rect 4713 6453 4727 6467
rect 6013 6453 6027 6467
rect 6073 6453 6087 6467
rect 6373 6453 6387 6467
rect 6473 6453 6487 6467
rect 2853 6433 2867 6447
rect 2893 6433 2907 6447
rect 3173 6433 3187 6447
rect 3213 6433 3227 6447
rect 3313 6433 3327 6447
rect 3373 6433 3387 6447
rect 4993 6433 5007 6447
rect 133 6413 147 6427
rect 213 6413 227 6427
rect 393 6413 407 6427
rect 673 6413 687 6427
rect 733 6413 747 6427
rect 814 6413 828 6427
rect 933 6413 947 6427
rect 1053 6413 1067 6427
rect 1273 6413 1287 6427
rect 1373 6413 1387 6427
rect 1533 6413 1547 6427
rect 1693 6413 1707 6427
rect 1733 6413 1747 6427
rect 1893 6413 1907 6427
rect 2093 6413 2107 6427
rect 2513 6413 2527 6427
rect 2673 6413 2687 6427
rect 2753 6413 2767 6427
rect 3053 6413 3067 6427
rect 3413 6413 3427 6427
rect 3533 6413 3547 6427
rect 3573 6413 3587 6427
rect 3713 6413 3727 6427
rect 3813 6413 3827 6427
rect 3993 6413 4007 6427
rect 4093 6413 4107 6427
rect 4433 6413 4447 6427
rect 4713 6413 4727 6427
rect 4753 6413 4767 6427
rect 4793 6413 4807 6427
rect 5933 6433 5947 6447
rect 6213 6433 6227 6447
rect 6253 6433 6267 6447
rect 5553 6413 5567 6427
rect 5693 6413 5707 6427
rect 5833 6413 5847 6427
rect 6053 6413 6067 6427
rect 6153 6413 6167 6427
rect 6373 6413 6387 6427
rect 6453 6413 6467 6427
rect 4993 6393 5007 6407
rect 5053 6393 5067 6407
rect 5113 6393 5127 6407
rect 5253 6393 5267 6407
rect 5393 6393 5407 6407
rect 2353 6373 2367 6387
rect 2773 6373 2787 6387
rect 3153 6373 3167 6387
rect 3233 6373 3247 6387
rect 4013 6373 4027 6387
rect 4253 6373 4267 6387
rect 4313 6373 4327 6387
rect 4413 6373 4427 6387
rect 4553 6373 4567 6387
rect 4613 6373 4627 6387
rect 6013 6373 6027 6387
rect 6193 6373 6207 6387
rect 193 6353 207 6367
rect 233 6353 247 6367
rect 273 6353 287 6367
rect 373 6353 387 6367
rect 413 6353 427 6367
rect 573 6353 587 6367
rect 613 6353 627 6367
rect 713 6353 727 6367
rect 753 6353 767 6367
rect 913 6353 927 6367
rect 953 6353 967 6367
rect 993 6353 1007 6367
rect 1153 6353 1167 6367
rect 1193 6353 1207 6367
rect 1313 6353 1327 6367
rect 1353 6353 1367 6367
rect 1473 6353 1487 6367
rect 1513 6353 1527 6367
rect 1673 6353 1687 6367
rect 1713 6353 1727 6367
rect 1833 6353 1847 6367
rect 1873 6353 1887 6367
rect 1953 6353 1967 6367
rect 1993 6353 2007 6367
rect 2113 6353 2127 6367
rect 2393 6353 2407 6367
rect 2433 6353 2447 6367
rect 2533 6353 2547 6367
rect 2573 6353 2587 6367
rect 2693 6353 2707 6367
rect 2733 6353 2747 6367
rect 2933 6353 2947 6367
rect 3193 6353 3207 6367
rect 2513 6333 2527 6347
rect 2833 6333 2847 6347
rect 2893 6333 2907 6347
rect 3073 6333 3087 6347
rect 3213 6333 3227 6347
rect 3513 6353 3527 6367
rect 3553 6353 3567 6367
rect 3653 6353 3667 6367
rect 3693 6353 3707 6367
rect 3753 6353 3767 6367
rect 4113 6353 4127 6367
rect 4733 6353 4747 6367
rect 4773 6353 4787 6367
rect 4893 6353 4907 6367
rect 4933 6353 4947 6367
rect 5553 6353 5567 6367
rect 5673 6353 5687 6367
rect 5713 6353 5727 6367
rect 5833 6353 5847 6367
rect 6033 6353 6047 6367
rect 6073 6353 6087 6367
rect 6173 6353 6187 6367
rect 6353 6353 6367 6367
rect 6393 6353 6407 6367
rect 3373 6333 3387 6347
rect 3413 6333 3427 6347
rect 6053 6333 6067 6347
rect 6113 6333 6127 6347
rect 133 6313 147 6327
rect 373 6313 387 6327
rect 513 6313 527 6327
rect 1273 6313 1287 6327
rect 1473 6313 1487 6327
rect 1673 6313 1687 6327
rect 1833 6313 1847 6327
rect 2493 6313 2507 6327
rect 2533 6313 2547 6327
rect 2712 6313 2726 6327
rect 2734 6313 2748 6327
rect 2773 6313 2787 6327
rect 3693 6313 3707 6327
rect 3993 6313 4007 6327
rect 4893 6313 4907 6327
rect 4953 6313 4967 6327
rect 5393 6313 5407 6327
rect 5553 6313 5567 6327
rect 5673 6313 5687 6327
rect 6153 6313 6167 6327
rect 913 6293 927 6307
rect 993 6293 1007 6307
rect 1093 6293 1107 6307
rect 1213 6293 1227 6307
rect 1373 6293 1387 6307
rect 1753 6293 1767 6307
rect 2813 6293 2827 6307
rect 3073 6293 3087 6307
rect 4013 6293 4027 6307
rect 4353 6293 4367 6307
rect 4733 6293 4747 6307
rect 4933 6293 4947 6307
rect 5093 6293 5107 6307
rect 5813 6293 5827 6307
rect 5933 6293 5947 6307
rect 733 6273 747 6287
rect 1193 6273 1207 6287
rect 2493 6273 2507 6287
rect 673 6253 687 6267
rect 1033 6253 1047 6267
rect 1333 6253 1347 6267
rect 1593 6253 1607 6267
rect 1873 6253 1887 6267
rect 1953 6253 1967 6267
rect 3193 6273 3207 6287
rect 4113 6273 4127 6287
rect 4473 6273 4487 6287
rect 4993 6273 5007 6287
rect 5213 6273 5227 6287
rect 5473 6273 5487 6287
rect 2813 6253 2827 6267
rect 3813 6253 3827 6267
rect 4233 6253 4247 6267
rect 4693 6253 4707 6267
rect 4873 6253 4887 6267
rect 5053 6253 5067 6267
rect 5653 6253 5667 6267
rect 5833 6253 5847 6267
rect 6253 6253 6267 6267
rect 6333 6253 6347 6267
rect 413 6233 427 6247
rect 473 6233 487 6247
rect 1153 6233 1167 6247
rect 1473 6233 1487 6247
rect 1553 6233 1567 6247
rect 1733 6233 1747 6247
rect 233 6213 247 6227
rect 1253 6213 1267 6227
rect 1353 6213 1367 6227
rect 1513 6213 1527 6227
rect 2693 6233 2707 6247
rect 2753 6233 2767 6247
rect 2873 6233 2887 6247
rect 3173 6233 3187 6247
rect 4433 6233 4447 6247
rect 4953 6233 4967 6247
rect 4993 6233 5007 6247
rect 5113 6233 5127 6247
rect 5173 6234 5187 6248
rect 5913 6233 5927 6247
rect 6313 6233 6327 6247
rect 1773 6213 1787 6227
rect 2512 6213 2526 6227
rect 2573 6213 2587 6227
rect 2833 6213 2847 6227
rect 3153 6213 3167 6227
rect 3633 6213 3647 6227
rect 3773 6213 3787 6227
rect 4093 6213 4107 6227
rect 4413 6213 4427 6227
rect 4593 6213 4607 6227
rect 4873 6213 4887 6227
rect 5033 6213 5047 6227
rect 5148 6213 5162 6227
rect 5193 6213 5207 6227
rect 5233 6213 5247 6227
rect 5293 6213 5307 6227
rect 5393 6213 5407 6227
rect 273 6193 287 6207
rect 613 6193 627 6207
rect 1213 6193 1227 6207
rect 1553 6193 1567 6207
rect 1953 6193 1967 6207
rect 2013 6193 2027 6207
rect 2353 6193 2367 6207
rect 2993 6193 3007 6207
rect 3373 6193 3387 6207
rect 3413 6193 3427 6207
rect 3473 6193 3487 6207
rect 3853 6193 3867 6207
rect 3913 6193 3927 6207
rect 4073 6187 4087 6201
rect 5333 6193 5347 6207
rect 5873 6193 5887 6207
rect 6193 6193 6207 6207
rect 353 6173 367 6187
rect 393 6173 407 6187
rect 1253 6173 1267 6187
rect 1293 6173 1307 6187
rect 1393 6173 1407 6187
rect 1513 6173 1527 6187
rect 1713 6173 1727 6187
rect 1833 6173 1847 6187
rect 1993 6173 2007 6187
rect 2553 6173 2567 6187
rect 273 6153 287 6167
rect 673 6153 687 6167
rect 2613 6173 2627 6187
rect 2733 6173 2747 6187
rect 3053 6173 3067 6187
rect 3313 6173 3327 6187
rect 3453 6173 3467 6187
rect 3573 6173 3587 6187
rect 3692 6173 3706 6187
rect 3714 6173 3728 6187
rect 3873 6173 3887 6187
rect 4033 6173 4047 6187
rect 4573 6173 4587 6187
rect 153 6133 167 6147
rect 4093 6153 4107 6167
rect 4233 6153 4247 6167
rect 6093 6173 6107 6187
rect 473 6133 487 6147
rect 513 6133 527 6147
rect 593 6133 607 6147
rect 633 6133 647 6147
rect 913 6133 927 6147
rect 953 6133 967 6147
rect 1053 6133 1067 6147
rect 1093 6133 1107 6147
rect 1213 6133 1227 6147
rect 1253 6133 1267 6147
rect 1513 6133 1527 6147
rect 1553 6133 1567 6147
rect 1833 6133 1847 6147
rect 1873 6133 1887 6147
rect 1993 6133 2007 6147
rect 2033 6133 2047 6147
rect 2073 6133 2087 6147
rect 2373 6133 2387 6147
rect 2613 6133 2627 6147
rect 2653 6133 2667 6147
rect 2773 6133 2787 6147
rect 2813 6133 2827 6147
rect 2933 6133 2947 6147
rect 3053 6133 3067 6147
rect 3233 6133 3247 6147
rect 3273 6133 3287 6147
rect 3373 6133 3387 6147
rect 3413 6133 3427 6147
rect 3493 6133 3507 6147
rect 3573 6133 3587 6147
rect 3613 6133 3627 6147
rect 3853 6133 3867 6147
rect 3893 6133 3907 6147
rect 3993 6133 4007 6147
rect 4033 6133 4047 6147
rect 4573 6133 4587 6147
rect 4613 6133 4627 6147
rect 4713 6133 4727 6147
rect 4753 6133 4767 6147
rect 5233 6133 5247 6147
rect 5293 6133 5307 6147
rect 5873 6133 5887 6147
rect 5913 6133 5927 6147
rect 6053 6133 6067 6147
rect 6153 6153 6167 6167
rect 6233 6153 6247 6167
rect 293 6113 307 6127
rect 853 6113 867 6127
rect 1293 6113 1307 6127
rect 1433 6113 1447 6127
rect 1593 6113 1607 6127
rect 2093 6113 2107 6127
rect 2413 6113 2427 6127
rect 2453 6113 2467 6127
rect 3193 6113 3207 6127
rect 4373 6113 4387 6127
rect 4433 6113 4447 6127
rect 6153 6113 6167 6127
rect 6233 6113 6247 6127
rect 1473 6093 1487 6107
rect 1573 6093 1587 6107
rect 1653 6093 1667 6107
rect 1733 6093 1747 6107
rect 4813 6093 4827 6107
rect 4873 6093 4887 6107
rect 5073 6093 5087 6107
rect 5173 6093 5187 6107
rect 5333 6093 5347 6107
rect 5453 6093 5467 6107
rect 5653 6093 5667 6107
rect 113 6073 127 6087
rect 233 6073 247 6087
rect 373 6073 387 6087
rect 573 6073 587 6087
rect 613 6073 627 6087
rect 673 6073 687 6087
rect 933 6073 947 6087
rect 973 6073 987 6087
rect 1013 6073 1027 6087
rect 1113 6073 1127 6087
rect 1213 6073 1227 6087
rect 1273 6073 1287 6087
rect 1393 6073 1407 6087
rect 1893 6073 1907 6087
rect 1953 6073 1967 6087
rect 2053 6073 2067 6087
rect 2293 6073 2307 6087
rect 2573 6073 2587 6087
rect 2673 6073 2687 6087
rect 2733 6073 2747 6087
rect 2833 6073 2847 6087
rect 2953 6073 2967 6087
rect 3073 6073 3087 6087
rect 3293 6073 3307 6087
rect 3433 6073 3447 6087
rect 3473 6073 3487 6087
rect 3593 6073 3607 6087
rect 3713 6073 3727 6087
rect 3813 6073 3827 6087
rect 3873 6073 3887 6087
rect 3913 6073 3927 6087
rect 4053 6073 4067 6087
rect 4193 6073 4207 6087
rect 4253 6073 4267 6087
rect 4473 6073 4487 6087
rect 4633 6073 4647 6087
rect 773 6053 787 6067
rect 813 6053 827 6067
rect 1433 6053 1447 6067
rect 1493 6053 1507 6067
rect 113 6033 127 6047
rect 353 6033 367 6047
rect 773 6013 787 6027
rect 913 6013 927 6027
rect 973 6033 987 6047
rect 1033 6033 1047 6047
rect 1393 6033 1407 6047
rect 1673 6053 1687 6067
rect 1713 6053 1727 6067
rect 2133 6053 2147 6067
rect 2173 6053 2187 6067
rect 1893 6033 1907 6047
rect 2093 6033 2107 6047
rect 2433 6053 2447 6067
rect 2493 6053 2507 6067
rect 2393 6033 2407 6047
rect 2753 6033 2767 6047
rect 2953 6033 2967 6047
rect 4433 6053 4447 6067
rect 3773 6033 3787 6047
rect 3853 6033 3867 6047
rect 3893 6033 3907 6047
rect 4053 6033 4067 6047
rect 4233 6033 4247 6047
rect 5173 6053 5187 6067
rect 5333 6053 5347 6067
rect 5593 6053 5607 6067
rect 5853 6073 5867 6087
rect 5933 6073 5947 6087
rect 6013 6073 6027 6087
rect 6313 6073 6327 6087
rect 6513 6073 6527 6087
rect 5633 6033 5647 6047
rect 6173 6053 6187 6067
rect 6213 6053 6227 6067
rect 673 5993 687 6007
rect 873 5993 887 6007
rect 933 5993 947 6007
rect 1313 6013 1327 6027
rect 3213 6013 3227 6027
rect 3393 6013 3407 6027
rect 3933 6013 3947 6027
rect 4013 6013 4027 6027
rect 5193 6013 5207 6027
rect 5293 6013 5307 6027
rect 5933 6013 5947 6027
rect 6213 6013 6227 6027
rect 993 5993 1007 6007
rect 1293 5993 1307 6007
rect 1673 5993 1687 6007
rect 1793 5993 1807 6007
rect 2053 5993 2067 6007
rect 2153 5993 2167 6007
rect 2213 5993 2227 6007
rect 2313 5993 2327 6007
rect 2373 5993 2387 6007
rect 2433 5993 2447 6007
rect 2513 5993 2527 6007
rect 3273 5993 3287 6007
rect 853 5973 867 5987
rect 1093 5973 1107 5987
rect 1213 5973 1227 5987
rect 2013 5973 2027 5987
rect 2133 5973 2147 5987
rect 2293 5973 2307 5987
rect 173 5953 187 5967
rect 233 5953 247 5967
rect 1772 5953 1786 5967
rect 1794 5953 1808 5967
rect 2113 5953 2127 5967
rect 2193 5953 2207 5967
rect 2393 5953 2407 5967
rect 2493 5973 2507 5987
rect 2573 5973 2587 5987
rect 2713 5953 2727 5967
rect 3253 5973 3267 5987
rect 4473 5993 4487 6007
rect 4753 5993 4767 6007
rect 5173 5993 5187 6007
rect 5853 5993 5867 6007
rect 6013 5993 6027 6007
rect 3133 5953 3147 5967
rect 4193 5973 4207 5987
rect 4853 5973 4867 5987
rect 4133 5953 4147 5967
rect 4253 5953 4267 5967
rect 4473 5953 4487 5967
rect 4993 5973 5007 5987
rect 5033 5973 5047 5987
rect 5073 5973 5087 5987
rect 5113 5973 5127 5987
rect 5153 5973 5167 5987
rect 5293 5973 5307 5987
rect 5453 5973 5467 5987
rect 5893 5973 5907 5987
rect 6173 5973 6187 5987
rect 6313 5973 6327 5987
rect 4953 5954 4967 5968
rect 5193 5953 5207 5967
rect 5433 5953 5447 5967
rect 5553 5953 5567 5967
rect 5593 5953 5607 5967
rect 5773 5953 5787 5967
rect 6053 5953 6067 5967
rect 473 5933 487 5947
rect 673 5933 687 5947
rect 813 5933 827 5947
rect 973 5933 987 5947
rect 1053 5933 1067 5947
rect 1253 5933 1267 5947
rect 1353 5933 1367 5947
rect 1093 5913 1107 5927
rect 1133 5913 1147 5927
rect 1753 5933 1767 5947
rect 2353 5933 2367 5947
rect 2813 5933 2827 5947
rect 2033 5913 2047 5927
rect 2073 5913 2087 5927
rect 2193 5913 2207 5927
rect 2253 5913 2267 5927
rect 2393 5913 2407 5927
rect 2553 5913 2567 5927
rect 3033 5933 3047 5947
rect 3173 5933 3187 5947
rect 3433 5933 3447 5947
rect 3473 5933 3487 5947
rect 3513 5933 3527 5947
rect 3313 5913 3327 5927
rect 3353 5913 3367 5927
rect 3633 5913 3647 5927
rect 3833 5913 3847 5927
rect 3893 5913 3907 5927
rect 4233 5933 4247 5947
rect 4273 5933 4287 5947
rect 4513 5933 4527 5947
rect 4573 5933 4587 5947
rect 4953 5932 4967 5946
rect 4253 5913 4267 5927
rect 5133 5933 5147 5947
rect 5253 5933 5267 5947
rect 5573 5933 5587 5947
rect 5633 5933 5647 5947
rect 6013 5933 6027 5947
rect 6113 5933 6127 5947
rect 6213 5933 6227 5947
rect 5393 5913 5407 5927
rect 5433 5913 5447 5927
rect 6293 5913 6307 5927
rect 6333 5913 6347 5927
rect 153 5893 167 5907
rect 253 5893 267 5907
rect 353 5893 367 5907
rect 473 5893 487 5907
rect 593 5893 607 5907
rect 673 5893 687 5907
rect 833 5893 847 5907
rect 933 5893 947 5907
rect 1033 5893 1047 5907
rect 1253 5893 1267 5907
rect 1293 5893 1307 5907
rect 1413 5893 1427 5907
rect 1573 5893 1587 5907
rect 1613 5893 1627 5907
rect 1713 5893 1727 5907
rect 1833 5893 1847 5907
rect 2353 5893 2367 5907
rect 2513 5893 2527 5907
rect 2713 5893 2727 5907
rect 2753 5893 2767 5907
rect 2853 5893 2867 5907
rect 3053 5893 3067 5907
rect 3133 5893 3147 5907
rect 3553 5893 3567 5907
rect 3673 5893 3687 5907
rect 3713 5893 3727 5907
rect 3913 5893 3927 5907
rect 3993 5893 4007 5907
rect 4213 5893 4227 5907
rect 4373 5893 4387 5907
rect 4513 5893 4527 5907
rect 4633 5893 4647 5907
rect 4753 5893 4767 5907
rect 5093 5893 5107 5907
rect 5253 5893 5267 5907
rect 5573 5893 5587 5907
rect 5613 5893 5627 5907
rect 5773 5893 5787 5907
rect 5853 5893 5867 5907
rect 5893 5893 5907 5907
rect 6013 5893 6027 5907
rect 6053 5893 6067 5907
rect 6213 5893 6227 5907
rect 1073 5873 1087 5887
rect 3573 5873 3587 5887
rect 433 5853 447 5867
rect 1113 5853 1127 5867
rect 2073 5853 2087 5867
rect 2113 5853 2127 5867
rect 2273 5853 2287 5867
rect 2313 5853 2327 5867
rect 3153 5853 3167 5867
rect 3273 5853 3287 5867
rect 4912 5853 4926 5867
rect 4934 5853 4948 5867
rect 5173 5853 5187 5867
rect 5313 5853 5327 5867
rect 5533 5853 5547 5867
rect 133 5833 147 5847
rect 173 5833 187 5847
rect 293 5833 307 5847
rect 333 5833 347 5847
rect 493 5833 507 5847
rect 653 5833 667 5847
rect 693 5833 707 5847
rect 773 5833 787 5847
rect 813 5833 827 5847
rect 913 5833 927 5847
rect 953 5833 967 5847
rect 993 5813 1007 5827
rect 1353 5833 1367 5847
rect 1393 5833 1407 5847
rect 1433 5833 1447 5847
rect 1513 5833 1527 5847
rect 1553 5833 1567 5847
rect 1693 5833 1707 5847
rect 1733 5833 1747 5847
rect 1853 5833 1867 5847
rect 1893 5833 1907 5847
rect 2373 5833 2387 5847
rect 2413 5833 2427 5847
rect 2533 5833 2547 5847
rect 2573 5833 2587 5847
rect 2613 5833 2627 5847
rect 2833 5833 2847 5847
rect 2873 5833 2887 5847
rect 2993 5833 3007 5847
rect 3033 5833 3047 5847
rect 3473 5833 3487 5847
rect 3513 5833 3527 5847
rect 3613 5833 3627 5847
rect 3653 5833 3667 5847
rect 3753 5833 3767 5847
rect 3793 5833 3807 5847
rect 3833 5833 3847 5847
rect 3893 5833 3907 5847
rect 3933 5833 3947 5847
rect 4073 5833 4087 5847
rect 4113 5833 4127 5847
rect 4233 5833 4247 5847
rect 4273 5833 4287 5847
rect 4393 5833 4407 5847
rect 4453 5833 4467 5847
rect 4653 5833 4667 5847
rect 4693 5833 4707 5847
rect 5233 5833 5247 5847
rect 5273 5833 5287 5847
rect 5593 5833 5607 5847
rect 5713 5833 5727 5847
rect 5753 5833 5767 5847
rect 5873 5833 5887 5847
rect 5913 5833 5927 5847
rect 6073 5833 6087 5847
rect 6153 5833 6167 5847
rect 6193 5833 6207 5847
rect 2053 5813 2067 5827
rect 2093 5813 2107 5827
rect 2273 5813 2287 5827
rect 2453 5813 2467 5827
rect 4853 5813 4867 5827
rect 253 5793 267 5807
rect 433 5793 447 5807
rect 733 5793 747 5807
rect 913 5793 927 5807
rect 953 5793 967 5807
rect 1353 5793 1367 5807
rect 1413 5793 1427 5807
rect 1553 5793 1567 5807
rect 1613 5793 1627 5807
rect 1893 5793 1907 5807
rect 2373 5793 2387 5807
rect 2653 5793 2667 5807
rect 2993 5793 3007 5807
rect 3653 5793 3667 5807
rect 3713 5793 3727 5807
rect 3933 5793 3947 5807
rect 4193 5793 4207 5807
rect 4433 5793 4447 5807
rect 4572 5793 4586 5807
rect 4993 5793 5007 5807
rect 5033 5793 5047 5807
rect 5533 5813 5547 5827
rect 5813 5813 5827 5827
rect 5853 5813 5867 5827
rect 6253 5813 6267 5827
rect 6473 5813 6487 5827
rect 5433 5793 5447 5807
rect 5472 5793 5486 5807
rect 5573 5793 5587 5807
rect 5833 5793 5847 5807
rect 6013 5793 6027 5807
rect 6193 5793 6207 5807
rect 1113 5773 1127 5787
rect 1233 5773 1247 5787
rect 1753 5773 1767 5787
rect 1853 5773 1867 5787
rect 2233 5773 2247 5787
rect 2292 5773 2306 5787
rect 2353 5773 2367 5787
rect 2532 5773 2546 5787
rect 2554 5773 2568 5787
rect 2673 5773 2687 5787
rect 2733 5773 2747 5787
rect 2873 5773 2887 5787
rect 3093 5773 3107 5787
rect 3153 5773 3167 5787
rect 3213 5773 3227 5787
rect 93 5753 107 5767
rect 133 5753 147 5767
rect 833 5753 847 5767
rect 953 5753 967 5767
rect 13 5733 27 5747
rect 1313 5753 1327 5767
rect 1693 5753 1707 5767
rect 2153 5753 2167 5767
rect 2333 5753 2347 5767
rect 2613 5753 2627 5767
rect 2774 5753 2788 5767
rect 3233 5753 3247 5767
rect 3433 5753 3447 5767
rect 3513 5773 3527 5787
rect 4153 5773 4167 5787
rect 4833 5773 4847 5787
rect 1013 5733 1027 5747
rect 2233 5733 2247 5747
rect 2293 5733 2307 5747
rect 2493 5733 2507 5747
rect 2533 5733 2547 5747
rect 2893 5733 2907 5747
rect 2973 5733 2987 5747
rect 3253 5733 3267 5747
rect 3353 5733 3367 5747
rect 3553 5733 3567 5747
rect 3793 5753 3807 5767
rect 3873 5753 3887 5767
rect 3913 5753 3927 5767
rect 4213 5753 4227 5767
rect 4614 5753 4628 5767
rect 4653 5754 4667 5768
rect 4773 5753 4787 5767
rect 5113 5753 5127 5767
rect 6513 5773 6527 5787
rect 5233 5753 5247 5767
rect 5292 5753 5306 5767
rect 5353 5753 5367 5767
rect 5713 5753 5727 5767
rect 5873 5753 5887 5767
rect 6053 5753 6067 5767
rect 6093 5754 6107 5768
rect 6173 5753 6187 5767
rect 693 5713 707 5727
rect 853 5693 867 5707
rect 973 5693 987 5707
rect 1353 5693 1367 5707
rect 1513 5693 1527 5707
rect 2173 5713 2187 5727
rect 2573 5713 2587 5727
rect 3193 5713 3207 5727
rect 3513 5713 3527 5727
rect 3933 5713 3947 5727
rect 2593 5693 2607 5707
rect 353 5673 367 5687
rect 1213 5673 1227 5687
rect 1573 5673 1587 5687
rect 1733 5673 1747 5687
rect 1813 5673 1827 5687
rect 1993 5673 2007 5687
rect 2053 5673 2067 5687
rect 2353 5673 2367 5687
rect 2913 5693 2927 5707
rect 3173 5693 3187 5707
rect 3433 5693 3447 5707
rect 3673 5693 3687 5707
rect 413 5653 427 5667
rect 653 5653 667 5667
rect 1053 5653 1067 5667
rect 1113 5633 1127 5647
rect 1473 5653 1487 5667
rect 1613 5653 1627 5667
rect 1693 5653 1707 5667
rect 2093 5653 2107 5667
rect 2833 5673 2847 5687
rect 2573 5653 2587 5667
rect 2873 5653 2887 5667
rect 3153 5673 3167 5687
rect 3313 5674 3327 5688
rect 3853 5693 3867 5707
rect 3913 5693 3927 5707
rect 3973 5733 3987 5747
rect 4133 5733 4147 5747
rect 4453 5733 4467 5747
rect 4592 5733 4606 5747
rect 4653 5732 4667 5746
rect 4813 5733 4827 5747
rect 4873 5733 4887 5747
rect 4253 5713 4267 5727
rect 4833 5713 4847 5727
rect 4273 5693 4287 5707
rect 4753 5693 4767 5707
rect 5093 5713 5107 5727
rect 5213 5733 5227 5747
rect 5913 5733 5927 5747
rect 6093 5732 6107 5746
rect 5233 5713 5247 5727
rect 5353 5713 5367 5727
rect 6513 5713 6527 5727
rect 5333 5693 5347 5707
rect 5753 5693 5767 5707
rect 6373 5693 6387 5707
rect 6413 5693 6427 5707
rect 3313 5652 3327 5666
rect 4553 5673 4567 5687
rect 4673 5673 4687 5687
rect 4853 5673 4867 5687
rect 4913 5673 4927 5687
rect 3753 5653 3767 5667
rect 3893 5653 3907 5667
rect 4493 5653 4507 5667
rect 4613 5653 4627 5667
rect 4713 5653 4727 5667
rect 4873 5653 4887 5667
rect 4953 5653 4967 5667
rect 5033 5653 5047 5667
rect 2073 5633 2087 5647
rect 2173 5633 2187 5647
rect 3333 5633 3347 5647
rect 3553 5633 3567 5647
rect 3793 5633 3807 5647
rect 4053 5633 4067 5647
rect 4173 5633 4187 5647
rect 4393 5633 4407 5647
rect 4473 5633 4487 5647
rect 5413 5653 5427 5667
rect 5453 5653 5467 5667
rect 5653 5653 5667 5667
rect 5713 5653 5727 5667
rect 6213 5653 6227 5667
rect 6353 5653 6367 5667
rect 6453 5653 6467 5667
rect 6393 5633 6407 5647
rect 113 5613 127 5627
rect 153 5613 167 5627
rect 253 5613 267 5627
rect 293 5613 307 5627
rect 333 5613 347 5627
rect 373 5613 387 5627
rect 413 5613 427 5627
rect 453 5613 467 5627
rect 553 5613 567 5627
rect 593 5613 607 5627
rect 673 5613 687 5627
rect 713 5613 727 5627
rect 753 5613 767 5627
rect 793 5613 807 5627
rect 933 5613 947 5627
rect 973 5613 987 5627
rect 1013 5613 1027 5627
rect 1133 5613 1147 5627
rect 1173 5613 1187 5627
rect 1413 5613 1427 5627
rect 1453 5613 1467 5627
rect 1573 5613 1587 5627
rect 1613 5613 1627 5627
rect 1773 5613 1787 5627
rect 1813 5613 1827 5627
rect 1853 5613 1867 5627
rect 1913 5613 1927 5627
rect 1953 5613 1967 5627
rect 2213 5613 2227 5627
rect 2253 5613 2267 5627
rect 2513 5613 2527 5627
rect 2553 5613 2567 5627
rect 2653 5613 2667 5627
rect 2693 5613 2707 5627
rect 2793 5613 2807 5627
rect 2833 5613 2847 5627
rect 2953 5613 2967 5627
rect 2993 5613 3007 5627
rect 3133 5613 3147 5627
rect 3173 5613 3187 5627
rect 3393 5613 3407 5627
rect 3433 5613 3447 5627
rect 3653 5613 3667 5627
rect 3693 5613 3707 5627
rect 3733 5613 3747 5627
rect 3893 5613 3907 5627
rect 3933 5613 3947 5627
rect 3973 5613 3987 5627
rect 4513 5613 4527 5627
rect 4553 5613 4567 5627
rect 4673 5613 4687 5627
rect 4713 5613 4727 5627
rect 4813 5613 4827 5627
rect 4853 5613 4867 5627
rect 4993 5613 5007 5627
rect 5013 5613 5027 5627
rect 5453 5613 5467 5627
rect 5493 5613 5507 5627
rect 5613 5613 5627 5627
rect 5653 5613 5667 5627
rect 5793 5613 5807 5627
rect 5833 5613 5847 5627
rect 5973 5613 5987 5627
rect 6013 5613 6027 5627
rect 6333 5613 6347 5627
rect 6413 5613 6427 5627
rect 6453 5613 6467 5627
rect 1053 5593 1067 5607
rect 1093 5593 1107 5607
rect 1873 5593 1887 5607
rect 2353 5593 2367 5607
rect 4093 5593 4107 5607
rect 4173 5593 4187 5607
rect 4333 5593 4347 5607
rect 4393 5593 4407 5607
rect 4433 5593 4447 5607
rect 5053 5593 5067 5607
rect 5113 5593 5127 5607
rect 6093 5593 6107 5607
rect 6193 5593 6207 5607
rect 6373 5593 6387 5607
rect 6513 5593 6527 5607
rect 93 5553 107 5567
rect 133 5553 147 5567
rect 374 5553 388 5567
rect 433 5553 447 5567
rect 533 5553 547 5567
rect 613 5553 627 5567
rect 753 5553 767 5567
rect 833 5553 847 5567
rect 1033 5553 1047 5567
rect 1113 5553 1127 5567
rect 1313 5553 1327 5567
rect 1473 5553 1487 5567
rect 1553 5553 1567 5567
rect 1633 5553 1647 5567
rect 1694 5553 1708 5567
rect 1793 5553 1807 5567
rect 1973 5553 1987 5567
rect 2273 5553 2287 5567
rect 2333 5553 2347 5567
rect 2493 5553 2507 5567
rect 2533 5553 2547 5567
rect 2713 5553 2727 5567
rect 2933 5573 2947 5587
rect 3393 5573 3407 5587
rect 3873 5573 3887 5587
rect 2873 5553 2887 5567
rect 3013 5553 3027 5567
rect 3053 5553 3067 5567
rect 3193 5553 3207 5567
rect 3313 5553 3327 5567
rect 3573 5553 3587 5567
rect 3633 5553 3647 5567
rect 3713 5553 3727 5567
rect 3993 5553 4007 5567
rect 4053 5553 4067 5567
rect 4213 5553 4227 5567
rect 4413 5553 4427 5567
rect 4593 5553 4607 5567
rect 4653 5553 4667 5567
rect 4773 5553 4787 5567
rect 4973 5553 4987 5567
rect 5233 5553 5247 5567
rect 5373 5553 5387 5567
rect 5473 5553 5487 5567
rect 5633 5553 5647 5567
rect 5773 5553 5787 5567
rect 5953 5573 5967 5587
rect 5933 5553 5947 5567
rect 6033 5553 6047 5567
rect 6153 5553 6167 5567
rect 6273 5553 6287 5567
rect 6313 5553 6327 5567
rect 573 5533 587 5547
rect 133 5513 147 5527
rect 293 5513 307 5527
rect 473 5513 487 5527
rect 713 5513 727 5527
rect 1153 5533 1167 5547
rect 1313 5513 1327 5527
rect 1413 5513 1427 5527
rect 1773 5513 1787 5527
rect 2053 5533 2067 5547
rect 2093 5533 2107 5547
rect 1993 5513 2007 5527
rect 2233 5513 2247 5527
rect 2433 5513 2447 5527
rect 2513 5513 2527 5527
rect 3413 5533 3427 5547
rect 3453 5533 3467 5547
rect 3673 5533 3687 5547
rect 4093 5533 4107 5547
rect 4153 5533 4167 5547
rect 2693 5513 2707 5527
rect 3073 5513 3087 5527
rect 153 5493 167 5507
rect 253 5493 267 5507
rect 333 5493 347 5507
rect 613 5493 627 5507
rect 833 5493 847 5507
rect 1173 5493 1187 5507
rect 1333 5493 1347 5507
rect 1853 5493 1867 5507
rect 2093 5493 2107 5507
rect 2533 5493 2547 5507
rect 3033 5493 3047 5507
rect 3333 5493 3347 5507
rect 3373 5493 3387 5507
rect 3693 5513 3707 5527
rect 4053 5513 4067 5527
rect 4513 5513 4527 5527
rect 4633 5513 4647 5527
rect 3613 5493 3627 5507
rect 3893 5493 3907 5507
rect 4093 5494 4107 5508
rect 4193 5493 4207 5507
rect 4613 5493 4627 5507
rect 4654 5493 4668 5507
rect 4713 5493 4727 5507
rect 113 5473 127 5487
rect 573 5473 587 5487
rect 993 5473 1007 5487
rect 1433 5473 1447 5487
rect 1473 5473 1487 5487
rect 1533 5473 1547 5487
rect 1633 5473 1647 5487
rect 1993 5473 2007 5487
rect 2333 5473 2347 5487
rect 2393 5473 2407 5487
rect 2433 5473 2447 5487
rect 2733 5473 2747 5487
rect 3113 5473 3127 5487
rect 3393 5473 3407 5487
rect 3453 5473 3467 5487
rect 3493 5473 3507 5487
rect 3573 5473 3587 5487
rect 3693 5473 3707 5487
rect 3873 5473 3887 5487
rect 4093 5472 4107 5486
rect 4333 5473 4347 5487
rect 4413 5473 4427 5487
rect 4453 5473 4467 5487
rect 4853 5513 4867 5527
rect 5373 5513 5387 5527
rect 5433 5513 5447 5527
rect 5573 5513 5587 5527
rect 5633 5513 5647 5527
rect 5773 5513 5787 5527
rect 6033 5514 6047 5528
rect 6073 5513 6087 5527
rect 6133 5513 6147 5527
rect 6393 5513 6407 5527
rect 4753 5493 4767 5507
rect 5113 5493 5127 5507
rect 4793 5473 4807 5487
rect 5473 5493 5487 5507
rect 5513 5493 5527 5507
rect 5613 5493 5627 5507
rect 5793 5493 5807 5507
rect 6033 5492 6047 5506
rect 6513 5493 6527 5507
rect 5293 5473 5307 5487
rect 5773 5473 5787 5487
rect 5973 5473 5987 5487
rect 6093 5473 6107 5487
rect 6333 5473 6347 5487
rect 493 5453 507 5467
rect 553 5453 567 5467
rect 1793 5453 1807 5467
rect 1953 5453 1967 5467
rect 2133 5453 2147 5467
rect 2533 5453 2547 5467
rect 2593 5453 2607 5467
rect 2793 5453 2807 5467
rect 2853 5453 2867 5467
rect 3273 5453 3287 5467
rect 3633 5453 3647 5467
rect 3833 5453 3847 5467
rect 3993 5453 4007 5467
rect 4033 5453 4047 5467
rect 4253 5453 4267 5467
rect 4473 5453 4487 5467
rect 4613 5453 4627 5467
rect 4673 5453 4687 5467
rect 4833 5453 4847 5467
rect 4953 5453 4967 5467
rect 5053 5453 5067 5467
rect 5133 5453 5147 5467
rect 5273 5453 5287 5467
rect 5333 5453 5347 5467
rect 5372 5453 5386 5467
rect 5394 5453 5408 5467
rect 5713 5453 5727 5467
rect 5893 5453 5907 5467
rect 6073 5453 6087 5467
rect 6253 5453 6267 5467
rect 6453 5453 6467 5467
rect 333 5433 347 5447
rect 673 5433 687 5447
rect 853 5433 867 5447
rect 893 5433 907 5447
rect 1153 5433 1167 5447
rect 1673 5433 1687 5447
rect 2033 5433 2047 5447
rect 2633 5433 2647 5447
rect 2673 5433 2687 5447
rect 3113 5433 3127 5447
rect 3173 5433 3187 5447
rect 3334 5433 3348 5447
rect 3413 5433 3427 5447
rect 3473 5433 3487 5447
rect 3713 5433 3727 5447
rect 3913 5433 3927 5447
rect 4093 5433 4107 5447
rect 4753 5433 4767 5447
rect 4993 5433 5007 5447
rect 5353 5433 5367 5447
rect 5493 5433 5507 5447
rect 5552 5433 5566 5447
rect 5593 5433 5607 5447
rect 5933 5433 5947 5447
rect 6273 5433 6287 5447
rect 6313 5434 6327 5448
rect 433 5413 447 5427
rect 493 5413 507 5427
rect 653 5413 667 5427
rect 1293 5413 1307 5427
rect 1233 5393 1247 5407
rect 1333 5393 1347 5407
rect 1713 5413 1727 5427
rect 2273 5413 2287 5427
rect 2413 5413 2427 5427
rect 2133 5393 2147 5407
rect 2173 5393 2187 5407
rect 2453 5393 2467 5407
rect 2493 5393 2507 5407
rect 2633 5393 2647 5407
rect 2912 5413 2926 5427
rect 2934 5413 2948 5427
rect 2973 5413 2987 5427
rect 3273 5413 3287 5427
rect 3313 5413 3327 5427
rect 3353 5413 3367 5427
rect 3433 5413 3447 5427
rect 3793 5413 3807 5427
rect 3834 5413 3848 5427
rect 3893 5413 3907 5427
rect 4173 5413 4187 5427
rect 4213 5413 4227 5427
rect 4493 5413 4507 5427
rect 4573 5413 4587 5427
rect 4633 5413 4647 5427
rect 4713 5413 4727 5427
rect 5013 5413 5027 5427
rect 5053 5413 5067 5427
rect 5213 5413 5227 5427
rect 5393 5413 5407 5427
rect 5613 5413 5627 5427
rect 5693 5413 5707 5427
rect 6153 5413 6167 5427
rect 6313 5412 6327 5426
rect 6373 5413 6387 5427
rect 6433 5413 6447 5427
rect 3073 5393 3087 5407
rect 3113 5393 3127 5407
rect 3233 5393 3247 5407
rect 3673 5393 3687 5407
rect 3713 5393 3727 5407
rect 73 5373 87 5387
rect 273 5373 287 5387
rect 393 5373 407 5387
rect 493 5373 507 5387
rect 553 5373 567 5387
rect 673 5373 687 5387
rect 733 5373 747 5387
rect 873 5373 887 5387
rect 973 5373 987 5387
rect 1133 5373 1147 5387
rect 1213 5373 1227 5387
rect 1373 5373 1387 5387
rect 1533 5373 1547 5387
rect 1573 5373 1587 5387
rect 1693 5373 1707 5387
rect 1793 5373 1807 5387
rect 1873 5373 1887 5387
rect 2033 5373 2047 5387
rect 2373 5373 2387 5387
rect 2593 5373 2607 5387
rect 2753 5373 2767 5387
rect 2953 5373 2967 5387
rect 2993 5373 3007 5387
rect 3033 5373 3047 5387
rect 3433 5373 3447 5387
rect 3473 5373 3487 5387
rect 3633 5373 3647 5387
rect 3753 5373 3767 5387
rect 3993 5373 4007 5387
rect 5333 5393 5347 5407
rect 5493 5393 5507 5407
rect 5533 5393 5547 5407
rect 5933 5393 5947 5407
rect 5973 5393 5987 5407
rect 6173 5393 6187 5407
rect 6513 5393 6527 5407
rect 4453 5373 4467 5387
rect 4633 5373 4647 5387
rect 4673 5373 4687 5387
rect 4733 5373 4747 5387
rect 4773 5373 4787 5387
rect 5053 5373 5067 5387
rect 5093 5373 5107 5387
rect 5273 5373 5287 5387
rect 5393 5373 5407 5387
rect 5633 5373 5647 5387
rect 5713 5373 5727 5387
rect 5753 5373 5767 5387
rect 5893 5373 5907 5387
rect 6133 5373 6147 5387
rect 6293 5373 6307 5387
rect 6433 5373 6447 5387
rect 6473 5373 6487 5387
rect 793 5353 807 5367
rect 833 5353 847 5367
rect 1453 5353 1467 5367
rect 2113 5333 2127 5347
rect 2193 5333 2207 5347
rect 3053 5333 3067 5347
rect 3133 5333 3147 5347
rect 3333 5333 3347 5347
rect 3653 5333 3667 5347
rect 3693 5333 3707 5347
rect 3733 5333 3747 5347
rect 4073 5333 4087 5347
rect 4273 5333 4287 5347
rect 4353 5333 4367 5347
rect 4393 5333 4407 5347
rect 4833 5333 4847 5347
rect 4953 5333 4967 5347
rect 5213 5333 5227 5347
rect 5333 5333 5347 5347
rect 5913 5333 5927 5347
rect 5993 5333 6007 5347
rect 113 5313 127 5327
rect 153 5313 167 5327
rect 293 5313 307 5327
rect 333 5313 347 5327
rect 473 5313 487 5327
rect 513 5313 527 5327
rect 653 5313 667 5327
rect 693 5313 707 5327
rect 753 5313 767 5327
rect 813 5313 827 5327
rect 853 5313 867 5327
rect 893 5313 907 5327
rect 1013 5313 1027 5327
rect 1053 5313 1067 5327
rect 1153 5313 1167 5327
rect 1193 5313 1207 5327
rect 1313 5313 1327 5327
rect 1353 5313 1367 5327
rect 1393 5313 1407 5327
rect 1473 5313 1487 5327
rect 1513 5313 1527 5327
rect 1673 5313 1687 5327
rect 1713 5313 1727 5327
rect 1813 5313 1827 5327
rect 1853 5313 1867 5327
rect 1973 5313 1987 5327
rect 2013 5313 2027 5327
rect 1373 5293 1387 5307
rect 1533 5293 1547 5307
rect 1573 5293 1587 5307
rect 2033 5293 2047 5307
rect 2333 5313 2347 5327
rect 2473 5313 2487 5327
rect 2613 5313 2627 5327
rect 2653 5313 2667 5327
rect 2773 5313 2787 5327
rect 2893 5313 2907 5327
rect 2933 5313 2947 5327
rect 2293 5293 2307 5307
rect 393 5273 407 5287
rect 513 5273 527 5287
rect 1053 5273 1067 5287
rect 1093 5273 1107 5287
rect 2493 5273 2507 5287
rect 3013 5293 3027 5307
rect 3213 5313 3227 5327
rect 3413 5313 3427 5327
rect 3453 5313 3467 5327
rect 3493 5313 3507 5327
rect 3533 5313 3547 5327
rect 3133 5293 3147 5307
rect 3173 5293 3187 5307
rect 3653 5293 3667 5307
rect 3853 5313 3867 5327
rect 3893 5313 3907 5327
rect 4013 5313 4027 5327
rect 4513 5313 4527 5327
rect 4553 5313 4567 5327
rect 4673 5313 4687 5327
rect 4713 5313 4727 5327
rect 5073 5313 5087 5327
rect 5113 5313 5127 5327
rect 5373 5313 5387 5327
rect 5653 5313 5667 5327
rect 5773 5313 5787 5327
rect 5813 5313 5827 5327
rect 5953 5313 5967 5327
rect 6113 5313 6127 5327
rect 6153 5313 6167 5327
rect 6313 5313 6327 5327
rect 6413 5313 6427 5327
rect 6453 5313 6467 5327
rect 4473 5293 4487 5307
rect 4953 5293 4967 5307
rect 5053 5293 5067 5307
rect 5993 5293 6007 5307
rect 2833 5273 2847 5287
rect 2913 5273 2927 5287
rect 2953 5273 2967 5287
rect 3053 5273 3067 5287
rect 3093 5273 3107 5287
rect 3193 5274 3207 5288
rect 473 5253 487 5267
rect 693 5253 707 5267
rect 1313 5253 1327 5267
rect 1473 5253 1487 5267
rect 1713 5253 1727 5267
rect 2113 5253 2127 5267
rect 3153 5253 3167 5267
rect 3193 5252 3207 5266
rect 3393 5273 3407 5287
rect 3573 5273 3587 5287
rect 3973 5273 3987 5287
rect 4013 5273 4027 5287
rect 4293 5273 4307 5287
rect 3433 5253 3447 5267
rect 3693 5253 3707 5267
rect 3733 5253 3747 5267
rect 4053 5253 4067 5267
rect 4653 5273 4667 5287
rect 5073 5273 5087 5287
rect 5213 5273 5227 5287
rect 5273 5273 5287 5287
rect 5653 5273 5667 5287
rect 5813 5273 5827 5287
rect 5953 5274 5967 5288
rect 6393 5273 6407 5287
rect 6453 5273 6467 5287
rect 4973 5253 4987 5267
rect 5713 5253 5727 5267
rect 5953 5252 5967 5266
rect 6073 5253 6087 5267
rect 6313 5253 6327 5267
rect 813 5233 827 5247
rect 1233 5233 1247 5247
rect 1413 5233 1427 5247
rect 1533 5233 1547 5247
rect 1793 5233 1807 5247
rect 1913 5233 1927 5247
rect 2073 5233 2087 5247
rect 2393 5233 2407 5247
rect 2493 5233 2507 5247
rect 2933 5233 2947 5247
rect 3233 5233 3247 5247
rect 3373 5233 3387 5247
rect 3453 5233 3467 5247
rect 3532 5233 3546 5247
rect 3554 5233 3568 5247
rect 3873 5233 3887 5247
rect 4553 5233 4567 5247
rect 1193 5213 1207 5227
rect 1393 5213 1407 5227
rect 1853 5213 1867 5227
rect 1973 5213 1987 5227
rect 2153 5213 2167 5227
rect 2693 5213 2707 5227
rect 3073 5213 3087 5227
rect 3353 5213 3367 5227
rect 4773 5233 4787 5247
rect 4813 5233 4827 5247
rect 4073 5213 4087 5227
rect 4193 5213 4207 5227
rect 293 5193 307 5207
rect 413 5193 427 5207
rect 1293 5193 1307 5207
rect 1813 5193 1827 5207
rect 2133 5193 2147 5207
rect 2413 5193 2427 5207
rect 2653 5193 2667 5207
rect 3193 5193 3207 5207
rect 113 5173 127 5187
rect 313 5173 327 5187
rect 593 5173 607 5187
rect 733 5173 747 5187
rect 933 5173 947 5187
rect 973 5173 987 5187
rect 1053 5173 1067 5187
rect 1093 5173 1107 5187
rect 1433 5173 1447 5187
rect 1533 5173 1547 5187
rect 1913 5173 1927 5187
rect 2013 5173 2027 5187
rect 2253 5173 2267 5187
rect 2333 5173 2347 5187
rect 2573 5173 2587 5187
rect 2993 5173 3007 5187
rect 3293 5173 3307 5187
rect 3453 5173 3467 5187
rect 3713 5173 3727 5187
rect 3773 5173 3787 5187
rect 3933 5173 3947 5187
rect 3973 5174 3987 5188
rect 4573 5193 4587 5207
rect 4633 5193 4647 5207
rect 4713 5213 4727 5227
rect 5073 5213 5087 5227
rect 5193 5233 5207 5247
rect 5553 5233 5567 5247
rect 5533 5213 5547 5227
rect 5693 5213 5707 5227
rect 5773 5213 5787 5227
rect 5873 5213 5887 5227
rect 5913 5213 5927 5227
rect 6293 5213 6307 5227
rect 6473 5213 6487 5227
rect 4993 5193 5007 5207
rect 6233 5193 6247 5207
rect 6413 5193 6427 5207
rect 6453 5193 6467 5207
rect 6153 5174 6167 5188
rect 6373 5173 6387 5187
rect 6473 5173 6487 5187
rect 273 5153 287 5167
rect 633 5153 647 5167
rect 1153 5153 1167 5167
rect 2233 5153 2247 5167
rect 2773 5153 2787 5167
rect 3093 5153 3107 5167
rect 3552 5153 3566 5167
rect 3574 5153 3588 5167
rect 3633 5153 3647 5167
rect 3693 5153 3707 5167
rect 3813 5153 3827 5167
rect 3973 5152 3987 5166
rect 73 5133 87 5147
rect 113 5133 127 5147
rect 153 5133 167 5147
rect 233 5133 247 5147
rect 533 5133 547 5147
rect 1113 5133 1127 5147
rect 1193 5133 1207 5147
rect 1372 5133 1386 5147
rect 1394 5133 1408 5147
rect 1513 5133 1527 5147
rect 1873 5133 1887 5147
rect 2093 5133 2107 5147
rect 2193 5133 2207 5147
rect 2433 5133 2447 5147
rect 2533 5133 2547 5147
rect 2612 5133 2626 5147
rect 3293 5133 3307 5147
rect 3333 5133 3347 5147
rect 3513 5133 3527 5147
rect 493 5113 507 5127
rect 2673 5113 2687 5127
rect 2733 5113 2747 5127
rect 2774 5113 2788 5127
rect 113 5093 127 5107
rect 153 5093 167 5107
rect 233 5093 247 5107
rect 273 5093 287 5107
rect 313 5093 327 5107
rect 433 5093 447 5107
rect 473 5093 487 5107
rect 593 5093 607 5107
rect 633 5093 647 5107
rect 873 5093 887 5107
rect 913 5093 927 5107
rect 953 5093 967 5107
rect 993 5093 1007 5107
rect 1033 5093 1047 5107
rect 1073 5093 1087 5107
rect 1193 5093 1207 5107
rect 1233 5093 1247 5107
rect 1353 5093 1367 5107
rect 1393 5093 1407 5107
rect 1513 5093 1527 5107
rect 1553 5093 1567 5107
rect 1693 5093 1707 5107
rect 1733 5093 1747 5107
rect 1873 5093 1887 5107
rect 1913 5093 1927 5107
rect 2033 5093 2047 5107
rect 2073 5093 2087 5107
rect 2213 5093 2227 5107
rect 2253 5093 2267 5107
rect 2353 5093 2367 5107
rect 2393 5093 2407 5107
rect 2533 5093 2547 5107
rect 2573 5093 2587 5107
rect 2913 5093 2927 5107
rect 3493 5113 3507 5127
rect 3653 5133 3667 5147
rect 3914 5133 3928 5147
rect 4252 5153 4266 5167
rect 4274 5153 4288 5167
rect 4773 5153 4787 5167
rect 4853 5153 4867 5167
rect 5913 5153 5927 5167
rect 6153 5152 6167 5166
rect 6253 5153 6267 5167
rect 4173 5133 4187 5147
rect 4373 5133 4387 5147
rect 4413 5133 4427 5147
rect 4813 5133 4827 5147
rect 3153 5093 3167 5107
rect 3293 5093 3307 5107
rect 3333 5093 3347 5107
rect 3433 5093 3447 5107
rect 3473 5093 3487 5107
rect 3673 5113 3687 5127
rect 4073 5113 4087 5127
rect 3773 5093 3787 5107
rect 3813 5093 3827 5107
rect 3873 5093 3887 5107
rect 3933 5093 3947 5107
rect 3973 5093 3987 5107
rect 4253 5093 4267 5107
rect 4293 5093 4307 5107
rect 4393 5093 4407 5107
rect 4693 5113 4707 5127
rect 4793 5113 4807 5127
rect 5633 5133 5647 5147
rect 6233 5133 6247 5147
rect 5613 5113 5627 5127
rect 5653 5112 5667 5126
rect 5714 5113 5728 5127
rect 5753 5113 5767 5127
rect 5793 5113 5807 5127
rect 5013 5093 5027 5107
rect 5173 5093 5187 5107
rect 5213 5093 5227 5107
rect 5473 5093 5487 5107
rect 5513 5093 5527 5107
rect 5913 5093 5927 5107
rect 5953 5093 5967 5107
rect 6033 5093 6047 5107
rect 6073 5093 6087 5107
rect 6193 5093 6207 5107
rect 6233 5093 6247 5107
rect 13 5073 27 5087
rect 2613 5073 2627 5087
rect 2733 5073 2747 5087
rect 3573 5073 3587 5087
rect 3653 5073 3667 5087
rect 4013 5073 4027 5087
rect 4753 5073 4767 5087
rect 4813 5073 4827 5087
rect 5073 5073 5087 5087
rect 5653 5073 5667 5087
rect 5773 5073 5787 5087
rect 2593 5053 2607 5067
rect 73 5033 87 5047
rect 133 5033 147 5047
rect 253 5033 267 5047
rect 393 5033 407 5047
rect 493 5033 507 5047
rect 573 5033 587 5047
rect 733 5033 747 5047
rect 793 5033 807 5047
rect 933 5033 947 5047
rect 1053 5033 1067 5047
rect 1253 5033 1267 5047
rect 1333 5033 1347 5047
rect 1373 5033 1387 5047
rect 1413 5033 1427 5047
rect 1573 5033 1587 5047
rect 1753 5033 1767 5047
rect 1893 5033 1907 5047
rect 2013 5033 2027 5047
rect 2093 5033 2107 5047
rect 2173 5033 2187 5047
rect 2233 5033 2247 5047
rect 2333 5033 2347 5047
rect 2433 5033 2447 5047
rect 2693 5033 2707 5047
rect 3213 5033 3227 5047
rect 3413 5053 3427 5067
rect 3373 5033 3387 5047
rect 3493 5033 3507 5047
rect 3673 5033 3687 5047
rect 3833 5033 3847 5047
rect 3912 5033 3926 5047
rect 4213 5033 4227 5047
rect 4393 5033 4407 5047
rect 4553 5033 4567 5047
rect 4713 5033 4727 5047
rect 4853 5033 4867 5047
rect 4893 5033 4907 5047
rect 5113 5033 5127 5047
rect 5293 5033 5307 5047
rect 5433 5033 5447 5047
rect 5533 5033 5547 5047
rect 6013 5033 6027 5047
rect 6053 5033 6067 5047
rect 6113 5033 6127 5047
rect 6313 5033 6327 5047
rect 293 5013 307 5027
rect 613 5013 627 5027
rect 893 5013 907 5027
rect 1493 5013 1507 5027
rect 133 4993 147 5007
rect 253 4993 267 5007
rect 313 4993 327 5007
rect 493 4993 507 5007
rect 573 4993 587 5007
rect 1213 4993 1227 5007
rect 1253 4993 1267 5007
rect 1293 4993 1307 5007
rect 1333 4993 1347 5007
rect 1553 4993 1567 5007
rect 1713 4993 1727 5007
rect 553 4973 567 4987
rect 1453 4973 1467 4987
rect 1633 4973 1647 4987
rect 1753 4973 1767 4987
rect 1793 4973 1807 4987
rect 1893 4993 1907 5007
rect 2033 4993 2047 5007
rect 2073 4993 2087 5007
rect 2133 4993 2147 5007
rect 2793 5013 2807 5027
rect 2892 5013 2906 5027
rect 2973 5013 2987 5027
rect 3033 5013 3047 5027
rect 3593 5013 3607 5027
rect 3633 5013 3647 5027
rect 4073 5013 4087 5027
rect 4113 5013 4127 5027
rect 5233 5013 5247 5027
rect 5313 5013 5327 5027
rect 5633 5013 5647 5027
rect 5673 5013 5687 5027
rect 5753 5013 5767 5027
rect 5793 5013 5807 5027
rect 5873 5013 5887 5027
rect 6353 5013 6367 5027
rect 6513 5013 6527 5027
rect 2513 4993 2527 5007
rect 2553 4993 2567 5007
rect 2693 4993 2707 5007
rect 2873 4993 2887 5007
rect 2912 4993 2926 5007
rect 2953 4993 2967 5007
rect 1873 4973 1887 4987
rect 2313 4973 2327 4987
rect 2633 4973 2647 4987
rect 3073 4993 3087 5007
rect 3233 4993 3247 5007
rect 3333 4994 3347 5008
rect 3673 4993 3687 5007
rect 3853 4993 3867 5007
rect 3913 4993 3927 5007
rect 4033 4993 4047 5007
rect 4193 4993 4207 5007
rect 4693 4993 4707 5007
rect 5153 4993 5167 5007
rect 5253 4993 5267 5007
rect 5473 4993 5487 5007
rect 5973 4993 5987 5007
rect 6073 4993 6087 5007
rect 3153 4973 3167 4987
rect 3333 4972 3347 4986
rect 3933 4973 3947 4987
rect 4073 4973 4087 4987
rect 4113 4973 4127 4987
rect 4513 4973 4527 4987
rect 4633 4973 4647 4987
rect 4733 4973 4747 4987
rect 5093 4973 5107 4987
rect 5333 4973 5347 4987
rect 5413 4973 5427 4987
rect 5673 4973 5687 4987
rect 5713 4973 5727 4987
rect 5893 4973 5907 4987
rect 6113 4973 6127 4987
rect 893 4953 907 4967
rect 1673 4953 1687 4967
rect 2033 4953 2047 4967
rect 2413 4953 2427 4967
rect 2833 4953 2847 4967
rect 2953 4953 2967 4967
rect 3033 4953 3047 4967
rect 3573 4953 3587 4967
rect 3613 4953 3627 4967
rect 4033 4953 4047 4967
rect 4233 4953 4247 4967
rect 4413 4953 4427 4967
rect 173 4933 187 4947
rect 393 4933 407 4947
rect 973 4933 987 4947
rect 1233 4933 1247 4947
rect 1453 4933 1467 4947
rect 1533 4933 1547 4947
rect 1573 4933 1587 4947
rect 1693 4933 1707 4947
rect 2193 4933 2207 4947
rect 2233 4933 2247 4947
rect 2373 4933 2387 4947
rect 2913 4933 2927 4947
rect 3053 4933 3067 4947
rect 3233 4933 3247 4947
rect 3293 4933 3307 4947
rect 3633 4933 3647 4947
rect 3953 4933 3967 4947
rect 4113 4933 4127 4947
rect 4313 4933 4327 4947
rect 293 4913 307 4927
rect 473 4913 487 4927
rect 653 4913 667 4927
rect 853 4913 867 4927
rect 1013 4913 1027 4927
rect 1733 4913 1747 4927
rect 2153 4913 2167 4927
rect 2313 4913 2327 4927
rect 93 4893 107 4907
rect 153 4893 167 4907
rect 413 4893 427 4907
rect 613 4893 627 4907
rect 713 4893 727 4907
rect 1293 4893 1307 4907
rect 1514 4893 1528 4907
rect 1613 4893 1627 4907
rect 2113 4893 2127 4907
rect 2232 4893 2246 4907
rect 2254 4893 2268 4907
rect 2733 4893 2747 4907
rect 2873 4893 2887 4907
rect 2973 4913 2987 4927
rect 3013 4913 3027 4927
rect 3133 4913 3147 4927
rect 2993 4893 3007 4907
rect 3073 4893 3087 4907
rect 3533 4913 3547 4927
rect 4233 4913 4247 4927
rect 4613 4953 4627 4967
rect 4813 4953 4827 4967
rect 5053 4953 5067 4967
rect 5313 4953 5327 4967
rect 5433 4953 5447 4967
rect 5613 4953 5627 4967
rect 6093 4953 6107 4967
rect 6253 4953 6267 4967
rect 6313 4953 6327 4967
rect 4473 4933 4487 4947
rect 4693 4933 4707 4947
rect 5293 4933 5307 4947
rect 6053 4933 6067 4947
rect 4553 4913 4567 4927
rect 4733 4913 4747 4927
rect 4833 4913 4847 4927
rect 4933 4913 4947 4927
rect 3692 4893 3706 4907
rect 453 4873 467 4887
rect 493 4873 507 4887
rect 813 4873 827 4887
rect 853 4873 867 4887
rect 933 4873 947 4887
rect 973 4873 987 4887
rect 1673 4873 1687 4887
rect 1713 4873 1727 4887
rect 1853 4873 1867 4887
rect 2273 4873 2287 4887
rect 2393 4873 2407 4887
rect 2453 4873 2467 4887
rect 2533 4873 2547 4887
rect 2693 4873 2707 4887
rect 93 4853 107 4867
rect 253 4853 267 4867
rect 293 4853 307 4867
rect 373 4853 387 4867
rect 433 4853 447 4867
rect 533 4853 547 4867
rect 673 4853 687 4867
rect 1013 4853 1027 4867
rect 1133 4853 1147 4867
rect 1233 4853 1247 4867
rect 1453 4853 1467 4867
rect 1973 4853 1987 4867
rect 2093 4853 2107 4867
rect 2133 4853 2147 4867
rect 2192 4853 2206 4867
rect 2214 4853 2228 4867
rect 2493 4853 2507 4867
rect 2733 4853 2747 4867
rect 3113 4873 3127 4887
rect 3153 4873 3167 4887
rect 3293 4873 3307 4887
rect 3333 4873 3347 4887
rect 3573 4873 3587 4887
rect 3893 4893 3907 4907
rect 4133 4893 4147 4907
rect 4593 4893 4607 4907
rect 4633 4893 4647 4907
rect 4713 4893 4727 4907
rect 4893 4893 4907 4907
rect 5013 4893 5027 4907
rect 5093 4893 5107 4907
rect 5133 4893 5147 4907
rect 5433 4913 5447 4927
rect 5473 4913 5487 4927
rect 5652 4913 5666 4927
rect 5713 4913 5727 4927
rect 5773 4913 5787 4927
rect 6273 4913 6287 4927
rect 6493 4913 6507 4927
rect 5733 4893 5747 4907
rect 5852 4893 5866 4907
rect 5874 4893 5888 4907
rect 3833 4873 3847 4887
rect 5253 4873 5267 4887
rect 5293 4873 5307 4887
rect 5573 4873 5587 4887
rect 5613 4873 5627 4887
rect 6213 4873 6227 4887
rect 6253 4873 6267 4887
rect 6373 4873 6387 4887
rect 6413 4873 6427 4887
rect 2913 4853 2927 4867
rect 3033 4853 3047 4867
rect 3453 4853 3467 4867
rect 3533 4853 3547 4867
rect 3613 4853 3627 4867
rect 3713 4853 3727 4867
rect 3893 4853 3907 4867
rect 3953 4853 3967 4867
rect 4033 4853 4047 4867
rect 4133 4853 4147 4867
rect 4233 4853 4247 4867
rect 4433 4853 4447 4867
rect 4793 4853 4807 4867
rect 4933 4853 4947 4867
rect 4993 4853 5007 4867
rect 5173 4853 5187 4867
rect 5213 4853 5227 4867
rect 5333 4853 5347 4867
rect 5473 4853 5487 4867
rect 5653 4853 5667 4867
rect 5753 4853 5767 4867
rect 5873 4853 5887 4867
rect 5913 4853 5927 4867
rect 6113 4853 6127 4867
rect 1173 4833 1187 4847
rect 1733 4833 1747 4847
rect 1793 4833 1807 4847
rect 2853 4833 2867 4847
rect 873 4813 887 4827
rect 2453 4813 2467 4827
rect 2513 4813 2527 4827
rect 2753 4813 2767 4827
rect 3233 4813 3247 4827
rect 3273 4813 3287 4827
rect 3353 4813 3367 4827
rect 3853 4813 3867 4827
rect 4253 4813 4267 4827
rect 4313 4813 4327 4827
rect 4893 4813 4907 4827
rect 4973 4813 4987 4827
rect 5193 4813 5207 4827
rect 5233 4813 5247 4827
rect 5313 4813 5327 4827
rect 5693 4813 5707 4827
rect 6173 4813 6187 4827
rect 6273 4813 6287 4827
rect 73 4793 87 4807
rect 113 4793 127 4807
rect 153 4793 167 4807
rect 413 4793 427 4807
rect 453 4793 467 4807
rect 573 4793 587 4807
rect 653 4793 667 4807
rect 693 4793 707 4807
rect 1113 4793 1127 4807
rect 1153 4793 1167 4807
rect 1193 4793 1207 4807
rect 1253 4793 1267 4807
rect 1293 4793 1307 4807
rect 1533 4793 1547 4807
rect 1573 4793 1587 4807
rect 1833 4793 1847 4807
rect 1873 4793 1887 4807
rect 1993 4793 2007 4807
rect 2033 4793 2047 4807
rect 2153 4793 2167 4807
rect 2193 4793 2207 4807
rect 2313 4793 2327 4807
rect 2353 4793 2367 4807
rect 2793 4793 2807 4807
rect 2833 4793 2847 4807
rect 3013 4793 3027 4807
rect 3313 4793 3327 4807
rect 3473 4793 3487 4807
rect 3593 4793 3607 4807
rect 3633 4793 3647 4807
rect 3733 4793 3747 4807
rect 4073 4793 4087 4807
rect 4193 4793 4207 4807
rect 4453 4793 4467 4807
rect 4533 4793 4547 4807
rect 4573 4793 4587 4807
rect 4613 4793 4627 4807
rect 4733 4793 4747 4807
rect 4773 4793 4787 4807
rect 5053 4793 5067 4807
rect 5093 4793 5107 4807
rect 973 4773 987 4787
rect 1053 4773 1067 4787
rect 113 4753 127 4767
rect 173 4753 187 4767
rect 293 4753 307 4767
rect 493 4753 507 4767
rect 1153 4753 1167 4767
rect 1213 4753 1227 4767
rect 1253 4753 1267 4767
rect 2433 4773 2447 4787
rect 2633 4773 2647 4787
rect 3053 4773 3067 4787
rect 3873 4773 3887 4787
rect 4793 4773 4807 4787
rect 5013 4773 5027 4787
rect 5273 4793 5287 4807
rect 5413 4793 5427 4807
rect 5453 4793 5467 4807
rect 5733 4793 5747 4807
rect 5773 4793 5787 4807
rect 5853 4793 5867 4807
rect 5893 4793 5907 4807
rect 6053 4793 6067 4807
rect 6093 4793 6107 4807
rect 5253 4773 5267 4787
rect 5313 4773 5327 4787
rect 5493 4773 5507 4787
rect 5553 4773 5567 4787
rect 5693 4773 5707 4787
rect 6133 4773 6147 4787
rect 6213 4773 6227 4787
rect 1612 4753 1626 4767
rect 1634 4753 1648 4767
rect 2073 4753 2087 4767
rect 2193 4753 2207 4767
rect 2353 4753 2367 4767
rect 2453 4753 2467 4767
rect 2753 4753 2767 4767
rect 3112 4753 3126 4767
rect 3134 4753 3148 4767
rect 3353 4753 3367 4767
rect 3813 4753 3827 4767
rect 3853 4753 3867 4767
rect 3893 4753 3907 4767
rect 3933 4753 3947 4767
rect 4073 4753 4087 4767
rect 4173 4753 4187 4767
rect 4453 4753 4467 4767
rect 4533 4753 4547 4767
rect 5333 4753 5347 4767
rect 5393 4753 5407 4767
rect 5453 4753 5467 4767
rect 1513 4733 1527 4747
rect 1673 4733 1687 4747
rect 1713 4733 1727 4747
rect 2373 4733 2387 4747
rect 733 4713 747 4727
rect 853 4713 867 4727
rect 913 4713 927 4727
rect 1533 4713 1547 4727
rect 2292 4713 2306 4727
rect 2314 4713 2328 4727
rect 2553 4733 2567 4747
rect 2413 4713 2427 4727
rect 2733 4733 2747 4747
rect 2793 4713 2807 4727
rect 2873 4713 2887 4727
rect 2953 4733 2967 4747
rect 3033 4713 3047 4727
rect 3173 4733 3187 4747
rect 3452 4733 3466 4747
rect 3474 4733 3488 4747
rect 3352 4713 3366 4727
rect 3553 4713 3567 4727
rect 3633 4733 3647 4747
rect 3674 4733 3688 4747
rect 4213 4733 4227 4747
rect 4793 4734 4807 4748
rect 6373 4753 6387 4767
rect 4833 4733 4847 4747
rect 4973 4733 4987 4747
rect 5613 4733 5627 4747
rect 5673 4733 5687 4747
rect 5713 4733 5727 4747
rect 6133 4733 6147 4747
rect 1053 4693 1067 4707
rect 1393 4693 1407 4707
rect 1833 4693 1847 4707
rect 2033 4693 2047 4707
rect 2393 4693 2407 4707
rect 2693 4693 2707 4707
rect 2893 4693 2907 4707
rect 3833 4713 3847 4727
rect 3873 4713 3887 4727
rect 4693 4713 4707 4727
rect 4793 4712 4807 4726
rect 5153 4713 5167 4727
rect 5573 4713 5587 4727
rect 793 4673 807 4687
rect 833 4673 847 4687
rect 1213 4673 1227 4687
rect 1533 4673 1547 4687
rect 1973 4673 1987 4687
rect 2053 4673 2067 4687
rect 2453 4673 2467 4687
rect 3133 4674 3147 4688
rect 3353 4673 3367 4687
rect 3432 4673 3446 4687
rect 3454 4674 3468 4688
rect 3773 4673 3787 4687
rect 3813 4693 3827 4707
rect 4273 4693 4287 4707
rect 4313 4693 4327 4707
rect 4493 4693 4507 4707
rect 4733 4693 4747 4707
rect 4893 4693 4907 4707
rect 4993 4693 5007 4707
rect 5373 4693 5387 4707
rect 5913 4693 5927 4707
rect 5133 4673 5147 4687
rect 5433 4673 5447 4687
rect 6153 4673 6167 4687
rect 673 4653 687 4667
rect 733 4653 747 4667
rect 1253 4653 1267 4667
rect 1592 4653 1606 4667
rect 1614 4653 1628 4667
rect 1953 4653 1967 4667
rect 1993 4653 2007 4667
rect 2252 4653 2266 4667
rect 2274 4653 2288 4667
rect 2353 4653 2367 4667
rect 2873 4653 2887 4667
rect 2972 4653 2986 4667
rect 2994 4653 3008 4667
rect 253 4633 267 4647
rect 433 4633 447 4647
rect 813 4633 827 4647
rect 993 4633 1007 4647
rect 1693 4633 1707 4647
rect 3133 4652 3147 4666
rect 3193 4653 3207 4667
rect 3313 4653 3327 4667
rect 3453 4652 3467 4666
rect 2713 4633 2727 4647
rect 2853 4633 2867 4647
rect 2893 4633 2907 4647
rect 3053 4633 3067 4647
rect 3433 4633 3447 4647
rect 3633 4633 3647 4647
rect 3733 4654 3747 4668
rect 3793 4653 3807 4667
rect 3853 4653 3867 4667
rect 4013 4653 4027 4667
rect 4633 4653 4647 4667
rect 4872 4653 4886 4667
rect 4894 4653 4908 4667
rect 5193 4653 5207 4667
rect 5273 4653 5287 4667
rect 5713 4653 5727 4667
rect 5833 4653 5847 4667
rect 5973 4653 5987 4667
rect 3733 4632 3747 4646
rect 3773 4633 3787 4647
rect 3913 4633 3927 4647
rect 3953 4633 3967 4647
rect 4053 4633 4067 4647
rect 4373 4633 4387 4647
rect 4833 4633 4847 4647
rect 5233 4633 5247 4647
rect 5453 4633 5467 4647
rect 5533 4633 5547 4647
rect 5733 4633 5747 4647
rect 6053 4633 6067 4647
rect 6233 4633 6247 4647
rect 6313 4633 6327 4647
rect 313 4613 327 4627
rect 373 4613 387 4627
rect 573 4613 587 4627
rect 773 4613 787 4627
rect 833 4613 847 4627
rect 933 4613 947 4627
rect 1213 4613 1227 4627
rect 1273 4613 1287 4627
rect 1553 4613 1567 4627
rect 1953 4613 1967 4627
rect 2033 4613 2047 4627
rect 2753 4613 2767 4627
rect 3173 4613 3187 4627
rect 3233 4613 3247 4627
rect 3333 4613 3347 4627
rect 4273 4613 4287 4627
rect 4533 4613 4547 4627
rect 5013 4613 5027 4627
rect 5093 4613 5107 4627
rect 5293 4613 5307 4627
rect 5393 4613 5407 4627
rect 6133 4613 6147 4627
rect 6293 4613 6307 4627
rect 1113 4593 1127 4607
rect 1513 4593 1527 4607
rect 1693 4593 1707 4607
rect 1873 4593 1887 4607
rect 2153 4593 2167 4607
rect 73 4573 87 4587
rect 113 4573 127 4587
rect 393 4573 407 4587
rect 433 4573 447 4587
rect 473 4573 487 4587
rect 533 4573 547 4587
rect 573 4573 587 4587
rect 733 4573 747 4587
rect 773 4573 787 4587
rect 1053 4573 1067 4587
rect 1093 4573 1107 4587
rect 1213 4573 1227 4587
rect 1253 4573 1267 4587
rect 1393 4573 1407 4587
rect 1553 4573 1567 4587
rect 1593 4573 1607 4587
rect 2033 4573 2047 4587
rect 2073 4573 2087 4587
rect 2853 4593 2867 4607
rect 3553 4593 3567 4607
rect 3633 4593 3647 4607
rect 3753 4593 3767 4607
rect 3813 4593 3827 4607
rect 4253 4593 4267 4607
rect 4333 4593 4347 4607
rect 6113 4593 6127 4607
rect 2353 4573 2367 4587
rect 2713 4573 2727 4587
rect 2773 4573 2787 4587
rect 2893 4573 2907 4587
rect 2933 4573 2947 4587
rect 3033 4573 3047 4587
rect 3073 4573 3087 4587
rect 3133 4573 3147 4587
rect 3293 4573 3307 4587
rect 3333 4573 3347 4587
rect 3693 4573 3707 4587
rect 3733 4573 3747 4587
rect 3773 4573 3787 4587
rect 3853 4573 3867 4587
rect 3893 4573 3907 4587
rect 3973 4573 3987 4587
rect 4013 4573 4027 4587
rect 4373 4573 4387 4587
rect 4413 4573 4427 4587
rect 4513 4573 4527 4587
rect 4553 4573 4567 4587
rect 4793 4573 4807 4587
rect 4833 4573 4847 4587
rect 4953 4573 4967 4587
rect 4993 4573 5007 4587
rect 5093 4573 5107 4587
rect 5133 4573 5147 4587
rect 5253 4573 5267 4587
rect 5293 4573 5307 4587
rect 5513 4573 5527 4587
rect 5553 4573 5567 4587
rect 5673 4573 5687 4587
rect 5713 4573 5727 4587
rect 5893 4573 5907 4587
rect 5973 4573 5987 4587
rect 6133 4573 6147 4587
rect 6173 4573 6187 4587
rect 13 4553 27 4567
rect 193 4553 207 4567
rect 313 4553 327 4567
rect 813 4553 827 4567
rect 1353 4553 1367 4567
rect 1433 4553 1447 4567
rect 1773 4553 1787 4567
rect 1853 4553 1867 4567
rect 2173 4553 2187 4567
rect 2253 4553 2267 4567
rect 2533 4553 2547 4567
rect 2593 4553 2607 4567
rect 3193 4553 3207 4567
rect 3253 4553 3267 4567
rect 3493 4553 3507 4567
rect 3553 4553 3567 4567
rect 4193 4553 4207 4567
rect 4253 4553 4267 4567
rect 6293 4553 6307 4567
rect 6353 4553 6367 4567
rect 6413 4553 6427 4567
rect 33 4533 47 4547
rect 1613 4533 1627 4547
rect 2093 4533 2107 4547
rect 4573 4533 4587 4547
rect 233 4513 247 4527
rect 273 4513 287 4527
rect 553 4513 567 4527
rect 633 4513 647 4527
rect 753 4513 767 4527
rect 933 4513 947 4527
rect 1033 4513 1047 4527
rect 1113 4513 1127 4527
rect 1213 4513 1227 4527
rect 1273 4513 1287 4527
rect 1453 4513 1467 4527
rect 1733 4513 1747 4527
rect 1893 4513 1907 4527
rect 1933 4513 1947 4527
rect 1993 4513 2007 4527
rect 2153 4513 2167 4527
rect 2293 4513 2307 4527
rect 2773 4513 2787 4527
rect 3333 4513 3347 4527
rect 3373 4513 3387 4527
rect 3573 4513 3587 4527
rect 3793 4513 3807 4527
rect 3833 4513 3847 4527
rect 4073 4513 4087 4527
rect 4433 4513 4447 4527
rect 4713 4513 4727 4527
rect 4773 4513 4787 4527
rect 5153 4513 5167 4527
rect 5273 4513 5287 4527
rect 5373 4513 5387 4527
rect 5533 4513 5547 4527
rect 5653 4513 5667 4527
rect 5733 4513 5747 4527
rect 5953 4513 5967 4527
rect 6033 4513 6047 4527
rect 6113 4513 6127 4527
rect 6153 4513 6167 4527
rect 6313 4513 6327 4527
rect 13 4473 27 4487
rect 513 4473 527 4487
rect 753 4473 767 4487
rect 893 4473 907 4487
rect 1373 4493 1387 4507
rect 1413 4493 1427 4507
rect 1773 4493 1787 4507
rect 1853 4493 1867 4507
rect 1152 4473 1166 4487
rect 1813 4473 1827 4487
rect 1873 4473 1887 4487
rect 2033 4473 2047 4487
rect 2193 4493 2207 4507
rect 2233 4493 2247 4507
rect 2733 4493 2747 4507
rect 2913 4493 2927 4507
rect 3013 4493 3027 4507
rect 3593 4493 3607 4507
rect 3673 4493 3687 4507
rect 2653 4473 2667 4487
rect 3273 4473 3287 4487
rect 3353 4474 3367 4488
rect 3453 4473 3467 4487
rect 3493 4474 3507 4488
rect 1093 4453 1107 4467
rect 1253 4453 1267 4467
rect 1413 4453 1427 4467
rect 1473 4453 1487 4467
rect 1633 4453 1647 4467
rect 2173 4453 2187 4467
rect 2233 4453 2247 4467
rect 2313 4453 2327 4467
rect 2613 4453 2627 4467
rect 2913 4453 2927 4467
rect 2953 4453 2967 4467
rect 3193 4453 3207 4467
rect 3233 4453 3247 4467
rect 3353 4452 3367 4466
rect 3433 4453 3447 4467
rect 3493 4452 3507 4466
rect 3573 4453 3587 4467
rect 3693 4453 3707 4467
rect 3733 4473 3747 4487
rect 4353 4493 4367 4507
rect 4273 4473 4287 4487
rect 3873 4453 3887 4467
rect 3973 4453 3987 4467
rect 4033 4453 4047 4467
rect 4293 4453 4307 4467
rect 4693 4473 4707 4487
rect 4773 4473 4787 4487
rect 4833 4473 4847 4487
rect 4953 4473 4967 4487
rect 5693 4493 5707 4507
rect 5993 4493 6007 4507
rect 5133 4473 5147 4487
rect 5293 4473 5307 4487
rect 5533 4473 5547 4487
rect 5953 4473 5967 4487
rect 6113 4473 6127 4487
rect 4473 4453 4487 4467
rect 4613 4453 4627 4467
rect 4713 4453 4727 4467
rect 4933 4453 4947 4467
rect 5093 4453 5107 4467
rect 5253 4453 5267 4467
rect 5333 4453 5347 4467
rect 5573 4453 5587 4467
rect 5753 4453 5767 4467
rect 5993 4453 6007 4467
rect 1033 4433 1047 4447
rect 1213 4433 1227 4447
rect 1353 4433 1367 4447
rect 1493 4433 1507 4447
rect 1613 4433 1627 4447
rect 1893 4433 1907 4447
rect 1953 4433 1967 4447
rect 133 4413 147 4427
rect 2273 4413 2287 4427
rect 2333 4413 2347 4427
rect 2433 4413 2447 4427
rect 2533 4433 2547 4447
rect 2733 4434 2747 4448
rect 2853 4433 2867 4447
rect 3113 4433 3127 4447
rect 3253 4433 3267 4447
rect 3333 4433 3347 4447
rect 3393 4433 3407 4447
rect 4653 4433 4667 4447
rect 4833 4433 4847 4447
rect 5013 4433 5027 4447
rect 2733 4412 2747 4426
rect 3153 4413 3167 4427
rect 3293 4413 3307 4427
rect 3413 4413 3427 4427
rect 693 4393 707 4407
rect 773 4393 787 4407
rect 1113 4393 1127 4407
rect 1173 4393 1187 4407
rect 1373 4393 1387 4407
rect 1733 4393 1747 4407
rect 1853 4393 1867 4407
rect 1953 4393 1967 4407
rect 1993 4393 2007 4407
rect 2173 4393 2187 4407
rect 2253 4393 2267 4407
rect 2513 4393 2527 4407
rect 2673 4393 2687 4407
rect 2993 4393 3007 4407
rect 3313 4393 3327 4407
rect 3353 4394 3367 4408
rect 3472 4413 3486 4427
rect 3494 4413 3508 4427
rect 3552 4413 3566 4427
rect 3574 4413 3588 4427
rect 3773 4413 3787 4427
rect 4133 4413 4147 4427
rect 5053 4413 5067 4427
rect 5153 4413 5167 4427
rect 5793 4413 5807 4427
rect 3693 4393 3707 4407
rect 4173 4393 4187 4407
rect 4233 4393 4247 4407
rect 4293 4393 4307 4407
rect 4353 4393 4367 4407
rect 5653 4393 5667 4407
rect 233 4373 247 4387
rect 333 4373 347 4387
rect 733 4373 747 4387
rect 853 4373 867 4387
rect 933 4373 947 4387
rect 1312 4373 1326 4387
rect 1334 4373 1348 4387
rect 1673 4373 1687 4387
rect 1752 4373 1766 4387
rect 1774 4373 1788 4387
rect 1833 4373 1847 4387
rect 2213 4373 2227 4387
rect 3213 4373 3227 4387
rect 3353 4372 3367 4386
rect 3893 4373 3907 4387
rect 4073 4373 4087 4387
rect 4513 4373 4527 4387
rect 4753 4373 4767 4387
rect 4813 4373 4827 4387
rect 5213 4373 5227 4387
rect 5513 4373 5527 4387
rect 5553 4373 5567 4387
rect 5753 4373 5767 4387
rect 5793 4373 5807 4387
rect 1413 4353 1427 4367
rect 1453 4353 1467 4367
rect 1933 4353 1947 4367
rect 1973 4353 1987 4367
rect 2493 4353 2507 4367
rect 2613 4353 2627 4367
rect 2653 4353 2667 4367
rect 3773 4353 3787 4367
rect 3953 4353 3967 4367
rect 4193 4353 4207 4367
rect 4933 4353 4947 4367
rect 6293 4393 6307 4407
rect 6353 4393 6367 4407
rect 6193 4353 6207 4367
rect 6313 4373 6327 4387
rect 6373 4373 6387 4387
rect 6433 4373 6447 4387
rect 133 4333 147 4347
rect 313 4333 327 4347
rect 353 4333 367 4347
rect 393 4333 407 4347
rect 533 4333 547 4347
rect 573 4333 587 4347
rect 733 4333 747 4347
rect 933 4333 947 4347
rect 1213 4333 1227 4347
rect 1293 4333 1307 4347
rect 1513 4333 1527 4347
rect 1653 4333 1667 4347
rect 1833 4333 1847 4347
rect 2113 4333 2127 4347
rect 2273 4333 2287 4347
rect 2313 4333 2327 4347
rect 2733 4333 2747 4347
rect 3112 4333 3126 4347
rect 3134 4333 3148 4347
rect 3413 4333 3427 4347
rect 3453 4333 3467 4347
rect 3673 4333 3687 4347
rect 3733 4333 3747 4347
rect 4233 4333 4247 4347
rect 4353 4333 4367 4347
rect 4453 4333 4467 4347
rect 4573 4333 4587 4347
rect 4653 4333 4667 4347
rect 4813 4333 4827 4347
rect 4973 4333 4987 4347
rect 5113 4333 5127 4347
rect 5213 4333 5227 4347
rect 5292 4333 5306 4347
rect 5493 4333 5507 4347
rect 5553 4333 5567 4347
rect 5633 4333 5647 4347
rect 5733 4333 5747 4347
rect 5773 4333 5787 4347
rect 5893 4333 5907 4347
rect 5932 4333 5946 4347
rect 5973 4333 5987 4347
rect 6013 4333 6027 4347
rect 6313 4333 6327 4347
rect 6393 4333 6407 4347
rect 6473 4333 6487 4347
rect 433 4313 447 4327
rect 473 4313 487 4327
rect 33 4293 47 4307
rect 1393 4293 1407 4307
rect 1473 4293 1487 4307
rect 1673 4293 1687 4307
rect 1913 4293 1927 4307
rect 1993 4293 2007 4307
rect 2433 4293 2447 4307
rect 2493 4293 2507 4307
rect 2593 4293 2607 4307
rect 2673 4293 2687 4307
rect 2853 4293 2867 4307
rect 2913 4293 2927 4307
rect 2933 4293 2947 4307
rect 3573 4293 3587 4307
rect 3633 4293 3647 4307
rect 4073 4293 4087 4307
rect 4153 4293 4167 4307
rect 6073 4293 6087 4307
rect 6353 4293 6367 4307
rect 233 4273 247 4287
rect 273 4273 287 4287
rect 373 4273 387 4287
rect 413 4273 427 4287
rect 513 4273 527 4287
rect 553 4273 567 4287
rect 673 4273 687 4287
rect 713 4273 727 4287
rect 913 4273 927 4287
rect 1053 4273 1067 4287
rect 1093 4273 1107 4287
rect 1133 4273 1147 4287
rect 1233 4273 1247 4287
rect 1273 4273 1287 4287
rect 1433 4273 1447 4287
rect 1593 4273 1607 4287
rect 1633 4273 1647 4287
rect 1773 4273 1787 4287
rect 1813 4273 1827 4287
rect 1953 4273 1967 4287
rect 2133 4273 2147 4287
rect 2293 4273 2307 4287
rect 2633 4273 2647 4287
rect 3053 4273 3067 4287
rect 3093 4273 3107 4287
rect 3193 4273 3207 4287
rect 3233 4273 3247 4287
rect 3353 4273 3367 4287
rect 3393 4273 3407 4287
rect 3753 4273 3767 4287
rect 3793 4273 3807 4287
rect 4333 4273 4347 4287
rect 4373 4273 4387 4287
rect 4473 4273 4487 4287
rect 4513 4273 4527 4287
rect 4653 4273 4667 4287
rect 4693 4273 4707 4287
rect 4993 4273 5007 4287
rect 5233 4273 5247 4287
rect 5273 4273 5287 4287
rect 5473 4273 5487 4287
rect 5533 4273 5547 4287
rect 5573 4273 5587 4287
rect 5713 4273 5727 4287
rect 5753 4273 5767 4287
rect 5913 4273 5927 4287
rect 5993 4273 6007 4287
rect 6033 4273 6047 4287
rect 6293 4273 6307 4287
rect 993 4253 1007 4267
rect 1393 4253 1407 4267
rect 1453 4253 1467 4267
rect 1493 4253 1507 4267
rect 193 4233 207 4247
rect 233 4233 247 4247
rect 373 4233 387 4247
rect 573 4233 587 4247
rect 713 4233 727 4247
rect 933 4233 947 4247
rect 973 4233 987 4247
rect 2093 4253 2107 4267
rect 2493 4253 2507 4267
rect 2573 4253 2587 4267
rect 2713 4253 2727 4267
rect 2913 4253 2927 4267
rect 2993 4253 3007 4267
rect 3413 4253 3427 4267
rect 4073 4253 4087 4267
rect 4113 4253 4127 4267
rect 4413 4253 4427 4267
rect 4453 4253 4467 4267
rect 313 4213 327 4227
rect 553 4213 567 4227
rect 1133 4213 1147 4227
rect 1233 4213 1247 4227
rect 1353 4213 1367 4227
rect 1773 4213 1787 4227
rect 1813 4213 1827 4227
rect 1973 4233 1987 4247
rect 2133 4233 2147 4247
rect 2633 4233 2647 4247
rect 3233 4233 3247 4247
rect 3373 4233 3387 4247
rect 3653 4233 3667 4247
rect 3893 4233 3907 4247
rect 1913 4213 1927 4227
rect 2073 4213 2087 4227
rect 2153 4213 2167 4227
rect 1253 4193 1267 4207
rect 1313 4193 1327 4207
rect 2173 4193 2187 4207
rect 2293 4193 2307 4207
rect 2593 4213 2607 4227
rect 2793 4213 2807 4227
rect 2533 4193 2547 4207
rect 2833 4193 2847 4207
rect 2953 4214 2967 4228
rect 3053 4214 3067 4228
rect 3193 4213 3207 4227
rect 3253 4213 3267 4227
rect 3413 4213 3427 4227
rect 4373 4233 4387 4247
rect 4433 4233 4447 4247
rect 4513 4233 4527 4247
rect 4653 4233 4667 4247
rect 4713 4233 4727 4247
rect 4773 4233 4787 4247
rect 4813 4233 4827 4247
rect 5173 4253 5187 4267
rect 5213 4253 5227 4267
rect 5233 4233 5247 4247
rect 5273 4233 5287 4247
rect 5873 4253 5887 4267
rect 6313 4233 6327 4247
rect 4353 4213 4367 4227
rect 4413 4213 4427 4227
rect 4973 4213 4987 4227
rect 5113 4213 5127 4227
rect 5553 4213 5567 4227
rect 5753 4213 5767 4227
rect 5873 4213 5887 4227
rect 6173 4213 6187 4227
rect 6353 4213 6367 4227
rect 273 4173 287 4187
rect 393 4173 407 4187
rect 1813 4173 1827 4187
rect 1873 4179 1887 4193
rect 2953 4192 2967 4206
rect 3053 4192 3067 4206
rect 3292 4193 3306 4207
rect 3314 4193 3328 4207
rect 3432 4193 3446 4207
rect 3454 4193 3468 4207
rect 3573 4193 3587 4207
rect 3714 4193 3728 4207
rect 2113 4173 2127 4187
rect 3153 4173 3167 4187
rect 3193 4173 3207 4187
rect 3233 4173 3247 4187
rect 3493 4173 3507 4187
rect 3753 4173 3767 4187
rect 4153 4173 4167 4187
rect 4193 4193 4207 4207
rect 4553 4193 4567 4207
rect 4913 4193 4927 4207
rect 5013 4193 5027 4207
rect 5313 4193 5326 4207
rect 5326 4193 5327 4207
rect 4273 4173 4287 4187
rect 4633 4173 4647 4187
rect 4693 4173 4707 4187
rect 5053 4173 5067 4187
rect 5454 4193 5468 4207
rect 5494 4193 5508 4207
rect 5533 4193 5547 4207
rect 5573 4193 5587 4207
rect 5693 4193 5707 4207
rect 5733 4193 5747 4207
rect 5913 4193 5927 4207
rect 5373 4173 5387 4187
rect 5553 4173 5567 4187
rect 853 4153 867 4167
rect 1313 4153 1327 4167
rect 1453 4153 1467 4167
rect 1913 4153 1927 4167
rect 2053 4153 2067 4167
rect 533 4133 547 4147
rect 1173 4133 1187 4147
rect 1293 4133 1307 4147
rect 1433 4133 1447 4147
rect 1473 4133 1487 4147
rect 1633 4133 1647 4147
rect 1953 4133 1967 4147
rect 1993 4133 2007 4147
rect 2113 4133 2127 4147
rect 2153 4133 2167 4147
rect 2253 4153 2267 4167
rect 2452 4153 2466 4167
rect 2474 4153 2488 4167
rect 2933 4153 2947 4167
rect 3033 4153 3047 4167
rect 3112 4153 3126 4167
rect 3134 4153 3148 4167
rect 3313 4153 3327 4167
rect 3373 4153 3387 4167
rect 2533 4133 2547 4147
rect 2613 4133 2627 4147
rect 2652 4133 2666 4147
rect 2674 4133 2688 4147
rect 2792 4133 2806 4147
rect 2814 4133 2828 4147
rect 2973 4133 2987 4147
rect 3053 4133 3067 4147
rect 3093 4133 3107 4147
rect 3193 4133 3207 4147
rect 3273 4133 3287 4147
rect 4053 4153 4067 4167
rect 4113 4153 4127 4167
rect 4373 4153 4387 4167
rect 4413 4153 4427 4167
rect 4873 4153 4887 4167
rect 5013 4153 5027 4167
rect 6193 4153 6207 4167
rect 3673 4133 3687 4147
rect 933 4113 947 4127
rect 1653 4113 1667 4127
rect 1693 4113 1707 4127
rect 1773 4113 1787 4127
rect 1933 4113 1947 4127
rect 1973 4113 1987 4127
rect 2073 4113 2087 4127
rect 353 4093 367 4107
rect 453 4093 467 4107
rect 553 4093 567 4107
rect 813 4093 827 4107
rect 1393 4093 1407 4107
rect 1533 4093 1547 4107
rect 1853 4093 1867 4107
rect 1913 4093 1927 4107
rect 2013 4093 2027 4107
rect 2173 4093 2187 4107
rect 2513 4093 2527 4107
rect 2873 4113 2887 4127
rect 3132 4114 3146 4128
rect 3013 4093 3027 4107
rect 3052 4093 3066 4107
rect 3074 4093 3088 4107
rect 913 4073 927 4087
rect 1033 4073 1047 4087
rect 1093 4073 1107 4087
rect 2333 4073 2347 4087
rect 2993 4073 3007 4087
rect 3133 4092 3147 4106
rect 3293 4093 3307 4107
rect 3333 4113 3347 4127
rect 3493 4113 3507 4127
rect 4593 4133 4607 4147
rect 4793 4133 4807 4147
rect 5173 4133 5187 4147
rect 5833 4133 5847 4147
rect 6113 4133 6127 4147
rect 4173 4113 4187 4127
rect 4753 4113 4767 4127
rect 4913 4113 4927 4127
rect 5053 4113 5067 4127
rect 5453 4113 5467 4127
rect 5493 4113 5507 4127
rect 5633 4113 5647 4127
rect 5853 4113 5867 4127
rect 6153 4114 6167 4128
rect 4233 4093 4247 4107
rect 4793 4093 4807 4107
rect 4873 4093 4887 4107
rect 4973 4093 4987 4107
rect 5133 4093 5147 4107
rect 5193 4093 5207 4107
rect 5253 4093 5267 4107
rect 5953 4093 5967 4107
rect 6153 4092 6167 4106
rect 3413 4073 3427 4087
rect 3453 4073 3467 4087
rect 153 4053 167 4067
rect 193 4053 207 4067
rect 233 4053 247 4067
rect 273 4053 287 4067
rect 313 4053 327 4067
rect 353 4053 367 4067
rect 393 4053 407 4067
rect 513 4053 527 4067
rect 553 4053 567 4067
rect 733 4053 747 4067
rect 793 4053 807 4067
rect 813 4053 827 4067
rect 853 4053 867 4067
rect 1293 4053 1307 4067
rect 1353 4053 1367 4067
rect 1393 4053 1407 4067
rect 1433 4053 1447 4067
rect 1493 4053 1507 4067
rect 1533 4053 1547 4067
rect 1653 4053 1667 4067
rect 1693 4053 1707 4067
rect 1973 4053 1987 4067
rect 2013 4053 2027 4067
rect 2353 4053 2367 4067
rect 2433 4053 2447 4067
rect 2513 4053 2527 4067
rect 2553 4053 2567 4067
rect 2593 4053 2607 4067
rect 2713 4053 2727 4067
rect 2753 4053 2767 4067
rect 2873 4053 2887 4067
rect 2913 4053 2927 4067
rect 3053 4053 3067 4067
rect 3093 4053 3107 4067
rect 3213 4053 3227 4067
rect 3333 4053 3347 4067
rect 3373 4053 3387 4067
rect 3493 4053 3507 4067
rect 3533 4053 3547 4067
rect 3773 4073 3787 4087
rect 4213 4073 4227 4087
rect 4313 4073 4327 4087
rect 4633 4073 4647 4087
rect 4893 4073 4907 4087
rect 5373 4073 5387 4087
rect 3673 4053 3687 4067
rect 3713 4053 3727 4067
rect 3793 4053 3807 4067
rect 3833 4053 3847 4067
rect 3953 4053 3967 4067
rect 3993 4053 4007 4067
rect 4113 4053 4127 4067
rect 4153 4053 4167 4067
rect 4613 4053 4627 4067
rect 4873 4053 4887 4067
rect 5053 4053 5067 4067
rect 5093 4053 5107 4067
rect 5133 4053 5147 4067
rect 5233 4053 5247 4067
rect 5493 4053 5507 4067
rect 5533 4053 5547 4067
rect 5633 4053 5647 4067
rect 5673 4053 5687 4067
rect 5793 4053 5807 4067
rect 5833 4053 5847 4067
rect 5873 4053 5887 4067
rect 5913 4053 5927 4067
rect 5953 4053 5967 4067
rect 5993 4053 6007 4067
rect 6113 4053 6127 4067
rect 6153 4053 6167 4067
rect 6293 4053 6307 4067
rect 6333 4053 6347 4067
rect 993 4033 1007 4047
rect 1873 4033 1887 4047
rect 2073 4033 2087 4047
rect 2173 4033 2187 4047
rect 2233 4033 2247 4047
rect 4293 4033 4307 4047
rect 4433 4033 4447 4047
rect 4713 4033 4727 4047
rect 4753 4033 4767 4047
rect 4793 4033 4807 4047
rect 2853 4013 2867 4027
rect 113 3993 127 4007
rect 213 3993 227 4007
rect 313 3993 327 4007
rect 413 3993 427 4007
rect 693 3993 707 4007
rect 833 3993 847 4007
rect 1173 3993 1187 4007
rect 1333 3993 1347 4007
rect 1413 3993 1427 4007
rect 1594 3993 1608 4007
rect 1833 3993 1847 4007
rect 2133 3993 2147 4007
rect 2213 3993 2227 4007
rect 2313 3993 2327 4007
rect 2474 3993 2488 4007
rect 2533 3993 2547 4007
rect 2573 3993 2587 4007
rect 4093 4013 4107 4027
rect 2893 3993 2907 4007
rect 2933 3993 2947 4007
rect 3113 3993 3127 4007
rect 3193 3993 3207 4007
rect 3233 3993 3247 4007
rect 3293 3993 3307 4007
rect 193 3953 207 3967
rect 933 3973 947 3987
rect 973 3973 987 3987
rect 1093 3973 1107 3987
rect 1133 3973 1147 3987
rect 2613 3973 2627 3987
rect 2773 3973 2787 3987
rect 2853 3973 2867 3987
rect 3073 3973 3087 3987
rect 3413 3993 3427 4007
rect 3553 3993 3567 4007
rect 3613 3993 3627 4007
rect 3673 3993 3687 4007
rect 3773 3993 3787 4007
rect 3813 3993 3827 4007
rect 4133 3993 4147 4007
rect 4173 3993 4187 4007
rect 4273 3993 4287 4007
rect 4413 3993 4427 4007
rect 4613 3993 4627 4007
rect 5053 3993 5067 4007
rect 5153 3993 5167 4007
rect 5273 3993 5287 4007
rect 5353 3993 5367 4007
rect 5473 3993 5487 4007
rect 5613 3993 5627 4007
rect 5653 3993 5667 4007
rect 5773 3993 5787 4007
rect 5853 3993 5867 4007
rect 6053 3993 6067 4007
rect 6273 3993 6287 4007
rect 6433 3993 6447 4007
rect 3473 3973 3487 3987
rect 4013 3973 4027 3987
rect 4093 3973 4107 3987
rect 4733 3973 4747 3987
rect 693 3953 707 3967
rect 833 3953 847 3967
rect 893 3953 907 3967
rect 1193 3953 1207 3967
rect 1473 3953 1487 3967
rect 1693 3953 1707 3967
rect 1733 3953 1747 3967
rect 2333 3953 2347 3967
rect 2493 3953 2507 3967
rect 3313 3953 3327 3967
rect 3453 3953 3467 3967
rect 3513 3953 3527 3967
rect 3573 3953 3587 3967
rect 3733 3953 3747 3967
rect 3913 3953 3927 3967
rect 3953 3954 3967 3968
rect 3993 3953 4007 3967
rect 4413 3953 4427 3967
rect 113 3933 127 3947
rect 153 3933 167 3947
rect 1093 3933 1107 3947
rect 1252 3933 1266 3947
rect 2353 3933 2367 3947
rect 2753 3934 2767 3948
rect 2913 3933 2927 3947
rect 3333 3933 3347 3947
rect 3653 3933 3667 3947
rect 3853 3933 3867 3947
rect 3953 3932 3967 3946
rect 4033 3933 4047 3947
rect 4072 3933 4086 3947
rect 4094 3933 4108 3947
rect 4153 3933 4167 3947
rect 4293 3933 4307 3947
rect 4433 3933 4447 3947
rect 4694 3933 4708 3947
rect 5553 3973 5567 3987
rect 5073 3953 5087 3967
rect 5353 3953 5367 3967
rect 5573 3953 5587 3967
rect 5613 3953 5627 3967
rect 4793 3934 4807 3948
rect 5093 3933 5107 3947
rect 5153 3933 5167 3947
rect 5273 3933 5287 3947
rect 5413 3933 5427 3947
rect 5553 3933 5567 3947
rect 5653 3933 5667 3947
rect 5713 3953 5727 3967
rect 5853 3953 5867 3967
rect 6013 3973 6027 3987
rect 6133 3953 6147 3967
rect 6213 3953 6227 3967
rect 6373 3953 6387 3967
rect 6453 3953 6467 3967
rect 5752 3933 5766 3947
rect 5793 3933 5807 3947
rect 5933 3933 5947 3947
rect 513 3913 527 3927
rect 613 3913 627 3927
rect 1113 3913 1127 3927
rect 233 3893 247 3907
rect 453 3893 467 3907
rect 913 3893 927 3907
rect 953 3893 967 3907
rect 993 3893 1007 3907
rect 1033 3893 1047 3907
rect 2292 3913 2306 3927
rect 2314 3913 2328 3927
rect 2453 3913 2467 3927
rect 2493 3913 2507 3927
rect 2612 3913 2626 3927
rect 2634 3913 2648 3927
rect 2713 3913 2727 3927
rect 2753 3912 2767 3926
rect 2993 3913 3007 3927
rect 3313 3913 3327 3927
rect 1293 3893 1307 3907
rect 2372 3893 2386 3907
rect 2394 3893 2408 3907
rect 2553 3893 2567 3907
rect 2593 3893 2607 3907
rect 2653 3893 2667 3907
rect 793 3873 807 3887
rect 873 3873 887 3887
rect 1393 3873 1407 3887
rect 1833 3873 1847 3887
rect 2053 3873 2067 3887
rect 2293 3873 2307 3887
rect 2334 3873 2348 3887
rect 2633 3873 2647 3887
rect 2733 3893 2747 3907
rect 2812 3893 2826 3907
rect 2834 3893 2848 3907
rect 2893 3893 2907 3907
rect 3213 3893 3227 3907
rect 3333 3893 3347 3907
rect 3373 3893 3387 3907
rect 3433 3913 3447 3927
rect 3553 3913 3567 3927
rect 3913 3913 3927 3927
rect 3973 3913 3987 3927
rect 4473 3913 4487 3927
rect 4753 3913 4767 3927
rect 4793 3912 4807 3926
rect 5013 3913 5027 3927
rect 5053 3913 5067 3927
rect 5253 3913 5267 3927
rect 5313 3914 5327 3928
rect 5393 3913 5407 3927
rect 3793 3893 3807 3907
rect 2753 3873 2767 3887
rect 3253 3873 3267 3887
rect 3293 3873 3307 3887
rect 4233 3893 4247 3907
rect 4593 3893 4607 3907
rect 4973 3893 4987 3907
rect 5233 3893 5247 3907
rect 5313 3892 5327 3906
rect 5613 3893 5627 3907
rect 5753 3893 5767 3907
rect 6113 3893 6127 3907
rect 4513 3873 4527 3887
rect 4653 3873 4667 3887
rect 4693 3873 4707 3887
rect 4833 3873 4847 3887
rect 4892 3873 4906 3887
rect 4953 3873 4967 3887
rect 5033 3873 5047 3887
rect 5253 3873 5267 3887
rect 5633 3872 5647 3886
rect 5813 3873 5827 3887
rect 6053 3873 6067 3887
rect 6393 3873 6407 3887
rect 553 3853 567 3867
rect 1933 3853 1947 3867
rect 673 3833 687 3847
rect 733 3833 747 3847
rect 773 3833 787 3847
rect 913 3833 927 3847
rect 1053 3833 1067 3847
rect 1093 3833 1107 3847
rect 2473 3853 2487 3867
rect 2513 3853 2527 3867
rect 3192 3853 3206 3867
rect 3214 3853 3228 3867
rect 3333 3853 3347 3867
rect 4673 3853 4687 3867
rect 4793 3853 4807 3867
rect 5193 3853 5207 3867
rect 5273 3853 5287 3867
rect 5473 3853 5487 3867
rect 5652 3853 5666 3867
rect 6013 3853 6027 3867
rect 3073 3833 3087 3847
rect 3133 3833 3147 3847
rect 4953 3833 4967 3847
rect 4993 3833 5007 3847
rect 6252 3853 6266 3867
rect 6274 3853 6288 3867
rect 6313 3853 6327 3867
rect 53 3813 67 3827
rect 153 3813 167 3827
rect 373 3813 387 3827
rect 514 3813 528 3827
rect 613 3813 627 3827
rect 873 3813 887 3827
rect 953 3813 967 3827
rect 1133 3813 1147 3827
rect 1253 3813 1267 3827
rect 1493 3813 1507 3827
rect 1553 3813 1567 3827
rect 1813 3813 1827 3827
rect 2013 3813 2027 3827
rect 2213 3813 2227 3827
rect 2373 3813 2387 3827
rect 2413 3813 2427 3827
rect 2653 3813 2667 3827
rect 2893 3813 2907 3827
rect 3213 3813 3227 3827
rect 3253 3813 3267 3827
rect 3293 3813 3307 3827
rect 3613 3813 3627 3827
rect 3673 3813 3687 3827
rect 3913 3813 3927 3827
rect 4473 3813 4487 3827
rect 4513 3813 4527 3827
rect 4673 3813 4687 3827
rect 4793 3813 4807 3827
rect 5073 3813 5087 3827
rect 5193 3813 5207 3827
rect 653 3793 667 3807
rect 4553 3793 4567 3807
rect 5173 3793 5187 3807
rect 5313 3813 5327 3827
rect 5413 3813 5427 3827
rect 5613 3813 5627 3827
rect 5773 3813 5787 3827
rect 5853 3813 5867 3827
rect 5933 3813 5947 3827
rect 5993 3813 6007 3827
rect 6093 3813 6107 3827
rect 6253 3814 6267 3828
rect 6293 3813 6307 3827
rect 6313 3814 6327 3828
rect 5693 3793 5707 3807
rect 853 3773 867 3787
rect 1113 3773 1127 3787
rect 1733 3773 1747 3787
rect 1813 3773 1827 3787
rect 1973 3773 1987 3787
rect 2473 3773 2487 3787
rect 2513 3773 2527 3787
rect 2773 3773 2787 3787
rect 2833 3773 2847 3787
rect 3073 3773 3087 3787
rect 3433 3773 3447 3787
rect 3493 3773 3507 3787
rect 3793 3773 3807 3787
rect 3853 3773 3867 3787
rect 4033 3773 4047 3787
rect 4093 3773 4107 3787
rect 4293 3773 4307 3787
rect 4353 3773 4367 3787
rect 4933 3773 4947 3787
rect 6373 3773 6387 3787
rect 6433 3773 6447 3787
rect 93 3753 107 3767
rect 133 3753 147 3767
rect 233 3753 247 3767
rect 273 3753 287 3767
rect 393 3753 407 3767
rect 433 3753 447 3767
rect 593 3753 607 3767
rect 633 3753 647 3767
rect 893 3753 907 3767
rect 933 3753 947 3767
rect 1173 3753 1187 3767
rect 1193 3753 1207 3767
rect 1233 3753 1247 3767
rect 1273 3753 1287 3767
rect 1353 3753 1367 3767
rect 1393 3753 1407 3767
rect 1533 3753 1547 3767
rect 1853 3753 1867 3767
rect 2193 3753 2207 3767
rect 2233 3753 2247 3767
rect 2273 3753 2287 3767
rect 2393 3753 2407 3767
rect 2433 3753 2447 3767
rect 2533 3753 2547 3767
rect 2553 3753 2567 3767
rect 2593 3753 2607 3767
rect 3013 3753 3027 3767
rect 3193 3753 3207 3767
rect 3233 3753 3247 3767
rect 3333 3753 3347 3767
rect 3373 3753 3387 3767
rect 733 3733 747 3747
rect 773 3733 787 3747
rect 973 3733 987 3747
rect 1053 3733 1067 3747
rect 2633 3733 2647 3747
rect 3073 3733 3087 3747
rect 4093 3733 4107 3747
rect 4493 3753 4507 3767
rect 4533 3753 4547 3767
rect 4653 3753 4667 3767
rect 4693 3753 4707 3767
rect 5093 3753 5107 3767
rect 5133 3753 5147 3767
rect 5253 3753 5267 3767
rect 5293 3753 5307 3767
rect 5333 3753 5347 3767
rect 5433 3753 5447 3767
rect 5473 3753 5487 3767
rect 5593 3753 5607 3767
rect 5633 3753 5647 3767
rect 5673 3753 5687 3767
rect 5753 3753 5767 3767
rect 5793 3753 5807 3767
rect 5913 3753 5927 3767
rect 5953 3753 5967 3767
rect 6073 3753 6087 3767
rect 6113 3753 6127 3767
rect 6293 3753 6307 3767
rect 6393 3733 6407 3747
rect 133 3713 147 3727
rect 313 3713 327 3727
rect 453 3713 467 3727
rect 593 3713 607 3727
rect 853 3713 867 3727
rect 893 3713 907 3727
rect 933 3713 947 3727
rect 1093 3713 1107 3727
rect 1133 3713 1147 3727
rect 1193 3713 1207 3727
rect 1233 3713 1247 3727
rect 1453 3713 1467 3727
rect 1733 3713 1747 3727
rect 1913 3713 1927 3727
rect 1973 3713 1987 3727
rect 2133 3713 2147 3727
rect 2233 3713 2247 3727
rect 2393 3713 2407 3727
rect 2433 3713 2447 3727
rect 3193 3713 3207 3727
rect 3293 3713 3307 3727
rect 4433 3713 4447 3727
rect 4493 3713 4507 3727
rect 4553 3713 4567 3727
rect 4614 3713 4628 3727
rect 4693 3713 4707 3727
rect 4753 3713 4767 3727
rect 4833 3713 4847 3727
rect 4933 3713 4947 3727
rect 5133 3713 5147 3727
rect 5293 3713 5307 3727
rect 5433 3713 5447 3727
rect 5733 3713 5747 3727
rect 5913 3713 5927 3727
rect 53 3693 67 3707
rect 233 3693 247 3707
rect 1493 3693 1507 3707
rect 2273 3693 2287 3707
rect 2313 3693 2327 3707
rect 3233 3693 3247 3707
rect 3373 3693 3387 3707
rect 4793 3693 4807 3707
rect 5333 3693 5347 3707
rect 5473 3693 5487 3707
rect 5753 3693 5767 3707
rect 5953 3693 5967 3707
rect 6013 3693 6027 3707
rect 273 3673 287 3687
rect 393 3673 407 3687
rect 1053 3673 1067 3687
rect 1153 3673 1167 3687
rect 2253 3673 2267 3687
rect 2413 3673 2427 3687
rect 2553 3673 2567 3687
rect 2733 3673 2747 3687
rect 2833 3673 2847 3687
rect 3113 3673 3127 3687
rect 3433 3673 3447 3687
rect 3853 3673 3867 3687
rect 4093 3673 4107 3687
rect 4153 3673 4167 3687
rect 4594 3673 4608 3687
rect 93 3653 107 3667
rect 553 3653 567 3667
rect 1473 3653 1487 3667
rect 1513 3653 1527 3667
rect 1853 3653 1867 3667
rect 253 3633 267 3647
rect 473 3633 487 3647
rect 773 3633 787 3647
rect 933 3633 947 3647
rect 2273 3633 2287 3647
rect 2533 3653 2547 3667
rect 2853 3653 2867 3667
rect 3153 3653 3167 3667
rect 3573 3653 3587 3667
rect 3673 3653 3687 3667
rect 3913 3653 3927 3667
rect 3993 3653 4007 3667
rect 2353 3633 2367 3647
rect 2473 3633 2487 3647
rect 733 3613 747 3627
rect 1253 3613 1267 3627
rect 2713 3633 2727 3647
rect 2893 3633 2907 3647
rect 3033 3633 3047 3647
rect 2513 3613 2527 3627
rect 3613 3633 3627 3647
rect 3933 3633 3947 3647
rect 4013 3633 4027 3647
rect 4653 3653 4667 3667
rect 5273 3673 5287 3687
rect 5553 3673 5567 3687
rect 5653 3673 5667 3687
rect 5813 3673 5827 3687
rect 5893 3673 5907 3687
rect 6473 3673 6487 3687
rect 5833 3653 5847 3667
rect 6073 3653 6087 3667
rect 6453 3653 6467 3667
rect 6493 3653 6507 3667
rect 4113 3633 4127 3647
rect 4693 3633 4707 3647
rect 4893 3633 4907 3647
rect 4933 3633 4947 3647
rect 5093 3633 5107 3647
rect 3133 3613 3147 3627
rect 3653 3613 3667 3627
rect 4353 3613 4367 3627
rect 4493 3613 4507 3627
rect 4613 3613 4627 3627
rect 4653 3613 4667 3627
rect 4993 3613 5007 3627
rect 5753 3613 5767 3627
rect 5933 3613 5947 3627
rect 6013 3613 6027 3627
rect 6213 3613 6227 3627
rect 6273 3613 6287 3627
rect 73 3573 87 3587
rect 193 3573 207 3587
rect 313 3573 327 3587
rect 413 3573 427 3587
rect 513 3573 527 3587
rect 593 3573 607 3587
rect 1373 3593 1387 3607
rect 1413 3593 1427 3607
rect 1533 3593 1547 3607
rect 1653 3593 1667 3607
rect 1813 3593 1827 3607
rect 3413 3593 3427 3607
rect 3513 3593 3527 3607
rect 4053 3593 4067 3607
rect 4253 3593 4267 3607
rect 893 3573 907 3587
rect 973 3573 987 3587
rect 1253 3573 1267 3587
rect 1553 3573 1567 3587
rect 1833 3573 1847 3587
rect 2333 3573 2347 3587
rect 2393 3573 2407 3587
rect 2493 3573 2507 3587
rect 2753 3573 2767 3587
rect 2853 3573 2867 3587
rect 3173 3573 3187 3587
rect 3253 3573 3267 3587
rect 3453 3573 3467 3587
rect 3553 3573 3567 3587
rect 3593 3573 3607 3587
rect 4033 3573 4047 3587
rect 4433 3573 4447 3587
rect 4573 3593 4587 3607
rect 5712 3593 5726 3607
rect 5893 3593 5907 3607
rect 5033 3573 5047 3587
rect 5333 3573 5347 3587
rect 5493 3573 5507 3587
rect 5833 3573 5847 3587
rect 5993 3573 6007 3587
rect 6073 3573 6087 3587
rect 6212 3573 6226 3587
rect 6234 3573 6248 3587
rect 6513 3573 6527 3587
rect 2813 3553 2827 3567
rect 73 3533 87 3547
rect 273 3533 287 3547
rect 313 3533 327 3547
rect 393 3533 407 3547
rect 593 3533 607 3547
rect 633 3533 647 3547
rect 733 3533 747 3547
rect 773 3533 787 3547
rect 893 3533 907 3547
rect 933 3533 947 3547
rect 1213 3533 1227 3547
rect 1253 3533 1267 3547
rect 1373 3533 1387 3547
rect 1413 3533 1427 3547
rect 1533 3533 1547 3547
rect 1573 3533 1587 3547
rect 1653 3533 1667 3547
rect 1833 3533 1847 3547
rect 1873 3533 1887 3547
rect 1913 3533 1927 3547
rect 1953 3533 1967 3547
rect 1993 3533 2007 3547
rect 2033 3533 2047 3547
rect 2193 3533 2207 3547
rect 2373 3533 2387 3547
rect 2413 3533 2427 3547
rect 2453 3533 2467 3547
rect 2493 3533 2507 3547
rect 2553 3533 2567 3547
rect 2593 3533 2607 3547
rect 3033 3553 3047 3567
rect 3093 3553 3107 3567
rect 4733 3553 4747 3567
rect 4833 3553 4847 3567
rect 4893 3553 4907 3567
rect 5553 3553 5567 3567
rect 3293 3533 3307 3547
rect 3473 3533 3487 3547
rect 3513 3533 3527 3547
rect 3613 3533 3627 3547
rect 3653 3533 3667 3547
rect 3993 3533 4007 3547
rect 4033 3533 4047 3547
rect 4393 3533 4407 3547
rect 4433 3533 4447 3547
rect 4573 3533 4587 3547
rect 4613 3533 4627 3547
rect 4693 3533 4707 3547
rect 4993 3533 5007 3547
rect 5093 3534 5107 3548
rect 5333 3533 5347 3547
rect 5373 3533 5387 3547
rect 5493 3533 5507 3547
rect 5533 3533 5547 3547
rect 5653 3533 5667 3547
rect 5693 3533 5707 3547
rect 5853 3533 5867 3547
rect 5893 3533 5907 3547
rect 5993 3533 6007 3547
rect 6033 3533 6047 3547
rect 6173 3533 6187 3547
rect 6213 3533 6227 3547
rect 6313 3533 6327 3547
rect 233 3513 247 3527
rect 433 3513 447 3527
rect 1173 3513 1187 3527
rect 1793 3513 1807 3527
rect 2733 3513 2747 3527
rect 2773 3513 2787 3527
rect 2813 3513 2827 3527
rect 3093 3513 3107 3527
rect 3153 3513 3167 3527
rect 3813 3513 3827 3527
rect 3893 3513 3907 3527
rect 4073 3513 4087 3527
rect 4293 3513 4307 3527
rect 4953 3513 4967 3527
rect 5093 3512 5107 3526
rect 5573 3513 5587 3527
rect 5613 3513 5627 3527
rect 953 3493 967 3507
rect 2473 3493 2487 3507
rect 2533 3493 2547 3507
rect 4893 3493 4907 3507
rect 4973 3493 4987 3507
rect 5713 3494 5727 3508
rect 5753 3493 5767 3507
rect 93 3473 107 3487
rect 373 3473 387 3487
rect 413 3473 427 3487
rect 553 3473 567 3487
rect 713 3473 727 3487
rect 793 3473 807 3487
rect 1273 3473 1287 3487
rect 1373 3473 1387 3487
rect 1433 3473 1447 3487
rect 1673 3473 1687 3487
rect 1873 3473 1887 3487
rect 1973 3473 1987 3487
rect 2153 3473 2167 3487
rect 2293 3473 2307 3487
rect 2453 3473 2467 3487
rect 2573 3473 2587 3487
rect 2713 3473 2727 3487
rect 2853 3473 2867 3487
rect 2933 3473 2947 3487
rect 2973 3473 2987 3487
rect 3173 3473 3187 3487
rect 3233 3473 3247 3487
rect 3273 3473 3287 3487
rect 3493 3473 3507 3487
rect 3533 3473 3547 3487
rect 3673 3473 3687 3487
rect 3713 3473 3727 3487
rect 3953 3473 3967 3487
rect 4533 3473 4547 3487
rect 4613 3473 4627 3487
rect 4793 3473 4807 3487
rect 4913 3473 4927 3487
rect 5153 3473 5167 3487
rect 5273 3473 5287 3487
rect 5313 3473 5327 3487
rect 5473 3473 5487 3487
rect 5553 3473 5567 3487
rect 5633 3473 5647 3487
rect 633 3433 647 3447
rect 1033 3453 1047 3467
rect 1073 3453 1087 3467
rect 813 3433 827 3447
rect 873 3433 887 3447
rect 2533 3453 2547 3467
rect 2753 3453 2767 3467
rect 2793 3453 2807 3467
rect 913 3413 927 3427
rect 1413 3433 1427 3447
rect 1573 3433 1587 3447
rect 1673 3434 1687 3448
rect 1813 3433 1827 3447
rect 2233 3433 2247 3447
rect 2573 3433 2587 3447
rect 2893 3433 2907 3447
rect 2953 3433 2967 3447
rect 3033 3433 3047 3447
rect 3093 3433 3107 3447
rect 3273 3433 3287 3447
rect 5713 3472 5727 3486
rect 5813 3473 5827 3487
rect 5873 3473 5887 3487
rect 6013 3473 6027 3487
rect 6093 3473 6107 3487
rect 6153 3473 6167 3487
rect 6193 3473 6207 3487
rect 6293 3473 6307 3487
rect 6333 3473 6347 3487
rect 4833 3453 4847 3467
rect 4873 3453 4887 3467
rect 5513 3453 5527 3467
rect 3333 3433 3347 3447
rect 3593 3433 3607 3447
rect 4033 3433 4047 3447
rect 4393 3433 4407 3447
rect 4513 3433 4527 3447
rect 4633 3433 4647 3447
rect 4673 3433 4687 3447
rect 5153 3433 5167 3447
rect 5313 3433 5327 3447
rect 5553 3433 5567 3447
rect 5873 3433 5887 3447
rect 6013 3433 6027 3447
rect 6113 3433 6127 3447
rect 6193 3433 6207 3447
rect 1093 3413 1107 3427
rect 1673 3412 1687 3426
rect 2033 3414 2047 3428
rect 2373 3413 2387 3427
rect 2633 3413 2647 3427
rect 593 3393 607 3407
rect 1313 3393 1327 3407
rect 1913 3393 1927 3407
rect 2033 3392 2047 3406
rect 2273 3393 2287 3407
rect 2513 3393 2527 3407
rect 2553 3393 2567 3407
rect 2673 3393 2687 3407
rect 2773 3413 2787 3427
rect 2793 3393 2807 3407
rect 2992 3393 3006 3407
rect 3014 3393 3028 3407
rect 3453 3413 3467 3427
rect 3493 3413 3507 3427
rect 3933 3413 3947 3427
rect 4173 3413 4187 3427
rect 4293 3413 4307 3427
rect 4453 3413 4467 3427
rect 4613 3413 4627 3427
rect 4873 3413 4887 3427
rect 5033 3413 5047 3427
rect 5173 3413 5187 3427
rect 5513 3413 5527 3427
rect 5673 3413 5687 3427
rect 6213 3413 6227 3427
rect 6272 3413 6286 3427
rect 6333 3413 6347 3427
rect 3293 3393 3307 3407
rect 3393 3393 3407 3407
rect 4633 3393 4647 3407
rect 4813 3393 4827 3407
rect 4993 3393 5007 3407
rect 5053 3393 5067 3407
rect 5613 3393 5627 3407
rect 5893 3394 5907 3408
rect 5993 3393 6007 3407
rect 713 3373 727 3387
rect 773 3373 787 3387
rect 1033 3373 1047 3387
rect 1093 3373 1107 3387
rect 1253 3373 1267 3387
rect 1333 3373 1347 3387
rect 1813 3373 1827 3387
rect 1873 3373 1887 3387
rect 2013 3373 2027 3387
rect 2153 3373 2167 3387
rect 2194 3373 2208 3387
rect 2333 3373 2347 3387
rect 2713 3374 2727 3388
rect 3313 3373 3327 3387
rect 3833 3373 3847 3387
rect 453 3353 467 3367
rect 733 3353 747 3367
rect 1153 3353 1167 3367
rect 1273 3353 1287 3367
rect 1373 3353 1387 3367
rect 1973 3353 1987 3367
rect 2113 3353 2127 3367
rect 2453 3353 2467 3367
rect 2572 3353 2586 3367
rect 2594 3353 2608 3367
rect 2713 3352 2727 3366
rect 2913 3353 2927 3367
rect 3013 3353 3027 3367
rect 3273 3353 3287 3367
rect 3353 3353 3367 3367
rect 3393 3353 3407 3367
rect 3473 3353 3487 3367
rect 3533 3353 3547 3367
rect 3713 3353 3727 3367
rect 3752 3353 3766 3367
rect 4113 3353 4127 3367
rect 4153 3353 4167 3367
rect 4213 3373 4227 3387
rect 4413 3373 4427 3387
rect 4793 3373 4807 3387
rect 4953 3373 4967 3387
rect 5093 3374 5107 3388
rect 5153 3373 5167 3387
rect 5193 3373 5207 3387
rect 5413 3373 5427 3387
rect 5893 3372 5907 3386
rect 4513 3353 4527 3367
rect 93 3333 107 3347
rect 193 3333 207 3347
rect 253 3333 267 3347
rect 433 3333 447 3347
rect 533 3333 547 3347
rect 1013 3333 1027 3347
rect 1353 3333 1367 3347
rect 1873 3333 1887 3347
rect 1933 3333 1947 3347
rect 2093 3333 2107 3347
rect 2253 3333 2267 3347
rect 2333 3333 2347 3347
rect 2493 3333 2507 3347
rect 2633 3333 2647 3347
rect 2753 3333 2767 3347
rect 593 3313 607 3327
rect 873 3313 887 3327
rect 913 3313 927 3327
rect 1333 3313 1347 3327
rect 1533 3313 1547 3327
rect 1613 3313 1627 3327
rect 2313 3313 2327 3327
rect 2393 3313 2407 3327
rect 2593 3313 2607 3327
rect 3633 3333 3647 3347
rect 3833 3333 3847 3347
rect 3893 3333 3907 3347
rect 4073 3333 4087 3347
rect 4133 3333 4147 3347
rect 4573 3353 4587 3367
rect 4673 3353 4687 3367
rect 4833 3353 4847 3367
rect 4933 3353 4947 3367
rect 4973 3353 4987 3367
rect 5094 3352 5108 3366
rect 5293 3353 5307 3367
rect 5373 3353 5387 3367
rect 5633 3353 5647 3367
rect 5953 3353 5967 3367
rect 6173 3353 6187 3367
rect 6273 3353 6287 3367
rect 6393 3353 6407 3367
rect 2933 3313 2947 3327
rect 2973 3313 2987 3327
rect 3113 3313 3127 3327
rect 3153 3313 3167 3327
rect 3353 3313 3367 3327
rect 3393 3313 3407 3327
rect 4553 3333 4567 3347
rect 4593 3333 4607 3347
rect 4693 3333 4707 3347
rect 4753 3333 4767 3347
rect 5133 3333 5147 3347
rect 5733 3333 5747 3347
rect 5773 3333 5787 3347
rect 6013 3333 6027 3347
rect 6093 3333 6107 3347
rect 6253 3333 6267 3347
rect 6293 3333 6307 3347
rect 4253 3313 4267 3327
rect 4293 3313 4307 3327
rect 5953 3313 5967 3327
rect 5993 3313 6007 3327
rect 53 3293 67 3307
rect 253 3293 267 3307
rect 313 3293 327 3307
rect 473 3293 487 3307
rect 553 3293 567 3307
rect 633 3293 647 3307
rect 793 3293 807 3307
rect 1013 3293 1027 3307
rect 1073 3293 1087 3307
rect 1473 3293 1487 3307
rect 1653 3293 1667 3307
rect 1693 3293 1707 3307
rect 1733 3293 1747 3307
rect 1813 3293 1827 3307
rect 1933 3293 1947 3307
rect 2033 3293 2047 3307
rect 2093 3293 2107 3307
rect 2193 3293 2207 3307
rect 2233 3293 2247 3307
rect 2413 3293 2427 3307
rect 2633 3293 2647 3307
rect 2753 3293 2767 3307
rect 3033 3293 3047 3307
rect 3233 3293 3247 3307
rect 3273 3293 3287 3307
rect 3433 3293 3447 3307
rect 3473 3293 3487 3307
rect 3513 3293 3527 3307
rect 3553 3293 3567 3307
rect 3693 3293 3707 3307
rect 3893 3293 3907 3307
rect 3933 3293 3947 3307
rect 4213 3293 4227 3307
rect 4413 3293 4427 3307
rect 4553 3293 4567 3307
rect 4693 3293 4707 3307
rect 4873 3293 4887 3307
rect 4953 3293 4967 3307
rect 5093 3293 5107 3307
rect 5133 3293 5147 3307
rect 5193 3293 5207 3307
rect 5293 3293 5307 3307
rect 5413 3293 5427 3307
rect 5453 3293 5467 3307
rect 5573 3293 5587 3307
rect 5633 3293 5647 3307
rect 5773 3293 5787 3307
rect 6093 3293 6107 3307
rect 6172 3293 6186 3307
rect 6333 3293 6347 3307
rect 6413 3293 6427 3307
rect 6453 3293 6467 3307
rect 2013 3273 2027 3287
rect 2053 3273 2067 3287
rect 5033 3273 5047 3287
rect 5073 3273 5087 3287
rect 973 3253 987 3267
rect 1573 3253 1587 3267
rect 1613 3253 1627 3267
rect 1733 3253 1747 3267
rect 2193 3253 2207 3267
rect 2913 3253 2927 3267
rect 2953 3253 2967 3267
rect 2993 3253 3007 3267
rect 3153 3253 3167 3267
rect 3213 3253 3227 3267
rect 3333 3253 3347 3267
rect 3413 3253 3427 3267
rect 3633 3253 3647 3267
rect 3653 3253 3667 3267
rect 3713 3253 3727 3267
rect 4052 3253 4066 3267
rect 4074 3253 4088 3267
rect 4233 3253 4247 3267
rect 4313 3253 4327 3267
rect 4492 3253 4506 3267
rect 4533 3253 4547 3267
rect 5613 3253 5627 3267
rect 5673 3253 5687 3267
rect 5933 3253 5947 3267
rect 6013 3253 6027 3267
rect 6433 3253 6447 3267
rect 93 3233 107 3247
rect 133 3233 147 3247
rect 233 3233 247 3247
rect 273 3233 287 3247
rect 393 3233 407 3247
rect 433 3233 447 3247
rect 533 3233 547 3247
rect 573 3233 587 3247
rect 673 3233 687 3247
rect 733 3233 747 3247
rect 773 3233 787 3247
rect 1033 3233 1047 3247
rect 1153 3233 1167 3247
rect 1213 3233 1227 3247
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1453 3233 1467 3247
rect 1873 3233 1887 3247
rect 1913 3233 1927 3247
rect 1953 3233 1967 3247
rect 1993 3233 2007 3247
rect 2073 3233 2087 3247
rect 2113 3233 2127 3247
rect 2253 3233 2267 3247
rect 2293 3233 2307 3247
rect 2393 3233 2407 3247
rect 2433 3233 2447 3247
rect 2573 3233 2587 3247
rect 2613 3233 2627 3247
rect 2733 3233 2747 3247
rect 2773 3233 2787 3247
rect 993 3213 1007 3227
rect 2813 3213 2827 3227
rect 2853 3213 2867 3227
rect 3373 3233 3387 3247
rect 3493 3233 3507 3247
rect 3533 3233 3547 3247
rect 4273 3233 4287 3247
rect 2973 3213 2987 3227
rect 3453 3213 3467 3227
rect 3893 3213 3907 3227
rect 3973 3213 3987 3227
rect 4053 3213 4067 3227
rect 4233 3213 4247 3227
rect 4313 3213 4327 3227
rect 4553 3233 4567 3247
rect 4633 3234 4647 3248
rect 4673 3233 4687 3247
rect 4713 3233 4727 3247
rect 4753 3233 4767 3247
rect 4973 3233 4987 3247
rect 5013 3233 5027 3247
rect 5113 3233 5127 3247
rect 5153 3233 5167 3247
rect 5233 3233 5247 3247
rect 5273 3233 5287 3247
rect 5313 3233 5327 3247
rect 5433 3233 5447 3247
rect 5473 3233 5487 3247
rect 5753 3233 5767 3247
rect 5793 3233 5807 3247
rect 4633 3212 4647 3226
rect 6113 3233 6127 3247
rect 6153 3233 6167 3247
rect 6313 3233 6327 3247
rect 6353 3233 6367 3247
rect 6073 3213 6087 3227
rect 213 3193 227 3207
rect 273 3193 287 3207
rect 393 3193 407 3207
rect 533 3193 547 3207
rect 1153 3193 1167 3207
rect 1533 3193 1547 3207
rect 1913 3193 1927 3207
rect 2113 3193 2127 3207
rect 2293 3193 2307 3207
rect 2373 3193 2387 3207
rect 2413 3193 2427 3207
rect 2473 3193 2487 3207
rect 2913 3193 2927 3207
rect 3233 3193 3247 3207
rect 3273 3193 3287 3207
rect 4293 3193 4307 3207
rect 4693 3193 4707 3207
rect 4813 3193 4827 3207
rect 5113 3193 5127 3207
rect 5273 3193 5287 3207
rect 5653 3193 5667 3207
rect 5733 3193 5747 3207
rect 5933 3193 5947 3207
rect 6153 3193 6167 3207
rect 6413 3213 6427 3227
rect 6473 3213 6487 3227
rect 133 3173 147 3187
rect 233 3173 247 3187
rect 633 3173 647 3187
rect 773 3173 787 3187
rect 833 3173 847 3187
rect 1333 3173 1347 3187
rect 1453 3173 1467 3187
rect 2493 3173 2507 3187
rect 673 3153 687 3167
rect 913 3153 927 3167
rect 1153 3153 1167 3167
rect 1473 3153 1487 3167
rect 2013 3153 2027 3167
rect 2953 3173 2967 3187
rect 3293 3173 3307 3187
rect 3373 3173 3387 3187
rect 3453 3173 3467 3187
rect 3653 3173 3667 3187
rect 3193 3153 3207 3167
rect 3513 3153 3527 3167
rect 3593 3153 3607 3167
rect 4333 3173 4347 3187
rect 4373 3173 4387 3187
rect 4453 3173 4467 3187
rect 4573 3173 4587 3187
rect 4793 3173 4807 3187
rect 4973 3173 4987 3187
rect 5033 3173 5047 3187
rect 5253 3173 5267 3187
rect 5413 3173 5427 3187
rect 4113 3153 4127 3167
rect 4873 3153 4887 3167
rect 5013 3153 5027 3167
rect 5153 3153 5167 3167
rect 5393 3154 5407 3168
rect 5453 3153 5467 3167
rect 5573 3173 5587 3187
rect 5753 3173 5767 3187
rect 5673 3153 5687 3167
rect 5813 3153 5827 3167
rect 5993 3153 6007 3167
rect 6353 3153 6367 3167
rect 6513 3153 6527 3167
rect 2373 3133 2387 3147
rect 2453 3133 2467 3147
rect 2513 3133 2527 3147
rect 2893 3133 2907 3147
rect 2953 3133 2967 3147
rect 3753 3133 3767 3147
rect 3913 3133 3927 3147
rect 4353 3133 4367 3147
rect 1133 3113 1147 3127
rect 1353 3113 1367 3127
rect 2613 3113 2627 3127
rect 3793 3113 3807 3127
rect 3833 3113 3847 3127
rect 4053 3113 4067 3127
rect 4153 3113 4167 3127
rect 4593 3113 4607 3127
rect 4653 3113 4667 3127
rect 4693 3133 4707 3147
rect 4933 3133 4947 3147
rect 5053 3133 5067 3147
rect 5393 3132 5407 3146
rect 5773 3113 5787 3127
rect 5873 3113 5887 3127
rect 6033 3113 6047 3127
rect 6093 3113 6107 3127
rect 6233 3113 6247 3127
rect 573 3093 587 3107
rect 813 3093 827 3107
rect 1253 3093 1267 3107
rect 2253 3093 2267 3107
rect 2493 3093 2507 3107
rect 2534 3093 2548 3107
rect 2573 3093 2587 3107
rect 2813 3094 2827 3108
rect 2913 3093 2927 3107
rect 2953 3093 2967 3107
rect 4393 3093 4407 3107
rect 4913 3093 4927 3107
rect 5033 3093 5047 3107
rect 5813 3093 5827 3107
rect 6353 3093 6367 3107
rect 6472 3093 6486 3107
rect 6513 3093 6527 3107
rect 753 3073 767 3087
rect 1073 3073 1087 3087
rect 1473 3073 1487 3087
rect 1613 3073 1627 3087
rect 1653 3073 1667 3087
rect 1973 3073 1987 3087
rect 2433 3073 2447 3087
rect 2773 3073 2787 3087
rect 2813 3072 2827 3086
rect 2893 3073 2907 3087
rect 3213 3073 3227 3087
rect 3813 3073 3827 3087
rect 4113 3073 4127 3087
rect 4253 3073 4267 3087
rect 4433 3073 4447 3087
rect 4713 3073 4727 3087
rect 4933 3073 4947 3087
rect 5073 3073 5087 3087
rect 6013 3073 6027 3087
rect 6073 3073 6087 3087
rect 6213 3074 6227 3088
rect 53 3053 67 3067
rect 93 3053 107 3067
rect 833 3053 847 3067
rect 873 3053 887 3067
rect 933 3053 947 3067
rect 1393 3053 1407 3067
rect 1573 3053 1587 3067
rect 1693 3053 1707 3067
rect 1773 3053 1787 3067
rect 1913 3053 1927 3067
rect 2333 3053 2347 3067
rect 2373 3053 2387 3067
rect 2413 3053 2427 3067
rect 2452 3053 2466 3067
rect 2474 3053 2488 3067
rect 2513 3053 2527 3067
rect 2613 3053 2627 3067
rect 2653 3053 2667 3067
rect 2953 3053 2967 3067
rect 4053 3053 4067 3067
rect 4173 3053 4187 3067
rect 4213 3053 4227 3067
rect 4293 3053 4307 3067
rect 4453 3053 4467 3067
rect 5013 3053 5027 3067
rect 5193 3053 5207 3067
rect 5373 3053 5387 3067
rect 5533 3053 5547 3067
rect 5713 3053 5727 3067
rect 5873 3053 5887 3067
rect 5993 3053 6007 3067
rect 6213 3052 6227 3066
rect 6313 3053 6327 3067
rect 6373 3053 6387 3067
rect 93 3013 107 3027
rect 273 3013 287 3027
rect 313 3013 327 3027
rect 473 3013 487 3027
rect 513 3013 527 3027
rect 793 3013 807 3027
rect 833 3013 847 3027
rect 873 3013 887 3027
rect 1053 3013 1067 3027
rect 1173 3013 1187 3027
rect 1213 3013 1227 3027
rect 1253 3013 1267 3027
rect 1353 3013 1367 3027
rect 1493 3013 1507 3027
rect 1613 3013 1627 3027
rect 1653 3013 1667 3027
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 2073 3013 2087 3027
rect 2233 3034 2247 3048
rect 2233 3012 2247 3026
rect 2273 3013 2287 3027
rect 2313 3013 2327 3027
rect 2433 3013 2447 3027
rect 2473 3013 2487 3027
rect 2613 3013 2627 3027
rect 2653 3013 2667 3027
rect 2833 3033 2847 3047
rect 3013 3013 3027 3027
rect 3153 3013 3167 3027
rect 3433 3013 3447 3027
rect 3813 3013 3827 3027
rect 4033 3033 4047 3047
rect 4833 3033 4847 3047
rect 4013 3013 4027 3027
rect 4073 3014 4087 3028
rect 4113 3013 4127 3027
rect 4153 3013 4167 3027
rect 4253 3013 4267 3027
rect 4293 3013 4307 3027
rect 4433 3013 4447 3027
rect 4473 3013 4487 3027
rect 4513 3013 4527 3027
rect 4553 3013 4567 3027
rect 4593 3013 4607 3027
rect 4733 3013 4747 3027
rect 4773 3013 4787 3027
rect 4873 3013 4887 3027
rect 4913 3013 4927 3027
rect 5033 3013 5047 3027
rect 5073 3013 5087 3027
rect 5213 3013 5227 3027
rect 5253 3013 5267 3027
rect 5373 3013 5387 3027
rect 5413 3013 5427 3027
rect 5533 3013 5547 3027
rect 5573 3013 5587 3027
rect 5673 3013 5687 3027
rect 5713 3013 5727 3027
rect 5833 3013 5847 3027
rect 5873 3013 5887 3027
rect 6013 3013 6027 3027
rect 6053 3013 6067 3027
rect 6213 3013 6227 3027
rect 6253 3013 6267 3027
rect 6373 3013 6387 3027
rect 6413 3013 6427 3027
rect 6513 3013 6527 3027
rect 233 2993 247 3007
rect 573 2993 587 3007
rect 673 2993 687 3007
rect 1893 2993 1907 3007
rect 2753 2993 2767 3007
rect 2833 2993 2847 3007
rect 3233 2993 3247 3007
rect 3293 2993 3307 3007
rect 3673 2993 3687 3007
rect 3853 2993 3867 3007
rect 3913 2993 3927 3007
rect 4073 2992 4087 3006
rect 4953 2993 4967 3007
rect 4993 2993 5007 3007
rect 2493 2973 2507 2987
rect 2553 2973 2567 2987
rect 4853 2973 4867 2987
rect 6433 2973 6447 2987
rect 113 2953 127 2967
rect 333 2953 347 2967
rect 493 2953 507 2967
rect 633 2953 647 2967
rect 693 2953 707 2967
rect 853 2953 867 2967
rect 933 2953 947 2967
rect 973 2953 987 2967
rect 1073 2953 1087 2967
rect 1153 2953 1167 2967
rect 1333 2953 1347 2967
rect 1593 2953 1607 2967
rect 1633 2953 1647 2967
rect 1793 2953 1807 2967
rect 1993 2953 2007 2967
rect 2093 2953 2107 2967
rect 2293 2953 2307 2967
rect 2413 2953 2427 2967
rect 2453 2953 2467 2967
rect 2633 2953 2647 2967
rect 2853 2953 2867 2967
rect 2993 2953 3007 2967
rect 3053 2953 3067 2967
rect 3113 2953 3127 2967
rect 3413 2953 3427 2967
rect 3453 2953 3467 2967
rect 3653 2953 3667 2967
rect 3893 2953 3907 2967
rect 3933 2953 3947 2967
rect 4213 2953 4227 2967
rect 4313 2953 4327 2967
rect 4453 2953 4467 2967
rect 4573 2953 4587 2967
rect 4633 2953 4647 2967
rect 4753 2953 4767 2967
rect 4793 2953 4807 2967
rect 4893 2953 4907 2967
rect 5053 2953 5067 2967
rect 5193 2953 5207 2967
rect 5353 2953 5367 2967
rect 5513 2953 5527 2967
rect 5653 2953 5667 2967
rect 5693 2953 5707 2967
rect 5813 2953 5827 2967
rect 5853 2953 5867 2967
rect 5913 2953 5927 2967
rect 5973 2953 5987 2967
rect 6033 2953 6047 2967
rect 6113 2953 6127 2967
rect 6233 2953 6247 2967
rect 6273 2953 6287 2967
rect 6393 2953 6407 2967
rect 333 2913 347 2927
rect 393 2913 407 2927
rect 813 2913 827 2927
rect 853 2913 867 2927
rect 1093 2913 1107 2927
rect 1653 2913 1667 2927
rect 1733 2933 1747 2947
rect 1773 2933 1787 2947
rect 1813 2913 1827 2927
rect 2593 2933 2607 2947
rect 2773 2933 2787 2947
rect 2813 2933 2827 2947
rect 2733 2913 2747 2927
rect 3213 2913 3227 2927
rect 4273 2933 4287 2947
rect 3653 2913 3667 2927
rect 4833 2933 4847 2947
rect 4873 2933 4887 2947
rect 4533 2913 4547 2927
rect 4573 2913 4587 2927
rect 4732 2913 4746 2927
rect 4754 2913 4768 2927
rect 4993 2933 5007 2947
rect 5233 2933 5247 2947
rect 5933 2933 5947 2947
rect 5413 2913 5427 2927
rect 5473 2913 5487 2927
rect 5693 2913 5707 2927
rect 5853 2913 5867 2927
rect 6193 2933 6207 2947
rect 6033 2913 6047 2927
rect 6233 2913 6247 2927
rect 6273 2913 6287 2927
rect 6353 2914 6367 2928
rect 6393 2913 6407 2927
rect 253 2893 267 2907
rect 553 2893 567 2907
rect 793 2893 807 2907
rect 933 2893 947 2907
rect 1053 2893 1067 2907
rect 1113 2893 1127 2907
rect 2073 2893 2087 2907
rect 2453 2893 2467 2907
rect 2534 2893 2548 2907
rect 2973 2893 2987 2907
rect 3433 2893 3447 2907
rect 3493 2893 3507 2907
rect 3573 2893 3587 2907
rect 3613 2893 3627 2907
rect 3933 2893 3947 2907
rect 4253 2893 4267 2907
rect 4353 2893 4367 2907
rect 4553 2893 4567 2907
rect 4593 2893 4607 2907
rect 4813 2893 4827 2907
rect 4874 2893 4888 2907
rect 5073 2893 5087 2907
rect 5353 2893 5367 2907
rect 5513 2893 5527 2907
rect 5873 2893 5887 2907
rect 6132 2893 6146 2907
rect 6173 2893 6187 2907
rect 6253 2893 6267 2907
rect 453 2873 467 2887
rect 1013 2873 1027 2887
rect 1073 2873 1087 2887
rect 1333 2873 1347 2887
rect 1633 2873 1647 2887
rect 1733 2873 1747 2887
rect 2093 2873 2107 2887
rect 2253 2873 2267 2887
rect 2393 2873 2407 2887
rect 2513 2873 2527 2887
rect 2593 2873 2607 2887
rect 2773 2873 2787 2887
rect 2893 2873 2907 2887
rect 3153 2873 3167 2887
rect 3193 2873 3207 2887
rect 493 2853 507 2867
rect 1113 2853 1127 2867
rect 2353 2853 2367 2867
rect 2413 2853 2427 2867
rect 3033 2853 3047 2867
rect 3233 2853 3247 2867
rect 3273 2873 3287 2887
rect 3773 2873 3787 2887
rect 4073 2873 4087 2887
rect 4493 2873 4507 2887
rect 4533 2873 4547 2887
rect 6353 2892 6367 2906
rect 5053 2873 5067 2887
rect 5113 2873 5127 2887
rect 5193 2873 5207 2887
rect 5253 2873 5267 2887
rect 5433 2873 5447 2887
rect 5473 2873 5487 2887
rect 5573 2873 5587 2887
rect 5733 2873 5747 2887
rect 5973 2873 5987 2887
rect 6293 2873 6307 2887
rect 6413 2873 6427 2887
rect 3533 2853 3547 2867
rect 3573 2853 3587 2867
rect 3853 2853 3867 2867
rect 3893 2853 3907 2867
rect 173 2833 187 2847
rect 573 2833 587 2847
rect 893 2833 907 2847
rect 953 2833 967 2847
rect 1553 2833 1567 2847
rect 1593 2833 1607 2847
rect 1693 2833 1707 2847
rect 2073 2833 2087 2847
rect 2313 2834 2327 2848
rect 2373 2833 2387 2847
rect 2593 2833 2607 2847
rect 2733 2833 2747 2847
rect 3113 2833 3127 2847
rect 3273 2833 3287 2847
rect 3493 2833 3507 2847
rect 4393 2853 4407 2867
rect 4593 2853 4607 2867
rect 4693 2853 4707 2867
rect 4792 2853 4806 2867
rect 4814 2853 4828 2867
rect 4873 2853 4887 2867
rect 5073 2853 5087 2867
rect 5593 2853 5607 2867
rect 5993 2853 6007 2867
rect 6313 2853 6327 2867
rect 253 2813 267 2827
rect 313 2813 327 2827
rect 393 2813 407 2827
rect 753 2813 767 2827
rect 1773 2813 1787 2827
rect 1833 2813 1847 2827
rect 1973 2813 1987 2827
rect 2013 2813 2027 2827
rect 2133 2813 2147 2827
rect 2273 2813 2287 2827
rect 2312 2812 2326 2826
rect 2334 2813 2348 2827
rect 2453 2813 2467 2827
rect 93 2793 107 2807
rect 133 2793 147 2807
rect 1553 2793 1567 2807
rect 1693 2793 1707 2807
rect 1733 2793 1747 2807
rect 1993 2793 2007 2807
rect 2713 2813 2727 2827
rect 3713 2813 3727 2827
rect 3753 2813 3767 2827
rect 3853 2813 3867 2827
rect 4452 2833 4466 2847
rect 4913 2833 4927 2847
rect 4993 2833 5007 2847
rect 5153 2833 5167 2847
rect 5213 2833 5227 2847
rect 5573 2833 5587 2847
rect 5633 2833 5647 2847
rect 5833 2833 5847 2847
rect 5973 2833 5987 2847
rect 6193 2834 6207 2848
rect 6333 2833 6347 2847
rect 6393 2833 6407 2847
rect 4293 2813 4307 2827
rect 4573 2813 4587 2827
rect 4633 2813 4647 2827
rect 4673 2813 4687 2827
rect 4793 2813 4807 2827
rect 4953 2813 4967 2827
rect 3193 2793 3207 2807
rect 3233 2793 3247 2807
rect 4053 2793 4067 2807
rect 4133 2793 4147 2807
rect 4173 2793 4187 2807
rect 5133 2813 5147 2827
rect 5432 2813 5446 2827
rect 5454 2813 5468 2827
rect 6193 2812 6207 2826
rect 6313 2813 6327 2827
rect 6353 2813 6367 2827
rect 6173 2793 6187 2807
rect 253 2773 267 2787
rect 333 2773 347 2787
rect 453 2773 467 2787
rect 493 2773 507 2787
rect 553 2773 567 2787
rect 593 2773 607 2787
rect 693 2773 707 2787
rect 733 2773 747 2787
rect 873 2773 887 2787
rect 953 2773 967 2787
rect 1213 2773 1227 2787
rect 1493 2773 1507 2787
rect 1833 2773 1847 2787
rect 1913 2773 1927 2787
rect 2033 2773 2047 2787
rect 2153 2773 2167 2787
rect 2253 2773 2267 2787
rect 2313 2773 2327 2787
rect 2453 2773 2467 2787
rect 2653 2773 2667 2787
rect 2733 2773 2747 2787
rect 2813 2773 2827 2787
rect 2853 2773 2867 2787
rect 3473 2773 3487 2787
rect 3513 2773 3527 2787
rect 3633 2773 3647 2787
rect 3753 2773 3767 2787
rect 3853 2773 3867 2787
rect 4193 2773 4207 2787
rect 4353 2773 4367 2787
rect 4533 2773 4547 2787
rect 4653 2773 4667 2787
rect 4793 2773 4807 2787
rect 4953 2773 4967 2787
rect 5253 2773 5267 2787
rect 5313 2773 5327 2787
rect 5453 2773 5467 2787
rect 5553 2773 5567 2787
rect 5593 2773 5607 2787
rect 5673 2773 5687 2787
rect 5713 2773 5727 2787
rect 5833 2773 5847 2787
rect 5973 2773 5987 2787
rect 6033 2773 6047 2787
rect 6133 2773 6147 2787
rect 6333 2773 6347 2787
rect 6433 2773 6447 2787
rect 4693 2753 4707 2767
rect 4753 2753 4767 2767
rect 4913 2753 4927 2767
rect 5873 2753 5887 2767
rect 5933 2753 5947 2767
rect 193 2733 207 2747
rect 733 2733 747 2747
rect 1773 2733 1787 2747
rect 2973 2733 2987 2747
rect 3033 2733 3047 2747
rect 3173 2733 3187 2747
rect 3253 2733 3267 2747
rect 3293 2733 3307 2747
rect 3353 2733 3367 2747
rect 3653 2733 3667 2747
rect 3973 2733 3987 2747
rect 4013 2733 4027 2747
rect 4493 2733 4507 2747
rect 4633 2733 4647 2747
rect 5273 2733 5287 2747
rect 353 2713 367 2727
rect 393 2713 407 2727
rect 533 2713 547 2727
rect 573 2713 587 2727
rect 813 2713 827 2727
rect 853 2713 867 2727
rect 893 2713 907 2727
rect 1073 2713 1087 2727
rect 1113 2713 1127 2727
rect 1353 2713 1367 2727
rect 1393 2713 1407 2727
rect 1533 2713 1547 2727
rect 1573 2713 1587 2727
rect 1813 2713 1827 2727
rect 1853 2713 1867 2727
rect 2013 2713 2027 2727
rect 2053 2713 2067 2727
rect 2133 2713 2147 2727
rect 2173 2713 2187 2727
rect 2293 2713 2307 2727
rect 2333 2713 2347 2727
rect 2373 2713 2387 2727
rect 2593 2713 2607 2727
rect 2633 2713 2647 2727
rect 2753 2713 2767 2727
rect 2793 2713 2807 2727
rect 93 2693 107 2707
rect 133 2693 147 2707
rect 193 2673 207 2687
rect 333 2693 347 2707
rect 533 2673 547 2687
rect 633 2673 647 2687
rect 813 2673 827 2687
rect 1073 2673 1087 2687
rect 1213 2673 1227 2687
rect 2673 2693 2687 2707
rect 2733 2693 2747 2707
rect 3133 2693 3147 2707
rect 3533 2713 3547 2727
rect 4173 2713 4187 2727
rect 4213 2713 4227 2727
rect 4333 2713 4347 2727
rect 4773 2713 4787 2727
rect 4813 2713 4827 2727
rect 4933 2713 4947 2727
rect 4973 2713 4987 2727
rect 5113 2713 5127 2727
rect 5153 2713 5167 2727
rect 5433 2713 5447 2727
rect 5473 2713 5487 2727
rect 5613 2713 5627 2727
rect 5653 2713 5667 2727
rect 5813 2713 5827 2727
rect 5853 2713 5867 2727
rect 5953 2713 5967 2727
rect 5993 2713 6007 2727
rect 6153 2713 6167 2727
rect 6193 2713 6207 2727
rect 6313 2713 6327 2727
rect 6353 2713 6367 2727
rect 1393 2673 1407 2687
rect 1813 2673 1827 2687
rect 1973 2673 1987 2687
rect 2013 2673 2027 2687
rect 2113 2673 2127 2687
rect 2153 2673 2167 2687
rect 2293 2673 2307 2687
rect 1353 2653 1367 2667
rect 533 2633 547 2647
rect 1073 2633 1087 2647
rect 1193 2633 1207 2647
rect 1293 2633 1307 2647
rect 1933 2653 1947 2667
rect 2053 2653 2067 2667
rect 2193 2653 2207 2667
rect 2233 2653 2247 2667
rect 2513 2673 2527 2687
rect 2793 2673 2807 2687
rect 3293 2693 3307 2707
rect 3253 2673 3267 2687
rect 3493 2673 3507 2687
rect 3713 2673 3727 2687
rect 3813 2673 3827 2687
rect 3853 2673 3867 2687
rect 4113 2673 4127 2687
rect 4173 2674 4187 2688
rect 4233 2673 4247 2687
rect 2333 2653 2347 2667
rect 1413 2633 1427 2647
rect 1553 2633 1567 2647
rect 1853 2633 1867 2647
rect 1993 2633 2007 2647
rect 2113 2633 2127 2647
rect 2753 2633 2767 2647
rect 2833 2633 2847 2647
rect 3173 2653 3187 2667
rect 3093 2633 3107 2647
rect 3433 2633 3447 2647
rect 4053 2654 4067 2668
rect 4273 2674 4287 2688
rect 4432 2673 4446 2687
rect 4533 2673 4547 2687
rect 5093 2673 5107 2687
rect 5153 2673 5167 2687
rect 5273 2673 5287 2687
rect 5813 2673 5827 2687
rect 5993 2673 6007 2687
rect 6293 2673 6307 2687
rect 6353 2673 6367 2687
rect 4173 2652 4187 2666
rect 4213 2653 4227 2667
rect 4273 2652 4287 2666
rect 4553 2653 4567 2667
rect 4673 2653 4687 2667
rect 4933 2653 4947 2667
rect 5253 2653 5267 2667
rect 5653 2653 5667 2667
rect 5853 2653 5867 2667
rect 1053 2613 1067 2627
rect 1433 2613 1447 2627
rect 1873 2613 1887 2627
rect 1933 2613 1947 2627
rect 2393 2613 2407 2627
rect 2533 2613 2547 2627
rect 2573 2613 2587 2627
rect 2633 2613 2647 2627
rect 2692 2613 2706 2627
rect 2714 2613 2728 2627
rect 2893 2613 2907 2627
rect 3253 2613 3267 2627
rect 3313 2613 3327 2627
rect 3933 2633 3947 2647
rect 4013 2633 4027 2647
rect 4053 2632 4067 2646
rect 4132 2633 4146 2647
rect 4154 2633 4168 2647
rect 4233 2633 4247 2647
rect 4513 2633 4527 2647
rect 4613 2633 4627 2647
rect 5113 2633 5127 2647
rect 5313 2633 5327 2647
rect 5633 2633 5647 2647
rect 5713 2633 5727 2647
rect 6513 2633 6527 2647
rect 3673 2613 3687 2627
rect 1273 2593 1287 2607
rect 1533 2593 1547 2607
rect 1693 2593 1707 2607
rect 3093 2593 3107 2607
rect 3513 2593 3527 2607
rect 3653 2593 3667 2607
rect 4113 2613 4127 2627
rect 4193 2613 4207 2627
rect 4393 2613 4407 2627
rect 4473 2613 4487 2627
rect 4693 2613 4707 2627
rect 4733 2613 4747 2627
rect 4873 2613 4887 2627
rect 5393 2613 5407 2627
rect 5433 2613 5447 2627
rect 5953 2613 5967 2627
rect 6413 2613 6427 2627
rect 3793 2593 3807 2607
rect 4153 2593 4167 2607
rect 4293 2593 4307 2607
rect 4593 2593 4607 2607
rect 4773 2593 4787 2607
rect 4933 2593 4947 2607
rect 5313 2593 5327 2607
rect 5413 2593 5427 2607
rect 5773 2593 5787 2607
rect 5973 2593 5987 2607
rect 6093 2593 6107 2607
rect 6133 2593 6147 2607
rect 493 2573 507 2587
rect 893 2573 907 2587
rect 933 2573 947 2587
rect 1253 2573 1267 2587
rect 1333 2573 1347 2587
rect 1373 2573 1387 2587
rect 2412 2573 2426 2587
rect 2493 2573 2507 2587
rect 2793 2573 2807 2587
rect 133 2553 147 2567
rect 333 2553 347 2567
rect 793 2553 807 2567
rect 173 2533 187 2547
rect 293 2533 307 2547
rect 673 2533 687 2547
rect 773 2533 787 2547
rect 853 2533 867 2547
rect 933 2533 947 2547
rect 1193 2553 1207 2567
rect 1393 2553 1407 2567
rect 1433 2553 1447 2567
rect 2212 2553 2226 2567
rect 2234 2553 2248 2567
rect 2353 2553 2367 2567
rect 2393 2553 2407 2567
rect 2553 2553 2567 2567
rect 3153 2573 3167 2587
rect 3712 2573 3726 2587
rect 3773 2573 3787 2587
rect 3913 2573 3927 2587
rect 4113 2573 4127 2587
rect 4193 2573 4207 2587
rect 4553 2573 4567 2587
rect 4633 2573 4647 2587
rect 4813 2573 4827 2587
rect 5212 2573 5226 2587
rect 5234 2573 5248 2587
rect 5373 2573 5387 2587
rect 5573 2573 5587 2587
rect 6073 2573 6087 2587
rect 2853 2553 2867 2567
rect 1013 2533 1027 2547
rect 1153 2533 1167 2547
rect 1213 2533 1227 2547
rect 3053 2553 3067 2567
rect 3113 2553 3127 2567
rect 3753 2553 3767 2567
rect 3973 2553 3987 2567
rect 4073 2554 4087 2568
rect 4153 2553 4167 2567
rect 4613 2553 4627 2567
rect 4973 2553 4987 2567
rect 5193 2553 5207 2567
rect 5613 2553 5627 2567
rect 6213 2553 6227 2567
rect 1753 2533 1767 2547
rect 1973 2533 1987 2547
rect 2013 2533 2027 2547
rect 2053 2533 2067 2547
rect 2373 2533 2387 2547
rect 2413 2533 2427 2547
rect 2613 2533 2627 2547
rect 2653 2533 2667 2547
rect 2713 2533 2727 2547
rect 2813 2533 2827 2547
rect 2913 2533 2927 2547
rect 2953 2533 2967 2547
rect 3353 2533 3367 2547
rect 3532 2533 3546 2547
rect 3572 2533 3586 2547
rect 3853 2533 3867 2547
rect 3913 2533 3927 2547
rect 4073 2532 4087 2546
rect 4373 2533 4387 2547
rect 4413 2533 4427 2547
rect 4493 2533 4507 2547
rect 4633 2533 4647 2547
rect 4712 2533 4726 2547
rect 5173 2533 5187 2547
rect 1133 2513 1147 2527
rect 133 2493 147 2507
rect 173 2493 187 2507
rect 293 2493 307 2507
rect 333 2493 347 2507
rect 453 2493 467 2507
rect 493 2493 507 2507
rect 593 2493 607 2507
rect 633 2493 647 2507
rect 733 2493 747 2507
rect 773 2493 787 2507
rect 1013 2493 1027 2507
rect 1053 2493 1067 2507
rect 1313 2513 1327 2527
rect 1553 2493 1567 2507
rect 1593 2493 1607 2507
rect 1713 2493 1727 2507
rect 1753 2493 1767 2507
rect 2013 2493 2027 2507
rect 2053 2493 2067 2507
rect 2433 2513 2447 2527
rect 2533 2513 2547 2527
rect 3633 2514 3647 2528
rect 4913 2513 4927 2527
rect 4993 2513 5007 2527
rect 5093 2514 5107 2528
rect 5513 2533 5527 2547
rect 5633 2533 5647 2547
rect 5793 2533 5807 2547
rect 5913 2533 5927 2547
rect 6033 2533 6047 2547
rect 6233 2533 6247 2547
rect 5733 2513 5747 2527
rect 2373 2493 2387 2507
rect 2473 2493 2487 2507
rect 2513 2493 2527 2507
rect 2613 2493 2627 2507
rect 2653 2493 2667 2507
rect 2893 2493 2907 2507
rect 2933 2493 2947 2507
rect 3073 2493 3087 2507
rect 3113 2493 3127 2507
rect 3432 2493 3446 2507
rect 3533 2493 3547 2507
rect 3633 2492 3647 2506
rect 3733 2493 3747 2507
rect 3793 2493 3807 2507
rect 3833 2493 3847 2507
rect 3913 2493 3927 2507
rect 3933 2493 3947 2507
rect 3973 2493 3987 2507
rect 4093 2493 4107 2507
rect 4133 2493 4147 2507
rect 4193 2493 4207 2507
rect 4373 2493 4387 2507
rect 4413 2493 4427 2507
rect 4673 2493 4687 2507
rect 4713 2493 4727 2507
rect 4793 2493 4807 2507
rect 4833 2493 4847 2507
rect 4873 2493 4887 2507
rect 5013 2493 5027 2507
rect 5053 2493 5067 2507
rect 5093 2492 5107 2506
rect 5133 2493 5147 2507
rect 5173 2493 5187 2507
rect 5213 2493 5227 2507
rect 5313 2493 5327 2507
rect 5353 2493 5367 2507
rect 5773 2493 5787 2507
rect 5813 2493 5827 2507
rect 5853 2493 5867 2507
rect 6033 2493 6047 2507
rect 6073 2493 6087 2507
rect 6213 2493 6227 2507
rect 6253 2493 6267 2507
rect 6313 2493 6327 2507
rect 1153 2473 1167 2487
rect 1233 2473 1247 2487
rect 1353 2473 1367 2487
rect 1433 2473 1447 2487
rect 1513 2473 1527 2487
rect 1853 2473 1867 2487
rect 1973 2473 1987 2487
rect 2093 2473 2107 2487
rect 2233 2473 2247 2487
rect 2273 2473 2287 2487
rect 2773 2473 2787 2487
rect 3153 2473 3167 2487
rect 3293 2473 3307 2487
rect 3653 2473 3667 2487
rect 4493 2473 4507 2487
rect 4633 2473 4647 2487
rect 5453 2473 5467 2487
rect 5513 2473 5527 2487
rect 5633 2473 5647 2487
rect 2453 2453 2467 2467
rect 93 2433 107 2447
rect 153 2433 167 2447
rect 193 2433 207 2447
rect 313 2433 327 2447
rect 473 2433 487 2447
rect 673 2433 687 2447
rect 713 2433 727 2447
rect 793 2433 807 2447
rect 1013 2433 1027 2447
rect 1593 2433 1607 2447
rect 1693 2433 1707 2447
rect 1893 2433 1907 2447
rect 2013 2433 2027 2447
rect 2093 2433 2107 2447
rect 2153 2433 2167 2447
rect 2193 2433 2207 2447
rect 2373 2433 2387 2447
rect 2533 2433 2547 2447
rect 2613 2433 2627 2447
rect 2813 2433 2827 2447
rect 2913 2433 2927 2447
rect 3053 2433 3067 2447
rect 3253 2433 3267 2447
rect 3413 2433 3427 2447
rect 3614 2433 3628 2447
rect 3873 2433 3887 2447
rect 3933 2433 3947 2447
rect 4073 2433 4087 2447
rect 4133 2433 4147 2447
rect 4273 2433 4287 2447
rect 4413 2433 4427 2447
rect 4533 2433 4547 2447
rect 4653 2433 4667 2447
rect 4773 2433 4787 2447
rect 4933 2433 4947 2447
rect 4993 2433 5007 2447
rect 5493 2433 5507 2447
rect 5793 2433 5807 2447
rect 5893 2433 5907 2447
rect 5913 2433 5927 2447
rect 5973 2433 5987 2447
rect 113 2413 127 2427
rect 893 2413 907 2427
rect 933 2413 947 2427
rect 1173 2413 1187 2427
rect 1213 2413 1227 2427
rect 1373 2413 1387 2427
rect 1413 2413 1427 2427
rect 1733 2413 1747 2427
rect 2953 2413 2967 2427
rect 6193 2430 6207 2444
rect 6413 2433 6427 2447
rect 3093 2413 3107 2427
rect 3773 2413 3787 2427
rect 4813 2413 4827 2427
rect 4892 2413 4906 2427
rect 153 2393 167 2407
rect 313 2393 327 2407
rect 374 2393 388 2407
rect 453 2393 467 2407
rect 573 2393 587 2407
rect 1453 2393 1467 2407
rect 1853 2393 1867 2407
rect 1913 2393 1927 2407
rect 1993 2393 2007 2407
rect 2133 2393 2147 2407
rect 2193 2393 2207 2407
rect 2273 2393 2287 2407
rect 2313 2393 2327 2407
rect 2473 2393 2487 2407
rect 3293 2393 3307 2407
rect 3433 2393 3447 2407
rect 3513 2393 3527 2407
rect 3594 2393 3608 2407
rect 4053 2393 4067 2407
rect 4333 2393 4347 2407
rect 4473 2393 4487 2407
rect 4613 2393 4627 2407
rect 4713 2393 4727 2407
rect 4753 2393 4767 2407
rect 4833 2393 4847 2407
rect 5093 2413 5107 2427
rect 5293 2413 5307 2427
rect 5613 2413 5627 2427
rect 5653 2413 5667 2427
rect 4913 2393 4927 2407
rect 4953 2393 4967 2407
rect 5033 2393 5047 2407
rect 5113 2393 5127 2407
rect 5353 2393 5367 2407
rect 5493 2393 5507 2407
rect 5533 2393 5547 2407
rect 5713 2393 5727 2407
rect 5773 2393 5787 2407
rect 6113 2390 6127 2404
rect 6193 2390 6207 2404
rect 473 2373 487 2387
rect 533 2373 547 2387
rect 413 2353 427 2367
rect 593 2353 607 2367
rect 1753 2373 1767 2387
rect 1813 2373 1827 2387
rect 1093 2353 1107 2367
rect 1273 2353 1287 2367
rect 1553 2353 1567 2367
rect 2413 2373 2427 2387
rect 2533 2373 2547 2387
rect 2573 2373 2587 2387
rect 2653 2373 2667 2387
rect 2833 2373 2847 2387
rect 2892 2373 2906 2387
rect 2914 2373 2928 2387
rect 3093 2374 3107 2388
rect 3153 2373 3167 2387
rect 3553 2373 3567 2387
rect 3713 2373 3727 2387
rect 4113 2373 4127 2387
rect 4253 2373 4267 2387
rect 4293 2373 4307 2387
rect 4653 2373 4667 2387
rect 4693 2373 4707 2387
rect 5433 2373 5447 2387
rect 5793 2373 5807 2387
rect 5853 2373 5867 2387
rect 6213 2373 6227 2387
rect 2253 2353 2267 2367
rect 2433 2353 2447 2367
rect 2613 2353 2627 2367
rect 793 2333 807 2347
rect 893 2333 907 2347
rect 1013 2334 1027 2348
rect 1193 2333 1207 2347
rect 1373 2333 1387 2347
rect 1833 2333 1847 2347
rect 2193 2333 2207 2347
rect 2413 2333 2427 2347
rect 2553 2333 2567 2347
rect 3093 2352 3107 2366
rect 773 2313 787 2327
rect 853 2313 867 2327
rect 933 2313 947 2327
rect 1013 2312 1027 2326
rect 1053 2313 1067 2327
rect 1233 2313 1247 2327
rect 1493 2313 1507 2327
rect 1692 2313 1706 2327
rect 1714 2313 1728 2327
rect 1793 2313 1807 2327
rect 1893 2313 1907 2327
rect 2332 2313 2346 2327
rect 2354 2313 2368 2327
rect 2473 2313 2487 2327
rect 2593 2313 2607 2327
rect 2733 2313 2747 2327
rect 2813 2313 2827 2327
rect 3153 2334 3167 2348
rect 3653 2353 3667 2367
rect 4013 2353 4027 2367
rect 4073 2353 4087 2367
rect 4193 2353 4207 2367
rect 3193 2333 3207 2347
rect 3313 2333 3327 2347
rect 3713 2333 3727 2347
rect 4533 2353 4547 2367
rect 4973 2353 4987 2367
rect 5153 2353 5167 2367
rect 5293 2353 5307 2367
rect 5453 2353 5467 2367
rect 5613 2353 5627 2367
rect 5833 2353 5847 2367
rect 6033 2353 6047 2367
rect 4333 2333 4347 2347
rect 4373 2333 4387 2347
rect 4413 2333 4427 2347
rect 5113 2333 5127 2347
rect 5313 2333 5327 2347
rect 5593 2333 5607 2347
rect 5653 2333 5667 2347
rect 2993 2314 3007 2328
rect 6213 2333 6227 2347
rect 3153 2312 3167 2326
rect 3253 2313 3267 2327
rect 3373 2313 3387 2327
rect 3413 2313 3427 2327
rect 3593 2313 3607 2327
rect 3913 2313 3927 2327
rect 4233 2313 4247 2327
rect 4433 2313 4447 2327
rect 4593 2313 4607 2327
rect 4813 2313 4827 2327
rect 4853 2313 4867 2327
rect 4993 2313 5007 2327
rect 5093 2313 5107 2327
rect 5173 2313 5187 2327
rect 5213 2313 5227 2327
rect 5253 2313 5267 2327
rect 5333 2313 5347 2327
rect 5433 2313 5447 2327
rect 5713 2313 5727 2327
rect 5753 2313 5767 2327
rect 5893 2313 5907 2327
rect 6033 2313 6047 2327
rect 6233 2313 6247 2327
rect 6313 2313 6327 2327
rect 553 2293 567 2307
rect 1213 2293 1227 2307
rect 1353 2293 1367 2307
rect 1473 2293 1487 2307
rect 1593 2293 1607 2307
rect 1633 2293 1647 2307
rect 1733 2293 1747 2307
rect 853 2273 867 2287
rect 893 2273 907 2287
rect 2173 2273 2187 2287
rect 2293 2293 2307 2307
rect 2633 2293 2647 2307
rect 2713 2293 2727 2307
rect 2793 2292 2807 2306
rect 2833 2293 2847 2307
rect 2873 2293 2887 2307
rect 2993 2292 3007 2306
rect 3053 2293 3067 2307
rect 3113 2293 3127 2307
rect 3773 2293 3787 2307
rect 4333 2293 4347 2307
rect 4513 2293 4527 2307
rect 4933 2293 4947 2307
rect 5193 2293 5207 2307
rect 5233 2293 5247 2307
rect 5373 2293 5387 2307
rect 5673 2293 5687 2307
rect 5873 2293 5887 2307
rect 2853 2273 2867 2287
rect 3333 2273 3347 2287
rect 3373 2273 3387 2287
rect 3553 2273 3567 2287
rect 3593 2273 3607 2287
rect 3633 2273 3647 2287
rect 3693 2273 3707 2287
rect 3893 2273 3907 2287
rect 3933 2273 3947 2287
rect 5833 2273 5847 2287
rect 6173 2293 6187 2307
rect 6273 2293 6287 2307
rect 6373 2293 6387 2307
rect 6433 2293 6447 2307
rect 6213 2273 6227 2287
rect 133 2253 147 2267
rect 153 2253 167 2267
rect 273 2253 287 2267
rect 413 2253 427 2267
rect 493 2253 507 2267
rect 633 2253 647 2267
rect 693 2253 707 2267
rect 773 2253 787 2267
rect 933 2253 947 2267
rect 1173 2253 1187 2267
rect 1213 2253 1227 2267
rect 1353 2253 1367 2267
rect 1393 2253 1407 2267
rect 1493 2253 1507 2267
rect 1533 2253 1547 2267
rect 1633 2253 1647 2267
rect 1813 2253 1827 2267
rect 1953 2253 1967 2267
rect 2053 2253 2067 2267
rect 2113 2253 2127 2267
rect 2253 2253 2267 2267
rect 2293 2253 2307 2267
rect 2433 2253 2447 2267
rect 2553 2253 2567 2267
rect 2653 2253 2667 2267
rect 2713 2253 2727 2267
rect 2813 2253 2827 2267
rect 2913 2253 2927 2267
rect 3193 2253 3207 2267
rect 3253 2253 3267 2267
rect 3293 2253 3307 2267
rect 3513 2253 3527 2267
rect 3733 2253 3747 2267
rect 4053 2253 4067 2267
rect 4253 2253 4267 2267
rect 4413 2253 4427 2267
rect 4573 2253 4587 2267
rect 4653 2253 4667 2267
rect 4813 2253 4827 2267
rect 4993 2253 5007 2267
rect 5033 2253 5047 2267
rect 5153 2253 5167 2267
rect 5193 2253 5207 2267
rect 5333 2253 5347 2267
rect 5373 2253 5387 2267
rect 5493 2253 5507 2267
rect 5533 2253 5547 2267
rect 5613 2253 5627 2267
rect 5733 2253 5747 2267
rect 5873 2253 5887 2267
rect 6033 2253 6047 2267
rect 6173 2253 6187 2267
rect 6373 2253 6387 2267
rect 4733 2233 4747 2247
rect 4773 2233 4787 2247
rect 373 2213 387 2227
rect 813 2213 827 2227
rect 3233 2213 3247 2227
rect 3313 2213 3327 2227
rect 3393 2213 3407 2227
rect 3533 2213 3547 2227
rect 3613 2213 3627 2227
rect 3693 2213 3707 2227
rect 3833 2213 3847 2227
rect 4013 2213 4027 2227
rect 4693 2213 4707 2227
rect 213 2193 227 2207
rect 433 2193 447 2207
rect 553 2193 567 2207
rect 593 2193 607 2207
rect 713 2193 727 2207
rect 753 2193 767 2207
rect 1013 2193 1027 2207
rect 1053 2193 1067 2207
rect 1153 2193 1167 2207
rect 1193 2193 1207 2207
rect 1293 2193 1307 2207
rect 1473 2193 1487 2207
rect 1513 2193 1527 2207
rect 1613 2193 1627 2207
rect 1653 2193 1667 2207
rect 1693 2193 1707 2207
rect 1833 2193 1847 2207
rect 2033 2193 2047 2207
rect 2073 2193 2087 2207
rect 2113 2193 2127 2207
rect 2333 2193 2347 2207
rect 2373 2193 2387 2207
rect 2413 2193 2427 2207
rect 2633 2193 2647 2207
rect 2693 2193 2707 2207
rect 2733 2193 2747 2207
rect 2833 2193 2847 2207
rect 2873 2193 2887 2207
rect 3013 2193 3027 2207
rect 3053 2193 3067 2207
rect 253 2173 267 2187
rect 3093 2173 3107 2187
rect 3393 2173 3407 2187
rect 3433 2173 3447 2187
rect 3533 2173 3547 2187
rect 3753 2193 3767 2207
rect 4193 2193 4207 2207
rect 4233 2193 4247 2207
rect 4333 2193 4347 2207
rect 4373 2193 4387 2207
rect 4513 2193 4527 2207
rect 4633 2193 4647 2207
rect 4793 2193 4807 2207
rect 4833 2193 4847 2207
rect 4933 2193 4947 2207
rect 4973 2193 4987 2207
rect 5093 2193 5107 2207
rect 5133 2193 5147 2207
rect 5253 2193 5267 2207
rect 5293 2193 5307 2207
rect 5393 2193 5407 2207
rect 5433 2193 5447 2207
rect 5673 2193 5687 2207
rect 5713 2193 5727 2207
rect 5853 2193 5867 2207
rect 5893 2193 5907 2207
rect 6013 2193 6027 2207
rect 6053 2193 6067 2207
rect 6153 2193 6167 2207
rect 6193 2193 6207 2207
rect 6353 2193 6367 2207
rect 6393 2193 6407 2207
rect 3673 2173 3687 2187
rect 3793 2173 3807 2187
rect 5333 2173 5347 2187
rect 5373 2173 5387 2187
rect 433 2153 447 2167
rect 553 2153 567 2167
rect 613 2153 627 2167
rect 713 2153 727 2167
rect 1133 2153 1147 2167
rect 1193 2153 1207 2167
rect 1313 2153 1327 2167
rect 1693 2153 1707 2167
rect 1813 2153 1827 2167
rect 1953 2153 1967 2167
rect 2133 2153 2147 2167
rect 2433 2153 2447 2167
rect 1033 2133 1047 2147
rect 1473 2133 1487 2147
rect 2113 2133 2127 2147
rect 2352 2133 2366 2147
rect 2374 2133 2388 2147
rect 2693 2153 2707 2167
rect 2913 2153 2927 2167
rect 2993 2153 3007 2167
rect 3353 2153 3367 2167
rect 3933 2153 3947 2167
rect 4353 2153 4367 2167
rect 4493 2153 4507 2167
rect 4973 2153 4987 2167
rect 5193 2153 5207 2167
rect 5533 2154 5547 2168
rect 6153 2153 6167 2167
rect 6293 2153 6307 2167
rect 6393 2153 6407 2167
rect 6513 2153 6527 2167
rect 2653 2133 2667 2147
rect 2853 2133 2867 2147
rect 2893 2133 2907 2147
rect 3013 2133 3027 2147
rect 3193 2133 3207 2147
rect 713 2113 727 2127
rect 913 2113 927 2127
rect 1433 2113 1447 2127
rect 2053 2113 2067 2127
rect 273 2093 287 2107
rect 573 2093 587 2107
rect 813 2093 827 2107
rect 893 2093 907 2107
rect 1693 2093 1707 2107
rect 2393 2113 2407 2127
rect 2613 2113 2627 2127
rect 2673 2113 2687 2127
rect 2833 2113 2847 2127
rect 2333 2093 2347 2107
rect 2733 2093 2747 2107
rect 2793 2093 2807 2107
rect 873 2073 887 2087
rect 972 2074 986 2088
rect 994 2073 1008 2087
rect 973 2052 987 2066
rect 1093 2053 1107 2067
rect 1653 2073 1667 2087
rect 2313 2073 2327 2087
rect 2353 2073 2367 2087
rect 2533 2073 2547 2087
rect 2633 2073 2647 2087
rect 2693 2073 2707 2087
rect 2773 2073 2787 2087
rect 2973 2093 2987 2107
rect 3053 2093 3067 2107
rect 3153 2113 3167 2127
rect 3233 2113 3247 2127
rect 3273 2133 3287 2147
rect 3513 2133 3527 2147
rect 4053 2133 4067 2147
rect 4193 2133 4207 2147
rect 4313 2133 4327 2147
rect 4553 2133 4567 2147
rect 4633 2133 4647 2147
rect 4833 2133 4847 2147
rect 4913 2133 4927 2147
rect 5093 2133 5107 2147
rect 3474 2113 3488 2127
rect 3553 2113 3567 2127
rect 3653 2113 3667 2127
rect 3753 2113 3767 2127
rect 3893 2113 3907 2127
rect 4033 2113 4047 2127
rect 4233 2113 4247 2127
rect 4492 2113 4506 2127
rect 4514 2113 4528 2127
rect 4613 2113 4627 2127
rect 4673 2113 4687 2127
rect 4733 2113 4747 2127
rect 4973 2113 4987 2127
rect 5013 2113 5027 2127
rect 5433 2133 5447 2147
rect 5493 2133 5507 2147
rect 5533 2132 5547 2146
rect 5893 2133 5907 2147
rect 5953 2133 5967 2147
rect 6013 2133 6027 2147
rect 5133 2113 5147 2127
rect 5693 2113 5707 2127
rect 6053 2113 6067 2127
rect 6173 2113 6187 2127
rect 6233 2113 6247 2127
rect 3533 2093 3547 2107
rect 4593 2093 4607 2107
rect 4713 2093 4727 2107
rect 4933 2093 4947 2107
rect 5253 2093 5267 2107
rect 5373 2093 5387 2107
rect 5593 2093 5607 2107
rect 3413 2073 3427 2087
rect 3453 2073 3467 2087
rect 3613 2073 3627 2087
rect 3713 2073 3727 2087
rect 3833 2073 3847 2087
rect 4173 2073 4187 2087
rect 4353 2073 4367 2087
rect 5013 2073 5027 2087
rect 5433 2073 5447 2087
rect 5513 2073 5527 2087
rect 5613 2073 5627 2087
rect 5733 2073 5747 2087
rect 2673 2053 2687 2067
rect 2754 2053 2768 2067
rect 2813 2053 2827 2067
rect 3013 2053 3027 2067
rect 3213 2053 3227 2067
rect 3493 2053 3507 2067
rect 3633 2053 3647 2067
rect 3773 2053 3787 2067
rect 4432 2053 4446 2067
rect 4454 2053 4468 2067
rect 4733 2053 4747 2067
rect 4813 2053 4827 2067
rect 5094 2053 5108 2067
rect 5193 2053 5207 2067
rect 5233 2053 5247 2067
rect 5413 2053 5427 2067
rect 5553 2053 5567 2067
rect 5713 2053 5727 2067
rect 5793 2053 5807 2067
rect 5853 2053 5867 2067
rect 113 2033 127 2047
rect 613 2033 627 2047
rect 1133 2033 1147 2047
rect 1253 2033 1267 2047
rect 2013 2033 2027 2047
rect 2053 2033 2067 2047
rect 433 2013 447 2027
rect 533 2013 547 2027
rect 673 2013 687 2027
rect 793 2013 807 2027
rect 933 2013 947 2027
rect 1172 2013 1186 2027
rect 1194 2013 1208 2027
rect 1293 2013 1307 2027
rect 1673 2013 1687 2027
rect 1813 2013 1827 2027
rect 1953 2013 1967 2027
rect 2033 2013 2047 2027
rect 2213 2013 2227 2027
rect 2293 2013 2307 2027
rect 2573 2013 2587 2027
rect 2693 2013 2707 2027
rect 2833 2033 2847 2047
rect 2913 2033 2927 2047
rect 3933 2033 3947 2047
rect 4113 2033 4127 2047
rect 4193 2033 4207 2047
rect 4513 2033 4527 2047
rect 4653 2033 4667 2047
rect 4774 2033 4788 2047
rect 4853 2033 4867 2047
rect 4953 2033 4967 2047
rect 5813 2033 5827 2047
rect 6353 2033 6367 2047
rect 6433 2033 6447 2047
rect 3313 2013 3327 2027
rect 3353 2013 3367 2027
rect 3393 2013 3407 2027
rect 3433 2013 3447 2027
rect 3513 2013 3527 2027
rect 4133 2013 4147 2027
rect 4253 2013 4267 2027
rect 4373 2013 4387 2027
rect 4413 2013 4427 2027
rect 4453 2013 4467 2027
rect 4493 2013 4507 2027
rect 4613 2013 4627 2027
rect 2173 1993 2187 2007
rect 2233 1993 2247 2007
rect 2473 1993 2487 2007
rect 3133 1993 3147 2007
rect 253 1973 267 1987
rect 293 1973 307 1987
rect 333 1973 347 1987
rect 533 1973 547 1987
rect 573 1973 587 1987
rect 853 1973 867 1987
rect 893 1973 907 1987
rect 1093 1973 1107 1987
rect 1133 1973 1147 1987
rect 1173 1973 1187 1987
rect 1253 1973 1267 1987
rect 1293 1973 1307 1987
rect 1473 1973 1487 1987
rect 1513 1973 1527 1987
rect 1813 1973 1827 1987
rect 1993 1973 2007 1987
rect 2033 1973 2047 1987
rect 2313 1973 2327 1987
rect 2353 1973 2367 1987
rect 2633 1973 2647 1987
rect 2673 1973 2687 1987
rect 2773 1973 2787 1987
rect 2813 1973 2827 1987
rect 3253 1993 3267 2007
rect 4853 1993 4867 2007
rect 4933 1993 4947 2007
rect 5113 2013 5127 2027
rect 5173 2013 5187 2027
rect 5293 2013 5307 2027
rect 5453 2013 5467 2027
rect 5653 2013 5667 2027
rect 5893 2010 5907 2024
rect 6113 2010 6127 2024
rect 6193 2013 6207 2027
rect 6273 2013 6287 2027
rect 6313 2013 6327 2027
rect 6413 2013 6427 2027
rect 5073 1993 5087 2007
rect 3313 1973 3327 1987
rect 3353 1973 3367 1987
rect 3453 1973 3467 1987
rect 3493 1973 3507 1987
rect 3613 1973 3627 1987
rect 3653 1973 3667 1987
rect 3753 1973 3767 1987
rect 3793 1973 3807 1987
rect 3913 1973 3927 1987
rect 3953 1973 3967 1987
rect 3993 1973 4007 1987
rect 4033 1973 4047 1987
rect 4073 1973 4087 1987
rect 4113 1973 4127 1987
rect 4433 1973 4447 1987
rect 4473 1973 4487 1987
rect 4513 1973 4527 1987
rect 4613 1973 4627 1987
rect 4653 1973 4667 1987
rect 4873 1973 4887 1987
rect 4953 1973 4967 1987
rect 5113 1973 5127 1987
rect 5153 1973 5167 1987
rect 5213 1973 5227 1987
rect 5293 1973 5307 1987
rect 5413 1973 5427 1987
rect 5453 1973 5467 1987
rect 5573 1973 5587 1987
rect 5613 1973 5627 1987
rect 5733 1973 5747 1987
rect 5773 1973 5787 1987
rect 5853 1973 5867 1987
rect 5893 1970 5907 1984
rect 6033 1973 6047 1987
rect 6073 1973 6087 1987
rect 6273 1973 6287 1987
rect 6413 1973 6427 1987
rect 6453 1973 6467 1987
rect 653 1953 667 1967
rect 1553 1953 1567 1967
rect 1893 1953 1907 1967
rect 2273 1953 2287 1967
rect 2433 1953 2447 1967
rect 2533 1953 2547 1967
rect 2953 1953 2967 1967
rect 3013 1953 3027 1967
rect 3093 1953 3107 1967
rect 3113 1953 3127 1967
rect 3193 1953 3207 1967
rect 4913 1953 4927 1967
rect 4993 1953 5007 1967
rect 1653 1933 1667 1947
rect 2753 1933 2767 1947
rect 3273 1934 3287 1948
rect 3733 1934 3747 1948
rect 4133 1933 4147 1947
rect 4793 1933 4807 1947
rect 5213 1933 5227 1947
rect 113 1913 127 1927
rect 273 1913 287 1927
rect 433 1913 447 1927
rect 593 1913 607 1927
rect 793 1913 807 1927
rect 1013 1913 1027 1927
rect 1153 1913 1167 1927
rect 1233 1913 1247 1927
rect 1273 1913 1287 1927
rect 1413 1913 1427 1927
rect 1493 1913 1507 1927
rect 233 1893 247 1907
rect 273 1873 287 1887
rect 433 1873 447 1887
rect 713 1893 727 1907
rect 753 1893 767 1907
rect 1773 1912 1787 1926
rect 1833 1912 1847 1926
rect 2013 1913 2027 1927
rect 2073 1913 2087 1927
rect 2293 1913 2307 1927
rect 2453 1913 2467 1927
rect 2493 1913 2507 1927
rect 2613 1913 2627 1927
rect 2693 1913 2707 1927
rect 2813 1913 2827 1927
rect 2993 1913 3007 1927
rect 3273 1912 3287 1926
rect 3593 1913 3607 1927
rect 1453 1893 1467 1907
rect 1593 1893 1607 1907
rect 1633 1893 1647 1907
rect 2153 1893 2167 1907
rect 2193 1893 2207 1907
rect 3133 1893 3147 1907
rect 3173 1893 3187 1907
rect 3213 1893 3227 1907
rect 3293 1893 3307 1907
rect 1493 1873 1507 1887
rect 2013 1873 2027 1887
rect 313 1853 327 1867
rect 473 1853 487 1867
rect 753 1853 767 1867
rect 1073 1853 1087 1867
rect 1593 1853 1607 1867
rect 1833 1853 1847 1867
rect 2293 1853 2307 1867
rect 2773 1854 2787 1868
rect 3233 1873 3247 1887
rect 3373 1873 3387 1887
rect 3733 1912 3747 1926
rect 3773 1913 3787 1927
rect 3893 1913 3907 1927
rect 4013 1913 4027 1927
rect 4173 1913 4187 1927
rect 4373 1913 4387 1927
rect 4453 1913 4467 1927
rect 4633 1913 4647 1927
rect 4693 1913 4707 1927
rect 4833 1913 4847 1927
rect 5133 1913 5147 1927
rect 5193 1913 5207 1927
rect 5273 1913 5287 1927
rect 5413 1913 5427 1927
rect 5513 1913 5527 1927
rect 5593 1913 5607 1927
rect 5653 1913 5667 1927
rect 5753 1913 5767 1927
rect 5873 1913 5887 1927
rect 5953 1913 5967 1927
rect 6093 1913 6107 1927
rect 6253 1912 6267 1926
rect 6313 1912 6327 1926
rect 6373 1913 6387 1927
rect 4213 1893 4227 1907
rect 4293 1893 4307 1907
rect 4933 1893 4947 1907
rect 4973 1893 4987 1907
rect 5913 1893 5927 1907
rect 3593 1873 3607 1887
rect 3833 1873 3847 1887
rect 3913 1873 3927 1887
rect 4073 1873 4087 1887
rect 4513 1873 4527 1887
rect 4573 1873 4587 1887
rect 4613 1873 4627 1887
rect 4833 1873 4847 1887
rect 5153 1873 5167 1887
rect 5233 1873 5247 1887
rect 5273 1873 5287 1887
rect 5453 1873 5467 1887
rect 5733 1873 5747 1887
rect 6133 1873 6147 1887
rect 6253 1873 6267 1887
rect 6413 1873 6427 1887
rect 6493 1873 6507 1887
rect 2853 1853 2867 1867
rect 2993 1853 3007 1867
rect 3133 1853 3147 1867
rect 3193 1853 3207 1867
rect 3413 1853 3427 1867
rect 3493 1853 3507 1867
rect 3633 1853 3647 1867
rect 3773 1853 3787 1867
rect 3813 1853 3827 1867
rect 4173 1853 4187 1867
rect 4292 1853 4306 1867
rect 4633 1853 4647 1867
rect 1273 1833 1287 1847
rect 1733 1833 1747 1847
rect 1773 1833 1787 1847
rect 1953 1833 1967 1847
rect 2013 1833 2027 1847
rect 2153 1833 2167 1847
rect 2533 1833 2547 1847
rect 2713 1833 2727 1847
rect 2773 1832 2787 1846
rect 2913 1833 2927 1847
rect 3093 1833 3107 1847
rect 3333 1833 3347 1847
rect 3513 1833 3527 1847
rect 233 1813 247 1827
rect 332 1813 346 1827
rect 354 1813 368 1827
rect 493 1813 507 1827
rect 613 1813 627 1827
rect 793 1813 807 1827
rect 933 1813 947 1827
rect 1213 1813 1227 1827
rect 1653 1813 1667 1827
rect 2173 1813 2187 1827
rect 2393 1813 2407 1827
rect 3033 1813 3047 1827
rect 3113 1813 3127 1827
rect 3813 1813 3827 1827
rect 213 1793 227 1807
rect 393 1793 407 1807
rect 1333 1793 1347 1807
rect 1533 1793 1547 1807
rect 1733 1793 1747 1807
rect 1913 1793 1927 1807
rect 2093 1793 2107 1807
rect 2953 1793 2967 1807
rect 3013 1793 3027 1807
rect 3053 1793 3067 1807
rect 3093 1793 3107 1807
rect 3134 1793 3148 1807
rect 3193 1793 3207 1807
rect 3233 1793 3247 1807
rect 3373 1793 3387 1807
rect 113 1773 127 1787
rect 193 1773 207 1787
rect 533 1773 547 1787
rect 653 1773 667 1787
rect 813 1773 827 1787
rect 1393 1773 1407 1787
rect 353 1753 367 1767
rect 393 1753 407 1767
rect 1273 1753 1287 1767
rect 1633 1773 1647 1787
rect 1692 1773 1706 1787
rect 1773 1773 1787 1787
rect 1813 1773 1827 1787
rect 1593 1753 1607 1767
rect 2033 1773 2047 1787
rect 2192 1773 2206 1787
rect 2233 1773 2247 1787
rect 2373 1773 2387 1787
rect 2573 1773 2587 1787
rect 2692 1773 2706 1787
rect 2714 1773 2728 1787
rect 2593 1753 2607 1767
rect 2753 1753 2767 1767
rect 3533 1793 3547 1807
rect 3673 1793 3687 1807
rect 3933 1833 3947 1847
rect 4273 1833 4287 1847
rect 4333 1833 4347 1847
rect 4933 1853 4947 1867
rect 5093 1853 5107 1867
rect 5253 1853 5267 1867
rect 5593 1853 5607 1867
rect 5793 1853 5807 1867
rect 6033 1853 6047 1867
rect 6313 1853 6327 1867
rect 4693 1833 4707 1847
rect 4833 1833 4847 1847
rect 4873 1833 4887 1847
rect 4973 1833 4987 1847
rect 5013 1833 5027 1847
rect 5313 1833 5327 1847
rect 5453 1833 5467 1847
rect 6093 1833 6107 1847
rect 6193 1833 6207 1847
rect 6293 1833 6307 1847
rect 6453 1834 6467 1848
rect 3893 1813 3907 1827
rect 4033 1813 4047 1827
rect 4073 1813 4087 1827
rect 4213 1813 4227 1827
rect 4473 1813 4487 1827
rect 4773 1813 4787 1827
rect 5373 1813 5387 1827
rect 5573 1813 5587 1827
rect 5753 1813 5767 1827
rect 6153 1813 6167 1827
rect 6453 1812 6467 1826
rect 3873 1793 3887 1807
rect 4333 1793 4347 1807
rect 4693 1793 4707 1807
rect 4793 1793 4807 1807
rect 4833 1793 4847 1807
rect 5013 1793 5027 1807
rect 5133 1793 5147 1807
rect 5193 1793 5207 1807
rect 5353 1793 5367 1807
rect 5493 1793 5507 1807
rect 5793 1793 5807 1807
rect 6473 1793 6487 1807
rect 3473 1773 3487 1787
rect 3693 1773 3707 1787
rect 3053 1753 3067 1767
rect 3093 1753 3107 1767
rect 3433 1753 3447 1767
rect 3633 1753 3647 1767
rect 3673 1753 3687 1767
rect 3933 1773 3947 1787
rect 4373 1773 4387 1787
rect 4433 1773 4447 1787
rect 4593 1773 4607 1787
rect 3913 1753 3927 1767
rect 4113 1753 4127 1767
rect 4153 1753 4167 1767
rect 4413 1753 4427 1767
rect 4453 1753 4467 1767
rect 4753 1773 4767 1787
rect 113 1733 127 1747
rect 313 1733 327 1747
rect 573 1733 587 1747
rect 653 1733 667 1747
rect 813 1733 827 1747
rect 913 1733 927 1747
rect 1133 1733 1147 1747
rect 1313 1733 1327 1747
rect 1413 1733 1427 1747
rect 1493 1733 1507 1747
rect 1633 1733 1647 1747
rect 1733 1733 1747 1747
rect 1813 1733 1827 1747
rect 1993 1733 2007 1747
rect 2033 1733 2047 1747
rect 2173 1733 2187 1747
rect 2293 1733 2307 1747
rect 2493 1733 2507 1747
rect 2553 1733 2567 1747
rect 3173 1733 3187 1747
rect 3313 1733 3327 1747
rect 3373 1733 3387 1747
rect 3513 1733 3527 1747
rect 4073 1733 4087 1747
rect 4373 1733 4387 1747
rect 4973 1773 4987 1787
rect 5053 1773 5067 1787
rect 5093 1773 5107 1787
rect 5473 1773 5487 1787
rect 5573 1773 5587 1787
rect 5733 1773 5747 1787
rect 5613 1753 5627 1767
rect 5653 1753 5667 1767
rect 6233 1773 6247 1787
rect 6313 1773 6327 1787
rect 6413 1773 6427 1787
rect 6453 1753 6467 1767
rect 4473 1733 4487 1747
rect 4554 1733 4568 1747
rect 4693 1733 4707 1747
rect 4793 1733 4807 1747
rect 4973 1733 4987 1747
rect 5013 1733 5027 1747
rect 5133 1733 5147 1747
rect 5173 1733 5187 1747
rect 5493 1733 5507 1747
rect 5533 1733 5547 1747
rect 5753 1733 5767 1747
rect 5833 1733 5847 1747
rect 5973 1733 5987 1747
rect 6153 1733 6167 1747
rect 6413 1733 6427 1747
rect 193 1713 207 1727
rect 2653 1713 2667 1727
rect 2713 1713 2727 1727
rect 2853 1713 2867 1727
rect 3353 1713 3367 1727
rect 3393 1713 3407 1727
rect 453 1693 467 1707
rect 613 1693 627 1707
rect 733 1693 747 1707
rect 893 1693 907 1707
rect 1533 1693 1547 1707
rect 1573 1693 1587 1707
rect 2013 1693 2027 1707
rect 2053 1693 2067 1707
rect 2173 1693 2187 1707
rect 2233 1694 2247 1708
rect 3053 1693 3067 1707
rect 3193 1693 3207 1707
rect 3613 1693 3627 1707
rect 3693 1693 3707 1707
rect 4033 1693 4047 1707
rect 4093 1693 4107 1707
rect 4173 1693 4187 1707
rect 5453 1693 5467 1707
rect 5573 1693 5587 1707
rect 73 1673 87 1687
rect 213 1673 227 1687
rect 253 1673 267 1687
rect 493 1673 507 1687
rect 533 1673 547 1687
rect 793 1673 807 1687
rect 973 1673 987 1687
rect 1013 1673 1027 1687
rect 1213 1673 1227 1687
rect 1253 1673 1267 1687
rect 1293 1673 1307 1687
rect 1433 1673 1447 1687
rect 1473 1673 1487 1687
rect 1553 1673 1567 1687
rect 1613 1673 1627 1687
rect 1753 1673 1767 1687
rect 1793 1673 1807 1687
rect 1833 1673 1847 1687
rect 1893 1673 1907 1687
rect 1933 1673 1947 1687
rect 1973 1673 1987 1687
rect 2093 1673 2107 1687
rect 2133 1673 2147 1687
rect 2233 1672 2247 1686
rect 2273 1673 2287 1687
rect 2313 1673 2327 1687
rect 2413 1673 2427 1687
rect 2453 1673 2467 1687
rect 2533 1673 2547 1687
rect 2573 1673 2587 1687
rect 2733 1673 2747 1687
rect 2773 1673 2787 1687
rect 2893 1673 2907 1687
rect 2933 1673 2947 1687
rect 3413 1673 3427 1687
rect 3453 1673 3467 1687
rect 3493 1673 3507 1687
rect 3653 1673 3667 1687
rect 3813 1673 3827 1687
rect 3853 1673 3867 1687
rect 3953 1673 3967 1687
rect 3993 1673 4007 1687
rect 1313 1653 1327 1667
rect 1493 1653 1507 1667
rect 1573 1653 1587 1667
rect 2613 1653 2627 1667
rect 2693 1653 2707 1667
rect 3073 1653 3087 1667
rect 3173 1653 3187 1667
rect 3533 1653 3547 1667
rect 3733 1653 3747 1667
rect 253 1633 267 1647
rect 353 1633 367 1647
rect 1133 1633 1147 1647
rect 1273 1633 1287 1647
rect 1333 1633 1347 1647
rect 1433 1633 1447 1647
rect 1473 1633 1487 1647
rect 1713 1633 1727 1647
rect 1793 1633 1807 1647
rect 2194 1633 2208 1647
rect 2813 1633 2827 1647
rect 2893 1633 2907 1647
rect 2953 1633 2967 1647
rect 3113 1633 3127 1647
rect 3253 1633 3267 1647
rect 3312 1633 3326 1647
rect 3334 1633 3348 1647
rect 3493 1633 3507 1647
rect 3573 1633 3587 1647
rect 1493 1613 1507 1627
rect 2053 1613 2067 1627
rect 2173 1613 2187 1627
rect 2653 1614 2667 1628
rect 2693 1613 2707 1627
rect 2733 1613 2747 1627
rect 2873 1613 2887 1627
rect 2913 1613 2927 1627
rect 3193 1613 3207 1627
rect 3513 1613 3527 1627
rect 3613 1614 3627 1628
rect 3693 1633 3707 1647
rect 3853 1633 3867 1647
rect 3893 1633 3907 1647
rect 3933 1634 3947 1648
rect 4053 1653 4067 1667
rect 4093 1653 4107 1667
rect 4313 1673 4327 1687
rect 4353 1673 4367 1687
rect 4453 1673 4467 1687
rect 4493 1673 4507 1687
rect 4633 1673 4647 1687
rect 4673 1673 4687 1687
rect 4813 1673 4827 1687
rect 4853 1673 4867 1687
rect 4953 1673 4967 1687
rect 4993 1673 5007 1687
rect 5113 1673 5127 1687
rect 5153 1673 5167 1687
rect 5313 1673 5327 1687
rect 5353 1673 5367 1687
rect 5513 1673 5527 1687
rect 5773 1673 5787 1687
rect 5873 1673 5887 1687
rect 5913 1673 5927 1687
rect 5953 1673 5967 1687
rect 6053 1673 6067 1687
rect 6093 1673 6107 1687
rect 6133 1673 6147 1687
rect 6273 1673 6287 1687
rect 6313 1673 6327 1687
rect 6393 1673 6407 1687
rect 6433 1673 6447 1687
rect 4373 1653 4387 1667
rect 4333 1633 4347 1647
rect 4633 1634 4647 1648
rect 4753 1633 4767 1647
rect 4953 1633 4967 1647
rect 5053 1633 5067 1647
rect 5112 1633 5126 1647
rect 5134 1633 5148 1647
rect 5173 1633 5187 1647
rect 5993 1633 6007 1647
rect 6093 1633 6107 1647
rect 6133 1633 6147 1647
rect 6353 1633 6367 1647
rect 6413 1633 6427 1647
rect 6453 1633 6467 1647
rect 3873 1613 3887 1627
rect 3933 1612 3947 1626
rect 3973 1613 3987 1627
rect 4012 1613 4026 1627
rect 4034 1613 4048 1627
rect 4133 1613 4147 1627
rect 4253 1613 4267 1627
rect 4453 1613 4467 1627
rect 4513 1613 4527 1627
rect 1293 1593 1307 1607
rect 1553 1593 1567 1607
rect 1593 1593 1607 1607
rect 1633 1593 1647 1607
rect 1693 1593 1707 1607
rect 1933 1593 1947 1607
rect 2073 1593 2087 1607
rect 2133 1593 2147 1607
rect 2313 1593 2327 1607
rect 2453 1593 2467 1607
rect 2493 1593 2507 1607
rect 973 1573 987 1587
rect 1573 1573 1587 1587
rect 1713 1573 1727 1587
rect 2193 1573 2207 1587
rect 2233 1573 2247 1587
rect 2332 1573 2346 1587
rect 2354 1573 2368 1587
rect 2553 1573 2567 1587
rect 2654 1592 2668 1606
rect 2713 1573 2727 1587
rect 2813 1573 2827 1587
rect 3333 1593 3347 1607
rect 3393 1593 3407 1607
rect 3553 1593 3567 1607
rect 3612 1592 3626 1606
rect 3634 1593 3648 1607
rect 3773 1593 3787 1607
rect 3953 1593 3967 1607
rect 4633 1612 4647 1626
rect 4713 1613 4727 1627
rect 4993 1613 5007 1627
rect 5153 1613 5167 1627
rect 5193 1613 5207 1627
rect 5393 1613 5407 1627
rect 4153 1593 4167 1607
rect 4593 1593 4607 1607
rect 4853 1593 4867 1607
rect 4953 1593 4967 1607
rect 5653 1613 5667 1627
rect 5533 1593 5547 1607
rect 6193 1593 6207 1607
rect 6353 1593 6367 1607
rect 6473 1593 6487 1607
rect 3073 1573 3087 1587
rect 3133 1573 3147 1587
rect 3173 1573 3187 1587
rect 3453 1573 3467 1587
rect 3513 1573 3527 1587
rect 3733 1573 3747 1587
rect 73 1553 87 1567
rect 273 1553 287 1567
rect 1013 1553 1027 1567
rect 1533 1553 1547 1567
rect 1673 1553 1687 1567
rect 192 1533 206 1547
rect 1593 1533 1607 1547
rect 1633 1534 1647 1548
rect 1793 1553 1807 1567
rect 2053 1553 2067 1567
rect 2173 1533 2187 1547
rect 2273 1553 2287 1567
rect 2413 1553 2427 1567
rect 5833 1573 5847 1587
rect 6213 1573 6227 1587
rect 6293 1573 6307 1587
rect 3773 1553 3787 1567
rect 3993 1553 4007 1567
rect 4173 1553 4187 1567
rect 4273 1553 4287 1567
rect 4353 1553 4367 1567
rect 4673 1553 4687 1567
rect 4813 1553 4827 1567
rect 5033 1553 5047 1567
rect 5133 1553 5147 1567
rect 2773 1533 2787 1547
rect 3033 1533 3047 1547
rect 3353 1533 3367 1547
rect 3493 1533 3507 1547
rect 3593 1533 3607 1547
rect 3653 1533 3667 1547
rect 3733 1533 3747 1547
rect 3913 1533 3927 1547
rect 4153 1533 4167 1547
rect 4313 1533 4327 1547
rect 4413 1533 4427 1547
rect 4453 1533 4467 1547
rect 4552 1533 4566 1547
rect 4574 1533 4588 1547
rect 4634 1533 4648 1547
rect 5193 1553 5207 1567
rect 5233 1553 5247 1567
rect 5313 1553 5327 1567
rect 5213 1533 5227 1547
rect 5413 1533 5427 1547
rect 5713 1533 5727 1547
rect 6233 1533 6247 1547
rect 6273 1533 6287 1547
rect 6393 1533 6407 1547
rect 214 1513 228 1527
rect 573 1513 587 1527
rect 953 1513 967 1527
rect 1633 1512 1647 1526
rect 173 1493 187 1507
rect 453 1493 467 1507
rect 612 1493 626 1507
rect 634 1493 648 1507
rect 793 1493 807 1507
rect 913 1493 927 1507
rect 1033 1493 1047 1507
rect 1073 1493 1087 1507
rect 1773 1493 1787 1507
rect 1853 1493 1867 1507
rect 2213 1513 2227 1527
rect 2393 1513 2407 1527
rect 2473 1513 2487 1527
rect 2893 1513 2907 1527
rect 3093 1513 3107 1527
rect 3133 1513 3147 1527
rect 3253 1513 3267 1527
rect 3553 1513 3567 1527
rect 3674 1513 3688 1527
rect 4193 1513 4207 1527
rect 4253 1513 4267 1527
rect 4393 1513 4407 1527
rect 4513 1513 4527 1527
rect 4733 1513 4747 1527
rect 5173 1513 5187 1527
rect 5353 1513 5367 1527
rect 5533 1513 5547 1527
rect 6293 1513 6307 1527
rect 6493 1513 6507 1527
rect 1493 1473 1507 1487
rect 73 1453 87 1467
rect 113 1453 127 1467
rect 153 1453 167 1467
rect 193 1453 207 1467
rect 233 1453 247 1467
rect 273 1453 287 1467
rect 433 1453 447 1467
rect 473 1453 487 1467
rect 573 1453 587 1467
rect 613 1453 627 1467
rect 713 1453 727 1467
rect 753 1453 767 1467
rect 793 1453 807 1467
rect 933 1453 947 1467
rect 973 1453 987 1467
rect 1013 1453 1027 1467
rect 1193 1453 1207 1467
rect 1233 1453 1247 1467
rect 1333 1453 1347 1467
rect 1373 1453 1387 1467
rect 1593 1453 1607 1467
rect 1633 1453 1647 1467
rect 1773 1453 1787 1467
rect 1813 1453 1827 1467
rect 1933 1453 1947 1467
rect 2073 1453 2087 1467
rect 2213 1453 2227 1467
rect 2253 1453 2267 1467
rect 2393 1453 2407 1467
rect 2433 1453 2447 1467
rect 2873 1493 2887 1507
rect 3293 1493 3307 1507
rect 3692 1493 3706 1507
rect 3714 1493 3728 1507
rect 3913 1493 3927 1507
rect 3973 1493 3987 1507
rect 4073 1493 4087 1507
rect 4293 1493 4307 1507
rect 4753 1493 4767 1507
rect 4793 1493 4807 1507
rect 5153 1493 5167 1507
rect 5193 1493 5207 1507
rect 5253 1493 5267 1507
rect 5613 1493 5627 1507
rect 5693 1493 5707 1507
rect 6253 1493 6267 1507
rect 6393 1493 6407 1507
rect 3093 1453 3107 1467
rect 3133 1453 3147 1467
rect 3293 1453 3307 1467
rect 3333 1453 3347 1467
rect 3553 1453 3567 1467
rect 3693 1453 3707 1467
rect 3733 1453 3747 1467
rect 3873 1453 3887 1467
rect 3913 1453 3927 1467
rect 4073 1453 4087 1467
rect 4113 1453 4127 1467
rect 4153 1453 4167 1467
rect 4193 1453 4207 1467
rect 4233 1453 4247 1467
rect 4273 1453 4287 1467
rect 4353 1453 4367 1467
rect 4393 1453 4407 1467
rect 4433 1453 4447 1467
rect 4513 1453 4527 1467
rect 4553 1453 4567 1467
rect 4713 1453 4727 1467
rect 4753 1453 4767 1467
rect 4873 1453 4887 1467
rect 4913 1453 4927 1467
rect 5053 1453 5067 1467
rect 5093 1453 5107 1467
rect 5193 1453 5207 1467
rect 5233 1453 5247 1467
rect 5353 1453 5367 1467
rect 5393 1453 5407 1467
rect 5533 1453 5547 1467
rect 5573 1453 5587 1467
rect 5633 1453 5647 1467
rect 5673 1453 5687 1467
rect 5833 1473 5847 1487
rect 5973 1473 5987 1487
rect 6313 1473 6327 1487
rect 6513 1473 6527 1487
rect 6013 1453 6027 1467
rect 6053 1453 6067 1467
rect 6133 1453 6147 1467
rect 6173 1453 6187 1467
rect 6353 1453 6367 1467
rect 2033 1433 2047 1447
rect 2113 1433 2127 1447
rect 2493 1433 2507 1447
rect 2593 1433 2607 1447
rect 2893 1433 2907 1447
rect 3833 1433 3847 1447
rect 4593 1433 4607 1447
rect 4673 1433 4687 1447
rect 4973 1433 4987 1447
rect 5013 1433 5027 1447
rect 5833 1433 5847 1447
rect 5933 1433 5947 1447
rect 6313 1433 6327 1447
rect 6393 1433 6407 1447
rect 3353 1413 3367 1427
rect 3673 1413 3687 1427
rect 5313 1413 5327 1427
rect 5653 1413 5667 1427
rect 93 1393 107 1407
rect 253 1393 267 1407
rect 352 1393 366 1407
rect 453 1393 467 1407
rect 493 1393 507 1407
rect 633 1393 647 1407
rect 733 1393 747 1407
rect 813 1393 827 1407
rect 953 1393 967 1407
rect 1053 1393 1067 1407
rect 1253 1393 1267 1407
rect 1293 1393 1307 1407
rect 1433 1393 1447 1407
rect 1473 1393 1487 1407
rect 1513 1393 1527 1407
rect 1733 1393 1747 1407
rect 1793 1393 1807 1407
rect 1853 1393 1867 1407
rect 1893 1393 1907 1407
rect 2133 1393 2147 1407
rect 2233 1393 2247 1407
rect 2333 1393 2347 1407
rect 2513 1393 2527 1407
rect 2553 1393 2567 1407
rect 2873 1393 2887 1407
rect 3113 1393 3127 1407
rect 3273 1393 3287 1407
rect 3373 1393 3387 1407
rect 3493 1393 3507 1407
rect 3573 1393 3587 1407
rect 3713 1393 3727 1407
rect 3813 1393 3827 1407
rect 3853 1393 3867 1407
rect 4093 1393 4107 1407
rect 4213 1393 4227 1407
rect 4273 1393 4287 1407
rect 4413 1393 4427 1407
rect 4533 1393 4547 1407
rect 4693 1393 4707 1407
rect 4813 1393 4827 1407
rect 4893 1393 4907 1407
rect 5033 1393 5047 1407
rect 5153 1393 5167 1407
rect 5213 1393 5227 1407
rect 5293 1393 5307 1407
rect 5373 1393 5387 1407
rect 5493 1393 5507 1407
rect 5693 1393 5707 1407
rect 5873 1393 5887 1407
rect 5973 1393 5987 1407
rect 6153 1393 6167 1407
rect 6293 1393 6307 1407
rect 6413 1393 6427 1407
rect 6493 1393 6507 1407
rect 133 1373 147 1387
rect 253 1353 267 1367
rect 313 1353 327 1367
rect 593 1373 607 1387
rect 773 1373 787 1387
rect 2053 1373 2067 1387
rect 2093 1373 2107 1387
rect 2593 1373 2607 1387
rect 2653 1373 2667 1387
rect 2673 1373 2687 1387
rect 2713 1373 2727 1387
rect 2953 1373 2967 1387
rect 2993 1373 3007 1387
rect 3153 1373 3167 1387
rect 3313 1373 3327 1387
rect 3613 1373 3627 1387
rect 3693 1373 3707 1387
rect 913 1353 927 1367
rect 1013 1353 1027 1367
rect 1233 1353 1247 1367
rect 1333 1353 1347 1367
rect 1813 1353 1827 1367
rect 2013 1353 2027 1367
rect 2253 1353 2267 1367
rect 2553 1353 2567 1367
rect 2613 1353 2627 1367
rect 2813 1353 2827 1367
rect 2873 1353 2887 1367
rect 3373 1353 3387 1367
rect 3493 1353 3507 1367
rect 3713 1353 3727 1367
rect 4053 1373 4067 1387
rect 4113 1373 4127 1387
rect 4173 1373 4187 1387
rect 4373 1373 4387 1387
rect 4733 1373 4747 1387
rect 5312 1373 5326 1387
rect 5353 1373 5367 1387
rect 6333 1373 6347 1387
rect 6373 1373 6387 1387
rect 4593 1353 4607 1367
rect 4713 1353 4727 1367
rect 4773 1353 4787 1367
rect 4893 1353 4907 1367
rect 4973 1353 4987 1367
rect 5153 1353 5167 1367
rect 5373 1353 5387 1367
rect 172 1333 186 1347
rect 213 1333 227 1347
rect 353 1333 367 1347
rect 453 1333 467 1347
rect 1373 1333 1387 1347
rect 1573 1333 1587 1347
rect 1693 1333 1707 1347
rect 1893 1333 1907 1347
rect 2093 1333 2107 1347
rect 2653 1333 2667 1347
rect 2693 1333 2707 1347
rect 2733 1333 2747 1347
rect 2773 1333 2787 1347
rect 2913 1333 2927 1347
rect 2953 1333 2967 1347
rect 3153 1333 3167 1347
rect 113 1313 127 1327
rect 413 1313 427 1327
rect 1173 1313 1187 1327
rect 1293 1313 1307 1327
rect 1433 1313 1447 1327
rect 1533 1313 1547 1327
rect 2013 1313 2027 1327
rect 2193 1313 2207 1327
rect 2293 1313 2307 1327
rect 2433 1313 2447 1327
rect 3053 1314 3067 1328
rect 3312 1334 3326 1348
rect 3334 1333 3348 1347
rect 3413 1333 3427 1347
rect 3633 1333 3647 1347
rect 3753 1333 3767 1347
rect 4053 1333 4067 1347
rect 4413 1333 4427 1347
rect 4473 1333 4487 1347
rect 4513 1333 4527 1347
rect 4573 1333 4587 1347
rect 4693 1333 4707 1347
rect 4873 1333 4887 1347
rect 4913 1333 4927 1347
rect 5013 1333 5027 1347
rect 5233 1333 5247 1347
rect 5513 1353 5527 1367
rect 5873 1353 5887 1367
rect 6053 1353 6067 1367
rect 5533 1333 5547 1347
rect 5653 1333 5667 1347
rect 5793 1333 5807 1347
rect 6173 1333 6187 1347
rect 6373 1333 6387 1347
rect 133 1293 147 1307
rect 453 1293 467 1307
rect 1793 1293 1807 1307
rect 2053 1293 2067 1307
rect 2133 1293 2147 1307
rect 2893 1293 2907 1307
rect 2953 1293 2967 1307
rect 2993 1293 3007 1307
rect 3053 1292 3067 1306
rect 3213 1313 3227 1327
rect 3273 1313 3287 1327
rect 3313 1312 3327 1326
rect 4213 1313 4227 1327
rect 4433 1313 4447 1327
rect 4813 1313 4827 1327
rect 4853 1313 4867 1327
rect 5093 1313 5107 1327
rect 5293 1313 5307 1327
rect 5893 1313 5907 1327
rect 5993 1313 6007 1327
rect 6133 1313 6147 1327
rect 6333 1313 6347 1327
rect 6493 1313 6507 1327
rect 4013 1293 4027 1307
rect 4073 1293 4087 1307
rect 4173 1293 4187 1307
rect 4333 1293 4347 1307
rect 4373 1293 4387 1307
rect 4793 1293 4807 1307
rect 5033 1293 5047 1307
rect 5173 1293 5187 1307
rect 5733 1293 5747 1307
rect 5933 1293 5947 1307
rect 6173 1293 6187 1307
rect 6233 1293 6247 1307
rect 6413 1293 6427 1307
rect 213 1273 227 1287
rect 393 1273 407 1287
rect 473 1273 487 1287
rect 1133 1273 1147 1287
rect 1313 1273 1327 1287
rect 1353 1273 1367 1287
rect 1393 1273 1407 1287
rect 1493 1273 1507 1287
rect 1553 1273 1567 1287
rect 1613 1273 1627 1287
rect 533 1253 547 1267
rect 733 1253 747 1267
rect 773 1253 787 1267
rect 1233 1253 1247 1267
rect 1593 1253 1607 1267
rect 2233 1273 2247 1287
rect 2273 1273 2287 1287
rect 2393 1273 2407 1287
rect 2833 1273 2847 1287
rect 3213 1273 3227 1287
rect 3673 1273 3687 1287
rect 3753 1273 3767 1287
rect 3893 1273 3907 1287
rect 3933 1273 3947 1287
rect 4233 1273 4247 1287
rect 4273 1273 4287 1287
rect 4733 1273 4747 1287
rect 4913 1273 4927 1287
rect 4972 1273 4986 1287
rect 4994 1273 5008 1287
rect 5373 1273 5387 1287
rect 5494 1273 5508 1287
rect 5833 1273 5847 1287
rect 6153 1273 6167 1287
rect 2373 1253 2387 1267
rect 2773 1253 2787 1267
rect 2873 1253 2887 1267
rect 3073 1253 3087 1267
rect 3113 1253 3127 1267
rect 3293 1253 3307 1267
rect 3333 1253 3347 1267
rect 3393 1253 3407 1267
rect 3553 1253 3567 1267
rect 1493 1233 1507 1247
rect 1533 1233 1547 1247
rect 2073 1233 2087 1247
rect 2153 1233 2167 1247
rect 2193 1233 2207 1247
rect 3713 1253 3727 1267
rect 3813 1253 3827 1267
rect 3993 1253 4007 1267
rect 4113 1253 4127 1267
rect 4193 1253 4207 1267
rect 4253 1253 4267 1267
rect 4293 1253 4307 1267
rect 4153 1233 4167 1247
rect 4233 1233 4247 1247
rect 4433 1233 4447 1247
rect 4473 1233 4487 1247
rect 4713 1233 4727 1247
rect 4753 1233 4767 1247
rect 4953 1253 4967 1267
rect 5073 1253 5087 1267
rect 5133 1253 5147 1267
rect 5353 1253 5367 1267
rect 5473 1253 5487 1267
rect 5753 1253 5767 1267
rect 5993 1253 6007 1267
rect 6433 1273 6447 1287
rect 6253 1253 6267 1267
rect 6193 1233 6207 1247
rect 113 1213 127 1227
rect 173 1213 187 1227
rect 213 1213 227 1227
rect 253 1213 267 1227
rect 393 1213 407 1227
rect 473 1213 487 1227
rect 573 1213 587 1227
rect 733 1213 747 1227
rect 1013 1213 1027 1227
rect 1133 1213 1147 1227
rect 1213 1213 1227 1227
rect 1293 1213 1307 1227
rect 1653 1213 1667 1227
rect 1733 1213 1747 1227
rect 1813 1213 1827 1227
rect 1893 1213 1907 1227
rect 2013 1213 2027 1227
rect 2293 1213 2307 1227
rect 2453 1213 2467 1227
rect 2533 1213 2547 1227
rect 2712 1213 2726 1227
rect 2812 1213 2826 1227
rect 3213 1213 3227 1227
rect 3313 1213 3327 1227
rect 3373 1213 3387 1227
rect 3513 1213 3527 1227
rect 3593 1213 3607 1227
rect 3673 1213 3687 1227
rect 3753 1213 3767 1227
rect 3913 1213 3927 1227
rect 3953 1213 3967 1227
rect 4113 1213 4127 1227
rect 4253 1213 4267 1227
rect 4334 1213 4348 1227
rect 4393 1213 4407 1227
rect 4513 1213 4527 1227
rect 4593 1213 4607 1227
rect 4873 1213 4887 1227
rect 4993 1213 5007 1227
rect 5033 1213 5047 1227
rect 5093 1213 5107 1227
rect 5173 1213 5187 1227
rect 5333 1213 5347 1227
rect 5373 1213 5387 1227
rect 5533 1213 5547 1227
rect 5733 1213 5747 1227
rect 5813 1213 5827 1227
rect 5913 1213 5927 1227
rect 6013 1213 6027 1227
rect 6233 1213 6247 1227
rect 6313 1213 6327 1227
rect 2733 1193 2747 1207
rect 633 1173 647 1187
rect 773 1173 787 1187
rect 1593 1173 1607 1187
rect 2053 1173 2067 1187
rect 2213 1173 2227 1187
rect 2393 1173 2407 1187
rect 4073 1173 4087 1187
rect 4313 1173 4327 1187
rect 4373 1173 4387 1187
rect 4413 1173 4427 1187
rect 4493 1173 4507 1187
rect 4813 1173 4827 1187
rect 113 1153 127 1167
rect 153 1153 167 1167
rect 273 1153 287 1167
rect 313 1153 327 1167
rect 453 1153 467 1167
rect 493 1153 507 1167
rect 873 1153 887 1167
rect 913 1153 927 1167
rect 993 1153 1007 1167
rect 1033 1153 1047 1167
rect 1193 1153 1207 1167
rect 1233 1153 1247 1167
rect 1313 1153 1327 1167
rect 1353 1153 1367 1167
rect 1473 1153 1487 1167
rect 1633 1153 1647 1167
rect 1673 1153 1687 1167
rect 1793 1153 1807 1167
rect 1833 1153 1847 1167
rect 1993 1153 2007 1167
rect 2273 1153 2287 1167
rect 2473 1153 2487 1167
rect 2513 1153 2527 1167
rect 2613 1153 2627 1167
rect 2653 1153 2667 1167
rect 2753 1153 2767 1167
rect 2793 1153 2807 1167
rect 2893 1153 2907 1167
rect 2933 1153 2947 1167
rect 3053 1153 3067 1167
rect 3093 1153 3107 1167
rect 3273 1153 3287 1167
rect 3353 1153 3367 1167
rect 3393 1153 3407 1167
rect 3573 1153 3587 1167
rect 3613 1153 3627 1167
rect 3653 1153 3667 1167
rect 3773 1153 3787 1167
rect 3813 1153 3827 1167
rect 3933 1153 3947 1167
rect 3973 1153 3987 1167
rect 4133 1153 4147 1167
rect 4233 1153 4247 1167
rect 4273 1153 4287 1167
rect 4453 1153 4467 1167
rect 4693 1153 4707 1167
rect 4853 1153 4867 1167
rect 4893 1153 4907 1167
rect 5013 1153 5027 1167
rect 5053 1153 5067 1167
rect 5153 1153 5167 1167
rect 5193 1153 5207 1167
rect 5233 1153 5247 1167
rect 5353 1153 5367 1167
rect 5393 1153 5407 1167
rect 5513 1153 5527 1167
rect 5553 1153 5567 1167
rect 5713 1153 5727 1167
rect 5753 1153 5767 1167
rect 5853 1153 5867 1167
rect 5893 1153 5907 1167
rect 5933 1153 5947 1167
rect 5993 1153 6007 1167
rect 6033 1153 6047 1167
rect 6173 1153 6187 1167
rect 6213 1153 6227 1167
rect 6333 1153 6347 1167
rect 6373 1153 6387 1167
rect 173 1133 187 1147
rect 253 1133 267 1147
rect 773 1133 787 1147
rect 813 1133 827 1147
rect 3753 1133 3767 1147
rect 4013 1133 4027 1147
rect 4153 1133 4167 1147
rect 4493 1133 4507 1147
rect 493 1113 507 1127
rect 534 1113 548 1127
rect 873 1113 887 1127
rect 993 1113 1007 1127
rect 1133 1113 1147 1127
rect 1353 1113 1367 1127
rect 1633 1113 1647 1127
rect 1793 1114 1807 1128
rect 1833 1113 1847 1127
rect 2532 1113 2546 1127
rect 2653 1113 2667 1127
rect 2733 1113 2747 1127
rect 2793 1113 2807 1127
rect 233 1093 247 1107
rect 313 1093 327 1107
rect 1193 1093 1207 1107
rect 1273 1093 1287 1107
rect 1313 1093 1327 1107
rect 1493 1093 1507 1107
rect 1533 1093 1547 1107
rect 1653 1093 1667 1107
rect 1813 1093 1827 1107
rect 2473 1093 2487 1107
rect 2813 1093 2827 1107
rect 2933 1113 2947 1127
rect 3053 1113 3067 1127
rect 3473 1113 3487 1127
rect 3533 1113 3547 1127
rect 3653 1113 3667 1127
rect 3693 1113 3707 1127
rect 3853 1113 3867 1127
rect 3913 1113 3927 1127
rect 4193 1113 4207 1127
rect 4312 1113 4326 1127
rect 4373 1113 4387 1127
rect 4893 1113 4907 1127
rect 5013 1113 5027 1127
rect 5193 1113 5207 1127
rect 5313 1113 5327 1127
rect 5353 1113 5367 1127
rect 5553 1113 5567 1127
rect 5853 1113 5867 1127
rect 6033 1113 6047 1127
rect 2913 1093 2927 1107
rect 3013 1093 3027 1107
rect 3093 1093 3107 1107
rect 3173 1093 3187 1107
rect 3333 1093 3347 1107
rect 3413 1093 3427 1107
rect 3833 1093 3847 1107
rect 3933 1093 3947 1107
rect 4073 1093 4087 1107
rect 4233 1093 4247 1107
rect 4273 1093 4287 1107
rect 973 1073 987 1087
rect 1033 1073 1047 1087
rect 1173 1073 1187 1087
rect 1333 1073 1347 1087
rect 1673 1073 1687 1087
rect 1833 1073 1847 1087
rect 1993 1073 2007 1087
rect 2253 1073 2267 1087
rect 2513 1073 2527 1087
rect 3432 1073 3446 1087
rect 3454 1073 3468 1087
rect 3692 1073 3706 1087
rect 3714 1073 3728 1087
rect 4053 1073 4067 1087
rect 4093 1073 4107 1087
rect 4753 1093 4767 1107
rect 5513 1093 5527 1107
rect 5313 1073 5327 1087
rect 5393 1073 5407 1087
rect 5474 1073 5488 1087
rect 5713 1093 5727 1107
rect 5893 1093 5907 1107
rect 6213 1093 6227 1107
rect 6333 1093 6347 1107
rect 6253 1073 6267 1087
rect 6293 1073 6307 1087
rect 613 1033 627 1047
rect 793 1033 807 1047
rect 1033 1033 1047 1047
rect 1393 1053 1407 1067
rect 1493 1053 1507 1067
rect 1633 1053 1647 1067
rect 1693 1053 1707 1067
rect 2853 1053 2867 1067
rect 1373 1033 1387 1047
rect 2873 1033 2887 1047
rect 3273 1033 3287 1047
rect 3393 1033 3407 1047
rect 3513 1033 3527 1047
rect 3953 1053 3967 1067
rect 4393 1053 4407 1067
rect 1733 1013 1747 1027
rect 2213 1013 2227 1027
rect 2373 1013 2387 1027
rect 2453 1013 2467 1027
rect 2493 1013 2507 1027
rect 2953 1013 2967 1027
rect 3033 1013 3047 1027
rect 3153 1013 3167 1027
rect 3413 1013 3427 1027
rect 3553 1013 3567 1027
rect 3593 1013 3607 1027
rect 4333 1033 4347 1047
rect 5133 1053 5147 1067
rect 5633 1053 5647 1067
rect 5673 1053 5687 1067
rect 5993 1053 6007 1067
rect 6153 1053 6167 1067
rect 4453 1033 4467 1047
rect 4553 1033 4567 1047
rect 4773 1033 4787 1047
rect 5473 1033 5487 1047
rect 6093 1033 6107 1047
rect 6253 1033 6267 1047
rect 3733 1013 3747 1027
rect 4013 1013 4027 1027
rect 4173 1013 4187 1027
rect 4293 1013 4307 1027
rect 5013 1013 5027 1027
rect 5093 1013 5107 1027
rect 593 993 607 1007
rect 773 993 787 1007
rect 1073 993 1087 1007
rect 1433 993 1447 1007
rect 1533 993 1547 1007
rect 2113 993 2127 1007
rect 2393 993 2407 1007
rect 2593 993 2607 1007
rect 2653 993 2667 1007
rect 2713 993 2727 1007
rect 2893 993 2907 1007
rect 3093 993 3107 1007
rect 3293 993 3307 1007
rect 153 973 167 987
rect 633 973 647 987
rect 733 973 747 987
rect 873 973 887 987
rect 1113 973 1127 987
rect 1193 973 1207 987
rect 1653 973 1667 987
rect 1813 973 1827 987
rect 2013 973 2027 987
rect 2133 973 2147 987
rect 2493 973 2507 987
rect 2633 973 2647 987
rect 2813 973 2827 987
rect 3013 973 3027 987
rect 3073 973 3087 987
rect 3193 973 3207 987
rect 3313 973 3327 987
rect 3393 993 3407 1007
rect 3693 993 3707 1007
rect 3893 993 3907 1007
rect 3933 993 3947 1007
rect 4133 994 4147 1008
rect 4234 993 4248 1007
rect 4473 993 4487 1007
rect 4733 993 4747 1007
rect 4773 993 4787 1007
rect 4833 993 4847 1007
rect 4933 993 4947 1007
rect 5073 993 5087 1007
rect 6013 993 6027 1007
rect 6053 993 6067 1007
rect 6293 993 6307 1007
rect 3453 973 3467 987
rect 4053 973 4067 987
rect 4133 972 4147 986
rect 4253 973 4267 987
rect 4393 973 4407 987
rect 4633 973 4647 987
rect 4713 973 4727 987
rect 4893 973 4907 987
rect 5093 973 5107 987
rect 5533 973 5547 987
rect 5593 973 5607 987
rect 5813 973 5827 987
rect 5893 973 5907 987
rect 6213 973 6227 987
rect 6473 973 6487 987
rect 3853 953 3867 967
rect 4093 953 4107 967
rect 113 933 127 947
rect 153 933 167 947
rect 273 933 287 947
rect 313 933 327 947
rect 373 933 387 947
rect 413 933 427 947
rect 453 933 467 947
rect 573 933 587 947
rect 613 933 627 947
rect 753 933 767 947
rect 793 933 807 947
rect 873 933 887 947
rect 913 933 927 947
rect 1033 933 1047 947
rect 1073 933 1087 947
rect 1193 933 1207 947
rect 1233 933 1247 947
rect 1493 933 1507 947
rect 1533 933 1547 947
rect 1613 933 1627 947
rect 1653 933 1667 947
rect 1773 933 1787 947
rect 1813 933 1827 947
rect 2093 933 2107 947
rect 2133 933 2147 947
rect 2253 933 2267 947
rect 2293 933 2307 947
rect 2413 933 2427 947
rect 2453 933 2467 947
rect 2533 933 2547 947
rect 2593 933 2607 947
rect 2633 933 2647 947
rect 2853 933 2867 947
rect 2893 933 2907 947
rect 3013 933 3027 947
rect 3053 933 3067 947
rect 3153 933 3167 947
rect 3193 933 3207 947
rect 3313 933 3327 947
rect 3353 933 3367 947
rect 3473 933 3487 947
rect 3513 933 3527 947
rect 3653 933 3667 947
rect 3693 933 3707 947
rect 3733 933 3747 947
rect 3773 933 3787 947
rect 3813 933 3827 947
rect 4133 933 4147 947
rect 4173 933 4187 947
rect 4253 933 4267 947
rect 4293 933 4307 947
rect 4333 933 4347 947
rect 4393 933 4407 947
rect 4433 933 4447 947
rect 4473 933 4487 947
rect 4593 933 4607 947
rect 4633 933 4647 947
rect 4733 933 4747 947
rect 4773 933 4787 947
rect 4893 933 4907 947
rect 4933 933 4947 947
rect 5053 933 5067 947
rect 5093 933 5107 947
rect 5133 933 5147 947
rect 5293 933 5307 947
rect 5393 933 5407 947
rect 5433 933 5447 947
rect 5533 933 5547 947
rect 5633 933 5647 947
rect 5693 933 5707 947
rect 5733 933 5747 947
rect 5773 933 5787 947
rect 5813 933 5827 947
rect 5853 933 5867 947
rect 5893 933 5907 947
rect 6033 933 6047 947
rect 6073 933 6087 947
rect 6173 933 6187 947
rect 6213 933 6227 947
rect 6333 933 6347 947
rect 6373 933 6387 947
rect 1873 913 1887 927
rect 2013 913 2027 927
rect 3973 913 3987 927
rect 4673 913 4687 927
rect 4373 893 4387 907
rect 4413 893 4427 907
rect 93 873 107 887
rect 133 873 147 887
rect 193 873 207 887
rect 293 873 307 887
rect 373 873 387 887
rect 534 873 548 887
rect 593 873 607 887
rect 713 873 727 887
rect 773 873 787 887
rect 833 873 847 887
rect 1013 873 1027 887
rect 1173 873 1187 887
rect 1393 873 1407 887
rect 1593 873 1607 887
rect 1793 873 1807 887
rect 1933 873 1947 887
rect 1973 873 1987 887
rect 2033 873 2047 887
rect 2233 873 2247 887
rect 2313 873 2327 887
rect 2393 873 2407 887
rect 2493 873 2507 887
rect 2613 873 2627 887
rect 2753 873 2767 887
rect 2973 873 2987 887
rect 3033 873 3047 887
rect 3173 873 3187 887
rect 3232 873 3246 887
rect 3453 873 3467 887
rect 3533 873 3547 887
rect 3673 873 3687 887
rect 3793 873 3807 887
rect 3933 873 3947 887
rect 4153 873 4167 887
rect 4273 873 4287 887
rect 4333 873 4347 887
rect 4393 873 4407 887
rect 4573 873 4587 887
rect 4713 873 4727 887
rect 4753 873 4767 887
rect 4853 873 4867 887
rect 4913 873 4927 887
rect 4973 873 4987 887
rect 5073 873 5087 887
rect 5173 873 5187 887
rect 5453 873 5467 887
rect 5553 873 5567 887
rect 5773 873 5787 887
rect 5873 873 5887 887
rect 5973 873 5987 887
rect 6013 873 6027 887
rect 6153 873 6167 887
rect 6193 873 6207 887
rect 6253 873 6267 887
rect 6353 873 6367 887
rect 6453 873 6467 887
rect 313 854 327 868
rect 1213 853 1227 867
rect 1633 853 1647 867
rect 2113 853 2127 867
rect 273 833 287 847
rect 313 832 327 846
rect 453 833 467 847
rect 572 833 586 847
rect 594 833 608 847
rect 813 833 827 847
rect 893 833 907 847
rect 1173 833 1187 847
rect 1733 833 1747 847
rect 1973 833 1987 847
rect 2093 833 2107 847
rect 2433 853 2447 867
rect 113 813 127 827
rect 353 813 367 827
rect 533 813 547 827
rect 753 814 767 828
rect 973 813 987 827
rect 1213 813 1227 827
rect 1393 813 1407 827
rect 1453 813 1467 827
rect 2313 813 2327 827
rect 2393 833 2407 847
rect 2753 833 2767 847
rect 3493 853 3507 867
rect 3013 833 3027 847
rect 3173 833 3187 847
rect 3213 833 3227 847
rect 2433 813 2447 827
rect 2533 813 2547 827
rect 2633 813 2647 827
rect 3033 813 3047 827
rect 3333 813 3347 827
rect 3373 833 3387 847
rect 3533 833 3547 847
rect 3573 833 3587 847
rect 3673 833 3687 847
rect 3793 833 3807 847
rect 4113 853 4127 867
rect 4653 853 4667 867
rect 4733 853 4747 867
rect 4153 833 4167 847
rect 4273 833 4287 847
rect 4353 833 4367 847
rect 4853 833 4867 847
rect 4913 833 4927 847
rect 5053 833 5067 847
rect 5413 853 5427 867
rect 5573 833 5587 847
rect 5833 853 5847 867
rect 6053 833 6067 847
rect 6353 833 6367 847
rect 3453 813 3467 827
rect 4553 813 4567 827
rect 4672 813 4686 827
rect 4713 813 4727 827
rect 5353 813 5367 827
rect 5873 813 5887 827
rect 5973 813 5987 827
rect 6033 813 6047 827
rect 193 793 207 807
rect 473 793 487 807
rect 673 793 687 807
rect 753 792 767 806
rect 853 793 867 807
rect 1833 793 1847 807
rect 2233 793 2247 807
rect 2793 793 2807 807
rect 2833 793 2847 807
rect 2993 793 3007 807
rect 3052 793 3066 807
rect 3074 793 3088 807
rect 3553 793 3567 807
rect 4353 793 4367 807
rect 4773 793 4787 807
rect 5253 793 5267 807
rect 5373 793 5387 807
rect 5413 793 5427 807
rect 5533 793 5547 807
rect 5693 793 5707 807
rect 5752 793 5766 807
rect 5774 793 5788 807
rect 6013 793 6027 807
rect 6113 793 6127 807
rect 293 773 307 787
rect 413 773 427 787
rect 833 773 847 787
rect 1813 773 1827 787
rect 1973 773 1987 787
rect 2032 773 2046 787
rect 2054 773 2068 787
rect 2553 773 2567 787
rect 2593 773 2607 787
rect 2693 773 2707 787
rect 2853 773 2867 787
rect 3273 773 3287 787
rect 3493 773 3507 787
rect 3773 773 3787 787
rect 3933 773 3947 787
rect 4113 773 4127 787
rect 4273 773 4287 787
rect 4673 773 4687 787
rect 4793 773 4807 787
rect 4913 773 4927 787
rect 5073 773 5087 787
rect 5173 773 5187 787
rect 5293 773 5307 787
rect 5433 773 5447 787
rect 5513 773 5527 787
rect 5553 773 5567 787
rect 5593 773 5607 787
rect 5813 773 5827 787
rect 113 753 127 767
rect 553 753 567 767
rect 713 753 727 767
rect 1173 753 1187 767
rect 1593 753 1607 767
rect 2193 753 2207 767
rect 2653 753 2667 767
rect 2713 753 2727 767
rect 2773 753 2787 767
rect 2913 753 2927 767
rect 3213 753 3227 767
rect 4413 753 4427 767
rect 4513 753 4527 767
rect 4653 753 4667 767
rect 4813 753 4827 767
rect 4873 753 4887 767
rect 4973 753 4987 767
rect 5393 753 5407 767
rect 5453 753 5467 767
rect 5613 753 5627 767
rect 5773 753 5787 767
rect 5873 753 5887 767
rect 153 733 167 747
rect 373 733 387 747
rect 873 733 887 747
rect 1033 733 1047 747
rect 1233 733 1247 747
rect 1273 733 1287 747
rect 1413 733 1427 747
rect 1693 733 1707 747
rect 1873 733 1887 747
rect 1933 733 1947 747
rect 1993 733 2007 747
rect 2393 733 2407 747
rect 2493 733 2507 747
rect 2633 733 2647 747
rect 2673 733 2687 747
rect 3073 733 3087 747
rect 3233 733 3247 747
rect 3713 733 3727 747
rect 3773 733 3787 747
rect 233 713 247 727
rect 713 713 727 727
rect 753 713 767 727
rect 2193 713 2207 727
rect 2233 713 2247 727
rect 2553 713 2567 727
rect 113 693 127 707
rect 273 693 287 707
rect 353 693 367 707
rect 533 693 547 707
rect 653 693 667 707
rect 873 693 887 707
rect 953 693 967 707
rect 1053 693 1067 707
rect 1113 693 1127 707
rect 1233 693 1247 707
rect 1333 693 1347 707
rect 1433 693 1447 707
rect 1493 693 1507 707
rect 1593 693 1607 707
rect 1753 693 1767 707
rect 1793 693 1807 707
rect 1833 693 1847 707
rect 1873 693 1887 707
rect 2053 693 2067 707
rect 2313 693 2327 707
rect 2393 693 2407 707
rect 2593 694 2607 708
rect 3053 713 3067 727
rect 3113 713 3127 727
rect 3153 713 3167 727
rect 3193 713 3207 727
rect 3333 713 3347 727
rect 3373 713 3387 727
rect 3793 713 3807 727
rect 2713 693 2727 707
rect 2793 693 2807 707
rect 2853 693 2867 707
rect 2953 693 2967 707
rect 2993 693 3007 707
rect 3233 693 3247 707
rect 3273 693 3287 707
rect 3493 693 3507 707
rect 3612 693 3626 707
rect 3693 693 3707 707
rect 3913 733 3927 747
rect 3973 733 3987 747
rect 4073 733 4087 747
rect 3953 713 3967 727
rect 4333 733 4347 747
rect 4593 733 4607 747
rect 4633 733 4647 747
rect 4913 733 4927 747
rect 4953 733 4967 747
rect 5053 733 5067 747
rect 5653 733 5667 747
rect 5733 733 5747 747
rect 5813 733 5827 747
rect 6013 733 6027 747
rect 6053 733 6067 747
rect 6413 733 6427 747
rect 3813 693 3827 707
rect 3873 693 3887 707
rect 3973 693 3987 707
rect 4033 693 4047 707
rect 4113 693 4127 707
rect 4193 693 4207 707
rect 4353 693 4367 707
rect 4513 693 4527 707
rect 4613 693 4627 707
rect 4793 693 4807 707
rect 4953 693 4967 707
rect 5113 693 5127 707
rect 5273 693 5287 707
rect 5353 693 5367 707
rect 5453 693 5467 707
rect 5553 693 5567 707
rect 5613 693 5627 707
rect 5813 693 5827 707
rect 5873 693 5887 707
rect 5933 693 5947 707
rect 6013 693 6027 707
rect 6113 693 6127 707
rect 6193 693 6207 707
rect 6333 693 6347 707
rect 2593 672 2607 686
rect 2633 673 2647 687
rect 3253 673 3267 687
rect 3313 673 3327 687
rect 693 653 707 667
rect 773 653 787 667
rect 2113 653 2127 667
rect 2913 653 2927 667
rect 3033 653 3047 667
rect 3133 653 3147 667
rect 3213 653 3227 667
rect 213 633 227 647
rect 253 633 267 647
rect 373 633 387 647
rect 413 633 427 647
rect 513 633 527 647
rect 553 633 567 647
rect 733 633 747 647
rect 853 633 867 647
rect 893 633 907 647
rect 1033 633 1047 647
rect 1073 633 1087 647
rect 1213 633 1227 647
rect 1253 633 1267 647
rect 1413 633 1427 647
rect 1453 633 1467 647
rect 1573 633 1587 647
rect 1613 633 1627 647
rect 1733 633 1747 647
rect 1773 633 1787 647
rect 1893 633 1907 647
rect 1933 633 1947 647
rect 2033 633 2047 647
rect 2073 633 2087 647
rect 2373 633 2387 647
rect 2413 633 2427 647
rect 2493 633 2507 647
rect 2533 633 2547 647
rect 2653 633 2667 647
rect 2693 633 2707 647
rect 2733 633 2747 647
rect 2833 633 2847 647
rect 2873 633 2887 647
rect 3173 633 3187 647
rect 3293 633 3307 647
rect 3393 633 3407 647
rect 3473 633 3487 647
rect 3513 633 3527 647
rect 3673 633 3687 647
rect 3713 633 3727 647
rect 3793 633 3807 647
rect 3833 633 3847 647
rect 3953 633 3967 647
rect 3993 633 4007 647
rect 4133 633 4147 647
rect 4173 633 4187 647
rect 4293 633 4307 647
rect 4333 633 4347 647
rect 4493 633 4507 647
rect 4533 633 4547 647
rect 4633 633 4647 647
rect 4673 633 4687 647
rect 4773 633 4787 647
rect 4813 633 4827 647
rect 4933 633 4947 647
rect 4973 633 4987 647
rect 5093 633 5107 647
rect 5133 633 5147 647
rect 5253 633 5267 647
rect 5293 633 5307 647
rect 5473 633 5487 647
rect 5513 633 5527 647
rect 5633 633 5647 647
rect 5673 633 5687 647
rect 5793 633 5807 647
rect 5833 633 5847 647
rect 5993 633 6007 647
rect 6033 633 6047 647
rect 6133 633 6147 647
rect 6173 633 6187 647
rect 6313 633 6327 647
rect 6353 633 6367 647
rect 353 613 367 627
rect 653 613 667 627
rect 1793 613 1807 627
rect 1833 613 1847 627
rect 2933 613 2947 627
rect 3033 613 3047 627
rect 3133 613 3147 627
rect 253 593 267 607
rect 853 593 867 607
rect 633 573 647 587
rect 993 593 1007 607
rect 1413 593 1427 607
rect 1573 593 1587 607
rect 1893 593 1907 607
rect 2113 593 2127 607
rect 2233 593 2247 607
rect 2533 593 2547 607
rect 2693 593 2707 607
rect 2973 593 2987 607
rect 3233 593 3247 607
rect 3753 593 3767 607
rect 4133 593 4147 607
rect 4533 593 4547 607
rect 4673 593 4687 607
rect 4833 593 4847 607
rect 4973 593 4987 607
rect 5013 593 5027 607
rect 5133 593 5147 607
rect 5273 593 5287 607
rect 5413 593 5427 607
rect 5593 593 5607 607
rect 5633 593 5647 607
rect 6033 593 6047 607
rect 6173 593 6187 607
rect 6353 593 6367 607
rect 1053 573 1067 587
rect 1213 573 1227 587
rect 1613 573 1627 587
rect 1693 573 1707 587
rect 2413 573 2427 587
rect 2613 573 2627 587
rect 2733 573 2747 587
rect 3093 573 3107 587
rect 3213 573 3227 587
rect 3793 573 3807 587
rect 3993 573 4007 587
rect 4813 573 4827 587
rect 5313 573 5327 587
rect 5373 573 5387 587
rect 5473 573 5487 587
rect 5673 573 5687 587
rect 5873 573 5887 587
rect 6313 573 6327 587
rect 6393 573 6407 587
rect 893 553 907 567
rect 933 553 947 567
rect 1493 553 1507 567
rect 473 533 487 547
rect 1333 533 1347 547
rect 1433 533 1447 547
rect 2053 553 2067 567
rect 2693 553 2707 567
rect 2833 553 2847 567
rect 3633 553 3647 567
rect 3673 553 3687 567
rect 3833 553 3847 567
rect 4173 553 4187 567
rect 4673 553 4687 567
rect 5233 553 5247 567
rect 5493 553 5507 567
rect 5973 553 5987 567
rect 6133 553 6147 567
rect 1573 533 1587 547
rect 1733 533 1747 547
rect 1993 533 2007 547
rect 2073 533 2087 547
rect 2553 533 2567 547
rect 3873 533 3887 547
rect 4193 533 4207 547
rect 4713 533 4727 547
rect 4933 533 4947 547
rect 5593 533 5607 547
rect 5653 533 5667 547
rect 6033 533 6047 547
rect 113 513 127 527
rect 233 513 247 527
rect 293 513 307 527
rect 1013 513 1027 527
rect 1093 513 1107 527
rect 1253 513 1267 527
rect 1753 513 1767 527
rect 2093 513 2107 527
rect 2493 513 2507 527
rect 3053 513 3067 527
rect 3433 513 3447 527
rect 733 493 747 507
rect 1393 493 1407 507
rect 2053 493 2067 507
rect 2373 493 2387 507
rect 2513 493 2527 507
rect 2553 493 2567 507
rect 3292 493 3306 507
rect 3553 513 3567 527
rect 5933 513 5947 527
rect 3913 493 3927 507
rect 3953 493 3967 507
rect 4012 493 4026 507
rect 4073 493 4087 507
rect 4133 493 4147 507
rect 5793 493 5807 507
rect 773 473 787 487
rect 1093 473 1107 487
rect 1233 473 1247 487
rect 1353 473 1367 487
rect 2933 473 2947 487
rect 3013 473 3027 487
rect 3173 473 3187 487
rect 3273 473 3287 487
rect 3713 473 3727 487
rect 4093 473 4107 487
rect 4192 473 4206 487
rect 4393 473 4407 487
rect 4753 473 4767 487
rect 5733 473 5747 487
rect 6193 473 6207 487
rect 6393 473 6407 487
rect 153 453 167 467
rect 273 453 287 467
rect 593 453 607 467
rect 952 453 966 467
rect 1173 453 1187 467
rect 1433 453 1447 467
rect 1513 453 1527 467
rect 1693 453 1707 467
rect 1873 453 1887 467
rect 3453 453 3467 467
rect 673 433 687 447
rect 713 433 727 447
rect 873 433 887 447
rect 1773 433 1787 447
rect 1813 433 1827 447
rect 2353 433 2367 447
rect 113 413 127 427
rect 153 413 167 427
rect 233 413 247 427
rect 393 413 407 427
rect 433 413 447 427
rect 593 413 607 427
rect 633 413 647 427
rect 733 413 747 427
rect 773 413 787 427
rect 893 413 907 427
rect 933 413 947 427
rect 1053 413 1067 427
rect 1093 413 1107 427
rect 1133 413 1147 427
rect 1173 413 1187 427
rect 1213 413 1227 427
rect 1353 413 1367 427
rect 1393 413 1407 427
rect 1533 413 1547 427
rect 1573 413 1587 427
rect 1653 413 1667 427
rect 1693 413 1707 427
rect 1833 413 1847 427
rect 1873 413 1887 427
rect 1993 413 2007 427
rect 2033 413 2047 427
rect 2153 413 2167 427
rect 2193 413 2207 427
rect 2373 413 2387 427
rect 2653 413 2667 427
rect 2693 413 2707 427
rect 2853 413 2867 427
rect 2893 413 2907 427
rect 3013 413 3027 427
rect 3053 413 3067 427
rect 3233 413 3247 427
rect 3433 413 3447 427
rect 3473 413 3487 427
rect 3533 453 3547 467
rect 4133 453 4147 467
rect 4253 453 4267 467
rect 4413 453 4427 467
rect 4613 453 4627 467
rect 4793 453 4807 467
rect 5113 453 5127 467
rect 5393 453 5407 467
rect 5433 453 5447 467
rect 5573 453 5587 467
rect 5753 453 5767 467
rect 6313 453 6327 467
rect 4193 433 4207 447
rect 3593 413 3607 427
rect 3633 413 3647 427
rect 3753 413 3767 427
rect 3793 413 3807 427
rect 3933 413 3947 427
rect 3973 413 3987 427
rect 4073 413 4087 427
rect 4113 413 4127 427
rect 5933 433 5947 447
rect 5973 433 5987 447
rect 4413 413 4427 427
rect 4453 413 4467 427
rect 4753 413 4767 427
rect 4793 413 4807 427
rect 5113 413 5127 427
rect 5253 413 5267 427
rect 5293 413 5307 427
rect 5393 413 5407 427
rect 5433 413 5447 427
rect 5533 413 5547 427
rect 5573 413 5587 427
rect 5713 413 5727 427
rect 5753 413 5767 427
rect 5833 413 5847 427
rect 5873 413 5887 427
rect 5913 413 5927 427
rect 6153 413 6167 427
rect 6193 413 6207 427
rect 6353 413 6367 427
rect 353 393 367 407
rect 1253 393 1267 407
rect 1313 393 1327 407
rect 2333 393 2347 407
rect 2413 393 2427 407
rect 4253 393 4267 407
rect 4333 393 4347 407
rect 4573 393 4587 407
rect 4673 393 4687 407
rect 4833 393 4847 407
rect 5053 393 5067 407
rect 6113 393 6127 407
rect 793 373 807 387
rect 3813 373 3827 387
rect 3873 374 3887 388
rect 3993 373 4007 387
rect 4053 373 4067 387
rect 253 353 267 367
rect 413 353 427 367
rect 533 353 547 367
rect 613 353 627 367
rect 713 353 727 367
rect 873 353 887 367
rect 993 353 1007 367
rect 1153 353 1167 367
rect 1193 353 1207 367
rect 1293 353 1307 367
rect 1333 353 1347 367
rect 1413 353 1427 367
rect 1453 353 1467 367
rect 1553 353 1567 367
rect 1593 353 1607 367
rect 1633 353 1647 367
rect 1673 353 1687 367
rect 1773 353 1787 367
rect 1813 353 1827 367
rect 2013 353 2027 367
rect 573 333 587 347
rect 753 333 767 347
rect 973 333 987 347
rect 1573 333 1587 347
rect 1613 333 1627 347
rect 413 313 427 327
rect 713 313 727 327
rect 853 313 867 327
rect 1413 313 1427 327
rect 1813 313 1827 327
rect 2173 353 2187 367
rect 2233 353 2247 367
rect 2633 353 2647 367
rect 2733 353 2747 367
rect 2873 353 2887 367
rect 2933 353 2947 367
rect 3033 353 3047 367
rect 2153 333 2167 347
rect 2353 333 2367 347
rect 2393 333 2407 347
rect 2493 333 2507 347
rect 2533 333 2547 347
rect 2013 313 2027 327
rect 2173 313 2187 327
rect 2313 313 2327 327
rect 2593 313 2607 327
rect 3213 352 3227 366
rect 3273 352 3287 366
rect 3453 353 3467 367
rect 3653 353 3667 367
rect 3733 353 3747 367
rect 3873 353 3887 367
rect 3953 353 3967 367
rect 4093 353 4107 367
rect 4613 353 4627 367
rect 4813 353 4827 367
rect 5093 353 5107 367
rect 5133 353 5147 367
rect 5273 353 5287 367
rect 5313 353 5327 367
rect 5453 353 5467 367
rect 5493 353 5507 367
rect 5593 353 5607 367
rect 5733 353 5747 367
rect 5793 353 5807 367
rect 5933 353 5947 367
rect 6113 353 6127 367
rect 6313 353 6327 367
rect 3413 333 3427 347
rect 2893 313 2907 327
rect 2993 313 3007 327
rect 3033 313 3047 327
rect 3493 313 3507 327
rect 3853 333 3867 347
rect 3973 333 3987 347
rect 4053 333 4067 347
rect 4133 333 4147 347
rect 4273 333 4287 347
rect 4313 333 4327 347
rect 4433 333 4447 347
rect 4233 313 4247 327
rect 4333 313 4347 327
rect 4613 313 4627 327
rect 4893 333 4907 347
rect 4933 333 4947 347
rect 5053 333 5067 347
rect 6033 333 6047 347
rect 6073 333 6087 347
rect 5393 313 5407 327
rect 5933 313 5947 327
rect 613 293 627 307
rect 753 293 767 307
rect 793 293 807 307
rect 1033 293 1047 307
rect 1193 293 1207 307
rect 1453 293 1467 307
rect 1793 293 1807 307
rect 2093 293 2107 307
rect 2133 293 2147 307
rect 2353 293 2367 307
rect 2393 293 2407 307
rect 2873 293 2887 307
rect 3133 293 3147 307
rect 3733 293 3747 307
rect 4273 293 4287 307
rect 93 273 107 287
rect 373 273 387 287
rect 573 273 587 287
rect 713 273 727 287
rect 893 273 907 287
rect 1873 273 1887 287
rect 1993 273 2007 287
rect 133 253 147 267
rect 433 253 447 267
rect 714 253 728 267
rect 833 253 847 267
rect 1093 253 1107 267
rect 1573 253 1587 267
rect 2013 253 2027 267
rect 2513 273 2527 287
rect 2653 273 2667 287
rect 2793 273 2807 287
rect 2833 273 2847 287
rect 3533 273 3547 287
rect 3593 273 3607 287
rect 3813 273 3827 287
rect 4673 293 4687 307
rect 4833 293 4847 307
rect 4893 293 4907 307
rect 5093 293 5107 307
rect 5513 293 5527 307
rect 5713 293 5727 307
rect 5973 293 5987 307
rect 4373 273 4387 287
rect 4453 273 4467 287
rect 4573 273 4587 287
rect 5153 273 5167 287
rect 5193 273 5207 287
rect 5433 273 5447 287
rect 6073 273 6087 287
rect 553 233 567 247
rect 692 233 706 247
rect 873 233 887 247
rect 1053 233 1067 247
rect 1353 233 1367 247
rect 1533 233 1547 247
rect 2133 233 2147 247
rect 2393 253 2407 267
rect 2853 253 2867 267
rect 2953 253 2967 267
rect 3053 253 3067 267
rect 3093 253 3107 267
rect 3273 253 3287 267
rect 3373 253 3387 267
rect 3693 253 3707 267
rect 3733 253 3747 267
rect 3893 253 3907 267
rect 2373 233 2387 247
rect 2413 233 2427 247
rect 2473 233 2487 247
rect 3173 233 3187 247
rect 3333 233 3347 247
rect 3413 233 3427 247
rect 3473 233 3487 247
rect 3633 233 3647 247
rect 3813 233 3827 247
rect 4153 253 4167 267
rect 5313 253 5327 267
rect 5473 253 5487 267
rect 5633 253 5647 267
rect 3993 233 4007 247
rect 4433 233 4447 247
rect 4593 233 4607 247
rect 4833 233 4847 247
rect 5013 233 5027 247
rect 5533 233 5547 247
rect 5753 233 5767 247
rect 5953 233 5967 247
rect 6112 233 6126 247
rect 6134 233 6148 247
rect 293 213 307 227
rect 433 213 447 227
rect 473 213 487 227
rect 653 213 667 227
rect 714 213 728 227
rect 832 213 846 227
rect 973 213 987 227
rect 1113 213 1127 227
rect 1293 213 1307 227
rect 1593 213 1607 227
rect 2033 213 2047 227
rect 2233 213 2247 227
rect 2293 213 2307 227
rect 2693 213 2707 227
rect 2753 213 2767 227
rect 3193 213 3207 227
rect 3433 213 3447 227
rect 3673 213 3687 227
rect 4093 213 4107 227
rect 4193 213 4207 227
rect 4373 213 4387 227
rect 4653 213 4667 227
rect 373 193 387 207
rect 1033 193 1047 207
rect 1373 193 1387 207
rect 1793 193 1807 207
rect 2193 193 2207 207
rect 2793 193 2807 207
rect 2993 193 3007 207
rect 3693 193 3707 207
rect 5133 213 5147 227
rect 5213 213 5227 227
rect 5353 213 5367 227
rect 5693 213 5707 227
rect 5973 213 5987 227
rect 234 173 248 187
rect 293 173 307 187
rect 433 173 447 187
rect 553 173 567 187
rect 333 153 347 167
rect 393 153 407 167
rect 653 173 667 187
rect 693 173 707 187
rect 793 173 807 187
rect 833 173 847 187
rect 933 173 947 187
rect 973 173 987 187
rect 1113 173 1127 187
rect 1273 173 1287 187
rect 1393 173 1407 187
rect 1533 173 1547 187
rect 1573 173 1587 187
rect 1713 173 1727 187
rect 1753 173 1767 187
rect 1833 173 1847 187
rect 1873 173 1887 187
rect 1913 173 1927 187
rect 1993 173 2007 187
rect 2093 173 2107 187
rect 2233 173 2247 187
rect 2313 173 2327 187
rect 2353 173 2367 187
rect 2413 173 2427 187
rect 2513 173 2527 187
rect 2633 173 2647 187
rect 2693 173 2707 187
rect 2833 173 2847 187
rect 2953 173 2967 187
rect 3113 173 3127 187
rect 3273 173 3287 187
rect 3333 173 3347 187
rect 3473 173 3487 187
rect 3533 173 3547 187
rect 3633 173 3647 187
rect 3813 173 3827 187
rect 3893 173 3907 187
rect 3993 173 4007 187
rect 4033 173 4047 187
rect 4073 173 4087 187
rect 4173 173 4187 187
rect 4273 173 4287 187
rect 4373 173 4387 187
rect 4453 173 4467 187
rect 4573 173 4587 187
rect 4693 173 4707 187
rect 4753 173 4767 187
rect 4953 173 4967 187
rect 5273 173 5287 187
rect 5353 173 5367 187
rect 5453 173 5467 187
rect 5533 173 5547 187
rect 5693 173 5707 187
rect 5833 173 5847 187
rect 5953 173 5967 187
rect 6093 173 6107 187
rect 6413 173 6427 187
rect 1013 153 1027 167
rect 1073 153 1087 167
rect 1313 153 1327 167
rect 1353 153 1367 167
rect 2873 153 2887 167
rect 2913 153 2927 167
rect 3073 153 3087 167
rect 3673 153 3687 167
rect 3713 153 3727 167
rect 3853 153 3867 167
rect 493 133 507 147
rect 693 133 707 147
rect 1133 133 1147 147
rect 1193 133 1207 147
rect 3013 133 3027 147
rect 3093 133 3107 147
rect 3293 133 3307 147
rect 3733 133 3747 147
rect 4433 133 4447 147
rect 93 113 107 127
rect 133 113 147 127
rect 273 113 287 127
rect 313 113 327 127
rect 373 113 387 127
rect 413 113 427 127
rect 453 113 467 127
rect 513 113 527 127
rect 593 113 607 127
rect 633 113 647 127
rect 673 113 687 127
rect 733 113 747 127
rect 773 113 787 127
rect 813 113 827 127
rect 953 113 967 127
rect 993 113 1007 127
rect 1033 113 1047 127
rect 1213 113 1227 127
rect 1253 113 1267 127
rect 1293 113 1307 127
rect 1373 113 1387 127
rect 1413 113 1427 127
rect 1553 113 1567 127
rect 1593 113 1607 127
rect 1733 113 1747 127
rect 1773 113 1787 127
rect 1893 113 1907 127
rect 1933 113 1947 127
rect 2173 113 2187 127
rect 2213 113 2227 127
rect 2253 113 2267 127
rect 2333 113 2347 127
rect 2373 113 2387 127
rect 2493 113 2507 127
rect 2533 113 2547 127
rect 2773 113 2787 127
rect 2813 113 2827 127
rect 2853 113 2867 127
rect 2933 113 2947 127
rect 2973 113 2987 127
rect 3133 113 3147 127
rect 3173 113 3187 127
rect 3453 113 3467 127
rect 3493 113 3507 127
rect 3613 113 3627 127
rect 3653 113 3667 127
rect 3793 113 3807 127
rect 3833 113 3847 127
rect 3933 113 3947 127
rect 3973 113 3987 127
rect 4093 113 4107 127
rect 4133 113 4147 127
rect 4313 113 4327 127
rect 4353 113 4367 127
rect 4393 113 4407 127
rect 4593 113 4607 127
rect 4693 113 4707 127
rect 4733 113 4747 127
rect 4853 113 4867 127
rect 4893 113 4907 127
rect 5013 113 5027 127
rect 5053 113 5067 127
rect 5173 113 5187 127
rect 5213 113 5227 127
rect 5333 113 5347 127
rect 5373 113 5387 127
rect 5473 113 5487 127
rect 5513 113 5527 127
rect 5673 113 5687 127
rect 5713 113 5727 127
rect 5753 113 5767 127
rect 5893 113 5907 127
rect 5933 113 5947 127
rect 5973 113 5987 127
rect 6113 113 6127 127
rect 6153 113 6167 127
rect 6253 113 6267 127
rect 6293 113 6307 127
rect 6333 113 6347 127
rect 3213 93 3227 107
rect 3373 93 3387 107
rect 3873 93 3887 107
rect 3993 93 4007 107
rect 4753 93 4767 107
rect 4813 93 4827 107
rect 6033 93 6047 107
rect 6093 93 6107 107
rect 6193 93 6207 107
rect 273 73 287 87
rect 633 73 647 87
rect 773 73 787 87
rect 813 73 827 87
rect 893 73 907 87
rect 953 73 967 87
rect 993 73 1007 87
rect 1253 73 1267 87
rect 1413 73 1427 87
rect 1453 73 1467 87
rect 1553 73 1567 87
rect 1893 73 1907 87
rect 2413 73 2427 87
rect 1733 53 1747 67
rect 1773 53 1787 67
rect 1933 53 1947 67
rect 3493 73 3507 87
rect 3653 73 3667 87
rect 3713 73 3727 87
rect 3833 73 3847 87
rect 3973 73 3987 87
rect 4593 73 4607 87
rect 4893 73 4907 87
rect 5053 73 5067 87
rect 5333 73 5347 87
rect 5673 73 5687 87
rect 2853 53 2867 67
rect 2973 53 2987 67
rect 3793 53 3807 67
rect 3933 53 3947 67
rect 5173 53 5187 67
rect 1033 33 1047 47
rect 1293 33 1307 47
rect 2053 33 2067 47
rect 2513 33 2527 47
rect 3054 33 3068 47
rect 4173 33 4187 47
rect 233 13 247 27
rect 853 13 867 27
rect 2093 13 2107 27
rect 2373 13 2387 27
rect 2533 13 2547 27
rect 2693 13 2707 27
rect 3112 13 3126 27
rect 3134 13 3148 27
rect 3533 13 3547 27
rect 3573 13 3587 27
rect 3673 13 3687 27
rect 3733 13 3747 27
rect 4953 13 4967 27
rect 5133 13 5147 27
rect 5173 13 5187 27
<< metal3 >>
rect 200 6424 213 6427
rect 196 6413 213 6424
rect 356 6416 393 6424
rect 136 6327 144 6413
rect 196 6367 204 6413
rect 236 6227 244 6353
rect 276 6207 284 6353
rect 276 6167 284 6193
rect 356 6187 364 6416
rect 556 6367 564 6473
rect 596 6367 604 6453
rect 556 6356 573 6367
rect 560 6353 573 6356
rect 596 6356 613 6367
rect 600 6353 613 6356
rect 376 6327 384 6353
rect 416 6247 424 6353
rect 116 6047 124 6073
rect 156 5907 164 6133
rect 236 5967 244 6073
rect 176 5847 184 5953
rect 136 5767 144 5833
rect 256 5807 264 5893
rect 296 5847 304 6113
rect 396 6087 404 6173
rect 476 6147 484 6233
rect 516 6147 524 6313
rect 676 6267 684 6413
rect 696 6367 704 6473
rect 736 6427 744 6453
rect 936 6427 944 6473
rect 696 6356 713 6367
rect 700 6353 713 6356
rect 816 6364 824 6413
rect 976 6367 984 6453
rect 1056 6427 1064 6513
rect 767 6356 824 6364
rect 967 6356 984 6367
rect 967 6353 980 6356
rect 916 6307 924 6353
rect 996 6307 1004 6353
rect 580 6144 593 6147
rect 576 6133 593 6144
rect 576 6087 584 6133
rect 616 6087 624 6193
rect 673 6144 687 6153
rect 647 6140 687 6144
rect 647 6136 684 6140
rect 387 6076 404 6087
rect 387 6073 400 6076
rect 356 5907 364 6033
rect 676 6007 684 6073
rect 476 5907 484 5933
rect 676 5907 684 5933
rect 16 5087 24 5733
rect 96 5567 104 5753
rect 336 5627 344 5833
rect 356 5687 364 5893
rect 436 5807 444 5853
rect 416 5627 424 5653
rect 467 5624 480 5627
rect 467 5613 484 5624
rect 116 5487 124 5613
rect 136 5527 144 5553
rect 156 5507 164 5613
rect 256 5507 264 5613
rect 296 5527 304 5613
rect 376 5567 384 5613
rect 76 5147 84 5373
rect 116 5327 124 5473
rect 156 5327 164 5493
rect 116 5147 124 5173
rect 276 5167 284 5373
rect 296 5327 304 5513
rect 336 5447 344 5493
rect 336 5327 344 5433
rect 436 5427 444 5553
rect 476 5527 484 5613
rect 496 5467 504 5833
rect 596 5627 604 5893
rect 656 5667 664 5833
rect 696 5727 704 5833
rect 736 5807 744 6273
rect 876 6136 913 6144
rect 776 6027 784 6053
rect 776 5847 784 6013
rect 816 5947 824 6053
rect 856 5987 864 6113
rect 876 6007 884 6136
rect 953 6124 967 6133
rect 953 6120 1024 6124
rect 956 6116 1024 6120
rect 1016 6087 1024 6116
rect 920 6084 933 6087
rect 916 6073 933 6084
rect 916 6027 924 6073
rect 976 6047 984 6073
rect 1036 6047 1044 6253
rect 1056 6147 1064 6413
rect 1096 6307 1104 6473
rect 1156 6247 1164 6353
rect 1196 6287 1204 6353
rect 1276 6327 1284 6413
rect 1316 6367 1324 6453
rect 1496 6447 1504 6493
rect 1536 6427 1544 6453
rect 1696 6427 1704 6493
rect 1856 6447 1864 6493
rect 2256 6487 2264 6564
rect 2296 6527 2304 6564
rect 2096 6427 2104 6473
rect 1216 6207 1224 6293
rect 1216 6147 1224 6193
rect 1256 6187 1264 6213
rect 1256 6147 1264 6173
rect 1107 6144 1120 6147
rect 1107 6133 1124 6144
rect 1016 6036 1033 6044
rect 816 5847 824 5933
rect 936 5907 944 5993
rect 836 5767 844 5893
rect 916 5807 924 5833
rect 956 5807 964 5833
rect 956 5767 964 5793
rect 976 5707 984 5933
rect 996 5827 1004 5993
rect 1016 5747 1024 6036
rect 1056 5947 1064 6133
rect 1116 6087 1124 6133
rect 1296 6127 1304 6173
rect 1336 6084 1344 6253
rect 1356 6227 1364 6353
rect 1376 6307 1384 6413
rect 1476 6327 1484 6353
rect 1396 6087 1404 6173
rect 1287 6076 1344 6084
rect 1216 5987 1224 6073
rect 1396 6047 1404 6073
rect 1436 6067 1444 6113
rect 1476 6107 1484 6233
rect 1516 6227 1524 6353
rect 1676 6327 1684 6353
rect 1556 6207 1564 6233
rect 1516 6147 1524 6173
rect 1536 6136 1553 6144
rect 1536 6064 1544 6136
rect 1567 6144 1580 6147
rect 1567 6133 1584 6144
rect 1576 6107 1584 6133
rect 1596 6127 1604 6253
rect 1716 6187 1724 6353
rect 1736 6247 1744 6413
rect 1896 6367 1904 6413
rect 2136 6367 2144 6433
rect 1887 6356 1904 6367
rect 1887 6353 1900 6356
rect 2127 6356 2144 6367
rect 2127 6353 2140 6356
rect 1836 6327 1844 6353
rect 1667 6096 1724 6104
rect 1716 6067 1724 6096
rect 1736 6067 1744 6093
rect 1507 6056 1544 6064
rect 1727 6056 1744 6067
rect 1727 6053 1740 6056
rect 1096 5927 1104 5973
rect 1120 5924 1133 5927
rect 1116 5913 1133 5924
rect 1116 5904 1124 5913
rect 1256 5907 1264 5933
rect 1296 5907 1304 5993
rect 1076 5900 1124 5904
rect 1073 5896 1124 5900
rect 687 5616 713 5624
rect 767 5616 793 5624
rect 556 5584 564 5613
rect 536 5580 564 5584
rect 533 5576 564 5580
rect 533 5567 547 5576
rect 576 5487 584 5533
rect 616 5507 624 5553
rect 556 5424 564 5453
rect 556 5416 584 5424
rect 496 5387 504 5413
rect 576 5404 584 5416
rect 576 5396 604 5404
rect 296 5207 304 5313
rect 396 5287 404 5373
rect 476 5267 484 5313
rect 516 5287 524 5313
rect 116 5107 124 5133
rect 156 5107 164 5133
rect 236 5107 244 5133
rect 316 5124 324 5173
rect 296 5116 324 5124
rect 296 5107 304 5116
rect 416 5107 424 5193
rect 556 5164 564 5373
rect 596 5187 604 5396
rect 656 5327 664 5413
rect 676 5387 684 5433
rect 716 5327 724 5513
rect 707 5316 724 5327
rect 707 5313 720 5316
rect 696 5267 704 5313
rect 736 5187 744 5373
rect 756 5327 764 5553
rect 836 5507 844 5553
rect 856 5447 864 5693
rect 1036 5627 1044 5893
rect 1073 5887 1087 5896
rect 1116 5787 1124 5853
rect 947 5616 973 5624
rect 1027 5616 1044 5627
rect 1027 5613 1040 5616
rect 1056 5607 1064 5653
rect 1113 5627 1127 5633
rect 1113 5620 1133 5627
rect 1116 5616 1133 5620
rect 1120 5613 1133 5616
rect 1056 5567 1064 5593
rect 1047 5556 1064 5567
rect 1096 5567 1104 5593
rect 1096 5556 1113 5567
rect 1047 5553 1060 5556
rect 1100 5553 1113 5556
rect 836 5380 873 5384
rect 833 5376 873 5380
rect 833 5367 847 5376
rect 556 5156 584 5164
rect 493 5107 507 5113
rect 287 5096 304 5107
rect 287 5093 300 5096
rect 416 5096 433 5107
rect 420 5093 433 5096
rect 487 5100 507 5107
rect 487 5096 504 5100
rect 487 5093 500 5096
rect 76 4807 84 5033
rect 136 5007 144 5033
rect 256 5007 264 5033
rect 96 4867 104 4893
rect 156 4807 164 4893
rect 76 4587 84 4793
rect 116 4767 124 4793
rect 176 4767 184 4933
rect 296 4927 304 5013
rect 316 5007 324 5093
rect 396 4947 404 5033
rect 496 5007 504 5033
rect 127 4756 144 4764
rect 136 4587 144 4756
rect 256 4647 264 4853
rect 296 4767 304 4853
rect 127 4576 144 4587
rect 127 4573 140 4576
rect 16 4487 24 4553
rect 36 4307 44 4533
rect 136 4347 144 4413
rect 196 4247 204 4553
rect 256 4527 264 4633
rect 376 4627 384 4853
rect 416 4807 424 4893
rect 453 4867 467 4873
rect 447 4860 467 4867
rect 447 4856 464 4860
rect 447 4853 460 4856
rect 476 4824 484 4913
rect 456 4820 484 4824
rect 453 4816 484 4820
rect 453 4807 467 4816
rect 496 4767 504 4873
rect 536 4867 544 5133
rect 576 5107 584 5156
rect 636 5107 644 5153
rect 576 5096 593 5107
rect 580 5093 593 5096
rect 796 5047 804 5353
rect 896 5327 904 5433
rect 827 5316 853 5324
rect 576 5007 584 5033
rect 556 4824 564 4973
rect 536 4816 564 4824
rect 316 4567 324 4613
rect 376 4587 384 4613
rect 436 4587 444 4633
rect 536 4587 544 4816
rect 576 4807 584 4993
rect 616 4907 624 5013
rect 656 4807 664 4913
rect 676 4667 684 4853
rect 716 4807 724 4893
rect 707 4796 724 4807
rect 707 4793 720 4796
rect 736 4727 744 5033
rect 816 4904 824 5233
rect 976 5187 984 5373
rect 996 5327 1004 5473
rect 1156 5447 1164 5533
rect 1176 5507 1184 5613
rect 1216 5387 1224 5673
rect 1236 5407 1244 5773
rect 1316 5767 1324 6013
rect 1676 6007 1684 6053
rect 1756 5947 1764 6293
rect 1956 6267 1964 6353
rect 1993 6344 2007 6353
rect 1993 6340 2024 6344
rect 1996 6336 2024 6340
rect 1776 5967 1784 6213
rect 1836 6147 1844 6173
rect 1876 6147 1884 6253
rect 2016 6207 2024 6336
rect 1956 6087 1964 6193
rect 1996 6147 2004 6173
rect 2047 6136 2073 6144
rect 1896 6047 1904 6073
rect 2056 6007 2064 6073
rect 2096 6047 2104 6113
rect 1796 5967 1804 5993
rect 2136 5987 2144 6053
rect 2176 6004 2184 6053
rect 2216 6007 2224 6453
rect 2296 6447 2304 6473
rect 2356 6207 2364 6373
rect 2396 6367 2404 6453
rect 2756 6427 2764 6493
rect 2500 6424 2513 6427
rect 2496 6413 2513 6424
rect 2447 6364 2460 6367
rect 2447 6353 2464 6364
rect 2167 5996 2184 6004
rect 1356 5847 1364 5933
rect 2016 5927 2024 5973
rect 2016 5916 2033 5927
rect 2020 5913 2033 5916
rect 2060 5924 2073 5927
rect 2056 5913 2073 5924
rect 1427 5904 1440 5907
rect 1427 5893 1444 5904
rect 1820 5904 1833 5907
rect 1727 5896 1764 5904
rect 1436 5847 1444 5893
rect 1407 5844 1420 5847
rect 1407 5833 1424 5844
rect 1416 5807 1424 5833
rect 1356 5707 1364 5793
rect 1516 5707 1524 5833
rect 1556 5807 1564 5833
rect 1576 5687 1584 5893
rect 1616 5807 1624 5893
rect 1696 5767 1704 5833
rect 1736 5687 1744 5833
rect 1756 5787 1764 5896
rect 1816 5893 1833 5904
rect 1816 5687 1824 5893
rect 1856 5787 1864 5833
rect 1896 5807 1904 5833
rect 2056 5827 2064 5913
rect 2116 5867 2124 5953
rect 2156 5884 2164 5993
rect 2296 5987 2304 6073
rect 2376 6007 2384 6133
rect 2456 6127 2464 6353
rect 2496 6327 2504 6413
rect 2676 6367 2684 6413
rect 2520 6364 2533 6367
rect 2516 6360 2533 6364
rect 2513 6353 2533 6360
rect 2676 6356 2693 6367
rect 2680 6353 2693 6356
rect 2513 6347 2527 6353
rect 2496 6287 2504 6313
rect 2400 6124 2413 6127
rect 2396 6113 2413 6124
rect 2396 6047 2404 6113
rect 2436 6007 2444 6053
rect 2196 5927 2204 5953
rect 2240 5924 2253 5927
rect 2236 5913 2253 5924
rect 2156 5876 2184 5884
rect 1907 5796 1924 5804
rect 1476 5627 1484 5653
rect 1616 5627 1624 5653
rect 1467 5616 1484 5627
rect 1560 5624 1573 5627
rect 1467 5613 1480 5616
rect 1556 5613 1573 5624
rect 1316 5527 1324 5553
rect 1416 5527 1424 5613
rect 1556 5567 1564 5613
rect 1696 5567 1704 5653
rect 1816 5627 1824 5673
rect 1916 5627 1924 5796
rect 1940 5624 1953 5627
rect 1936 5613 1953 5624
rect 1136 5344 1144 5373
rect 1116 5336 1144 5344
rect 996 5316 1013 5327
rect 1000 5313 1013 5316
rect 1056 5287 1064 5313
rect 1096 5187 1104 5273
rect 936 5107 944 5173
rect 887 5096 913 5104
rect 936 5096 953 5107
rect 940 5093 953 5096
rect 976 5044 984 5173
rect 1056 5107 1064 5173
rect 1116 5147 1124 5336
rect 1296 5327 1304 5413
rect 1336 5407 1344 5493
rect 1476 5487 1484 5553
rect 1636 5487 1644 5553
rect 1776 5527 1784 5613
rect 1387 5384 1400 5387
rect 1387 5373 1404 5384
rect 1396 5327 1404 5373
rect 1296 5316 1313 5327
rect 1300 5313 1313 5316
rect 1156 5167 1164 5313
rect 1196 5227 1204 5313
rect 1353 5307 1367 5313
rect 1353 5300 1373 5307
rect 1356 5296 1373 5300
rect 1360 5293 1373 5296
rect 1196 5107 1204 5133
rect 1236 5107 1244 5233
rect 1007 5096 1033 5104
rect 1056 5096 1073 5107
rect 1060 5093 1073 5096
rect 947 5036 984 5044
rect 896 4967 904 5013
rect 796 4896 824 4904
rect 796 4687 804 4896
rect 856 4887 864 4913
rect 827 4884 840 4887
rect 827 4873 844 4884
rect 836 4824 844 4873
rect 836 4816 873 4824
rect 576 4587 584 4613
rect 736 4587 744 4653
rect 776 4587 784 4613
rect 376 4576 393 4587
rect 380 4573 393 4576
rect 256 4516 273 4527
rect 260 4513 273 4516
rect 236 4387 244 4513
rect 336 4347 344 4373
rect 336 4336 353 4347
rect 340 4333 353 4336
rect 236 4247 244 4273
rect 276 4187 284 4273
rect 316 4227 324 4333
rect 376 4247 384 4273
rect 396 4187 404 4333
rect 476 4327 484 4573
rect 567 4516 633 4524
rect 756 4487 764 4513
rect 436 4287 444 4313
rect 516 4287 524 4473
rect 776 4407 784 4573
rect 816 4567 824 4633
rect 836 4627 844 4673
rect 427 4276 444 4287
rect 427 4273 440 4276
rect 536 4147 544 4333
rect 556 4227 564 4273
rect 576 4247 584 4333
rect 696 4287 704 4393
rect 856 4387 864 4713
rect 896 4487 904 4953
rect 976 4887 984 4933
rect 920 4884 933 4887
rect 916 4873 933 4884
rect 916 4727 924 4873
rect 1016 4867 1024 4913
rect 1056 4787 1064 5033
rect 1256 5007 1264 5033
rect 1296 5007 1304 5193
rect 1147 4856 1204 4864
rect 1173 4824 1187 4833
rect 1156 4820 1187 4824
rect 1153 4816 1184 4820
rect 1153 4807 1167 4816
rect 1196 4807 1204 4856
rect 916 4384 924 4713
rect 936 4527 944 4613
rect 916 4376 933 4384
rect 736 4347 744 4373
rect 936 4347 944 4373
rect 687 4276 704 4287
rect 687 4273 700 4276
rect 716 4247 724 4273
rect 356 4067 364 4093
rect 167 4056 193 4064
rect 247 4056 273 4064
rect 376 4056 393 4064
rect 313 4044 327 4053
rect 376 4044 384 4056
rect 407 4064 420 4067
rect 407 4053 424 4064
rect 313 4040 384 4044
rect 316 4036 384 4040
rect 416 4007 424 4053
rect 227 4004 240 4007
rect 227 3993 244 4004
rect 116 3947 124 3993
rect 156 3827 164 3933
rect 56 3707 64 3813
rect 96 3667 104 3753
rect 136 3727 144 3753
rect 107 3656 124 3664
rect 76 3547 84 3573
rect 116 3487 124 3656
rect 196 3587 204 3953
rect 236 3907 244 3993
rect 260 3764 273 3767
rect 256 3753 273 3764
rect 236 3707 244 3753
rect 256 3664 264 3753
rect 316 3727 324 3993
rect 456 3907 464 4093
rect 556 4067 564 4093
rect 816 4067 824 4093
rect 856 4067 864 4153
rect 916 4087 924 4273
rect 976 4247 984 4773
rect 996 4267 1004 4633
rect 1056 4587 1064 4693
rect 1116 4607 1124 4793
rect 1216 4767 1224 4993
rect 1236 4867 1244 4933
rect 1296 4807 1304 4893
rect 1256 4767 1264 4793
rect 1080 4584 1093 4587
rect 1076 4573 1093 4584
rect 1076 4564 1084 4573
rect 1056 4556 1084 4564
rect 1036 4447 1044 4513
rect 1056 4287 1064 4556
rect 1096 4287 1104 4453
rect 1116 4407 1124 4513
rect 1156 4487 1164 4753
rect 1216 4627 1224 4673
rect 1256 4587 1264 4653
rect 1200 4584 1213 4587
rect 1196 4573 1213 4584
rect 1196 4407 1204 4573
rect 1276 4527 1284 4613
rect 1260 4524 1273 4527
rect 1256 4513 1273 4524
rect 1216 4447 1224 4513
rect 1256 4467 1264 4513
rect 1187 4393 1204 4407
rect 936 4127 944 4233
rect 1096 4087 1104 4273
rect 1136 4227 1144 4273
rect 1196 4264 1204 4393
rect 1316 4387 1324 5253
rect 1396 5147 1404 5213
rect 1340 5104 1353 5107
rect 1336 5093 1353 5104
rect 1336 5047 1344 5093
rect 1376 5047 1384 5133
rect 1416 5107 1424 5233
rect 1436 5187 1444 5473
rect 1536 5387 1544 5473
rect 1467 5356 1524 5364
rect 1516 5327 1524 5356
rect 1527 5324 1540 5327
rect 1527 5320 1544 5324
rect 1527 5313 1547 5320
rect 1476 5267 1484 5313
rect 1533 5307 1547 5313
rect 1576 5307 1584 5373
rect 1536 5187 1544 5233
rect 1516 5107 1524 5133
rect 1407 5096 1424 5107
rect 1407 5093 1420 5096
rect 1427 5036 1464 5044
rect 1336 4387 1344 4993
rect 1456 4987 1464 5036
rect 1456 4867 1464 4933
rect 1396 4587 1404 4693
rect 1496 4584 1504 5013
rect 1556 5007 1564 5093
rect 1536 4996 1553 5004
rect 1536 4947 1544 4996
rect 1576 4947 1584 5033
rect 1636 4987 1644 5473
rect 1796 5467 1804 5553
rect 1856 5507 1864 5613
rect 1676 5404 1684 5433
rect 1656 5396 1684 5404
rect 1656 5344 1664 5396
rect 1716 5387 1724 5413
rect 1707 5376 1724 5387
rect 1707 5373 1720 5376
rect 1656 5340 1684 5344
rect 1656 5336 1687 5340
rect 1673 5327 1687 5336
rect 1716 5267 1724 5313
rect 1796 5247 1804 5373
rect 1856 5327 1864 5493
rect 1876 5387 1884 5593
rect 1936 5464 1944 5613
rect 1996 5567 2004 5673
rect 1987 5556 2004 5567
rect 1987 5553 2000 5556
rect 2056 5547 2064 5673
rect 2076 5647 2084 5853
rect 2096 5667 2104 5813
rect 1996 5487 2004 5513
rect 2096 5507 2104 5533
rect 2076 5496 2093 5504
rect 1936 5456 1953 5464
rect 1816 5207 1824 5313
rect 1616 4976 1633 4984
rect 1516 4807 1524 4893
rect 1576 4807 1584 4933
rect 1616 4907 1624 4976
rect 1676 4887 1684 4953
rect 1696 4947 1704 5093
rect 1733 5084 1747 5093
rect 1716 5080 1747 5084
rect 1716 5076 1744 5080
rect 1716 5007 1724 5076
rect 1716 4964 1724 4993
rect 1756 4987 1764 5033
rect 1716 4956 1744 4964
rect 1736 4927 1744 4956
rect 1516 4796 1533 4807
rect 1520 4793 1533 4796
rect 1516 4607 1524 4733
rect 1536 4687 1544 4713
rect 1616 4667 1624 4753
rect 1556 4587 1564 4613
rect 1596 4587 1604 4653
rect 1496 4576 1524 4584
rect 1447 4564 1460 4567
rect 1447 4553 1464 4564
rect 1356 4447 1364 4553
rect 1456 4527 1464 4553
rect 1376 4407 1384 4493
rect 1416 4467 1424 4493
rect 1476 4367 1484 4453
rect 1467 4356 1484 4367
rect 1467 4353 1480 4356
rect 1413 4344 1427 4353
rect 1307 4336 1344 4344
rect 1216 4287 1224 4333
rect 1216 4276 1233 4287
rect 1220 4273 1233 4276
rect 1287 4284 1300 4287
rect 1287 4273 1304 4284
rect 1196 4256 1244 4264
rect 1236 4227 1244 4256
rect 516 3927 524 4053
rect 556 3867 564 4053
rect 696 3967 704 3993
rect 616 3827 624 3913
rect 736 3847 744 4053
rect 796 3887 804 4053
rect 916 3996 984 4004
rect 836 3967 844 3993
rect 916 3967 924 3996
rect 976 3987 984 3996
rect 996 3987 1004 4033
rect 947 3984 960 3987
rect 947 3973 964 3984
rect 987 3976 1004 3987
rect 987 3973 1000 3976
rect 907 3956 924 3967
rect 907 3953 920 3956
rect 956 3907 964 3973
rect 1036 3907 1044 4073
rect 1176 4007 1184 4133
rect 1256 4084 1264 4193
rect 1296 4147 1304 4273
rect 1316 4167 1324 4193
rect 1256 4076 1284 4084
rect 1096 3947 1104 3973
rect 387 3816 424 3824
rect 396 3687 404 3753
rect 236 3660 264 3664
rect 236 3656 267 3660
rect 107 3476 124 3487
rect 107 3473 120 3476
rect 196 3347 204 3573
rect 236 3527 244 3656
rect 253 3647 267 3656
rect 276 3547 284 3673
rect 316 3547 324 3573
rect 396 3547 404 3673
rect 416 3587 424 3816
rect 447 3756 484 3764
rect 416 3487 424 3573
rect 56 3067 64 3293
rect 96 3247 104 3333
rect 256 3307 264 3333
rect 136 3187 144 3233
rect 96 3027 104 3053
rect 96 2807 104 3013
rect 127 2964 140 2967
rect 127 2953 144 2964
rect 136 2807 144 2953
rect 136 2707 144 2793
rect 96 2447 104 2693
rect 136 2507 144 2553
rect 176 2547 184 2833
rect 216 2764 224 3193
rect 236 3187 244 3233
rect 276 3207 284 3233
rect 316 3027 324 3293
rect 376 3247 384 3473
rect 436 3347 444 3513
rect 456 3367 464 3713
rect 476 3647 484 3756
rect 516 3587 524 3813
rect 640 3804 653 3807
rect 636 3793 653 3804
rect 636 3767 644 3793
rect 596 3727 604 3753
rect 556 3487 564 3653
rect 596 3547 604 3573
rect 636 3447 644 3533
rect 436 3247 444 3333
rect 536 3307 544 3333
rect 596 3327 604 3393
rect 536 3296 553 3307
rect 540 3293 553 3296
rect 376 3236 393 3247
rect 380 3233 393 3236
rect 396 3207 404 3233
rect 476 3027 484 3293
rect 536 3207 544 3233
rect 576 3107 584 3233
rect 636 3187 644 3293
rect 676 3247 684 3833
rect 776 3747 784 3833
rect 876 3827 884 3873
rect 916 3847 924 3893
rect 967 3824 980 3827
rect 967 3813 984 3824
rect 736 3627 744 3733
rect 856 3727 864 3773
rect 896 3727 904 3753
rect 936 3727 944 3753
rect 976 3747 984 3813
rect 936 3647 944 3713
rect 736 3547 744 3613
rect 776 3547 784 3633
rect 996 3584 1004 3893
rect 1056 3747 1064 3833
rect 1056 3687 1064 3733
rect 1096 3727 1104 3833
rect 1116 3787 1124 3913
rect 1136 3827 1144 3973
rect 1196 3804 1204 3953
rect 1256 3827 1264 3933
rect 1176 3796 1204 3804
rect 1176 3767 1184 3796
rect 1276 3767 1284 4076
rect 1296 3907 1304 4053
rect 1336 4007 1344 4336
rect 1376 4340 1427 4344
rect 1376 4336 1424 4340
rect 1356 4067 1364 4213
rect 1376 3884 1384 4336
rect 1396 4267 1404 4293
rect 1436 4147 1444 4273
rect 1456 4167 1464 4253
rect 1476 4147 1484 4293
rect 1496 4267 1504 4433
rect 1516 4347 1524 4576
rect 1607 4584 1620 4587
rect 1607 4573 1624 4584
rect 1616 4547 1624 4573
rect 1636 4467 1644 4753
rect 1716 4747 1724 4873
rect 1796 4847 1804 4973
rect 1856 4887 1864 5213
rect 1916 5187 1924 5233
rect 1876 5107 1884 5133
rect 1916 5107 1924 5173
rect 1956 5084 1964 5453
rect 2036 5387 2044 5433
rect 2027 5324 2040 5327
rect 2027 5320 2044 5324
rect 2027 5313 2047 5320
rect 1976 5227 1984 5313
rect 2033 5307 2047 5313
rect 2076 5247 2084 5496
rect 2156 5464 2164 5753
rect 2176 5727 2184 5876
rect 2236 5787 2244 5913
rect 2316 5867 2324 5993
rect 2496 5987 2504 6053
rect 2516 6007 2524 6213
rect 2356 5907 2364 5933
rect 2396 5927 2404 5953
rect 2536 5907 2544 6313
rect 2576 6227 2584 6353
rect 2696 6247 2704 6353
rect 2736 6327 2744 6353
rect 2776 6327 2784 6373
rect 2556 5927 2564 6173
rect 2616 6147 2624 6173
rect 2576 5987 2584 6073
rect 2527 5896 2544 5907
rect 2527 5893 2540 5896
rect 2356 5856 2424 5864
rect 2276 5827 2284 5853
rect 2356 5804 2364 5856
rect 2416 5847 2424 5856
rect 2427 5844 2440 5847
rect 2427 5833 2444 5844
rect 2376 5807 2384 5833
rect 2436 5827 2444 5833
rect 2436 5816 2453 5827
rect 2440 5813 2453 5816
rect 2336 5796 2364 5804
rect 2336 5784 2344 5796
rect 2536 5787 2544 5833
rect 2306 5776 2344 5784
rect 2173 5624 2187 5633
rect 2236 5627 2244 5733
rect 2173 5620 2213 5624
rect 2176 5616 2213 5620
rect 2236 5613 2253 5627
rect 2236 5527 2244 5613
rect 2147 5456 2164 5464
rect 2136 5407 2144 5453
rect 2276 5427 2284 5553
rect 2173 5384 2187 5393
rect 2156 5380 2187 5384
rect 2156 5376 2184 5380
rect 2116 5267 2124 5333
rect 1936 5076 1964 5084
rect 1896 5007 1904 5033
rect 1396 4067 1404 4093
rect 1536 4067 1544 4093
rect 1480 4064 1493 4067
rect 1476 4053 1493 4064
rect 1436 4007 1444 4053
rect 1427 3996 1444 4007
rect 1427 3993 1440 3996
rect 1476 3967 1484 4053
rect 1596 4007 1604 4273
rect 1376 3876 1393 3884
rect 1396 3767 1404 3873
rect 1196 3727 1204 3753
rect 1236 3727 1244 3753
rect 1096 3664 1104 3713
rect 987 3576 1004 3584
rect 1076 3656 1104 3664
rect 896 3547 904 3573
rect 947 3544 960 3547
rect 947 3533 964 3544
rect 956 3507 964 3533
rect 807 3484 820 3487
rect 807 3473 824 3484
rect 716 3387 724 3473
rect 816 3447 824 3473
rect 736 3247 744 3353
rect 776 3307 784 3373
rect 876 3327 884 3433
rect 916 3327 924 3413
rect 776 3296 793 3307
rect 780 3293 793 3296
rect 976 3267 984 3573
rect 1076 3467 1084 3656
rect 1036 3387 1044 3453
rect 1016 3307 1024 3333
rect 1036 3247 1044 3373
rect 1076 3307 1084 3453
rect 1096 3387 1104 3413
rect 776 3187 784 3233
rect 236 3020 273 3024
rect 233 3016 273 3020
rect 233 3007 247 3016
rect 256 2907 264 3016
rect 527 3024 540 3027
rect 527 3013 544 3024
rect 316 2827 324 3013
rect 336 2927 344 2953
rect 396 2827 404 2913
rect 256 2787 264 2813
rect 316 2787 324 2813
rect 316 2776 333 2787
rect 320 2773 333 2776
rect 216 2756 244 2764
rect 196 2687 204 2733
rect 176 2507 184 2533
rect 116 2267 124 2413
rect 156 2407 164 2433
rect 116 2256 133 2267
rect 120 2253 133 2256
rect 116 1927 124 2033
rect 116 1747 124 1773
rect 76 1567 84 1673
rect 76 1467 84 1553
rect 156 1467 164 2253
rect 196 1787 204 2433
rect 236 2424 244 2756
rect 396 2727 404 2813
rect 456 2787 464 2873
rect 496 2867 504 2953
rect 536 2904 544 3013
rect 676 3007 684 3153
rect 536 2896 553 2904
rect 496 2787 504 2853
rect 556 2787 564 2893
rect 576 2847 584 2993
rect 647 2956 693 2964
rect 756 2827 764 3073
rect 796 2907 804 3013
rect 816 2927 824 3093
rect 836 3067 844 3173
rect 836 3027 844 3053
rect 876 3027 884 3053
rect 856 2927 864 2953
rect 896 2787 904 2833
rect 596 2727 604 2773
rect 693 2764 707 2773
rect 887 2776 904 2787
rect 887 2773 900 2776
rect 733 2764 747 2773
rect 693 2760 747 2764
rect 696 2756 744 2760
rect 340 2724 353 2727
rect 336 2720 353 2724
rect 333 2713 353 2720
rect 587 2716 604 2727
rect 587 2713 600 2716
rect 333 2707 347 2713
rect 536 2687 544 2713
rect 296 2507 304 2533
rect 336 2507 344 2553
rect 496 2507 504 2573
rect 216 2416 244 2424
rect 216 2207 224 2416
rect 316 2407 324 2433
rect 456 2407 464 2493
rect 487 2444 500 2447
rect 487 2433 504 2444
rect 216 1807 224 2193
rect 256 1987 264 2173
rect 276 2107 284 2253
rect 376 2227 384 2393
rect 416 2267 424 2353
rect 436 2167 444 2193
rect 307 1976 333 1984
rect 436 1927 444 2013
rect 236 1827 244 1893
rect 276 1887 284 1913
rect 176 1776 193 1784
rect 176 1507 184 1776
rect 316 1747 324 1853
rect 196 1547 204 1713
rect 216 1527 224 1673
rect 256 1647 264 1673
rect 276 1467 284 1553
rect 100 1464 113 1467
rect 96 1453 113 1464
rect 207 1456 233 1464
rect 96 1444 104 1453
rect 76 1436 104 1444
rect 76 1384 84 1436
rect 156 1404 164 1453
rect 107 1396 164 1404
rect 76 1376 104 1384
rect 96 1167 104 1376
rect 116 1227 124 1313
rect 136 1307 144 1373
rect 256 1367 264 1393
rect 176 1227 184 1333
rect 216 1287 224 1333
rect 227 1216 253 1224
rect 316 1167 324 1353
rect 96 1153 113 1167
rect 167 1164 180 1167
rect 260 1164 273 1167
rect 167 1160 184 1164
rect 256 1160 273 1164
rect 167 1153 187 1160
rect 96 887 104 1153
rect 173 1147 187 1153
rect 253 1153 273 1160
rect 253 1147 267 1153
rect 316 1107 324 1153
rect 156 947 164 973
rect 116 827 124 933
rect 136 764 144 873
rect 196 807 204 873
rect 127 756 144 764
rect 116 707 124 753
rect 116 427 124 513
rect 156 467 164 733
rect 196 647 204 793
rect 236 727 244 1093
rect 336 947 344 1813
rect 356 1767 364 1813
rect 396 1767 404 1793
rect 356 1407 364 1633
rect 436 1484 444 1873
rect 476 1867 484 2373
rect 496 2267 504 2433
rect 536 2387 544 2633
rect 636 2507 644 2673
rect 580 2504 593 2507
rect 576 2493 593 2504
rect 576 2407 584 2493
rect 556 2207 564 2293
rect 596 2207 604 2353
rect 636 2267 644 2493
rect 676 2447 684 2533
rect 736 2507 744 2733
rect 816 2687 824 2713
rect 776 2507 784 2533
rect 796 2447 804 2553
rect 856 2547 864 2713
rect 896 2587 904 2713
rect 916 2444 924 3153
rect 936 2967 944 3053
rect 936 2587 944 2893
rect 956 2787 964 2833
rect 896 2440 924 2444
rect 893 2436 924 2440
rect 713 2424 727 2433
rect 893 2427 907 2436
rect 936 2427 944 2533
rect 713 2420 744 2424
rect 716 2416 744 2420
rect 680 2264 693 2267
rect 676 2253 693 2264
rect 556 2167 564 2193
rect 536 1987 544 2013
rect 576 1987 584 2093
rect 616 2047 624 2153
rect 616 1927 624 2033
rect 676 2027 684 2253
rect 716 2167 724 2193
rect 736 2184 744 2416
rect 896 2364 904 2413
rect 896 2356 924 2364
rect 776 2267 784 2313
rect 796 2204 804 2333
rect 856 2287 864 2313
rect 896 2287 904 2333
rect 767 2196 804 2204
rect 736 2176 764 2184
rect 607 1916 624 1927
rect 607 1913 620 1916
rect 456 1507 464 1693
rect 496 1687 504 1813
rect 536 1687 544 1773
rect 576 1527 584 1733
rect 616 1707 624 1813
rect 656 1787 664 1953
rect 716 1907 724 2113
rect 756 1907 764 2176
rect 816 2107 824 2213
rect 916 2127 924 2356
rect 936 2267 944 2313
rect 796 1927 804 2013
rect 876 2004 884 2073
rect 856 2000 884 2004
rect 853 1996 884 2000
rect 853 1987 867 1996
rect 896 1987 904 2093
rect 976 2088 984 2953
rect 996 2507 1004 3213
rect 1076 3087 1084 3293
rect 1016 3016 1053 3024
rect 1016 2887 1024 3016
rect 1060 2964 1073 2967
rect 1056 2953 1073 2964
rect 1056 2907 1064 2953
rect 1096 2927 1104 3373
rect 1136 3127 1144 3713
rect 1156 3367 1164 3673
rect 1256 3587 1264 3613
rect 1256 3547 1264 3573
rect 1176 3540 1213 3544
rect 1173 3536 1213 3540
rect 1173 3527 1187 3536
rect 1276 3404 1284 3473
rect 1256 3400 1284 3404
rect 1253 3396 1284 3400
rect 1253 3387 1267 3396
rect 1156 3207 1164 3233
rect 1156 2967 1164 3153
rect 1216 3027 1224 3233
rect 1276 3184 1284 3353
rect 1316 3247 1324 3393
rect 1336 3327 1344 3373
rect 1356 3347 1364 3753
rect 1376 3547 1384 3593
rect 1376 3367 1384 3473
rect 1353 3224 1367 3233
rect 1336 3220 1367 3224
rect 1336 3216 1364 3220
rect 1336 3187 1344 3216
rect 1276 3176 1304 3184
rect 1256 3027 1264 3093
rect 1187 3024 1200 3027
rect 1187 3013 1204 3024
rect 1076 2727 1084 2873
rect 1116 2867 1124 2893
rect 1116 2727 1124 2853
rect 1196 2787 1204 3013
rect 1196 2773 1213 2787
rect 1216 2687 1224 2773
rect 1076 2647 1084 2673
rect 1296 2647 1304 3176
rect 1336 2967 1344 3173
rect 1356 3027 1364 3113
rect 1396 3067 1404 3753
rect 1416 3547 1424 3593
rect 1420 3484 1433 3487
rect 1416 3473 1433 3484
rect 1416 3447 1424 3473
rect 1456 3464 1464 3713
rect 1476 3667 1484 3953
rect 1496 3707 1504 3813
rect 1436 3456 1464 3464
rect 1407 3056 1424 3064
rect 1367 3024 1380 3027
rect 1367 3013 1384 3024
rect 1336 2887 1344 2953
rect 1356 2667 1364 2713
rect 1016 2507 1024 2533
rect 1056 2507 1064 2613
rect 1196 2567 1204 2633
rect 996 2493 1013 2507
rect 996 2087 1004 2493
rect 1016 2348 1024 2433
rect 1016 2207 1024 2312
rect 1056 2207 1064 2313
rect 756 1867 764 1893
rect 936 1827 944 2013
rect 656 1747 664 1773
rect 436 1476 464 1484
rect 420 1464 433 1467
rect 416 1453 433 1464
rect 356 1347 364 1393
rect 416 1327 424 1453
rect 456 1424 464 1476
rect 576 1467 584 1513
rect 616 1467 624 1493
rect 487 1464 500 1467
rect 487 1453 504 1464
rect 436 1416 464 1424
rect 396 1227 404 1273
rect 436 964 444 1416
rect 496 1407 504 1453
rect 636 1407 644 1493
rect 736 1467 744 1693
rect 796 1687 804 1813
rect 816 1747 824 1773
rect 796 1467 804 1493
rect 736 1456 753 1467
rect 740 1453 753 1456
rect 896 1464 904 1693
rect 916 1507 924 1733
rect 976 1687 984 2052
rect 1036 1927 1044 2133
rect 1096 2067 1104 2353
rect 1136 2167 1144 2513
rect 1156 2487 1164 2533
rect 1216 2504 1224 2533
rect 1196 2496 1224 2504
rect 1196 2444 1204 2496
rect 1256 2487 1264 2573
rect 1247 2476 1264 2487
rect 1247 2473 1260 2476
rect 1196 2440 1224 2444
rect 1196 2436 1227 2440
rect 1213 2427 1227 2436
rect 1187 2424 1200 2427
rect 1187 2413 1204 2424
rect 1196 2347 1204 2413
rect 1236 2327 1244 2473
rect 1276 2367 1284 2593
rect 1376 2587 1384 3013
rect 1396 2687 1404 2713
rect 1416 2647 1424 3056
rect 1436 2627 1444 3456
rect 1456 3187 1464 3233
rect 1476 3167 1484 3293
rect 1476 3087 1484 3153
rect 1496 2787 1504 3013
rect 1216 2267 1224 2293
rect 1156 2044 1164 2193
rect 1147 2036 1164 2044
rect 1136 1987 1144 2033
rect 1176 2027 1184 2253
rect 1196 2167 1204 2193
rect 1196 1987 1204 2013
rect 1256 1987 1264 2033
rect 1296 2027 1304 2193
rect 1316 2167 1324 2513
rect 1336 2487 1344 2573
rect 1436 2567 1444 2613
rect 1336 2476 1353 2487
rect 1340 2473 1353 2476
rect 1396 2427 1404 2553
rect 1516 2487 1524 3653
rect 1536 3607 1544 3753
rect 1536 3547 1544 3593
rect 1556 3587 1564 3813
rect 1576 3447 1584 3533
rect 1616 3327 1624 4433
rect 1676 4387 1684 4733
rect 1696 4607 1704 4633
rect 1667 4344 1680 4347
rect 1667 4333 1684 4344
rect 1676 4307 1684 4333
rect 1636 4147 1644 4273
rect 1696 4127 1704 4593
rect 1736 4527 1744 4833
rect 1876 4807 1884 4973
rect 1836 4744 1844 4793
rect 1816 4736 1844 4744
rect 1736 4407 1744 4513
rect 1776 4507 1784 4553
rect 1816 4487 1824 4736
rect 1656 4067 1664 4113
rect 1696 3967 1704 4053
rect 1736 3967 1744 4393
rect 1836 4387 1844 4693
rect 1876 4607 1884 4793
rect 1856 4507 1864 4553
rect 1936 4527 1944 5076
rect 2016 5047 2024 5173
rect 2076 5107 2084 5233
rect 2036 5007 2044 5093
rect 2096 5047 2104 5133
rect 1976 4687 1984 4853
rect 2036 4807 2044 4953
rect 1956 4680 1973 4684
rect 1953 4676 1973 4680
rect 1953 4667 1967 4676
rect 1996 4667 2004 4793
rect 2036 4707 2044 4793
rect 2076 4767 2084 4993
rect 2116 4907 2124 5253
rect 2156 5227 2164 5376
rect 2136 5007 2144 5193
rect 2196 5147 2204 5333
rect 2296 5307 2304 5733
rect 2336 5567 2344 5753
rect 2356 5687 2364 5773
rect 2536 5747 2544 5773
rect 2356 5607 2364 5673
rect 2496 5567 2504 5733
rect 2556 5627 2564 5773
rect 2576 5727 2584 5833
rect 2616 5767 2624 5833
rect 2656 5807 2664 6133
rect 2576 5667 2584 5713
rect 2336 5487 2344 5553
rect 2516 5527 2524 5613
rect 2436 5487 2444 5513
rect 2536 5507 2544 5553
rect 2396 5387 2404 5473
rect 2596 5467 2604 5693
rect 2656 5627 2664 5793
rect 2676 5787 2684 6073
rect 2716 5967 2724 6313
rect 2816 6307 2824 6473
rect 2856 6447 2864 6473
rect 2896 6347 2904 6433
rect 2936 6367 2944 6493
rect 3176 6447 3184 6473
rect 3067 6424 3080 6427
rect 3067 6413 3084 6424
rect 3076 6347 3084 6413
rect 2816 6267 2824 6293
rect 2736 6087 2744 6173
rect 2756 6147 2764 6233
rect 2816 6147 2824 6253
rect 2836 6227 2844 6333
rect 2756 6136 2773 6147
rect 2760 6133 2773 6136
rect 2836 6087 2844 6213
rect 2756 5907 2764 6033
rect 2727 5896 2753 5904
rect 2816 5847 2824 5933
rect 2876 5907 2884 6233
rect 2867 5896 2884 5907
rect 2867 5893 2880 5896
rect 2816 5836 2833 5847
rect 2820 5833 2833 5836
rect 2876 5787 2884 5833
rect 2696 5527 2704 5613
rect 2736 5567 2744 5773
rect 2776 5627 2784 5753
rect 2836 5627 2844 5673
rect 2776 5616 2793 5627
rect 2780 5613 2793 5616
rect 2876 5567 2884 5653
rect 2727 5556 2744 5567
rect 2727 5553 2740 5556
rect 2413 5404 2427 5413
rect 2413 5400 2453 5404
rect 2416 5396 2453 5400
rect 2387 5376 2404 5387
rect 2387 5373 2400 5376
rect 2336 5187 2344 5313
rect 2236 5107 2244 5153
rect 2256 5107 2264 5173
rect 2227 5096 2244 5107
rect 2227 5093 2240 5096
rect 2336 5047 2344 5173
rect 2396 5107 2404 5233
rect 2353 5084 2367 5093
rect 2353 5080 2384 5084
rect 2356 5076 2384 5080
rect 2176 4964 2184 5033
rect 2156 4956 2184 4964
rect 2156 4927 2164 4956
rect 2236 4947 2244 5033
rect 2196 4867 2204 4933
rect 2316 4927 2324 4973
rect 2376 4947 2384 5076
rect 2416 4967 2424 5193
rect 2436 5047 2444 5133
rect 2107 4856 2133 4864
rect 2216 4807 2224 4853
rect 2207 4796 2224 4807
rect 2207 4793 2220 4796
rect 1856 4407 1864 4493
rect 1756 4204 1764 4373
rect 1776 4287 1784 4373
rect 1847 4344 1860 4347
rect 1876 4344 1884 4473
rect 1896 4447 1904 4513
rect 1956 4447 1964 4613
rect 2036 4587 2044 4613
rect 2056 4587 2064 4673
rect 2156 4607 2164 4793
rect 2056 4576 2073 4587
rect 2060 4573 2073 4576
rect 2160 4564 2173 4567
rect 2156 4553 2173 4564
rect 2080 4544 2093 4547
rect 2076 4533 2093 4544
rect 1996 4407 2004 4513
rect 1956 4367 1964 4393
rect 2036 4384 2044 4473
rect 1996 4376 2044 4384
rect 1996 4367 2004 4376
rect 1947 4356 1964 4367
rect 1947 4353 1960 4356
rect 1987 4356 2004 4367
rect 1987 4353 2000 4356
rect 1847 4336 1884 4344
rect 1847 4333 1864 4336
rect 1776 4227 1784 4273
rect 1816 4227 1824 4273
rect 1756 4196 1784 4204
rect 1776 4127 1784 4196
rect 1736 3787 1744 3953
rect 1816 3827 1824 4173
rect 1856 4107 1864 4333
rect 1916 4227 1924 4293
rect 1876 4047 1884 4179
rect 1916 4167 1924 4213
rect 1956 4147 1964 4273
rect 1976 4127 1984 4233
rect 1996 4147 2004 4293
rect 2076 4227 2084 4533
rect 2156 4527 2164 4553
rect 2196 4507 2204 4753
rect 2236 4567 2244 4893
rect 2256 4667 2264 4893
rect 2276 4667 2284 4873
rect 2316 4807 2324 4913
rect 2356 4767 2364 4793
rect 2396 4747 2404 4873
rect 2456 4827 2464 4873
rect 2476 4867 2484 5313
rect 2496 5287 2504 5393
rect 2536 5384 2544 5453
rect 2636 5407 2644 5433
rect 2516 5376 2544 5384
rect 2496 5247 2504 5273
rect 2516 5007 2524 5376
rect 2593 5364 2607 5373
rect 2576 5360 2607 5364
rect 2576 5356 2604 5360
rect 2576 5187 2584 5356
rect 2676 5344 2684 5433
rect 2736 5387 2744 5473
rect 2736 5376 2753 5387
rect 2740 5373 2753 5376
rect 2676 5336 2704 5344
rect 2616 5147 2624 5313
rect 2656 5207 2664 5313
rect 2696 5227 2704 5336
rect 2776 5167 2784 5313
rect 2536 5107 2544 5133
rect 2576 5067 2584 5093
rect 2616 5087 2624 5133
rect 2576 5056 2593 5067
rect 2580 5053 2593 5056
rect 2476 4856 2493 4867
rect 2480 4853 2493 4856
rect 2536 4827 2544 4873
rect 2527 4816 2544 4827
rect 2527 4813 2540 4816
rect 2387 4736 2404 4747
rect 2387 4733 2400 4736
rect 2236 4553 2253 4567
rect 2236 4524 2244 4553
rect 2296 4527 2304 4713
rect 2216 4516 2244 4524
rect 2176 4407 2184 4453
rect 2216 4387 2224 4516
rect 2247 4504 2260 4507
rect 2247 4493 2264 4504
rect 2100 4344 2113 4347
rect 2096 4333 2113 4344
rect 2096 4267 2104 4333
rect 2120 4284 2133 4287
rect 2116 4273 2133 4284
rect 2116 4187 2124 4273
rect 1836 3887 1844 3993
rect 1656 3547 1664 3593
rect 1676 3448 1684 3473
rect 1536 3207 1544 3313
rect 1676 3307 1684 3412
rect 1736 3307 1744 3713
rect 1816 3607 1824 3773
rect 1856 3667 1864 3753
rect 1916 3727 1924 4093
rect 1936 3867 1944 4113
rect 1976 4067 1984 4113
rect 2016 4067 2024 4093
rect 2056 3887 2064 4153
rect 2076 4047 2084 4113
rect 1976 3727 1984 3773
rect 1836 3547 1844 3573
rect 1860 3544 1873 3547
rect 1856 3533 1873 3544
rect 1967 3536 1993 3544
rect 1856 3524 1864 3533
rect 1807 3516 1864 3524
rect 1816 3387 1824 3433
rect 1876 3387 1884 3473
rect 1916 3407 1924 3533
rect 2016 3504 2024 3813
rect 1996 3496 2024 3504
rect 1816 3307 1824 3373
rect 1976 3367 1984 3473
rect 1667 3296 1684 3307
rect 1667 3293 1680 3296
rect 1587 3256 1613 3264
rect 1536 2727 1544 3193
rect 1556 2807 1564 2833
rect 1576 2727 1584 3053
rect 1616 3027 1624 3073
rect 1656 3027 1664 3073
rect 1696 3067 1704 3293
rect 1596 2847 1604 2953
rect 1636 2887 1644 2953
rect 1736 2947 1744 3253
rect 1876 3247 1884 3333
rect 1936 3307 1944 3333
rect 1996 3264 2004 3496
rect 2036 3428 2044 3533
rect 2016 3287 2024 3373
rect 2036 3307 2044 3392
rect 2116 3367 2124 4133
rect 2136 4007 2144 4233
rect 2156 4147 2164 4213
rect 2176 4107 2184 4193
rect 2176 4047 2184 4093
rect 2236 4047 2244 4453
rect 2256 4407 2264 4493
rect 2316 4467 2324 4713
rect 2356 4587 2364 4653
rect 2256 4167 2264 4393
rect 2276 4347 2284 4413
rect 2287 4336 2313 4344
rect 2296 4207 2304 4273
rect 2336 4087 2344 4413
rect 2136 3727 2144 3993
rect 2216 3844 2224 3993
rect 2316 3927 2324 3993
rect 2296 3887 2304 3913
rect 2336 3887 2344 3953
rect 2356 3947 2364 4053
rect 2396 3907 2404 4693
rect 2416 4067 2424 4713
rect 2436 4427 2444 4773
rect 2456 4687 2464 4753
rect 2556 4747 2564 4993
rect 2636 4787 2644 4973
rect 2607 4564 2620 4567
rect 2607 4553 2624 4564
rect 2536 4447 2544 4553
rect 2616 4467 2624 4553
rect 2493 4344 2507 4353
rect 2476 4340 2507 4344
rect 2476 4336 2504 4340
rect 2476 4324 2484 4336
rect 2456 4316 2484 4324
rect 2456 4307 2464 4316
rect 2447 4296 2464 4307
rect 2480 4304 2493 4307
rect 2447 4293 2460 4296
rect 2476 4293 2493 4304
rect 2476 4167 2484 4293
rect 2416 4056 2433 4067
rect 2420 4053 2433 4056
rect 2216 3836 2244 3844
rect 2200 3824 2213 3827
rect 2196 3813 2213 3824
rect 2196 3767 2204 3813
rect 2236 3767 2244 3836
rect 2376 3827 2384 3893
rect 2236 3727 2244 3753
rect 2276 3707 2284 3753
rect 2396 3727 2404 3753
rect 2416 3704 2424 3813
rect 2436 3784 2444 4053
rect 2456 4024 2464 4153
rect 2496 4044 2504 4253
rect 2516 4107 2524 4393
rect 2656 4367 2664 4473
rect 2676 4407 2684 5113
rect 2736 5087 2744 5113
rect 2696 5007 2704 5033
rect 2720 4904 2733 4907
rect 2716 4893 2733 4904
rect 2716 4887 2724 4893
rect 2707 4876 2724 4887
rect 2707 4873 2720 4876
rect 2696 4707 2704 4873
rect 2736 4747 2744 4853
rect 2776 4844 2784 5113
rect 2796 5027 2804 5453
rect 2836 4967 2844 5273
rect 2856 4847 2864 5453
rect 2896 5327 2904 5733
rect 2936 5724 2944 6133
rect 2956 6047 2964 6073
rect 2996 5984 3004 6193
rect 3056 6147 3064 6173
rect 3076 6087 3084 6293
rect 3156 6227 3164 6373
rect 3196 6287 3204 6353
rect 3216 6347 3224 6433
rect 3256 6387 3264 6493
rect 3316 6447 3324 6564
rect 3247 6376 3264 6387
rect 3247 6373 3260 6376
rect 2976 5976 3004 5984
rect 2976 5747 2984 5976
rect 3036 5847 3044 5933
rect 3136 5907 3144 5953
rect 3176 5947 3184 6233
rect 3316 6187 3324 6433
rect 3376 6347 3384 6433
rect 3416 6427 3424 6493
rect 3416 6207 3424 6333
rect 3376 6147 3384 6193
rect 3416 6147 3424 6193
rect 3196 6140 3233 6144
rect 3193 6136 3233 6140
rect 3193 6127 3207 6136
rect 3287 6144 3300 6147
rect 3287 6133 3304 6144
rect 3296 6087 3304 6133
rect 3456 6104 3464 6173
rect 3436 6100 3464 6104
rect 3433 6096 3464 6100
rect 3433 6087 3447 6096
rect 3476 6087 3484 6193
rect 3496 6147 3504 6564
rect 3976 6527 3984 6564
rect 3536 6427 3544 6453
rect 3576 6427 3584 6473
rect 3656 6367 3664 6453
rect 3067 5896 3104 5904
rect 2996 5807 3004 5833
rect 3096 5787 3104 5896
rect 3156 5787 3164 5853
rect 3216 5787 3224 6013
rect 3256 5844 3264 5973
rect 3276 5867 3284 5993
rect 3256 5836 3284 5844
rect 2916 5716 2944 5724
rect 2916 5707 2924 5716
rect 2916 5427 2924 5693
rect 3156 5627 3164 5673
rect 3176 5627 3184 5693
rect 2940 5624 2953 5627
rect 2936 5613 2953 5624
rect 3007 5616 3064 5624
rect 2936 5587 2944 5613
rect 3056 5567 3064 5616
rect 3147 5613 3164 5627
rect 2936 5327 2944 5413
rect 2896 5027 2904 5313
rect 2956 5287 2964 5373
rect 2916 5107 2924 5273
rect 2876 4907 2884 4993
rect 2916 4947 2924 4993
rect 2776 4836 2804 4844
rect 2796 4824 2804 4836
rect 2796 4816 2824 4824
rect 2756 4767 2764 4813
rect 2816 4807 2824 4816
rect 2816 4796 2833 4807
rect 2820 4793 2833 4796
rect 2796 4727 2804 4793
rect 2876 4667 2884 4713
rect 2896 4647 2904 4693
rect 2716 4587 2724 4633
rect 2736 4448 2744 4493
rect 2536 4147 2544 4193
rect 2576 4084 2584 4253
rect 2596 4227 2604 4293
rect 2616 4147 2624 4353
rect 2736 4347 2744 4412
rect 2756 4324 2764 4613
rect 2856 4607 2864 4633
rect 2916 4587 2924 4853
rect 2936 4587 2944 5233
rect 2976 5027 2984 5413
rect 2996 5187 3004 5373
rect 3016 5307 3024 5553
rect 3036 5387 3044 5493
rect 3076 5407 3084 5513
rect 3116 5447 3124 5473
rect 3116 5407 3124 5433
rect 3056 5287 3064 5333
rect 3076 5227 3084 5393
rect 3136 5307 3144 5333
rect 3096 5167 3104 5273
rect 3156 5267 3164 5613
rect 3196 5567 3204 5713
rect 3176 5307 3184 5433
rect 3196 5288 3204 5553
rect 3236 5424 3244 5753
rect 3216 5416 3244 5424
rect 3216 5327 3224 5416
rect 3256 5407 3264 5733
rect 3276 5467 3284 5836
rect 3316 5688 3324 5913
rect 3356 5747 3364 5913
rect 3313 5647 3327 5652
rect 3313 5640 3333 5647
rect 3316 5636 3333 5640
rect 3320 5633 3333 5636
rect 3396 5627 3404 6013
rect 3436 5947 3444 6073
rect 3516 5947 3524 6353
rect 3436 5767 3444 5933
rect 3476 5847 3484 5933
rect 3556 5907 3564 6353
rect 3696 6327 3704 6353
rect 3576 6147 3584 6173
rect 3556 5844 3564 5893
rect 3576 5887 3584 6133
rect 3616 6087 3624 6133
rect 3607 6076 3624 6087
rect 3607 6073 3620 6076
rect 3636 5927 3644 6213
rect 3696 6187 3704 6313
rect 3716 6187 3724 6413
rect 3756 6367 3764 6453
rect 3816 6267 3824 6413
rect 3716 6087 3724 6173
rect 3776 6047 3784 6213
rect 3816 6087 3824 6253
rect 3856 6147 3864 6193
rect 3876 6087 3884 6173
rect 3896 6047 3904 6133
rect 3916 6087 3924 6193
rect 3687 5904 3700 5907
rect 3687 5893 3704 5904
rect 3556 5836 3613 5844
rect 3516 5787 3524 5833
rect 3656 5807 3664 5833
rect 3696 5824 3704 5893
rect 3676 5816 3704 5824
rect 3516 5727 3524 5773
rect 3436 5627 3444 5693
rect 3556 5647 3564 5733
rect 3676 5707 3684 5816
rect 3716 5807 3724 5893
rect 3836 5847 3844 5913
rect 3756 5667 3764 5833
rect 3796 5767 3804 5833
rect 3856 5707 3864 6033
rect 3936 6027 3944 6513
rect 3996 6327 4004 6413
rect 4016 6387 4024 6513
rect 4093 6404 4107 6413
rect 4076 6400 4107 6404
rect 4076 6396 4104 6400
rect 3996 6147 4004 6313
rect 4016 6307 4024 6373
rect 4076 6201 4084 6396
rect 4256 6387 4264 6564
rect 4556 6476 4633 6484
rect 4116 6287 4124 6353
rect 4036 6147 4044 6173
rect 4096 6167 4104 6213
rect 4236 6167 4244 6253
rect 4236 6087 4244 6153
rect 4236 6076 4253 6087
rect 4240 6073 4253 6076
rect 4056 6047 4064 6073
rect 3893 5907 3907 5913
rect 3893 5900 3913 5907
rect 3896 5896 3913 5900
rect 3900 5893 3913 5896
rect 3996 5844 4004 5893
rect 3947 5836 4004 5844
rect 3640 5624 3653 5627
rect 3636 5613 3653 5624
rect 3707 5616 3733 5624
rect 3276 5427 3284 5453
rect 3316 5427 3324 5553
rect 3396 5547 3404 5573
rect 3636 5567 3644 5613
rect 3396 5536 3413 5547
rect 3400 5533 3413 5536
rect 3336 5447 3344 5493
rect 3247 5396 3264 5407
rect 3247 5393 3260 5396
rect 3196 5207 3204 5252
rect 3140 5104 3153 5107
rect 3136 5093 3153 5104
rect 3033 5004 3047 5013
rect 3033 5000 3064 5004
rect 3036 4996 3064 5000
rect 2953 4984 2967 4993
rect 2953 4980 2984 4984
rect 2956 4976 2984 4980
rect 2956 4747 2964 4953
rect 2976 4927 2984 4976
rect 2996 4667 3004 4893
rect 3016 4807 3024 4913
rect 3036 4867 3044 4953
rect 3056 4947 3064 4996
rect 3076 4907 3084 4993
rect 3136 4927 3144 5093
rect 3156 4887 3164 4973
rect 2907 4576 2924 4587
rect 2907 4573 2920 4576
rect 2776 4527 2784 4573
rect 2916 4467 2924 4493
rect 2716 4316 2764 4324
rect 2687 4304 2700 4307
rect 2687 4293 2704 4304
rect 2636 4247 2644 4273
rect 2576 4080 2604 4084
rect 2576 4076 2607 4080
rect 2593 4067 2607 4076
rect 2527 4056 2553 4064
rect 2496 4036 2524 4044
rect 2456 4016 2504 4024
rect 2456 3844 2464 3913
rect 2476 3867 2484 3993
rect 2496 3967 2504 4016
rect 2456 3836 2484 3844
rect 2476 3787 2484 3836
rect 2436 3776 2464 3784
rect 2436 3727 2444 3753
rect 2396 3696 2424 3704
rect 2156 3387 2164 3473
rect 2196 3387 2204 3533
rect 2096 3307 2104 3333
rect 2236 3307 2244 3433
rect 2256 3347 2264 3673
rect 2276 3407 2284 3633
rect 2316 3524 2324 3693
rect 2296 3516 2324 3524
rect 2296 3487 2304 3516
rect 2336 3387 2344 3573
rect 2276 3316 2313 3324
rect 2193 3284 2207 3293
rect 2276 3284 2284 3316
rect 2193 3280 2284 3284
rect 2196 3276 2284 3280
rect 1996 3256 2024 3264
rect 1967 3236 1993 3244
rect 1916 3207 1924 3233
rect 1916 3067 1924 3193
rect 2016 3167 2024 3256
rect 2056 3247 2064 3273
rect 2056 3236 2073 3247
rect 2060 3233 2073 3236
rect 2116 3207 2124 3233
rect 1776 3027 1784 3053
rect 1780 2964 1793 2967
rect 1776 2960 1793 2964
rect 1773 2953 1793 2960
rect 1773 2947 1787 2953
rect 1816 2927 1824 3013
rect 1536 2607 1544 2713
rect 1556 2507 1564 2633
rect 1576 2524 1584 2713
rect 1576 2520 1604 2524
rect 1576 2516 1607 2520
rect 1593 2507 1607 2516
rect 1396 2416 1413 2427
rect 1400 2413 1413 2416
rect 1376 2347 1384 2413
rect 1436 2407 1444 2473
rect 1436 2393 1453 2407
rect 1356 2267 1364 2293
rect 1296 1987 1304 2013
rect 1187 1976 1204 1987
rect 1187 1973 1200 1976
rect 1027 1916 1044 1927
rect 1096 1924 1104 1973
rect 1096 1916 1153 1924
rect 1027 1913 1040 1916
rect 1247 1916 1273 1924
rect 976 1587 984 1673
rect 1016 1567 1024 1673
rect 896 1456 933 1464
rect 716 1407 724 1453
rect 956 1407 964 1513
rect 1076 1507 1084 1853
rect 1136 1647 1144 1733
rect 1216 1687 1224 1813
rect 1276 1767 1284 1833
rect 1336 1747 1344 1793
rect 1396 1787 1404 2253
rect 1436 2127 1444 2393
rect 1556 2367 1564 2493
rect 1656 2444 1664 2913
rect 1696 2807 1704 2833
rect 1736 2807 1744 2873
rect 1776 2747 1784 2813
rect 1836 2787 1844 2813
rect 1896 2804 1904 2993
rect 1876 2796 1904 2804
rect 1816 2687 1824 2713
rect 1696 2507 1704 2593
rect 1756 2507 1764 2533
rect 1696 2496 1713 2507
rect 1700 2493 1713 2496
rect 1656 2436 1693 2444
rect 1476 2207 1484 2293
rect 1496 2267 1504 2313
rect 1596 2307 1604 2433
rect 1716 2327 1724 2493
rect 1536 2207 1544 2253
rect 1527 2196 1544 2207
rect 1596 2207 1604 2293
rect 1636 2267 1644 2293
rect 1696 2207 1704 2313
rect 1736 2307 1744 2413
rect 1816 2387 1824 2673
rect 1856 2647 1864 2713
rect 1876 2627 1884 2796
rect 1916 2787 1924 3053
rect 1976 2924 1984 3073
rect 2016 2984 2024 3153
rect 1996 2980 2024 2984
rect 1993 2976 2024 2980
rect 1993 2967 2007 2976
rect 1976 2916 2004 2924
rect 1976 2687 1984 2813
rect 1996 2807 2004 2916
rect 2076 2907 2084 3013
rect 2076 2847 2084 2893
rect 2096 2887 2104 2953
rect 2016 2787 2024 2813
rect 2136 2787 2144 2813
rect 2016 2776 2033 2787
rect 2020 2773 2033 2776
rect 2136 2776 2153 2787
rect 2140 2773 2153 2776
rect 2196 2764 2204 3253
rect 2256 3107 2264 3233
rect 2296 3207 2304 3233
rect 2336 3067 2344 3333
rect 2247 3044 2260 3047
rect 2247 3034 2264 3044
rect 2240 3033 2264 3034
rect 2256 3027 2264 3033
rect 2256 3016 2273 3027
rect 2260 3013 2273 3016
rect 2196 2756 2224 2764
rect 2120 2724 2133 2727
rect 2116 2713 2133 2724
rect 2187 2724 2200 2727
rect 2187 2713 2204 2724
rect 2016 2687 2024 2713
rect 1936 2627 1944 2653
rect 2016 2644 2024 2673
rect 2056 2667 2064 2713
rect 2116 2687 2124 2713
rect 2007 2636 2024 2644
rect 1856 2407 1864 2473
rect 1876 2447 1884 2613
rect 1976 2487 1984 2533
rect 1876 2436 1893 2447
rect 1880 2433 1893 2436
rect 1996 2407 2004 2633
rect 2056 2547 2064 2653
rect 2016 2507 2024 2533
rect 2067 2500 2104 2504
rect 2067 2496 2107 2500
rect 2093 2487 2107 2496
rect 1596 2196 1613 2207
rect 1527 2193 1540 2196
rect 1600 2193 1613 2196
rect 1476 1987 1484 2133
rect 1656 2087 1664 2193
rect 1696 2107 1704 2153
rect 1756 2144 1764 2373
rect 1796 2267 1804 2313
rect 1796 2256 1813 2267
rect 1800 2253 1813 2256
rect 1836 2207 1844 2333
rect 1736 2136 1764 2144
rect 1527 1980 1564 1984
rect 1527 1976 1567 1980
rect 1553 1967 1567 1976
rect 1416 1747 1424 1913
rect 1327 1733 1344 1747
rect 1307 1684 1320 1687
rect 1307 1680 1324 1684
rect 1307 1673 1327 1680
rect 987 1456 1013 1464
rect 1036 1407 1044 1493
rect 1180 1464 1193 1467
rect 1176 1453 1193 1464
rect 716 1396 733 1407
rect 720 1393 733 1396
rect 1036 1396 1053 1407
rect 1040 1393 1053 1396
rect 456 1347 464 1393
rect 456 1167 464 1293
rect 476 1227 484 1273
rect 496 1127 504 1153
rect 536 1127 544 1253
rect 596 1244 604 1373
rect 776 1267 784 1373
rect 576 1240 604 1244
rect 573 1236 604 1240
rect 573 1227 587 1236
rect 736 1227 744 1253
rect 436 960 464 964
rect 436 956 467 960
rect 453 947 467 956
rect 327 936 344 947
rect 327 933 340 936
rect 387 936 413 944
rect 276 847 284 933
rect 307 884 320 887
rect 307 880 324 884
rect 307 873 327 880
rect 313 868 327 873
rect 296 707 304 773
rect 287 696 304 707
rect 287 693 300 696
rect 316 684 324 832
rect 356 707 364 813
rect 376 747 384 873
rect 456 847 464 933
rect 536 827 544 873
rect 576 847 584 933
rect 596 887 604 993
rect 616 947 624 1033
rect 636 987 644 1173
rect 736 987 744 1213
rect 776 1147 784 1173
rect 816 1147 824 1393
rect 916 1167 924 1353
rect 1016 1227 1024 1353
rect 1176 1327 1184 1453
rect 1236 1367 1244 1453
rect 1256 1407 1264 1673
rect 1313 1667 1327 1673
rect 1336 1647 1344 1733
rect 1436 1647 1444 1673
rect 1136 1227 1144 1273
rect 1236 1267 1244 1353
rect 1176 1216 1213 1224
rect 296 676 324 684
rect 196 636 213 647
rect 200 633 213 636
rect 256 607 264 633
rect 296 527 304 676
rect 416 647 424 773
rect 360 644 373 647
rect 356 640 373 644
rect 353 633 373 640
rect 476 644 484 793
rect 556 707 564 753
rect 547 696 564 707
rect 547 693 560 696
rect 476 636 513 644
rect 596 644 604 833
rect 567 636 604 644
rect 353 627 367 633
rect 156 427 164 453
rect 236 427 244 513
rect 276 367 284 453
rect 416 444 424 633
rect 656 627 664 693
rect 676 667 684 793
rect 716 767 724 873
rect 756 828 764 933
rect 776 887 784 993
rect 796 947 804 1033
rect 816 847 824 1133
rect 876 1127 884 1153
rect 996 1127 1004 1153
rect 1036 1087 1044 1153
rect 876 947 884 973
rect 900 944 913 947
rect 896 933 913 944
rect 716 727 724 753
rect 756 727 764 792
rect 676 656 693 667
rect 680 653 693 656
rect 816 664 824 833
rect 836 787 844 873
rect 876 864 884 933
rect 856 856 884 864
rect 856 807 864 856
rect 896 847 904 933
rect 976 827 984 1073
rect 1036 947 1044 1033
rect 1076 947 1084 993
rect 876 707 884 733
rect 787 656 824 664
rect 416 440 444 444
rect 416 436 447 440
rect 433 427 447 436
rect 356 420 393 424
rect 353 416 393 420
rect 353 407 367 416
rect 267 356 284 367
rect 267 353 280 356
rect 416 327 424 353
rect 96 127 104 273
rect 136 127 144 253
rect 296 187 304 213
rect 376 207 384 273
rect 436 227 444 253
rect 476 227 484 533
rect 596 427 604 453
rect 636 427 644 573
rect 736 507 744 633
rect 856 607 864 633
rect 896 567 904 633
rect 660 444 673 447
rect 656 433 673 444
rect 656 404 664 433
rect 713 427 727 433
rect 776 427 784 473
rect 873 427 887 433
rect 936 427 944 553
rect 956 467 964 693
rect 713 420 733 427
rect 716 416 733 420
rect 720 413 733 416
rect 747 416 764 424
rect 536 396 664 404
rect 536 367 544 396
rect 756 384 764 416
rect 873 420 893 427
rect 876 416 893 420
rect 880 413 893 416
rect 756 376 793 384
rect 996 367 1004 593
rect 1016 527 1024 873
rect 1036 647 1044 733
rect 1116 707 1124 973
rect 1056 587 1064 693
rect 1087 644 1100 647
rect 1087 633 1104 644
rect 1096 527 1104 633
rect 1096 487 1104 513
rect 1136 427 1144 1113
rect 1176 1087 1184 1216
rect 1247 1164 1260 1167
rect 1247 1153 1264 1164
rect 1196 1107 1204 1153
rect 1196 947 1204 973
rect 1256 944 1264 1153
rect 1276 1107 1284 1633
rect 1296 1407 1304 1593
rect 1360 1464 1373 1467
rect 1356 1453 1373 1464
rect 1336 1367 1344 1453
rect 1296 1227 1304 1313
rect 1356 1287 1364 1453
rect 1316 1167 1324 1273
rect 1356 1127 1364 1153
rect 1247 936 1284 944
rect 1176 847 1184 873
rect 1176 767 1184 833
rect 1216 827 1224 853
rect 1276 747 1284 936
rect 1236 707 1244 733
rect 1216 587 1224 633
rect 1256 527 1264 633
rect 1176 427 1184 453
rect 1236 427 1244 473
rect 1227 416 1244 427
rect 1227 413 1240 416
rect 860 364 873 367
rect 856 353 873 364
rect 576 287 584 333
rect 616 307 624 353
rect 716 327 724 353
rect 756 307 764 333
rect 856 327 864 353
rect 713 267 727 273
rect 713 260 714 267
rect 706 233 707 240
rect 436 187 444 213
rect 556 187 564 233
rect 693 227 707 233
rect 693 220 714 227
rect 696 216 714 220
rect 700 213 714 216
rect 656 187 664 213
rect 796 187 804 293
rect 836 227 844 253
rect 236 27 244 173
rect 407 156 524 164
rect 336 127 344 153
rect 327 116 344 127
rect 327 113 340 116
rect 387 116 413 124
rect 493 124 507 133
rect 516 127 524 156
rect 696 147 704 173
rect 616 140 684 144
rect 616 136 687 140
rect 616 127 624 136
rect 673 127 687 136
rect 836 144 844 173
rect 876 164 884 233
rect 736 140 844 144
rect 733 136 844 140
rect 856 156 884 164
rect 467 120 507 124
rect 467 116 504 120
rect 607 116 624 127
rect 607 113 620 116
rect 733 127 747 136
rect 276 87 284 113
rect 636 87 644 113
rect 776 87 784 113
rect 816 87 824 113
rect 856 27 864 156
rect 896 87 904 273
rect 976 227 984 333
rect 976 187 984 213
rect 1036 207 1044 293
rect 1056 247 1064 413
rect 1096 267 1104 413
rect 1316 407 1324 1093
rect 1336 707 1344 1073
rect 1376 1047 1384 1333
rect 1436 1327 1444 1393
rect 1456 1284 1464 1893
rect 1496 1887 1504 1913
rect 1556 1896 1593 1904
rect 1476 1647 1484 1673
rect 1496 1667 1504 1733
rect 1536 1707 1544 1793
rect 1556 1687 1564 1896
rect 1620 1904 1633 1907
rect 1616 1893 1633 1904
rect 1596 1767 1604 1853
rect 1616 1724 1624 1893
rect 1656 1827 1664 1933
rect 1636 1747 1644 1773
rect 1616 1716 1644 1724
rect 1587 1704 1600 1707
rect 1587 1693 1604 1704
rect 1596 1687 1604 1693
rect 1596 1676 1613 1687
rect 1600 1673 1613 1676
rect 1587 1664 1600 1667
rect 1587 1653 1604 1664
rect 1496 1487 1504 1613
rect 1596 1607 1604 1653
rect 1636 1607 1644 1716
rect 1436 1276 1464 1284
rect 1396 1067 1404 1273
rect 1436 1007 1444 1276
rect 1476 1167 1484 1393
rect 1516 1344 1524 1393
rect 1496 1336 1524 1344
rect 1496 1287 1504 1336
rect 1536 1327 1544 1553
rect 1536 1247 1544 1313
rect 1556 1287 1564 1593
rect 1576 1347 1584 1573
rect 1636 1548 1644 1593
rect 1676 1567 1684 2013
rect 1736 1847 1744 2136
rect 1816 2027 1824 2153
rect 1816 1987 1824 2013
rect 1896 1967 1904 2313
rect 1776 1847 1784 1912
rect 1836 1867 1844 1912
rect 1696 1607 1704 1773
rect 1736 1747 1744 1793
rect 1776 1787 1784 1833
rect 1916 1807 1924 2393
rect 1956 2167 1964 2253
rect 2016 2047 2024 2433
rect 2040 2264 2053 2267
rect 2036 2253 2053 2264
rect 2036 2207 2044 2253
rect 2056 2047 2064 2113
rect 1956 1847 1964 2013
rect 2036 1987 2044 2013
rect 2007 1984 2020 1987
rect 2007 1973 2024 1984
rect 2016 1964 2024 1973
rect 2016 1956 2044 1964
rect 2016 1887 2024 1913
rect 2016 1847 2024 1873
rect 2036 1787 2044 1956
rect 2076 1927 2084 2193
rect 2096 1807 2104 2433
rect 2116 2267 2124 2633
rect 2156 2447 2164 2673
rect 2196 2667 2204 2713
rect 2216 2567 2224 2756
rect 2236 2667 2244 3012
rect 2256 2787 2264 2873
rect 2296 2824 2304 2953
rect 2316 2848 2324 3013
rect 2356 2867 2364 3633
rect 2396 3587 2404 3696
rect 2416 3547 2424 3673
rect 2456 3547 2464 3776
rect 2476 3647 2484 3773
rect 2496 3587 2504 3913
rect 2516 3867 2524 4036
rect 2547 3996 2573 4004
rect 2616 3927 2624 3973
rect 2516 3627 2524 3773
rect 2556 3767 2564 3893
rect 2596 3767 2604 3893
rect 2636 3887 2644 3913
rect 2656 3907 2664 4133
rect 2636 3827 2644 3873
rect 2636 3816 2653 3827
rect 2640 3813 2653 3816
rect 2536 3667 2544 3753
rect 2556 3547 2564 3673
rect 2580 3544 2593 3547
rect 2576 3533 2593 3544
rect 2376 3427 2384 3533
rect 2376 3247 2384 3413
rect 2456 3367 2464 3473
rect 2393 3307 2407 3313
rect 2393 3300 2413 3307
rect 2396 3296 2413 3300
rect 2400 3293 2413 3296
rect 2376 3236 2393 3247
rect 2380 3233 2393 3236
rect 2447 3244 2460 3247
rect 2447 3233 2464 3244
rect 2376 3147 2384 3193
rect 2416 3067 2424 3193
rect 2456 3147 2464 3233
rect 2476 3207 2484 3493
rect 2496 3347 2504 3533
rect 2576 3524 2584 3533
rect 2536 3520 2584 3524
rect 2533 3516 2584 3520
rect 2533 3507 2547 3516
rect 2496 3107 2504 3173
rect 2516 3147 2524 3393
rect 2376 2847 2384 3053
rect 2436 3027 2444 3073
rect 2516 3067 2524 3133
rect 2536 3107 2544 3453
rect 2576 3447 2584 3473
rect 2636 3427 2644 3733
rect 2676 3407 2684 4133
rect 2456 2967 2464 3053
rect 2476 3027 2484 3053
rect 2556 2987 2564 3393
rect 2576 3247 2584 3353
rect 2596 3327 2604 3353
rect 2636 3307 2644 3333
rect 2616 3127 2624 3233
rect 2696 3224 2704 4293
rect 2716 4267 2724 4316
rect 2856 4307 2864 4433
rect 2916 4307 2924 4453
rect 2876 4256 2913 4264
rect 2796 4147 2804 4213
rect 2716 3927 2724 4053
rect 2756 3948 2764 4053
rect 2736 3687 2744 3893
rect 2756 3887 2764 3912
rect 2776 3787 2784 3973
rect 2816 3907 2824 4133
rect 2836 3907 2844 4193
rect 2876 4127 2884 4256
rect 2936 4167 2944 4293
rect 2956 4228 2964 4453
rect 2860 4064 2873 4067
rect 2856 4053 2873 4064
rect 2856 4027 2864 4053
rect 2856 4000 2893 4004
rect 2853 3996 2893 4000
rect 2853 3987 2867 3996
rect 2916 3947 2924 4053
rect 2956 4007 2964 4192
rect 2976 4147 2984 4653
rect 3036 4587 3044 4713
rect 3056 4647 3064 4773
rect 3116 4767 3124 4873
rect 3136 4688 3144 4753
rect 3136 4587 3144 4652
rect 3176 4627 3184 4733
rect 3196 4667 3204 5193
rect 2996 4267 3004 4393
rect 3016 4107 3024 4493
rect 3036 4167 3044 4573
rect 3056 4228 3064 4273
rect 3056 4147 3064 4192
rect 3076 4164 3084 4573
rect 3196 4467 3204 4553
rect 3116 4347 3124 4433
rect 3136 4284 3144 4333
rect 3107 4276 3144 4284
rect 3156 4284 3164 4413
rect 3216 4387 3224 5033
rect 3236 5007 3244 5233
rect 3296 5147 3304 5173
rect 3336 5147 3344 5333
rect 3356 5227 3364 5413
rect 3376 5247 3384 5493
rect 3456 5487 3464 5533
rect 3576 5487 3584 5553
rect 3396 5287 3404 5473
rect 3416 5327 3424 5433
rect 3436 5387 3444 5413
rect 3476 5387 3484 5433
rect 3496 5327 3504 5473
rect 3616 5364 3624 5493
rect 3636 5387 3644 5453
rect 3676 5407 3684 5533
rect 3696 5487 3704 5513
rect 3716 5447 3724 5553
rect 3796 5427 3804 5633
rect 3876 5587 3884 5753
rect 3896 5667 3904 5833
rect 3916 5707 3924 5753
rect 3936 5727 3944 5793
rect 3907 5656 3924 5664
rect 3896 5507 3904 5613
rect 3916 5524 3924 5656
rect 3936 5627 3944 5713
rect 3976 5627 3984 5733
rect 4016 5584 4024 6013
rect 4056 5664 4064 6033
rect 4196 5987 4204 6073
rect 4136 5847 4144 5953
rect 4236 5947 4244 6033
rect 4256 5927 4264 5953
rect 4200 5904 4213 5907
rect 4087 5844 4100 5847
rect 4087 5833 4104 5844
rect 4127 5836 4144 5847
rect 4196 5893 4213 5904
rect 4127 5833 4140 5836
rect 4056 5656 4084 5664
rect 3976 5576 4024 5584
rect 3916 5516 3944 5524
rect 3836 5427 3844 5453
rect 3727 5400 3764 5404
rect 3727 5396 3767 5400
rect 3753 5387 3767 5396
rect 3616 5360 3704 5364
rect 3616 5356 3707 5360
rect 3693 5347 3707 5356
rect 3440 5324 3453 5327
rect 3436 5313 3453 5324
rect 3436 5267 3444 5313
rect 3536 5247 3544 5313
rect 3656 5307 3664 5333
rect 3456 5187 3464 5233
rect 3556 5167 3564 5233
rect 3576 5167 3584 5273
rect 3736 5267 3744 5333
rect 3876 5327 3884 5473
rect 3896 5327 3904 5413
rect 3867 5316 3884 5327
rect 3867 5313 3880 5316
rect 3696 5167 3704 5253
rect 3296 5107 3304 5133
rect 3493 5107 3507 5113
rect 3420 5104 3433 5107
rect 3416 5093 3433 5104
rect 3487 5100 3507 5107
rect 3487 5096 3504 5100
rect 3487 5093 3500 5096
rect 3336 5008 3344 5093
rect 3416 5067 3424 5093
rect 3516 5047 3524 5133
rect 3556 5087 3564 5153
rect 3556 5076 3573 5087
rect 3560 5073 3573 5076
rect 3507 5036 3524 5047
rect 3507 5033 3520 5036
rect 3236 4827 3244 4933
rect 3296 4887 3304 4933
rect 3336 4887 3344 4972
rect 3260 4824 3273 4827
rect 3256 4813 3273 4824
rect 3236 4467 3244 4613
rect 3256 4567 3264 4813
rect 3316 4667 3324 4793
rect 3356 4767 3364 4813
rect 3376 4727 3384 5033
rect 3636 5027 3644 5153
rect 3656 5087 3664 5133
rect 3676 5047 3684 5113
rect 3593 5004 3607 5013
rect 3593 5000 3644 5004
rect 3596 4996 3644 5000
rect 3536 4867 3544 4913
rect 3576 4887 3584 4953
rect 3616 4867 3624 4953
rect 3636 4947 3644 4996
rect 3676 4964 3684 4993
rect 3656 4956 3684 4964
rect 3440 4864 3453 4867
rect 3366 4716 3384 4727
rect 3436 4853 3453 4864
rect 3366 4713 3380 4716
rect 3436 4687 3444 4853
rect 3656 4824 3664 4956
rect 3696 4944 3704 5153
rect 3636 4820 3664 4824
rect 3633 4816 3664 4820
rect 3676 4936 3704 4944
rect 3633 4807 3647 4816
rect 3460 4804 3473 4807
rect 3456 4793 3473 4804
rect 3456 4747 3464 4793
rect 3456 4688 3464 4733
rect 3336 4587 3344 4613
rect 3156 4276 3193 4284
rect 3236 4247 3244 4273
rect 3196 4187 3204 4213
rect 3236 4187 3244 4233
rect 3256 4227 3264 4433
rect 3076 4156 3104 4164
rect 3093 4147 3104 4156
rect 3116 4107 3124 4153
rect 3136 4128 3144 4153
rect 3116 4106 3140 4107
rect 3116 4093 3133 4106
rect 2947 3996 2964 4007
rect 2947 3993 2960 3996
rect 2996 3927 3004 4073
rect 3056 4067 3064 4093
rect 3076 4067 3084 4093
rect 3076 4056 3093 4067
rect 3080 4053 3093 4056
rect 3116 4007 3124 4093
rect 2896 3827 2904 3893
rect 3076 3847 3084 3973
rect 3087 3776 3124 3784
rect 2836 3687 2844 3773
rect 3013 3744 3027 3753
rect 3013 3740 3073 3744
rect 3016 3736 3073 3740
rect 3116 3687 3124 3776
rect 2716 3527 2724 3633
rect 2856 3587 2864 3653
rect 2716 3516 2733 3527
rect 2720 3513 2733 3516
rect 2756 3484 2764 3573
rect 2816 3527 2824 3553
rect 2736 3476 2764 3484
rect 2716 3388 2724 3473
rect 2716 3247 2724 3352
rect 2736 3307 2744 3476
rect 2756 3347 2764 3453
rect 2776 3427 2784 3513
rect 2796 3407 2804 3453
rect 2736 3296 2753 3307
rect 2740 3293 2753 3296
rect 2796 3247 2804 3393
rect 2716 3236 2733 3247
rect 2720 3233 2733 3236
rect 2787 3236 2804 3247
rect 2787 3233 2800 3236
rect 2696 3216 2724 3224
rect 2576 3004 2584 3093
rect 2616 3027 2624 3053
rect 2656 3027 2664 3053
rect 2576 2996 2604 3004
rect 2400 2964 2413 2967
rect 2396 2953 2413 2964
rect 2396 2887 2404 2953
rect 2296 2816 2312 2824
rect 2276 2664 2284 2813
rect 2316 2787 2324 2812
rect 2336 2727 2344 2813
rect 2296 2687 2304 2713
rect 2276 2656 2304 2664
rect 2236 2487 2244 2553
rect 2196 2407 2204 2433
rect 2276 2407 2284 2473
rect 2116 2147 2124 2193
rect 2136 2167 2144 2393
rect 2196 2347 2204 2393
rect 2176 2007 2184 2273
rect 2256 2267 2264 2353
rect 2296 2307 2304 2656
rect 2296 2027 2304 2253
rect 2316 2087 2324 2393
rect 2336 2327 2344 2653
rect 2356 2327 2364 2553
rect 2376 2547 2384 2713
rect 2396 2567 2404 2613
rect 2416 2587 2424 2853
rect 2456 2827 2464 2893
rect 2456 2787 2464 2813
rect 2496 2587 2504 2973
rect 2596 2964 2604 2996
rect 2596 2956 2633 2964
rect 2516 2900 2524 2904
rect 2513 2887 2527 2900
rect 2516 2687 2524 2873
rect 2536 2627 2544 2893
rect 2596 2887 2604 2933
rect 2596 2727 2604 2833
rect 2716 2827 2724 3216
rect 2776 3087 2784 3233
rect 2856 3227 2864 3473
rect 2896 3447 2904 3633
rect 3036 3567 3044 3633
rect 3136 3627 3144 3833
rect 3156 3667 3164 4173
rect 3276 4147 3284 4473
rect 3296 4427 3304 4573
rect 3356 4564 3364 4673
rect 3420 4644 3433 4647
rect 3336 4556 3364 4564
rect 3416 4633 3433 4644
rect 3336 4527 3344 4556
rect 3336 4447 3344 4513
rect 3373 4504 3387 4513
rect 3356 4500 3387 4504
rect 3353 4496 3384 4500
rect 3353 4488 3367 4496
rect 3296 4207 3304 4413
rect 3356 4408 3364 4452
rect 3316 4207 3324 4393
rect 3356 4287 3364 4372
rect 3396 4287 3404 4433
rect 3416 4427 3424 4633
rect 3456 4487 3464 4652
rect 3436 4404 3444 4453
rect 3476 4427 3484 4733
rect 3556 4607 3564 4713
rect 3556 4567 3564 4593
rect 3507 4556 3544 4564
rect 3536 4544 3544 4556
rect 3536 4540 3584 4544
rect 3536 4536 3587 4540
rect 3573 4527 3587 4536
rect 3596 4507 3604 4793
rect 3676 4747 3684 4936
rect 3716 4904 3724 5173
rect 3776 5107 3784 5173
rect 3816 5107 3824 5153
rect 3706 4896 3724 4904
rect 3696 4867 3704 4893
rect 3836 4887 3844 5033
rect 3856 5007 3864 5313
rect 3876 5107 3884 5233
rect 3916 5147 3924 5433
rect 3936 5187 3944 5516
rect 3976 5387 3984 5576
rect 4056 5567 4064 5633
rect 3996 5467 4004 5553
rect 3976 5376 3993 5387
rect 3980 5373 3993 5376
rect 4016 5287 4024 5313
rect 3976 5188 3984 5273
rect 3976 5107 3984 5152
rect 3920 5104 3933 5107
rect 3916 5093 3933 5104
rect 3987 5100 4024 5104
rect 3987 5096 4027 5100
rect 3916 5047 3924 5093
rect 4013 5087 4027 5096
rect 4036 5007 4044 5453
rect 4056 5267 4064 5513
rect 4076 5347 4084 5656
rect 4096 5607 4104 5833
rect 4196 5807 4204 5893
rect 4276 5847 4284 5933
rect 4220 5844 4233 5847
rect 4216 5833 4233 5844
rect 4136 5547 4144 5733
rect 4156 5584 4164 5773
rect 4216 5767 4224 5833
rect 4176 5607 4184 5633
rect 4156 5576 4184 5584
rect 4136 5536 4153 5547
rect 4140 5533 4153 5536
rect 4096 5508 4104 5533
rect 4096 5447 4104 5472
rect 4176 5427 4184 5576
rect 3896 4867 3904 4893
rect 3696 4856 3713 4867
rect 3700 4853 3713 4856
rect 3840 4824 3853 4827
rect 3836 4813 3853 4824
rect 3636 4647 3644 4733
rect 3736 4668 3744 4793
rect 3816 4707 3824 4753
rect 3836 4727 3844 4813
rect 3856 4704 3864 4753
rect 3876 4727 3884 4773
rect 3896 4767 3904 4853
rect 3836 4696 3864 4704
rect 3836 4684 3844 4696
rect 3816 4676 3844 4684
rect 3776 4647 3784 4673
rect 3736 4607 3744 4632
rect 3736 4596 3753 4607
rect 3740 4593 3753 4596
rect 3507 4480 3584 4484
rect 3507 4476 3587 4480
rect 3573 4467 3587 4476
rect 3496 4427 3504 4452
rect 3596 4444 3604 4493
rect 3556 4440 3604 4444
rect 3553 4436 3604 4440
rect 3553 4427 3567 4436
rect 3566 4420 3567 4427
rect 3416 4396 3444 4404
rect 3416 4347 3424 4396
rect 3416 4267 3424 4333
rect 3376 4167 3384 4233
rect 3196 4007 3204 4133
rect 3316 4124 3324 4153
rect 3296 4120 3324 4124
rect 3293 4116 3324 4120
rect 3293 4107 3307 4116
rect 3336 4067 3344 4113
rect 3416 4087 3424 4213
rect 3456 4207 3464 4333
rect 3576 4307 3584 4413
rect 3636 4307 3644 4593
rect 3747 4576 3773 4584
rect 3693 4564 3707 4573
rect 3693 4560 3744 4564
rect 3696 4556 3744 4560
rect 3673 4484 3687 4493
rect 3736 4487 3744 4556
rect 3796 4527 3804 4653
rect 3816 4607 3824 4676
rect 3856 4587 3864 4653
rect 3916 4647 3924 4993
rect 4056 4984 4064 5253
rect 4076 5227 4084 5244
rect 4196 5227 4204 5493
rect 4216 5427 4224 5553
rect 4256 5467 4264 5713
rect 4276 5444 4284 5693
rect 4316 5444 4324 6373
rect 4356 5907 4364 6293
rect 4416 6227 4424 6373
rect 4436 6247 4444 6413
rect 4556 6387 4564 6476
rect 4716 6427 4724 6453
rect 4756 6427 4764 6473
rect 4600 6384 4613 6387
rect 4596 6373 4613 6384
rect 4416 6127 4424 6213
rect 4416 6116 4433 6127
rect 4420 6113 4433 6116
rect 4376 6064 4384 6113
rect 4476 6087 4484 6273
rect 4596 6227 4604 6373
rect 4796 6367 4804 6413
rect 4996 6407 5004 6433
rect 5256 6407 5264 6493
rect 5556 6427 5564 6564
rect 5696 6427 5704 6493
rect 5936 6487 5944 6564
rect 6176 6556 6204 6564
rect 5856 6427 5864 6473
rect 5847 6416 5864 6427
rect 5847 6413 5860 6416
rect 5127 6396 5204 6404
rect 4787 6356 4804 6367
rect 4787 6353 4800 6356
rect 4736 6307 4744 6353
rect 4896 6327 4904 6353
rect 4936 6307 4944 6353
rect 4576 6147 4584 6173
rect 4696 6147 4704 6253
rect 4876 6227 4884 6253
rect 4627 6144 4640 6147
rect 4627 6133 4644 6144
rect 4696 6136 4713 6147
rect 4700 6133 4713 6136
rect 4636 6087 4644 6133
rect 4376 6056 4433 6064
rect 4756 6007 4764 6133
rect 4876 6107 4884 6213
rect 4813 6084 4827 6093
rect 4813 6080 4844 6084
rect 4816 6076 4844 6080
rect 4476 5967 4484 5993
rect 4516 5907 4524 5933
rect 4356 5896 4373 5907
rect 4360 5893 4373 5896
rect 4396 5647 4404 5833
rect 4436 5607 4444 5793
rect 4456 5747 4464 5833
rect 4576 5807 4584 5933
rect 4336 5487 4344 5593
rect 4256 5436 4284 5444
rect 4296 5436 4324 5444
rect 4256 5324 4264 5436
rect 4296 5424 4304 5436
rect 4276 5416 4304 5424
rect 4276 5347 4284 5416
rect 4256 5316 4284 5324
rect 4076 5127 4084 5213
rect 4276 5167 4284 5316
rect 4076 5027 4084 5113
rect 4176 5084 4184 5133
rect 4256 5107 4264 5153
rect 4296 5107 4304 5273
rect 4156 5076 4184 5084
rect 4116 4987 4124 5013
rect 4036 4980 4064 4984
rect 4033 4976 4064 4980
rect 3936 4767 3944 4973
rect 4033 4967 4047 4976
rect 3956 4867 3964 4933
rect 4036 4744 4044 4853
rect 4076 4807 4084 4973
rect 4036 4736 4064 4744
rect 3673 4480 3724 4484
rect 3676 4476 3724 4480
rect 3696 4407 3704 4453
rect 3716 4347 3724 4476
rect 3776 4367 3784 4413
rect 3716 4336 3733 4347
rect 3720 4333 3733 4336
rect 3647 4304 3660 4307
rect 3647 4293 3664 4304
rect 3656 4247 3664 4293
rect 3227 4064 3240 4067
rect 3227 4053 3244 4064
rect 3387 4056 3424 4064
rect 3236 4007 3244 4053
rect 3416 4007 3424 4056
rect 3216 3867 3224 3893
rect 3296 3887 3304 3993
rect 3316 3927 3324 3953
rect 3336 3907 3344 3933
rect 3436 3927 3444 4193
rect 3496 4127 3504 4173
rect 3456 3967 3464 4073
rect 3496 4067 3504 4113
rect 3533 4044 3547 4053
rect 3533 4040 3564 4044
rect 3536 4036 3564 4040
rect 3556 4007 3564 4036
rect 3196 3827 3204 3853
rect 3256 3827 3264 3873
rect 3196 3816 3213 3827
rect 3200 3813 3213 3816
rect 3196 3727 3204 3753
rect 3236 3707 3244 3753
rect 3296 3727 3304 3813
rect 3336 3767 3344 3853
rect 3376 3767 3384 3893
rect 3476 3787 3484 3973
rect 3576 3967 3584 4193
rect 3676 4147 3684 4333
rect 3796 4304 3804 4513
rect 3776 4296 3804 4304
rect 3716 4067 3724 4193
rect 3756 4187 3764 4273
rect 3776 4104 3784 4296
rect 3836 4284 3844 4513
rect 3876 4364 3884 4453
rect 3896 4387 3904 4573
rect 3956 4367 3964 4633
rect 4016 4587 4024 4653
rect 4056 4647 4064 4736
rect 3976 4467 3984 4573
rect 4076 4527 4084 4753
rect 3876 4356 3904 4364
rect 3807 4276 3844 4284
rect 3896 4247 3904 4356
rect 4036 4304 4044 4453
rect 4076 4387 4084 4513
rect 4036 4296 4064 4304
rect 4056 4167 4064 4296
rect 4076 4267 4084 4293
rect 4116 4267 4124 4933
rect 4136 4867 4144 4893
rect 4136 4427 4144 4853
rect 4156 4384 4164 5076
rect 4196 4807 4204 4993
rect 4176 4407 4184 4753
rect 4216 4747 4224 5033
rect 4236 4927 4244 4953
rect 4316 4947 4324 5436
rect 4396 5347 4404 5593
rect 4416 5487 4424 5553
rect 4456 5387 4464 5473
rect 4476 5467 4484 5633
rect 4496 5427 4504 5653
rect 4556 5627 4564 5673
rect 4516 5527 4524 5613
rect 4596 5567 4604 5733
rect 4616 5667 4624 5753
rect 4636 5527 4644 5893
rect 4656 5768 4664 5833
rect 4656 5567 4664 5732
rect 4696 5684 4704 5833
rect 4756 5707 4764 5893
rect 4836 5787 4844 6076
rect 4856 5827 4864 5973
rect 4936 5867 4944 6293
rect 4956 6247 4964 6313
rect 4996 6247 5004 6273
rect 5056 6267 5064 6393
rect 5093 6284 5107 6293
rect 5196 6287 5204 6396
rect 5396 6327 5404 6393
rect 5556 6327 5564 6353
rect 5676 6327 5684 6353
rect 5093 6280 5124 6284
rect 5096 6276 5124 6280
rect 5196 6276 5213 6287
rect 5116 6264 5124 6276
rect 5200 6273 5213 6276
rect 5116 6260 5184 6264
rect 5116 6256 5187 6260
rect 5173 6248 5187 6256
rect 4956 5968 4964 6233
rect 4996 6216 5033 6224
rect 4996 5987 5004 6216
rect 5076 5987 5084 6093
rect 5116 5987 5124 6233
rect 5396 6227 5404 6313
rect 5180 6224 5193 6227
rect 5162 6213 5164 6224
rect 5156 6067 5164 6213
rect 5176 6213 5193 6224
rect 5176 6107 5184 6213
rect 5236 6147 5244 6213
rect 5296 6147 5304 6213
rect 5336 6107 5344 6193
rect 5156 6056 5173 6067
rect 5160 6053 5173 6056
rect 5156 6016 5193 6024
rect 5156 5987 5164 6016
rect 4687 5676 4704 5684
rect 4676 5627 4684 5673
rect 4716 5627 4724 5653
rect 4716 5507 4724 5613
rect 4776 5567 4784 5753
rect 4816 5627 4824 5733
rect 4836 5727 4844 5773
rect 4856 5627 4864 5673
rect 4876 5667 4884 5733
rect 4916 5687 4924 5853
rect 4956 5667 4964 5932
rect 5036 5807 5044 5973
rect 4996 5627 5004 5793
rect 5096 5727 5104 5893
rect 4973 5544 4987 5553
rect 4856 5540 4904 5544
rect 4973 5540 5004 5544
rect 4853 5536 4904 5540
rect 4976 5536 5004 5540
rect 4853 5527 4867 5536
rect 4896 5524 4904 5536
rect 4896 5516 4924 5524
rect 4613 5484 4627 5493
rect 4596 5480 4627 5484
rect 4596 5476 4624 5480
rect 4233 4844 4247 4853
rect 4233 4840 4284 4844
rect 4236 4836 4284 4840
rect 4276 4824 4284 4836
rect 4276 4816 4313 4824
rect 4256 4607 4264 4813
rect 4356 4784 4364 5333
rect 4476 5320 4513 5324
rect 4473 5316 4513 5320
rect 4473 5307 4487 5316
rect 4556 5247 4564 5313
rect 4576 5207 4584 5413
rect 4376 5107 4384 5133
rect 4376 5096 4393 5107
rect 4380 5093 4393 5096
rect 4396 4824 4404 5033
rect 4416 4967 4424 5133
rect 4476 4864 4484 4933
rect 4447 4856 4484 4864
rect 4396 4816 4444 4824
rect 4436 4807 4444 4816
rect 4436 4796 4453 4807
rect 4440 4793 4453 4796
rect 4516 4784 4524 4973
rect 4556 4927 4564 5033
rect 4596 4907 4604 5476
rect 4616 4967 4624 5453
rect 4636 5387 4644 5413
rect 4656 5287 4664 5493
rect 4756 5464 4764 5493
rect 4736 5456 4764 5464
rect 4676 5387 4684 5453
rect 4716 5344 4724 5413
rect 4736 5387 4744 5456
rect 4696 5336 4724 5344
rect 4696 5327 4704 5336
rect 4687 5316 4704 5327
rect 4687 5313 4700 5316
rect 4716 5227 4724 5313
rect 4636 4987 4644 5193
rect 4696 5064 4704 5113
rect 4756 5087 4764 5433
rect 4776 5247 4784 5373
rect 4776 5167 4784 5233
rect 4796 5127 4804 5473
rect 4836 5347 4844 5453
rect 4916 5264 4924 5516
rect 4956 5347 4964 5453
rect 4996 5447 5004 5536
rect 4956 5307 4964 5333
rect 4916 5256 4973 5264
rect 4816 5147 4824 5233
rect 4996 5207 5004 5433
rect 5016 5427 5024 5613
rect 5036 5607 5044 5653
rect 5036 5596 5053 5607
rect 5040 5593 5053 5596
rect 5056 5467 5064 5593
rect 5096 5507 5104 5713
rect 5116 5607 5124 5753
rect 5096 5496 5113 5507
rect 5100 5493 5113 5496
rect 5136 5467 5144 5933
rect 5176 5867 5184 5993
rect 5296 5987 5304 6013
rect 5056 5387 5064 5413
rect 5080 5384 5093 5387
rect 5076 5373 5093 5384
rect 5076 5364 5084 5373
rect 5016 5356 5084 5364
rect 4676 5056 4704 5064
rect 4676 4964 4684 5056
rect 4656 4956 4684 4964
rect 4636 4864 4644 4893
rect 4596 4856 4644 4864
rect 4547 4796 4573 4804
rect 4336 4776 4364 4784
rect 4496 4776 4524 4784
rect 4276 4627 4284 4693
rect 4256 4567 4264 4593
rect 4207 4556 4244 4564
rect 4236 4544 4244 4556
rect 4236 4536 4284 4544
rect 4276 4487 4284 4536
rect 4296 4407 4304 4453
rect 4156 4376 4184 4384
rect 4116 4167 4124 4253
rect 4156 4187 4164 4293
rect 3756 4096 3784 4104
rect 3676 4007 3684 4053
rect 3756 4007 3764 4096
rect 3773 4067 3787 4073
rect 3773 4060 3793 4067
rect 3776 4056 3793 4060
rect 3780 4053 3793 4056
rect 3847 4064 3860 4067
rect 3847 4053 3864 4064
rect 4007 4064 4020 4067
rect 4007 4053 4024 4064
rect 3756 3996 3773 4007
rect 3760 3993 3773 3996
rect 3476 3776 3493 3787
rect 3480 3773 3493 3776
rect 3156 3587 3164 3653
rect 3156 3576 3173 3587
rect 3160 3573 3173 3576
rect 3093 3544 3107 3553
rect 3093 3540 3124 3544
rect 3096 3536 3124 3540
rect 2947 3476 2973 3484
rect 3096 3447 3104 3513
rect 2996 3436 3033 3444
rect 2916 3327 2924 3353
rect 2916 3316 2933 3327
rect 2920 3313 2933 3316
rect 2956 3267 2964 3433
rect 2996 3407 3004 3436
rect 3016 3367 3024 3393
rect 3116 3327 3124 3536
rect 3153 3504 3167 3513
rect 3153 3500 3184 3504
rect 3156 3496 3187 3500
rect 3173 3487 3187 3496
rect 3256 3487 3264 3573
rect 3256 3476 3273 3487
rect 3260 3473 3273 3476
rect 2816 3108 2824 3213
rect 2916 3207 2924 3253
rect 2976 3227 2984 3313
rect 3033 3284 3047 3293
rect 3033 3280 3064 3284
rect 3036 3276 3064 3280
rect 3007 3264 3020 3267
rect 3007 3253 3024 3264
rect 2956 3147 2964 3173
rect 2896 3087 2904 3133
rect 2740 3004 2753 3007
rect 2736 2993 2753 3004
rect 2736 2927 2744 2993
rect 2816 2947 2824 3072
rect 2836 3007 2844 3033
rect 2776 2887 2784 2933
rect 2736 2787 2744 2833
rect 2856 2787 2864 2953
rect 2667 2784 2680 2787
rect 2667 2773 2684 2784
rect 2636 2627 2644 2713
rect 2676 2707 2684 2773
rect 2376 2447 2384 2493
rect 2416 2387 2424 2533
rect 2520 2524 2533 2527
rect 2516 2520 2533 2524
rect 2433 2504 2447 2513
rect 2513 2513 2533 2520
rect 2513 2507 2527 2513
rect 2433 2500 2473 2504
rect 2436 2496 2473 2500
rect 2416 2207 2424 2333
rect 2436 2267 2444 2353
rect 2336 2107 2344 2193
rect 2376 2147 2384 2193
rect 2356 2087 2364 2133
rect 2156 1847 2164 1893
rect 1816 1747 1824 1773
rect 2176 1747 2184 1813
rect 2196 1787 2204 1893
rect 1993 1724 2007 1733
rect 1993 1720 2024 1724
rect 1996 1716 2027 1720
rect 2013 1707 2027 1716
rect 1896 1700 1984 1704
rect 1893 1696 1984 1700
rect 1893 1687 1907 1696
rect 1976 1687 1984 1696
rect 1740 1684 1753 1687
rect 1736 1673 1753 1684
rect 1807 1676 1833 1684
rect 2036 1684 2044 1733
rect 2116 1696 2173 1704
rect 1987 1676 2044 1684
rect 1716 1587 1724 1633
rect 1596 1467 1604 1533
rect 1636 1467 1644 1512
rect 1736 1407 1744 1673
rect 1796 1567 1804 1633
rect 1936 1607 1944 1673
rect 2056 1627 2064 1693
rect 2116 1687 2124 1696
rect 2107 1676 2124 1687
rect 2107 1673 2120 1676
rect 1776 1467 1784 1493
rect 1496 1107 1504 1233
rect 1596 1187 1604 1253
rect 1616 1167 1624 1273
rect 1616 1156 1633 1167
rect 1620 1153 1633 1156
rect 1636 1127 1644 1153
rect 1496 947 1504 1053
rect 1536 1007 1544 1093
rect 1636 1067 1644 1113
rect 1656 1107 1664 1213
rect 1676 1087 1684 1153
rect 1696 1067 1704 1333
rect 1796 1307 1804 1393
rect 1816 1367 1824 1453
rect 1856 1407 1864 1493
rect 1936 1467 1944 1593
rect 2056 1567 2064 1613
rect 2136 1607 2144 1673
rect 2076 1467 2084 1593
rect 2176 1547 2184 1613
rect 2196 1587 2204 1633
rect 2216 1527 2224 2013
rect 2236 1787 2244 1993
rect 2356 1987 2364 2073
rect 2276 1980 2313 1984
rect 2273 1976 2313 1980
rect 2273 1967 2287 1976
rect 2296 1867 2304 1913
rect 2396 1827 2404 2113
rect 2436 1967 2444 2153
rect 2456 1927 2464 2453
rect 2556 2447 2564 2553
rect 2547 2436 2564 2447
rect 2547 2433 2560 2436
rect 2476 2327 2484 2393
rect 2576 2387 2584 2613
rect 2616 2507 2624 2533
rect 2656 2507 2664 2533
rect 2616 2484 2624 2493
rect 2696 2484 2704 2613
rect 2716 2547 2724 2613
rect 2616 2476 2644 2484
rect 2636 2464 2644 2476
rect 2676 2476 2704 2484
rect 2636 2456 2664 2464
rect 2476 2007 2484 2313
rect 2536 2087 2544 2373
rect 2616 2367 2624 2433
rect 2656 2387 2664 2456
rect 2556 2267 2564 2333
rect 2276 1736 2293 1744
rect 2276 1705 2284 1736
rect 2307 1736 2364 1744
rect 2247 1697 2284 1705
rect 2236 1587 2244 1672
rect 2276 1567 2284 1673
rect 2316 1607 2324 1673
rect 2356 1587 2364 1736
rect 2256 1556 2273 1564
rect 2256 1484 2264 1556
rect 2236 1476 2264 1484
rect 2236 1467 2244 1476
rect 2227 1456 2244 1467
rect 2227 1453 2240 1456
rect 2020 1444 2033 1447
rect 2016 1433 2033 1444
rect 2127 1444 2140 1447
rect 2127 1433 2144 1444
rect 1896 1347 1904 1393
rect 2016 1367 2024 1433
rect 2136 1407 2144 1433
rect 2016 1227 2024 1313
rect 2056 1307 2064 1373
rect 2093 1364 2107 1373
rect 2093 1356 2124 1364
rect 2093 1347 2107 1356
rect 1736 1027 1744 1213
rect 1796 1128 1804 1153
rect 1776 1116 1793 1124
rect 1536 947 1544 993
rect 1656 947 1664 973
rect 1776 947 1784 1116
rect 1816 1107 1824 1213
rect 1836 1127 1844 1153
rect 1796 1096 1813 1104
rect 1600 944 1613 947
rect 1596 933 1613 944
rect 1596 887 1604 933
rect 1796 887 1804 1096
rect 1836 1087 1844 1113
rect 1816 947 1824 973
rect 1827 944 1840 947
rect 1827 933 1844 944
rect 1396 827 1404 873
rect 1416 707 1424 733
rect 1416 696 1433 707
rect 1420 693 1433 696
rect 1336 547 1344 693
rect 1456 647 1464 813
rect 1596 767 1604 873
rect 1636 704 1644 853
rect 1607 696 1644 704
rect 1416 607 1424 633
rect 1496 567 1504 693
rect 1576 607 1584 633
rect 1616 587 1624 633
rect 1356 427 1364 473
rect 1396 427 1404 493
rect 1436 467 1444 533
rect 1516 427 1524 453
rect 1576 427 1584 533
rect 1636 427 1644 696
rect 1696 587 1704 733
rect 1736 647 1744 833
rect 1836 807 1844 933
rect 1816 707 1824 773
rect 1876 747 1884 913
rect 1896 707 1904 1213
rect 2076 1187 2084 1233
rect 2067 1176 2084 1187
rect 2067 1173 2080 1176
rect 1996 1087 2004 1153
rect 2116 1007 2124 1356
rect 2136 1247 2144 1293
rect 2196 1247 2204 1313
rect 2236 1287 2244 1393
rect 2256 1367 2264 1453
rect 2336 1407 2344 1573
rect 2136 1236 2153 1247
rect 2140 1233 2153 1236
rect 2216 1027 2224 1173
rect 2276 1167 2284 1273
rect 2296 1227 2304 1313
rect 2016 927 2024 973
rect 2136 947 2144 973
rect 1936 747 1944 873
rect 1976 847 1984 873
rect 2036 787 2044 873
rect 2096 847 2104 933
rect 2216 887 2224 1013
rect 2256 947 2264 1073
rect 2307 944 2320 947
rect 2307 933 2324 944
rect 2316 887 2324 933
rect 2216 876 2233 887
rect 2220 873 2233 876
rect 1807 696 1824 707
rect 1807 693 1820 696
rect 1887 696 1904 707
rect 1976 704 1984 773
rect 1956 696 1984 704
rect 1887 693 1900 696
rect 1696 467 1704 573
rect 1736 547 1744 633
rect 1756 527 1764 693
rect 1787 644 1800 647
rect 1787 640 1804 644
rect 1787 633 1807 640
rect 1793 627 1807 633
rect 1836 627 1844 693
rect 1956 647 1964 696
rect 1947 636 1964 647
rect 1996 644 2004 733
rect 2056 707 2064 773
rect 2116 684 2124 853
rect 2196 727 2204 753
rect 2236 727 2244 793
rect 2316 707 2324 813
rect 2096 676 2124 684
rect 2096 647 2104 676
rect 1996 636 2033 644
rect 1947 633 1960 636
rect 2087 636 2104 647
rect 2087 633 2100 636
rect 1896 607 1904 633
rect 2116 607 2124 653
rect 1696 427 1704 453
rect 1516 416 1533 427
rect 1520 413 1533 416
rect 1587 413 1604 427
rect 1636 424 1653 427
rect 1196 396 1253 404
rect 1196 384 1204 396
rect 1156 380 1204 384
rect 1153 376 1204 380
rect 1153 367 1167 376
rect 1596 367 1604 413
rect 1616 416 1653 424
rect 1567 364 1580 367
rect 1567 360 1584 364
rect 1567 353 1587 360
rect 1196 307 1204 353
rect 1296 227 1304 353
rect 1336 247 1344 353
rect 1416 327 1424 353
rect 1456 307 1464 353
rect 1573 347 1587 353
rect 1616 347 1624 416
rect 1640 413 1653 416
rect 1776 367 1784 433
rect 1813 427 1827 433
rect 1876 427 1884 453
rect 1996 427 2004 533
rect 2056 507 2064 553
rect 1813 420 1833 427
rect 1816 416 1833 420
rect 1820 413 1833 416
rect 1647 356 1673 364
rect 1816 327 1824 353
rect 1336 236 1353 247
rect 1340 233 1353 236
rect 1116 187 1124 213
rect 1373 187 1387 193
rect 1536 187 1544 233
rect 1576 187 1584 253
rect 1196 176 1273 184
rect 933 164 947 173
rect 933 160 1013 164
rect 936 156 1013 160
rect 1073 144 1087 153
rect 1196 147 1204 176
rect 1373 180 1393 187
rect 1376 176 1393 180
rect 1380 173 1393 176
rect 1216 156 1313 164
rect 1073 140 1133 144
rect 1076 136 1133 140
rect 1216 127 1224 156
rect 1356 127 1364 153
rect 1376 136 1444 144
rect 1376 127 1384 136
rect 1356 116 1373 127
rect 1360 113 1373 116
rect 956 87 964 113
rect 996 87 1004 113
rect 1036 47 1044 113
rect 1256 87 1264 113
rect 1296 47 1304 113
rect 1416 87 1424 113
rect 1436 104 1444 136
rect 1596 127 1604 213
rect 1796 207 1804 293
rect 1876 287 1884 413
rect 2016 327 2024 353
rect 1996 187 2004 273
rect 2016 267 2024 313
rect 2036 227 2044 413
rect 2076 204 2084 533
rect 2096 307 2104 513
rect 2140 424 2153 427
rect 2136 413 2153 424
rect 2207 424 2220 427
rect 2207 413 2224 424
rect 2136 307 2144 413
rect 2160 364 2173 367
rect 2156 360 2173 364
rect 2153 353 2173 360
rect 2153 347 2167 353
rect 2176 327 2184 353
rect 2216 304 2224 413
rect 2236 367 2244 593
rect 2356 447 2364 1573
rect 2376 1267 2384 1773
rect 2496 1747 2504 1913
rect 2536 1847 2544 1953
rect 2576 1787 2584 2013
rect 2596 1767 2604 2313
rect 2636 2207 2644 2293
rect 2656 2147 2664 2253
rect 2676 2127 2684 2476
rect 2736 2327 2744 2693
rect 2756 2647 2764 2713
rect 2796 2687 2804 2713
rect 2816 2704 2824 2773
rect 2816 2696 2844 2704
rect 2836 2647 2844 2696
rect 2856 2584 2864 2773
rect 2896 2627 2904 2873
rect 2856 2576 2884 2584
rect 2716 2267 2724 2293
rect 2696 2167 2704 2193
rect 2616 1927 2624 2113
rect 2736 2107 2744 2193
rect 2776 2087 2784 2473
rect 2796 2324 2804 2573
rect 2816 2447 2824 2533
rect 2796 2316 2813 2324
rect 2796 2107 2804 2292
rect 2816 2267 2824 2313
rect 2836 2307 2844 2373
rect 2856 2287 2864 2553
rect 2876 2307 2884 2576
rect 2916 2547 2924 3093
rect 2956 3067 2964 3093
rect 3016 3027 3024 3253
rect 3056 2967 3064 3276
rect 3156 3267 3164 3313
rect 3236 3307 3244 3473
rect 3276 3367 3284 3433
rect 3296 3407 3304 3533
rect 3336 3447 3344 3753
rect 3376 3707 3384 3753
rect 3436 3687 3444 3773
rect 3516 3607 3524 3953
rect 3236 3267 3244 3293
rect 3227 3256 3244 3267
rect 3227 3253 3240 3256
rect 3276 3207 3284 3293
rect 3316 3267 3324 3373
rect 3396 3367 3404 3393
rect 3416 3384 3424 3593
rect 3556 3587 3564 3913
rect 3616 3827 3624 3993
rect 3456 3427 3464 3573
rect 3527 3544 3540 3547
rect 3527 3533 3544 3544
rect 3416 3376 3444 3384
rect 3356 3327 3364 3353
rect 3396 3327 3404 3353
rect 3436 3307 3444 3376
rect 3476 3367 3484 3533
rect 3536 3487 3544 3533
rect 3496 3427 3504 3473
rect 3507 3416 3524 3424
rect 3516 3307 3524 3416
rect 3316 3256 3333 3267
rect 3320 3253 3333 3256
rect 2976 2747 2984 2893
rect 2956 2507 2964 2533
rect 2947 2496 2964 2507
rect 2947 2493 2960 2496
rect 2896 2387 2904 2493
rect 2916 2387 2924 2433
rect 2887 2204 2900 2207
rect 2887 2193 2904 2204
rect 2836 2127 2844 2193
rect 2896 2147 2904 2193
rect 2916 2167 2924 2253
rect 2816 2116 2833 2124
rect 2636 1987 2644 2073
rect 2676 1987 2684 2053
rect 2696 2027 2704 2073
rect 2816 2067 2824 2116
rect 2756 1964 2764 2053
rect 2836 1987 2844 2033
rect 2827 1976 2844 1987
rect 2827 1973 2840 1976
rect 2736 1956 2764 1964
rect 2696 1787 2704 1913
rect 2716 1787 2724 1833
rect 2736 1764 2744 1956
rect 2756 1767 2764 1933
rect 2776 1868 2784 1973
rect 2716 1756 2744 1764
rect 2567 1736 2624 1744
rect 2496 1684 2504 1733
rect 2496 1676 2533 1684
rect 2560 1684 2573 1687
rect 2556 1673 2573 1684
rect 2416 1567 2424 1673
rect 2456 1607 2464 1673
rect 2396 1467 2404 1513
rect 2396 1287 2404 1453
rect 2436 1327 2444 1453
rect 2376 944 2384 1013
rect 2396 1007 2404 1173
rect 2456 1124 2464 1213
rect 2476 1167 2484 1513
rect 2496 1447 2504 1593
rect 2556 1587 2564 1673
rect 2616 1667 2624 1736
rect 2716 1727 2724 1756
rect 2516 1184 2524 1393
rect 2556 1367 2564 1393
rect 2596 1387 2604 1433
rect 2616 1367 2624 1653
rect 2656 1628 2664 1713
rect 2776 1687 2784 1832
rect 2696 1627 2704 1653
rect 2736 1627 2744 1673
rect 2656 1387 2664 1592
rect 2716 1387 2724 1573
rect 2776 1547 2784 1673
rect 2816 1647 2824 1913
rect 2856 1884 2864 2133
rect 2956 2124 2964 2413
rect 2996 2328 3004 2953
rect 3036 2747 3044 2853
rect 3116 2847 3124 2953
rect 3156 2944 3164 3013
rect 3136 2936 3164 2944
rect 3096 2607 3104 2633
rect 3056 2447 3064 2553
rect 3096 2524 3104 2593
rect 3116 2567 3124 2833
rect 3136 2707 3144 2936
rect 3196 2924 3204 3153
rect 3236 3144 3244 3193
rect 3216 3136 3244 3144
rect 3216 3087 3224 3136
rect 3276 3004 3284 3193
rect 3376 3187 3384 3233
rect 3296 3007 3304 3173
rect 3416 3044 3424 3253
rect 3476 3247 3484 3293
rect 3536 3247 3544 3353
rect 3476 3236 3493 3247
rect 3480 3233 3493 3236
rect 3520 3244 3533 3247
rect 3516 3233 3533 3244
rect 3456 3187 3464 3213
rect 3516 3167 3524 3233
rect 3416 3040 3444 3044
rect 3416 3036 3447 3040
rect 3433 3027 3447 3036
rect 3247 2996 3284 3004
rect 3196 2916 3213 2924
rect 3156 2587 3164 2873
rect 3196 2807 3204 2873
rect 3216 2824 3224 2913
rect 3256 2884 3264 2996
rect 3276 2904 3284 2996
rect 3427 2956 3453 2964
rect 3276 2896 3304 2904
rect 3236 2880 3264 2884
rect 3233 2876 3264 2880
rect 3233 2867 3247 2876
rect 3276 2847 3284 2873
rect 3216 2820 3244 2824
rect 3216 2816 3247 2820
rect 3233 2807 3247 2816
rect 3296 2747 3304 2896
rect 3267 2744 3280 2747
rect 3267 2733 3284 2744
rect 3316 2736 3353 2744
rect 3176 2667 3184 2733
rect 3256 2627 3264 2673
rect 3276 2664 3284 2733
rect 3316 2724 3324 2736
rect 3296 2720 3324 2724
rect 3293 2716 3324 2720
rect 3293 2707 3307 2716
rect 3276 2656 3364 2664
rect 3076 2520 3104 2524
rect 3073 2516 3104 2520
rect 3073 2507 3087 2516
rect 3127 2500 3164 2504
rect 3127 2496 3167 2500
rect 3096 2388 3104 2413
rect 2996 2167 3004 2292
rect 3056 2207 3064 2293
rect 3016 2147 3024 2193
rect 3096 2187 3104 2352
rect 3116 2307 3124 2493
rect 3153 2487 3167 2496
rect 3156 2348 3164 2373
rect 3156 2127 3164 2312
rect 3196 2267 3204 2333
rect 3256 2327 3264 2433
rect 3296 2407 3304 2473
rect 3316 2364 3324 2613
rect 3356 2547 3364 2656
rect 3436 2647 3444 2893
rect 3496 2847 3504 2893
rect 3556 2884 3564 3293
rect 3576 2907 3584 3653
rect 3616 3647 3624 3813
rect 3656 3644 3664 3933
rect 3676 3667 3684 3813
rect 3656 3636 3684 3644
rect 3596 3547 3604 3573
rect 3656 3547 3664 3613
rect 3596 3536 3613 3547
rect 3600 3533 3613 3536
rect 3676 3487 3684 3636
rect 3596 3167 3604 3433
rect 3636 3267 3644 3333
rect 3676 3307 3684 3473
rect 3716 3367 3724 3473
rect 3676 3296 3693 3307
rect 3680 3293 3693 3296
rect 3656 3187 3664 3253
rect 3656 2927 3664 2953
rect 3536 2880 3564 2884
rect 3533 2876 3564 2880
rect 3533 2867 3547 2876
rect 3487 2776 3513 2784
rect 3436 2524 3444 2633
rect 3436 2516 3464 2524
rect 3436 2464 3444 2493
rect 3456 2484 3464 2516
rect 3456 2476 3484 2484
rect 3436 2456 3464 2464
rect 3296 2356 3324 2364
rect 3296 2267 3304 2356
rect 3316 2287 3324 2333
rect 3416 2327 3424 2433
rect 3376 2287 3384 2313
rect 3316 2276 3333 2287
rect 3320 2273 3333 2276
rect 3256 2227 3264 2253
rect 3247 2216 3264 2227
rect 3296 2227 3304 2253
rect 3296 2216 3313 2227
rect 3247 2213 3260 2216
rect 3300 2213 3313 2216
rect 2956 2120 2984 2124
rect 2956 2116 2987 2120
rect 2973 2107 2987 2116
rect 2836 1876 2864 1884
rect 2816 1587 2824 1633
rect 2687 1384 2700 1387
rect 2687 1373 2704 1384
rect 2727 1384 2740 1387
rect 2727 1373 2744 1384
rect 2696 1364 2704 1373
rect 2696 1356 2724 1364
rect 2496 1176 2524 1184
rect 2456 1120 2484 1124
rect 2456 1116 2487 1120
rect 2473 1107 2487 1116
rect 2496 1027 2504 1176
rect 2516 1087 2524 1153
rect 2536 1127 2544 1213
rect 2616 1167 2624 1353
rect 2656 1167 2664 1333
rect 2667 1164 2680 1167
rect 2667 1153 2684 1164
rect 2456 947 2464 1013
rect 2376 936 2413 944
rect 2496 887 2504 973
rect 2596 947 2604 993
rect 2396 847 2404 873
rect 2436 827 2444 853
rect 2536 827 2544 933
rect 2616 924 2624 1153
rect 2656 1007 2664 1113
rect 2636 947 2644 973
rect 2596 916 2624 924
rect 2596 864 2604 916
rect 2627 884 2640 887
rect 2627 873 2644 884
rect 2596 856 2624 864
rect 2396 707 2404 733
rect 2496 647 2504 733
rect 2556 727 2564 773
rect 2596 708 2604 773
rect 2376 507 2384 633
rect 2416 587 2424 633
rect 2496 527 2504 633
rect 2536 607 2544 633
rect 2556 507 2564 533
rect 2387 416 2444 424
rect 2320 404 2333 407
rect 2316 393 2333 404
rect 2316 327 2324 393
rect 2356 307 2364 333
rect 2396 307 2404 333
rect 2196 296 2224 304
rect 2136 247 2144 293
rect 2196 207 2204 296
rect 2396 267 2404 293
rect 2416 247 2424 393
rect 2436 344 2444 416
rect 2516 347 2524 493
rect 2436 336 2493 344
rect 2516 333 2533 347
rect 2516 287 2524 333
rect 2596 327 2604 672
rect 2616 587 2624 856
rect 2636 827 2644 873
rect 2636 687 2644 733
rect 2656 647 2664 753
rect 2676 747 2684 1153
rect 2696 787 2704 1333
rect 2716 1227 2724 1356
rect 2736 1347 2744 1373
rect 2816 1367 2824 1573
rect 2776 1267 2784 1333
rect 2836 1287 2844 1876
rect 2856 1727 2864 1853
rect 2916 1847 2924 2033
rect 3016 1967 3024 2053
rect 2916 1687 2924 1833
rect 2956 1807 2964 1953
rect 2996 1867 3004 1913
rect 2916 1676 2933 1687
rect 2920 1673 2933 1676
rect 2896 1647 2904 1673
rect 2956 1647 2964 1793
rect 2876 1507 2884 1613
rect 2896 1447 2904 1513
rect 2876 1367 2884 1393
rect 2916 1347 2924 1613
rect 2956 1347 2964 1373
rect 2956 1307 2964 1333
rect 2996 1307 3004 1373
rect 2736 1167 2744 1193
rect 2736 1156 2753 1167
rect 2740 1153 2753 1156
rect 2796 1127 2804 1153
rect 2716 767 2724 993
rect 2736 724 2744 1113
rect 2816 1107 2824 1213
rect 2816 987 2824 1093
rect 2756 847 2764 873
rect 2836 807 2844 1273
rect 2856 947 2864 1053
rect 2876 1047 2884 1253
rect 2896 1167 2904 1293
rect 2936 1127 2944 1153
rect 3016 1107 3024 1793
rect 3036 1767 3044 1813
rect 3056 1807 3064 2093
rect 3196 2044 3204 2133
rect 3136 2036 3204 2044
rect 3136 2007 3144 2036
rect 3136 1984 3144 1993
rect 3216 1984 3224 2053
rect 3116 1980 3144 1984
rect 3196 1980 3224 1984
rect 3113 1976 3144 1980
rect 3193 1976 3224 1980
rect 3113 1967 3127 1976
rect 3193 1967 3207 1976
rect 3096 1847 3104 1953
rect 3136 1867 3144 1893
rect 3173 1884 3187 1893
rect 3213 1884 3227 1893
rect 3236 1887 3244 2113
rect 3173 1880 3227 1884
rect 3176 1876 3224 1880
rect 3096 1767 3104 1793
rect 3036 1756 3053 1767
rect 3040 1753 3053 1756
rect 3056 1724 3064 1753
rect 3056 1716 3084 1724
rect 2916 1024 2924 1093
rect 3036 1027 3044 1533
rect 3056 1328 3064 1693
rect 3076 1667 3084 1716
rect 3116 1647 3124 1813
rect 3196 1807 3204 1853
rect 3056 1167 3064 1292
rect 3076 1267 3084 1573
rect 3096 1467 3104 1513
rect 3116 1407 3124 1633
rect 3136 1587 3144 1793
rect 3236 1744 3244 1793
rect 3187 1736 3244 1744
rect 3176 1587 3184 1653
rect 3196 1627 3204 1693
rect 3256 1647 3264 1993
rect 3276 1948 3284 2133
rect 3316 2027 3324 2213
rect 3396 2187 3404 2213
rect 3436 2187 3444 2393
rect 3356 2027 3364 2153
rect 3456 2087 3464 2456
rect 3476 2127 3484 2476
rect 3316 1987 3324 2013
rect 3340 1984 3353 1987
rect 3336 1973 3353 1984
rect 3256 1527 3264 1633
rect 3136 1467 3144 1513
rect 3276 1467 3284 1912
rect 3296 1507 3304 1893
rect 3336 1847 3344 1973
rect 3376 1807 3384 1873
rect 3316 1647 3324 1733
rect 3336 1607 3344 1633
rect 3356 1547 3364 1713
rect 3276 1456 3293 1467
rect 3280 1453 3293 1456
rect 3333 1444 3347 1453
rect 3333 1440 3364 1444
rect 3336 1436 3367 1440
rect 3353 1427 3367 1436
rect 3376 1407 3384 1733
rect 3396 1727 3404 2013
rect 3416 1867 3424 2073
rect 3496 2067 3504 2673
rect 3516 2507 3524 2593
rect 3536 2547 3544 2713
rect 3576 2547 3584 2853
rect 3516 2496 3533 2507
rect 3520 2493 3533 2496
rect 3616 2447 3624 2893
rect 3636 2528 3644 2773
rect 3656 2607 3664 2733
rect 3676 2627 3684 2993
rect 3716 2827 3724 3253
rect 3716 2587 3724 2673
rect 3516 2267 3524 2393
rect 3556 2287 3564 2373
rect 3596 2327 3604 2393
rect 3596 2287 3604 2313
rect 3636 2287 3644 2492
rect 3656 2367 3664 2473
rect 3716 2387 3724 2573
rect 3736 2507 3744 3953
rect 3796 3787 3804 3893
rect 3816 3527 3824 3993
rect 3856 3947 3864 4053
rect 3956 3968 3964 4053
rect 4016 3987 4024 4053
rect 3916 3927 3924 3953
rect 3916 3827 3924 3913
rect 3856 3687 3864 3773
rect 3756 3147 3764 3353
rect 3836 3347 3844 3373
rect 3896 3347 3904 3513
rect 3916 3304 3924 3653
rect 3936 3427 3944 3633
rect 3956 3487 3964 3932
rect 3907 3296 3933 3304
rect 3976 3227 3984 3913
rect 3996 3667 4004 3953
rect 4036 3787 4044 3933
rect 4013 3624 4027 3633
rect 3996 3620 4027 3624
rect 3996 3616 4024 3620
rect 3996 3547 4004 3616
rect 4056 3607 4064 4153
rect 4176 4127 4184 4376
rect 4196 4207 4204 4353
rect 4236 4347 4244 4393
rect 4316 4304 4324 4693
rect 4336 4607 4344 4776
rect 4376 4587 4384 4633
rect 4427 4584 4440 4587
rect 4427 4573 4444 4584
rect 4436 4527 4444 4573
rect 4456 4504 4464 4753
rect 4496 4707 4504 4776
rect 4536 4627 4544 4753
rect 4567 4584 4580 4587
rect 4567 4573 4584 4584
rect 4396 4496 4464 4504
rect 4356 4424 4364 4493
rect 4356 4416 4384 4424
rect 4356 4347 4364 4393
rect 4296 4296 4324 4304
rect 4376 4304 4384 4416
rect 4396 4304 4404 4496
rect 4476 4347 4484 4453
rect 4516 4387 4524 4573
rect 4576 4547 4584 4573
rect 4467 4336 4484 4347
rect 4467 4333 4480 4336
rect 4376 4296 4404 4304
rect 4296 4204 4304 4296
rect 4347 4284 4360 4287
rect 4347 4273 4364 4284
rect 4356 4227 4364 4273
rect 4376 4247 4384 4273
rect 4396 4267 4404 4296
rect 4396 4256 4413 4267
rect 4400 4253 4413 4256
rect 4296 4196 4324 4204
rect 4100 4064 4113 4067
rect 4096 4053 4113 4064
rect 4096 4027 4104 4053
rect 4076 3996 4133 4004
rect 4076 3947 4084 3996
rect 4096 3947 4104 3973
rect 4156 3947 4164 4053
rect 4176 4007 4184 4113
rect 4096 3747 4104 3773
rect 4096 3687 4104 3733
rect 4036 3547 4044 3573
rect 3756 2827 3764 3133
rect 3756 2787 3764 2813
rect 3776 2587 3784 2873
rect 3796 2607 3804 3113
rect 3816 3027 3824 3073
rect 3816 2687 3824 3013
rect 3656 2224 3664 2353
rect 3716 2347 3724 2373
rect 3696 2227 3704 2273
rect 3716 2267 3724 2333
rect 3756 2284 3764 2553
rect 3836 2507 3844 3113
rect 3856 2867 3864 2993
rect 3896 2967 3904 3213
rect 3916 3007 3924 3133
rect 3896 2867 3904 2953
rect 3936 2907 3944 2953
rect 3996 2864 4004 3533
rect 4036 3047 4044 3433
rect 4076 3347 4084 3513
rect 4116 3367 4124 3633
rect 4156 3367 4164 3673
rect 4056 3227 4064 3253
rect 4056 3127 4064 3213
rect 3976 2856 4004 2864
rect 3856 2787 3864 2813
rect 3976 2747 3984 2856
rect 4016 2747 4024 3013
rect 4056 2807 4064 3053
rect 4076 3028 4084 3253
rect 4116 3087 4124 3153
rect 4116 3027 4124 3073
rect 4076 2887 4084 2992
rect 4136 2807 4144 3333
rect 4156 3027 4164 3113
rect 4176 3067 4184 3413
rect 4216 3387 4224 4073
rect 4236 3907 4244 4093
rect 4276 4007 4284 4173
rect 4316 4087 4324 4196
rect 4416 4167 4424 4213
rect 4296 3947 4304 4033
rect 4376 3787 4384 4153
rect 4436 4047 4444 4233
rect 4416 3967 4424 3993
rect 4367 3776 4384 3787
rect 4367 3773 4380 3776
rect 4216 3307 4224 3373
rect 4256 3327 4264 3593
rect 4296 3527 4304 3773
rect 4436 3727 4444 3933
rect 4456 3827 4464 4253
rect 4476 3927 4484 4273
rect 4516 4247 4524 4273
rect 4516 3827 4524 3873
rect 4456 3816 4473 3827
rect 4460 3813 4473 3816
rect 4556 3807 4564 4193
rect 4496 3727 4504 3753
rect 4296 3327 4304 3413
rect 4236 3227 4244 3253
rect 4273 3224 4287 3233
rect 4316 3227 4324 3253
rect 4273 3220 4304 3224
rect 4276 3216 4304 3220
rect 4216 2967 4224 3053
rect 4236 2864 4244 3213
rect 4296 3207 4304 3216
rect 4296 3084 4304 3193
rect 4296 3076 4324 3084
rect 4256 3027 4264 3073
rect 4296 3027 4304 3053
rect 4256 2907 4264 3013
rect 4316 2967 4324 3076
rect 4236 2856 4264 2864
rect 3856 2547 3864 2673
rect 4016 2647 4024 2733
rect 4056 2668 4064 2793
rect 4067 2656 4084 2664
rect 3916 2547 3924 2573
rect 3936 2507 3944 2633
rect 3976 2507 3984 2553
rect 3776 2307 3784 2413
rect 3796 2324 3804 2493
rect 3796 2316 3824 2324
rect 3756 2276 3784 2284
rect 3716 2256 3733 2267
rect 3720 2253 3733 2256
rect 3627 2216 3664 2224
rect 3536 2187 3544 2213
rect 3476 2056 3493 2064
rect 3436 1767 3444 2013
rect 3456 1764 3464 1973
rect 3476 1787 3484 2056
rect 3516 2027 3524 2133
rect 3496 1867 3504 1973
rect 3456 1756 3484 1764
rect 3476 1704 3484 1756
rect 3516 1747 3524 1833
rect 3536 1807 3544 2093
rect 3556 1924 3564 2113
rect 3616 1987 3624 2073
rect 3556 1916 3593 1924
rect 3476 1696 3564 1704
rect 3427 1676 3453 1684
rect 3496 1647 3504 1673
rect 3156 1347 3164 1373
rect 3116 1167 3124 1253
rect 3107 1156 3124 1167
rect 3107 1153 3120 1156
rect 3056 1127 3064 1153
rect 2916 1016 2944 1024
rect 2896 947 2904 993
rect 2736 716 2764 724
rect 2727 704 2740 707
rect 2727 693 2744 704
rect 2736 647 2744 693
rect 2696 607 2704 633
rect 2696 427 2704 553
rect 2056 196 2084 204
rect 1727 176 1753 184
rect 1767 176 1833 184
rect 1887 176 1913 184
rect 1436 100 1464 104
rect 1436 96 1467 100
rect 1453 87 1467 96
rect 1556 87 1564 113
rect 1736 67 1744 113
rect 1776 67 1784 113
rect 1896 87 1904 113
rect 1936 67 1944 113
rect 2056 47 2064 196
rect 2236 187 2244 213
rect 2096 27 2104 173
rect 2296 144 2304 213
rect 2327 176 2353 184
rect 2256 140 2304 144
rect 2253 136 2304 140
rect 2253 127 2267 136
rect 2187 116 2213 124
rect 2296 124 2304 136
rect 2376 127 2384 233
rect 2296 116 2333 124
rect 2376 27 2384 113
rect 2416 87 2424 173
rect 2476 127 2484 233
rect 2636 187 2644 353
rect 2656 287 2664 413
rect 2736 367 2744 573
rect 2756 227 2764 716
rect 2696 187 2704 213
rect 2476 116 2493 127
rect 2480 113 2493 116
rect 2516 47 2524 173
rect 2536 27 2544 113
rect 2696 27 2704 173
rect 2776 144 2784 753
rect 2796 707 2804 793
rect 2856 707 2864 773
rect 2916 667 2924 753
rect 2913 644 2927 653
rect 2887 640 2927 644
rect 2887 636 2924 640
rect 2836 567 2844 633
rect 2936 627 2944 1016
rect 2956 707 2964 1013
rect 3096 1007 3104 1093
rect 3156 1027 3164 1333
rect 3276 1327 3284 1393
rect 3316 1348 3324 1373
rect 3216 1287 3224 1313
rect 3216 1227 3224 1273
rect 3016 947 3024 973
rect 3076 947 3084 973
rect 3176 947 3184 1093
rect 3276 1047 3284 1153
rect 3296 1007 3304 1253
rect 3316 1227 3324 1312
rect 3336 1267 3344 1333
rect 3376 1227 3384 1353
rect 3396 1267 3404 1593
rect 3516 1587 3524 1613
rect 3340 1164 3353 1167
rect 3336 1153 3353 1164
rect 3336 1107 3344 1153
rect 3396 1047 3404 1153
rect 3416 1107 3424 1333
rect 3456 1087 3464 1573
rect 3496 1407 3504 1533
rect 3496 1227 3504 1353
rect 3496 1216 3513 1227
rect 3500 1213 3513 1216
rect 3536 1127 3544 1653
rect 3556 1607 3564 1696
rect 3556 1467 3564 1513
rect 3576 1407 3584 1633
rect 3596 1547 3604 1873
rect 3636 1867 3644 2053
rect 3656 1987 3664 2113
rect 3636 1767 3644 1853
rect 3676 1807 3684 2173
rect 3756 2127 3764 2193
rect 3716 1804 3724 2073
rect 3776 2067 3784 2276
rect 3796 1987 3804 2173
rect 3816 2064 3824 2316
rect 3876 2287 3884 2433
rect 3916 2327 3924 2493
rect 3936 2287 3944 2433
rect 4056 2407 4064 2632
rect 4076 2568 4084 2656
rect 4116 2627 4124 2673
rect 4136 2647 4144 2793
rect 4173 2787 4187 2793
rect 4173 2780 4193 2787
rect 4176 2776 4193 2780
rect 4180 2773 4193 2776
rect 4176 2688 4184 2713
rect 4216 2667 4224 2713
rect 4256 2704 4264 2856
rect 4236 2700 4264 2704
rect 4233 2696 4264 2700
rect 4233 2687 4247 2696
rect 4276 2688 4284 2933
rect 4156 2607 4164 2633
rect 4076 2507 4084 2532
rect 4116 2507 4124 2573
rect 4076 2496 4093 2507
rect 4080 2493 4093 2496
rect 4116 2496 4133 2507
rect 4120 2493 4133 2496
rect 3876 2276 3893 2287
rect 3880 2273 3893 2276
rect 4016 2227 4024 2353
rect 4056 2267 4064 2393
rect 4076 2367 4084 2433
rect 3836 2087 3844 2213
rect 3816 2056 3844 2064
rect 3740 1984 3753 1987
rect 3736 1973 3753 1984
rect 3736 1948 3744 1973
rect 3747 1916 3773 1924
rect 3836 1887 3844 2056
rect 3896 1987 3904 2113
rect 3936 2047 3944 2153
rect 4036 1987 4044 2113
rect 3896 1984 3913 1987
rect 3876 1976 3913 1984
rect 3716 1796 3744 1804
rect 3693 1767 3707 1773
rect 3687 1764 3707 1767
rect 3687 1756 3724 1764
rect 3687 1753 3700 1756
rect 3616 1628 3624 1693
rect 3616 1387 3624 1592
rect 3636 1347 3644 1593
rect 3656 1564 3664 1673
rect 3696 1647 3704 1693
rect 3656 1556 3684 1564
rect 3656 1484 3664 1533
rect 3676 1527 3684 1556
rect 3716 1524 3724 1756
rect 3736 1667 3744 1796
rect 3776 1607 3784 1853
rect 3816 1827 3824 1853
rect 3816 1687 3824 1813
rect 3876 1807 3884 1976
rect 3900 1973 3913 1976
rect 3967 1976 3993 1984
rect 3896 1827 3904 1913
rect 3916 1767 3924 1873
rect 3936 1787 3944 1833
rect 3856 1647 3864 1673
rect 3907 1636 3933 1644
rect 3747 1584 3760 1587
rect 3747 1573 3764 1584
rect 3756 1567 3764 1573
rect 3756 1556 3773 1567
rect 3760 1553 3773 1556
rect 3696 1516 3724 1524
rect 3696 1507 3707 1516
rect 3706 1500 3707 1507
rect 3713 1493 3714 1500
rect 3713 1484 3727 1493
rect 3656 1480 3727 1484
rect 3656 1476 3724 1480
rect 3736 1467 3744 1533
rect 3876 1467 3884 1613
rect 3916 1507 3924 1533
rect 3916 1467 3924 1493
rect 3680 1464 3693 1467
rect 3676 1453 3693 1464
rect 3676 1427 3684 1453
rect 3696 1416 3744 1424
rect 3696 1387 3704 1416
rect 3716 1367 3724 1393
rect 3487 1116 3524 1124
rect 3396 1007 3404 1033
rect 3436 1027 3444 1073
rect 3516 1047 3524 1116
rect 3556 1027 3564 1253
rect 3676 1227 3684 1273
rect 3596 1167 3604 1213
rect 3596 1156 3613 1167
rect 3600 1153 3613 1156
rect 3427 1016 3444 1027
rect 3427 1013 3440 1016
rect 3196 947 3204 973
rect 3316 947 3324 973
rect 3456 947 3464 973
rect 3067 936 3084 947
rect 3067 933 3080 936
rect 3167 936 3184 947
rect 3167 933 3180 936
rect 3367 944 3380 947
rect 3367 933 3384 944
rect 3456 936 3473 947
rect 3460 933 3473 936
rect 3527 944 3540 947
rect 3527 933 3544 944
rect 2976 607 2984 873
rect 3016 847 3024 933
rect 3036 827 3044 873
rect 3176 847 3184 873
rect 2996 707 3004 793
rect 3056 727 3064 793
rect 3076 747 3084 793
rect 3216 767 3224 833
rect 3236 747 3244 873
rect 3376 847 3384 933
rect 3536 887 3544 933
rect 3467 876 3524 884
rect 3127 716 3153 724
rect 3207 716 3264 724
rect 3233 684 3247 693
rect 3256 687 3264 716
rect 3276 707 3284 773
rect 3336 727 3344 813
rect 3376 727 3384 833
rect 3216 680 3247 684
rect 3213 676 3244 680
rect 3213 667 3227 676
rect 3327 676 3404 684
rect 3036 627 3044 653
rect 3136 627 3144 653
rect 3396 647 3404 676
rect 3456 647 3464 813
rect 3496 787 3504 853
rect 3496 707 3504 773
rect 3516 647 3524 876
rect 3536 847 3544 873
rect 3576 847 3584 1153
rect 3656 1127 3664 1153
rect 3456 636 3473 647
rect 3460 633 3473 636
rect 2840 424 2853 427
rect 2836 413 2853 424
rect 2836 287 2844 413
rect 2876 307 2884 353
rect 2896 327 2904 413
rect 2936 367 2944 473
rect 3016 427 3024 473
rect 3056 427 3064 513
rect 3036 327 3044 353
rect 2796 207 2804 273
rect 2856 187 2864 253
rect 2956 187 2964 253
rect 2996 207 3004 313
rect 3096 267 3104 573
rect 3176 487 3184 633
rect 3216 366 3224 573
rect 3236 427 3244 593
rect 3296 507 3304 633
rect 3556 527 3564 793
rect 3276 366 3284 473
rect 3436 427 3444 513
rect 3456 367 3464 453
rect 3487 424 3500 427
rect 3487 413 3504 424
rect 2847 176 2864 187
rect 2847 173 2860 176
rect 2756 136 2784 144
rect 2816 156 2873 164
rect 2756 -16 2764 136
rect 2816 127 2824 156
rect 2916 127 2924 153
rect 2936 136 3013 144
rect 2936 127 2944 136
rect 2787 116 2813 124
rect 2916 116 2933 127
rect 2920 113 2933 116
rect 2856 67 2864 113
rect 2976 67 2984 113
rect 3056 47 3064 253
rect 3136 204 3144 293
rect 3076 196 3144 204
rect 3076 167 3084 196
rect 3100 184 3113 187
rect 3096 173 3113 184
rect 3096 147 3104 173
rect 3176 127 3184 233
rect 3136 27 3144 113
rect 3126 13 3127 20
rect 3113 4 3127 13
rect 3113 0 3184 4
rect 3116 -4 3184 0
rect 2756 -24 2784 -16
rect 3176 -36 3184 -4
rect 3196 -24 3204 213
rect 3276 187 3284 253
rect 3336 187 3344 233
rect 3216 -36 3224 93
rect 3296 -24 3304 133
rect 3376 107 3384 253
rect 3416 247 3424 333
rect 3496 327 3504 413
rect 3536 287 3544 453
rect 3596 444 3604 1013
rect 3656 947 3664 1113
rect 3696 1087 3704 1113
rect 3716 1087 3724 1253
rect 3736 1027 3744 1416
rect 3836 1407 3844 1433
rect 3836 1396 3853 1407
rect 3840 1393 3853 1396
rect 3756 1287 3764 1333
rect 3756 1227 3764 1273
rect 3816 1267 3824 1393
rect 3936 1287 3944 1612
rect 3956 1607 3964 1673
rect 3976 1507 3984 1613
rect 3996 1567 4004 1673
rect 4016 1627 4024 1913
rect 4036 1707 4044 1813
rect 4056 1667 4064 2133
rect 4116 2047 4124 2373
rect 4136 2027 4144 2433
rect 4127 1984 4140 1987
rect 4127 1973 4144 1984
rect 4076 1887 4084 1973
rect 4136 1947 4144 1973
rect 4076 1747 4084 1813
rect 4156 1767 4164 2553
rect 4176 2087 4184 2652
rect 4196 2587 4204 2613
rect 4196 2367 4204 2493
rect 4236 2327 4244 2633
rect 4276 2447 4284 2652
rect 4296 2607 4304 2813
rect 4336 2727 4344 3173
rect 4356 3147 4364 3613
rect 4436 3587 4444 3713
rect 4436 3547 4444 3573
rect 4396 3447 4404 3533
rect 4416 3307 4424 3373
rect 4456 3187 4464 3413
rect 4496 3267 4504 3613
rect 4536 3487 4544 3753
rect 4516 3367 4524 3433
rect 4556 3347 4564 3713
rect 4576 3607 4584 4333
rect 4596 4147 4604 4856
rect 4627 4804 4640 4807
rect 4627 4793 4644 4804
rect 4636 4667 4644 4793
rect 4656 4484 4664 4956
rect 4696 4947 4704 4993
rect 4716 4907 4724 5033
rect 4736 4927 4744 4973
rect 4816 4967 4824 5073
rect 4856 5047 4864 5153
rect 5016 5107 5024 5356
rect 5056 5087 5064 5293
rect 5076 5287 5084 5313
rect 5076 5227 5084 5273
rect 5056 5076 5073 5087
rect 5060 5073 5073 5076
rect 5116 5047 5124 5313
rect 5196 5247 5204 5953
rect 5256 5907 5264 5933
rect 5313 5844 5327 5853
rect 5287 5840 5327 5844
rect 5287 5836 5324 5840
rect 5236 5767 5244 5833
rect 5336 5784 5344 6053
rect 5456 5987 5464 6093
rect 5436 5927 5444 5953
rect 5393 5904 5407 5913
rect 5393 5900 5424 5904
rect 5396 5896 5424 5900
rect 5336 5780 5364 5784
rect 5336 5776 5367 5780
rect 5353 5767 5367 5776
rect 5216 5427 5224 5733
rect 5236 5567 5244 5713
rect 5233 5544 5247 5553
rect 5233 5540 5264 5544
rect 5236 5536 5264 5540
rect 5216 5287 5224 5333
rect 5216 5107 5224 5273
rect 5187 5104 5200 5107
rect 5187 5093 5204 5104
rect 4907 5044 4920 5047
rect 4907 5033 4924 5044
rect 4916 4984 4924 5033
rect 4896 4976 4924 4984
rect 4807 4864 4820 4867
rect 4836 4864 4844 4913
rect 4896 4907 4904 4976
rect 4936 4867 4944 4913
rect 4807 4853 4824 4864
rect 4836 4856 4864 4864
rect 4816 4804 4824 4853
rect 4816 4796 4844 4804
rect 4696 4527 4704 4713
rect 4736 4707 4744 4793
rect 4776 4527 4784 4793
rect 4796 4748 4804 4773
rect 4836 4747 4844 4796
rect 4796 4587 4804 4712
rect 4836 4587 4844 4633
rect 4696 4513 4713 4527
rect 4696 4487 4704 4513
rect 4636 4476 4664 4484
rect 4616 4067 4624 4453
rect 4636 4187 4644 4476
rect 4656 4347 4664 4433
rect 4656 4247 4664 4273
rect 4696 4187 4704 4273
rect 4716 4247 4724 4453
rect 4756 4127 4764 4373
rect 4776 4247 4784 4473
rect 4796 4147 4804 4573
rect 4836 4487 4844 4573
rect 4856 4444 4864 4856
rect 4996 4827 5004 4853
rect 4987 4816 5004 4827
rect 4987 4813 5000 4816
rect 4896 4744 4904 4813
rect 4976 4747 4984 4813
rect 5016 4787 5024 4893
rect 5056 4807 5064 4953
rect 5096 4907 5104 4973
rect 4876 4736 4904 4744
rect 4876 4667 4884 4736
rect 4896 4667 4904 4693
rect 4847 4436 4864 4444
rect 4816 4347 4824 4373
rect 4816 4104 4824 4233
rect 4807 4096 4824 4104
rect 4596 3687 4604 3893
rect 4616 3727 4624 3993
rect 4616 3627 4624 3713
rect 4616 3547 4624 3613
rect 4576 3367 4584 3533
rect 4616 3427 4624 3473
rect 4636 3447 4644 4073
rect 4796 4047 4804 4093
rect 4696 3887 4704 3933
rect 4656 3767 4664 3873
rect 4676 3827 4684 3853
rect 4716 3767 4724 4033
rect 4756 4004 4764 4033
rect 4756 3996 4784 4004
rect 4707 3753 4724 3767
rect 4696 3727 4704 3753
rect 4656 3627 4664 3653
rect 4696 3547 4704 3633
rect 4736 3567 4744 3973
rect 4776 3947 4784 3996
rect 4776 3937 4793 3947
rect 4780 3934 4793 3937
rect 4780 3933 4800 3934
rect 4756 3727 4764 3913
rect 4796 3867 4804 3912
rect 4836 3887 4844 4433
rect 4876 4107 4884 4153
rect 4876 4067 4884 4093
rect 4896 4087 4904 4653
rect 4996 4587 5004 4693
rect 5096 4627 5104 4793
rect 5136 4687 5144 4893
rect 5156 4727 5164 4993
rect 5176 4784 5184 4853
rect 5196 4827 5204 5093
rect 5220 5024 5233 5027
rect 5216 5013 5233 5024
rect 5216 4867 5224 5013
rect 5256 5007 5264 5536
rect 5296 5487 5304 5753
rect 5336 5467 5344 5693
rect 5276 5387 5284 5453
rect 5356 5447 5364 5713
rect 5416 5667 5424 5896
rect 5476 5807 5484 6273
rect 5656 6107 5664 6253
rect 5596 5967 5604 6053
rect 5536 5827 5544 5853
rect 5376 5527 5384 5553
rect 5436 5527 5444 5793
rect 5456 5627 5464 5653
rect 5507 5624 5520 5627
rect 5507 5613 5524 5624
rect 5336 5347 5344 5393
rect 5376 5327 5384 5453
rect 5396 5427 5404 5453
rect 5396 5387 5404 5413
rect 5276 4887 5284 5273
rect 5436 5047 5444 5513
rect 5476 5507 5484 5553
rect 5516 5507 5524 5613
rect 5556 5447 5564 5953
rect 5636 5947 5644 6033
rect 5716 6024 5724 6353
rect 5696 6016 5724 6024
rect 5576 5907 5584 5933
rect 5616 5847 5624 5893
rect 5607 5836 5624 5847
rect 5607 5833 5620 5836
rect 5576 5527 5584 5793
rect 5656 5627 5664 5653
rect 5600 5624 5613 5627
rect 5596 5613 5613 5624
rect 5596 5447 5604 5613
rect 5636 5527 5644 5553
rect 5496 5407 5504 5433
rect 5556 5424 5564 5433
rect 5616 5427 5624 5493
rect 5696 5427 5704 6016
rect 5776 5907 5784 5953
rect 5716 5767 5724 5833
rect 5756 5707 5764 5833
rect 5816 5827 5824 6293
rect 5836 6267 5844 6353
rect 5936 6307 5944 6433
rect 6016 6387 6024 6453
rect 6040 6424 6053 6427
rect 6036 6413 6053 6424
rect 6036 6367 6044 6413
rect 6076 6367 6084 6453
rect 5836 5907 5844 6253
rect 5876 6147 5884 6193
rect 5916 6147 5924 6233
rect 6056 6147 6064 6333
rect 5856 6007 5864 6073
rect 5936 6027 5944 6073
rect 6016 6007 6024 6073
rect 5896 5907 5904 5973
rect 6016 5907 6024 5933
rect 6056 5907 6064 5953
rect 5836 5896 5853 5907
rect 5840 5893 5853 5896
rect 5860 5844 5873 5847
rect 5856 5840 5873 5844
rect 5853 5833 5873 5840
rect 5853 5827 5867 5833
rect 5716 5467 5724 5653
rect 5836 5627 5844 5793
rect 5876 5704 5884 5753
rect 5916 5747 5924 5833
rect 6016 5807 6024 5893
rect 5876 5696 5904 5704
rect 5776 5527 5784 5553
rect 5796 5507 5804 5613
rect 5556 5416 5584 5424
rect 5536 5227 5544 5393
rect 5576 5384 5584 5416
rect 5776 5387 5784 5473
rect 5896 5467 5904 5696
rect 6056 5644 6064 5753
rect 6016 5640 6064 5644
rect 6013 5636 6064 5640
rect 6013 5627 6027 5636
rect 5960 5624 5973 5627
rect 5956 5613 5973 5624
rect 5956 5587 5964 5613
rect 5936 5447 5944 5553
rect 6036 5528 6044 5553
rect 6076 5527 6084 5833
rect 6096 5768 6104 6173
rect 6116 5947 6124 6333
rect 6156 6327 6164 6413
rect 6176 6367 6184 6556
rect 6196 6447 6204 6556
rect 6236 6527 6244 6564
rect 6196 6436 6213 6447
rect 6200 6433 6213 6436
rect 6196 6207 6204 6373
rect 6256 6267 6264 6433
rect 6156 6127 6164 6153
rect 6196 6084 6204 6193
rect 6236 6127 6244 6153
rect 6176 6080 6204 6084
rect 6173 6076 6204 6080
rect 6173 6067 6187 6076
rect 6216 6027 6224 6053
rect 6176 5864 6184 5973
rect 6216 5947 6224 6013
rect 6276 5927 6284 6513
rect 6376 6427 6384 6453
rect 6367 6364 6380 6367
rect 6367 6353 6384 6364
rect 6316 6087 6324 6233
rect 6313 5964 6327 5973
rect 6336 5964 6344 6253
rect 6313 5960 6344 5964
rect 6316 5956 6344 5960
rect 6316 5927 6324 5956
rect 6276 5924 6293 5927
rect 6256 5916 6293 5924
rect 6256 5904 6264 5916
rect 6227 5896 6264 5904
rect 6276 5913 6293 5916
rect 6316 5916 6333 5927
rect 6320 5913 6333 5916
rect 6156 5860 6184 5864
rect 6153 5856 6184 5860
rect 6153 5847 6167 5856
rect 6196 5807 6204 5833
rect 6096 5607 6104 5732
rect 6176 5607 6184 5753
rect 6176 5596 6193 5607
rect 6180 5593 6193 5596
rect 6167 5564 6180 5567
rect 6167 5553 6184 5564
rect 5976 5407 5984 5473
rect 5896 5400 5933 5404
rect 5576 5376 5633 5384
rect 5767 5376 5784 5387
rect 5893 5396 5933 5400
rect 5893 5387 5907 5396
rect 5767 5373 5780 5376
rect 5656 5287 5664 5313
rect 5296 4947 5304 5033
rect 5313 5004 5327 5013
rect 5476 5007 5484 5093
rect 5513 5084 5527 5093
rect 5556 5084 5564 5233
rect 5656 5144 5664 5273
rect 5716 5267 5724 5373
rect 5647 5136 5664 5144
rect 5513 5080 5564 5084
rect 5516 5076 5564 5080
rect 5313 5000 5344 5004
rect 5316 4996 5347 5000
rect 5333 4987 5347 4996
rect 5276 4876 5293 4887
rect 5280 4873 5293 4876
rect 5176 4776 5204 4784
rect 5196 4667 5204 4776
rect 5236 4647 5244 4813
rect 5256 4787 5264 4873
rect 5316 4827 5324 4953
rect 5276 4667 5284 4793
rect 4956 4487 4964 4573
rect 4936 4367 4944 4453
rect 5016 4447 5024 4613
rect 5296 4587 5304 4613
rect 5096 4467 5104 4573
rect 5136 4487 5144 4573
rect 5156 4427 5164 4513
rect 5256 4467 5264 4573
rect 5316 4544 5324 4773
rect 5336 4767 5344 4853
rect 5416 4807 5424 4973
rect 5436 4927 5444 4953
rect 5476 4867 5484 4913
rect 5456 4767 5464 4793
rect 5316 4536 5344 4544
rect 5287 4524 5300 4527
rect 5287 4513 5304 4524
rect 5296 4487 5304 4513
rect 4976 4227 4984 4333
rect 5007 4284 5020 4287
rect 5007 4273 5024 4284
rect 5016 4207 5024 4273
rect 4916 4127 4924 4193
rect 5056 4187 5064 4413
rect 5216 4347 5224 4373
rect 5296 4347 5304 4473
rect 5336 4467 5344 4536
rect 5376 4527 5384 4693
rect 5396 4627 5404 4753
rect 5496 4744 5504 4773
rect 5476 4736 5504 4744
rect 5116 4227 5124 4333
rect 5216 4267 5224 4333
rect 4976 3907 4984 4093
rect 5016 3927 5024 4153
rect 5176 4147 5184 4253
rect 5236 4247 5244 4273
rect 5276 4247 5284 4273
rect 5056 4067 5064 4113
rect 5136 4067 5144 4093
rect 5080 4064 5093 4067
rect 5076 4053 5093 4064
rect 5056 3927 5064 3993
rect 5076 3967 5084 4053
rect 4796 3707 4804 3813
rect 4796 3487 4804 3693
rect 4836 3567 4844 3713
rect 4896 3647 4904 3873
rect 4956 3847 4964 3873
rect 5016 3847 5024 3913
rect 5007 3836 5024 3847
rect 5007 3833 5020 3836
rect 4936 3727 4944 3773
rect 4896 3507 4904 3553
rect 4796 3464 4804 3473
rect 4796 3456 4833 3464
rect 4636 3407 4644 3433
rect 4676 3367 4684 3433
rect 4876 3427 4884 3453
rect 4540 3304 4553 3307
rect 4536 3293 4553 3304
rect 4536 3267 4544 3293
rect 4356 2787 4364 2893
rect 4336 2424 4344 2713
rect 4376 2547 4384 3173
rect 4396 2867 4404 3093
rect 4436 3027 4444 3073
rect 4456 2967 4464 3053
rect 4556 3027 4564 3233
rect 4576 3044 4584 3173
rect 4596 3127 4604 3333
rect 4696 3307 4704 3333
rect 4756 3247 4764 3333
rect 4647 3236 4673 3244
rect 4636 3144 4644 3212
rect 4696 3147 4704 3193
rect 4636 3140 4664 3144
rect 4636 3136 4667 3140
rect 4653 3127 4667 3136
rect 4607 3116 4624 3124
rect 4576 3040 4604 3044
rect 4576 3036 4607 3040
rect 4593 3027 4607 3036
rect 4487 3016 4513 3024
rect 4576 2927 4584 2953
rect 4536 2887 4544 2913
rect 4396 2524 4404 2613
rect 4376 2520 4404 2524
rect 4373 2516 4404 2520
rect 4373 2507 4387 2516
rect 4416 2507 4424 2533
rect 4316 2416 4344 2424
rect 4256 2267 4264 2373
rect 4196 2147 4204 2193
rect 4236 2127 4244 2193
rect 4176 1867 4184 1913
rect 4113 1744 4127 1753
rect 4113 1740 4144 1744
rect 4116 1736 4144 1740
rect 4096 1667 4104 1693
rect 4136 1627 4144 1736
rect 4036 1404 4044 1613
rect 4156 1547 4164 1593
rect 4176 1567 4184 1693
rect 4196 1544 4204 2033
rect 4216 1827 4224 1893
rect 4256 1627 4264 2013
rect 4296 1907 4304 2373
rect 4316 2147 4324 2416
rect 4336 2347 4344 2393
rect 4416 2347 4424 2433
rect 4436 2344 4444 2673
rect 4456 2364 4464 2833
rect 4496 2784 4504 2873
rect 4556 2804 4564 2893
rect 4596 2867 4604 2893
rect 4536 2800 4564 2804
rect 4476 2776 4504 2784
rect 4533 2796 4564 2800
rect 4533 2787 4547 2796
rect 4476 2747 4484 2776
rect 4476 2736 4493 2747
rect 4480 2733 4493 2736
rect 4476 2407 4484 2613
rect 4496 2547 4504 2733
rect 4536 2687 4544 2773
rect 4496 2487 4504 2533
rect 4456 2356 4484 2364
rect 4436 2336 4464 2344
rect 4336 2207 4344 2293
rect 4376 2207 4384 2333
rect 4356 2087 4364 2153
rect 4416 2027 4424 2253
rect 4436 2067 4444 2313
rect 4456 2067 4464 2336
rect 4476 2184 4484 2356
rect 4516 2307 4524 2633
rect 4556 2587 4564 2653
rect 4536 2367 4544 2433
rect 4576 2284 4584 2813
rect 4616 2647 4624 3116
rect 4636 2827 4644 2953
rect 4696 2867 4704 3133
rect 4716 3087 4724 3233
rect 4756 3027 4764 3233
rect 4796 3187 4804 3373
rect 4816 3207 4824 3393
rect 4796 3027 4804 3173
rect 4836 3047 4844 3353
rect 4876 3167 4884 3293
rect 4916 3107 4924 3473
rect 4936 3367 4944 3633
rect 4996 3547 5004 3613
rect 5036 3587 5044 3873
rect 5076 3827 5084 3953
rect 5156 3947 5164 3993
rect 5096 3767 5104 3933
rect 5196 3867 5204 4093
rect 5236 3907 5244 4053
rect 5256 3927 5264 4093
rect 5276 3947 5284 3993
rect 5316 3928 5324 4193
rect 5376 4087 5384 4173
rect 5356 3967 5364 3993
rect 5136 3727 5144 3753
rect 5096 3548 5104 3633
rect 4956 3387 4964 3513
rect 4976 3367 4984 3493
rect 4996 3407 5004 3533
rect 4940 3304 4953 3307
rect 4936 3293 4953 3304
rect 4936 3147 4944 3293
rect 5036 3287 5044 3413
rect 4976 3187 4984 3233
rect 5016 3167 5024 3233
rect 4936 3027 4944 3073
rect 5016 3067 5024 3153
rect 5036 3107 5044 3173
rect 5056 3147 5064 3393
rect 5096 3388 5104 3512
rect 5156 3447 5164 3473
rect 5176 3427 5184 3793
rect 5196 3387 5204 3813
rect 5256 3767 5264 3873
rect 5276 3784 5284 3853
rect 5316 3827 5324 3892
rect 5276 3780 5304 3784
rect 5276 3776 5307 3780
rect 5293 3767 5307 3776
rect 5296 3727 5304 3753
rect 5336 3707 5344 3753
rect 5276 3487 5284 3673
rect 5336 3547 5344 3573
rect 5316 3447 5324 3473
rect 5096 3307 5104 3352
rect 5136 3307 5144 3333
rect 5076 3087 5084 3273
rect 5096 3247 5104 3293
rect 5156 3247 5164 3373
rect 5376 3367 5384 3533
rect 5296 3307 5304 3353
rect 5096 3236 5113 3247
rect 5100 3233 5113 3236
rect 5076 3027 5084 3073
rect 4747 3016 4764 3027
rect 4747 3013 4760 3016
rect 4787 3016 4804 3027
rect 4860 3024 4873 3027
rect 4787 3013 4800 3016
rect 4856 3013 4873 3024
rect 4927 3016 4944 3027
rect 4996 3020 5033 3024
rect 4993 3016 5033 3020
rect 4927 3013 4940 3016
rect 4856 2987 4864 3013
rect 4993 3007 5007 3016
rect 4916 2996 4953 3004
rect 4756 2980 4844 2984
rect 4753 2976 4844 2980
rect 4753 2967 4767 2976
rect 4676 2787 4684 2813
rect 4667 2773 4684 2787
rect 4596 2327 4604 2593
rect 4636 2587 4644 2733
rect 4676 2667 4684 2773
rect 4696 2627 4704 2753
rect 4736 2627 4744 2913
rect 4756 2767 4764 2913
rect 4796 2867 4804 2953
rect 4836 2947 4844 2976
rect 4880 2964 4893 2967
rect 4876 2960 4893 2964
rect 4873 2953 4893 2960
rect 4916 2964 4924 2996
rect 4907 2956 4924 2964
rect 4873 2947 4887 2953
rect 4816 2867 4824 2893
rect 4876 2867 4884 2893
rect 4996 2847 5004 2933
rect 5056 2887 5064 2953
rect 5076 2867 5084 2893
rect 5116 2887 5124 3193
rect 5156 2847 5164 3153
rect 5196 3067 5204 3293
rect 5236 3260 5304 3264
rect 5233 3256 5304 3260
rect 5233 3247 5247 3256
rect 5296 3247 5304 3256
rect 5296 3236 5313 3247
rect 5300 3233 5313 3236
rect 5276 3207 5284 3233
rect 5196 3027 5204 3053
rect 5256 3027 5264 3173
rect 5396 3168 5404 3913
rect 5416 3827 5424 3933
rect 5436 3804 5444 4673
rect 5476 4664 5484 4736
rect 5456 4660 5484 4664
rect 5453 4656 5484 4660
rect 5453 4647 5467 4656
rect 5536 4647 5544 5033
rect 5556 4787 5564 5076
rect 5616 4967 5624 5113
rect 5636 5027 5644 5133
rect 5656 5087 5664 5112
rect 5696 5104 5704 5213
rect 5716 5127 5724 5253
rect 5776 5227 5784 5313
rect 5816 5287 5824 5313
rect 5916 5227 5924 5333
rect 5956 5288 5964 5313
rect 5996 5307 6004 5333
rect 5676 5096 5704 5104
rect 5676 5027 5684 5096
rect 5756 5027 5764 5113
rect 5796 5087 5804 5113
rect 5787 5076 5804 5087
rect 5787 5073 5800 5076
rect 5876 5027 5884 5213
rect 5916 5107 5924 5153
rect 5956 5107 5964 5252
rect 6036 5107 6044 5492
rect 6076 5267 6084 5453
rect 6096 5327 6104 5473
rect 6136 5387 6144 5513
rect 6156 5327 6164 5413
rect 6176 5407 6184 5553
rect 6096 5316 6113 5327
rect 6100 5313 6113 5316
rect 6156 5188 6164 5313
rect 6027 5036 6053 5044
rect 5676 4987 5684 5013
rect 5716 4927 5724 4973
rect 5576 4727 5584 4873
rect 5616 4747 5624 4873
rect 5656 4867 5664 4913
rect 5707 4824 5720 4827
rect 5707 4813 5724 4824
rect 5716 4807 5724 4813
rect 5736 4807 5744 4893
rect 5776 4867 5784 4913
rect 5767 4856 5784 4867
rect 5767 4853 5780 4856
rect 5716 4796 5733 4807
rect 5720 4793 5733 4796
rect 5760 4804 5773 4807
rect 5756 4793 5773 4804
rect 5756 4784 5764 4793
rect 5707 4776 5764 4784
rect 5676 4587 5684 4733
rect 5716 4667 5724 4733
rect 5716 4587 5724 4653
rect 5516 4387 5524 4573
rect 5553 4564 5567 4573
rect 5553 4560 5584 4564
rect 5556 4556 5584 4560
rect 5536 4487 5544 4513
rect 5576 4467 5584 4556
rect 5736 4527 5744 4633
rect 5656 4407 5664 4513
rect 5556 4347 5564 4373
rect 5456 4127 5464 4193
rect 5476 4007 5484 4273
rect 5496 4207 5504 4333
rect 5547 4284 5560 4287
rect 5547 4273 5564 4284
rect 5556 4227 5564 4273
rect 5576 4207 5584 4273
rect 5496 4067 5504 4113
rect 5536 4067 5544 4193
rect 5476 3904 5484 3993
rect 5556 3987 5564 4173
rect 5636 4127 5644 4333
rect 5696 4287 5704 4493
rect 5756 4387 5764 4453
rect 5796 4427 5804 5013
rect 6076 5007 6084 5093
rect 5856 4807 5864 4893
rect 5876 4867 5884 4893
rect 5896 4807 5904 4973
rect 5916 4707 5924 4853
rect 5976 4667 5984 4993
rect 6116 4987 6124 5033
rect 6056 4807 6064 4933
rect 6096 4807 6104 4953
rect 6127 4864 6140 4867
rect 6127 4853 6144 4864
rect 5756 4347 5764 4373
rect 5747 4336 5764 4347
rect 5747 4333 5760 4336
rect 5776 4287 5784 4333
rect 5696 4273 5713 4287
rect 5767 4276 5784 4287
rect 5767 4273 5780 4276
rect 5696 4207 5704 4273
rect 5756 4227 5764 4273
rect 5616 3967 5624 3993
rect 5476 3896 5504 3904
rect 5416 3796 5444 3804
rect 5416 3387 5424 3796
rect 5476 3767 5484 3853
rect 5436 3727 5444 3753
rect 5476 3707 5484 3753
rect 5496 3587 5504 3896
rect 5556 3687 5564 3933
rect 5576 3767 5584 3953
rect 5636 3904 5644 4053
rect 5656 3947 5664 3993
rect 5627 3896 5644 3904
rect 5616 3827 5624 3893
rect 5636 3767 5644 3872
rect 5656 3867 5664 3933
rect 5676 3767 5684 4053
rect 5716 3924 5724 3953
rect 5696 3916 5724 3924
rect 5696 3807 5704 3916
rect 5736 3904 5744 4193
rect 5796 4067 5804 4373
rect 5836 4147 5844 4653
rect 6056 4647 6064 4793
rect 6136 4787 6144 4853
rect 6136 4747 6144 4773
rect 6156 4687 6164 5152
rect 6180 5104 6193 5107
rect 6176 5093 6193 5104
rect 6176 4827 6184 5093
rect 6216 5084 6224 5653
rect 6256 5644 6264 5813
rect 6236 5636 6264 5644
rect 6236 5207 6244 5636
rect 6276 5567 6284 5913
rect 6376 5707 6384 6353
rect 6396 6144 6404 6353
rect 6396 6136 6424 6144
rect 6416 5707 6424 6136
rect 6456 5667 6464 6413
rect 6476 5827 6484 6453
rect 6516 5787 6524 6073
rect 6256 5167 6264 5453
rect 6316 5448 6324 5553
rect 6336 5487 6344 5613
rect 6236 5107 6244 5133
rect 6196 5076 6224 5084
rect 6196 4744 6204 5076
rect 6256 4887 6264 4953
rect 6276 4927 6284 5433
rect 6316 5387 6324 5412
rect 6307 5376 6324 5387
rect 6307 5373 6320 5376
rect 6316 5267 6324 5313
rect 6296 4944 6304 5213
rect 6316 4967 6324 5033
rect 6356 5027 6364 5653
rect 6393 5627 6407 5633
rect 6393 5620 6413 5627
rect 6396 5616 6413 5620
rect 6400 5613 6413 5616
rect 6376 5427 6384 5593
rect 6376 5187 6384 5413
rect 6396 5287 6404 5513
rect 6456 5467 6464 5613
rect 6516 5607 6524 5713
rect 6436 5387 6444 5413
rect 6516 5407 6524 5493
rect 6416 5207 6424 5313
rect 6456 5287 6464 5313
rect 6476 5227 6484 5373
rect 6296 4936 6324 4944
rect 6267 4884 6280 4887
rect 6267 4873 6284 4884
rect 6216 4787 6224 4873
rect 6276 4827 6284 4873
rect 6196 4736 6224 4744
rect 6113 4587 6127 4593
rect 6136 4587 6144 4613
rect 5960 4584 5973 4587
rect 5956 4573 5973 4584
rect 6113 4580 6133 4587
rect 6116 4576 6133 4580
rect 6120 4573 6133 4576
rect 6187 4584 6200 4587
rect 6187 4573 6204 4584
rect 5896 4347 5904 4573
rect 5956 4527 5964 4573
rect 5956 4487 5964 4513
rect 5996 4467 6004 4493
rect 5987 4336 6013 4344
rect 5936 4284 5944 4333
rect 6036 4287 6044 4513
rect 6116 4487 6124 4513
rect 5936 4276 5993 4284
rect 6073 4284 6087 4293
rect 6047 4280 6087 4284
rect 6047 4276 6084 4280
rect 5876 4227 5884 4253
rect 5916 4207 5924 4273
rect 5856 4084 5864 4113
rect 5836 4080 5864 4084
rect 5833 4076 5864 4080
rect 5833 4067 5847 4076
rect 5956 4067 5964 4093
rect 6116 4067 6124 4133
rect 6156 4128 6164 4513
rect 6196 4504 6204 4573
rect 6176 4496 6204 4504
rect 6176 4227 6184 4496
rect 6196 4167 6204 4353
rect 6156 4067 6164 4092
rect 5860 4064 5873 4067
rect 5856 4053 5873 4064
rect 5980 4064 5993 4067
rect 5976 4053 5993 4064
rect 5856 4044 5864 4053
rect 5776 4036 5864 4044
rect 5913 4044 5927 4053
rect 5976 4044 5984 4053
rect 5913 4040 5984 4044
rect 5916 4036 5984 4040
rect 5776 4007 5784 4036
rect 5856 3967 5864 3993
rect 5756 3907 5764 3933
rect 5716 3896 5744 3904
rect 5576 3756 5593 3767
rect 5580 3753 5593 3756
rect 5553 3547 5567 3553
rect 5656 3547 5664 3673
rect 5716 3607 5724 3896
rect 5736 3816 5773 3824
rect 5736 3727 5744 3816
rect 5796 3767 5804 3933
rect 5756 3707 5764 3753
rect 5816 3687 5824 3873
rect 5936 3827 5944 3933
rect 6016 3867 6024 3973
rect 6056 3887 6064 3993
rect 6216 3967 6224 4736
rect 6316 4647 6324 4936
rect 6376 4767 6384 4873
rect 5480 3544 5493 3547
rect 5476 3533 5493 3544
rect 5547 3540 5567 3547
rect 5547 3536 5564 3540
rect 5547 3533 5560 3536
rect 5707 3544 5720 3547
rect 5707 3533 5724 3544
rect 5476 3487 5484 3533
rect 5496 3524 5504 3533
rect 5496 3516 5573 3524
rect 5613 3504 5627 3513
rect 5716 3508 5724 3533
rect 5613 3500 5644 3504
rect 5616 3496 5647 3500
rect 5633 3487 5647 3496
rect 5756 3507 5764 3613
rect 5836 3587 5844 3653
rect 5856 3547 5864 3813
rect 5916 3727 5924 3753
rect 5956 3707 5964 3753
rect 5896 3607 5904 3673
rect 5516 3427 5524 3453
rect 5556 3447 5564 3473
rect 5427 3296 5453 3304
rect 5416 3187 5424 3293
rect 5376 3027 5384 3053
rect 5196 3016 5213 3027
rect 5200 3013 5213 3016
rect 5207 2956 5264 2964
rect 4796 2787 4804 2813
rect 4916 2767 4924 2833
rect 4956 2787 4964 2813
rect 5136 2727 5144 2813
rect 5136 2716 5153 2727
rect 5140 2713 5153 2716
rect 4776 2607 4784 2713
rect 4816 2587 4824 2713
rect 4936 2667 4944 2713
rect 4973 2704 4987 2713
rect 4956 2700 4987 2704
rect 4956 2696 4984 2700
rect 4616 2444 4624 2553
rect 4636 2487 4644 2533
rect 4716 2507 4724 2533
rect 4876 2507 4884 2613
rect 4900 2524 4913 2527
rect 4896 2513 4913 2524
rect 4687 2504 4700 2507
rect 4687 2493 4704 2504
rect 4696 2484 4704 2493
rect 4696 2476 4724 2484
rect 4616 2436 4653 2444
rect 4716 2407 4724 2476
rect 4576 2276 4604 2284
rect 4476 2176 4504 2184
rect 4496 2167 4504 2176
rect 4496 2127 4504 2153
rect 4516 2127 4524 2193
rect 4496 2027 4504 2113
rect 4516 2047 4524 2113
rect 4376 1927 4384 2013
rect 4196 1536 4224 1544
rect 4076 1467 4084 1493
rect 4196 1467 4204 1513
rect 4127 1456 4153 1464
rect 4216 1424 4224 1536
rect 4256 1527 4264 1613
rect 4276 1567 4284 1833
rect 4296 1704 4304 1853
rect 4336 1807 4344 1833
rect 4376 1747 4384 1773
rect 4416 1767 4424 2013
rect 4456 1987 4464 2013
rect 4456 1976 4473 1987
rect 4460 1973 4473 1976
rect 4556 1984 4564 2133
rect 4527 1976 4564 1984
rect 4576 1984 4584 2253
rect 4596 2107 4604 2276
rect 4616 2127 4624 2393
rect 4656 2267 4664 2373
rect 4636 2147 4644 2193
rect 4616 2027 4624 2113
rect 4656 2047 4664 2253
rect 4696 2227 4704 2373
rect 4736 2127 4744 2233
rect 4676 1987 4684 2113
rect 4576 1976 4613 1984
rect 4667 1976 4684 1987
rect 4667 1973 4680 1976
rect 4436 1787 4444 1973
rect 4467 1924 4480 1927
rect 4467 1913 4484 1924
rect 4476 1827 4484 1913
rect 4616 1887 4624 1973
rect 4453 1747 4467 1753
rect 4453 1740 4473 1747
rect 4456 1736 4473 1740
rect 4460 1733 4473 1736
rect 4296 1700 4324 1704
rect 4296 1696 4327 1700
rect 4296 1507 4304 1696
rect 4313 1687 4327 1696
rect 4416 1696 4484 1704
rect 4367 1684 4380 1687
rect 4367 1680 4384 1684
rect 4367 1673 4387 1680
rect 4316 1547 4324 1673
rect 4373 1667 4387 1673
rect 4247 1456 4273 1464
rect 4216 1416 4244 1424
rect 4016 1396 4044 1404
rect 4016 1307 4024 1396
rect 4107 1404 4120 1407
rect 4107 1400 4124 1404
rect 4176 1400 4213 1404
rect 4107 1393 4127 1400
rect 4113 1387 4127 1393
rect 4173 1396 4213 1400
rect 4173 1387 4187 1396
rect 4056 1347 4064 1373
rect 3760 1164 3773 1167
rect 3756 1160 3773 1164
rect 3753 1153 3773 1160
rect 3753 1147 3767 1153
rect 3813 1144 3827 1153
rect 3796 1140 3827 1144
rect 3796 1136 3824 1140
rect 3696 947 3704 993
rect 3747 936 3773 944
rect 3796 887 3804 1136
rect 3836 947 3844 1093
rect 3856 967 3864 1113
rect 3896 1007 3904 1273
rect 3916 1127 3924 1213
rect 3936 1107 3944 1153
rect 3956 1067 3964 1213
rect 3996 1167 4004 1253
rect 4076 1187 4084 1293
rect 4116 1227 4124 1253
rect 3987 1156 4004 1167
rect 3987 1153 4000 1156
rect 4016 1027 4024 1133
rect 4076 1107 4084 1173
rect 3827 936 3844 947
rect 3827 933 3840 936
rect 3936 887 3944 993
rect 4056 987 4064 1073
rect 4096 967 4104 1073
rect 4136 1008 4144 1153
rect 4156 1147 4164 1233
rect 4176 1027 4184 1293
rect 4196 1127 4204 1253
rect 4216 1167 4224 1313
rect 4236 1287 4244 1416
rect 4276 1287 4284 1393
rect 4296 1267 4304 1493
rect 4336 1307 4344 1633
rect 4356 1467 4364 1553
rect 4416 1547 4424 1696
rect 4476 1687 4484 1696
rect 4476 1676 4493 1687
rect 4480 1673 4493 1676
rect 4456 1627 4464 1673
rect 4516 1627 4524 1873
rect 4556 1547 4564 1733
rect 4576 1547 4584 1873
rect 4636 1867 4644 1913
rect 4696 1847 4704 1913
rect 4596 1607 4604 1773
rect 4696 1747 4704 1793
rect 4636 1648 4644 1673
rect 4636 1547 4644 1612
rect 4676 1567 4684 1673
rect 4716 1627 4724 2093
rect 4396 1467 4404 1513
rect 4456 1467 4464 1533
rect 4516 1467 4524 1513
rect 4556 1467 4564 1533
rect 4736 1527 4744 2053
rect 4756 1804 4764 2393
rect 4776 2247 4784 2433
rect 4796 2207 4804 2493
rect 4816 2327 4824 2413
rect 4836 2407 4844 2493
rect 4896 2427 4904 2513
rect 4936 2447 4944 2593
rect 4956 2407 4964 2696
rect 4816 2067 4824 2253
rect 4836 2147 4844 2193
rect 4856 2047 4864 2313
rect 4916 2147 4924 2393
rect 4976 2367 4984 2553
rect 5096 2528 5104 2673
rect 5116 2647 5124 2713
rect 5156 2687 5164 2713
rect 5196 2567 5204 2873
rect 5216 2587 5224 2833
rect 5236 2587 5244 2933
rect 5256 2887 5264 2956
rect 5356 2907 5364 2953
rect 5256 2787 5264 2873
rect 5276 2687 5284 2733
rect 4993 2507 5007 2513
rect 5176 2507 5184 2533
rect 4993 2500 5013 2507
rect 4996 2496 5013 2500
rect 5000 2493 5013 2496
rect 5067 2496 5093 2504
rect 5133 2484 5147 2493
rect 5213 2484 5227 2493
rect 5133 2480 5227 2484
rect 5136 2476 5224 2480
rect 4996 2327 5004 2433
rect 4936 2207 4944 2293
rect 4996 2267 5004 2313
rect 5036 2267 5044 2393
rect 5096 2327 5104 2413
rect 5116 2347 5124 2393
rect 5156 2267 5164 2353
rect 5256 2327 5264 2653
rect 5316 2647 5324 2773
rect 5316 2607 5324 2633
rect 5396 2627 5404 3132
rect 5436 3027 5444 3233
rect 5427 3013 5444 3027
rect 5416 2727 5424 2913
rect 5436 2887 5444 3013
rect 5456 2827 5464 3153
rect 5476 2927 5484 3233
rect 5576 3187 5584 3293
rect 5616 3267 5624 3393
rect 5636 3307 5644 3353
rect 5536 3027 5544 3053
rect 5516 2907 5524 2953
rect 5496 2896 5513 2904
rect 5436 2787 5444 2813
rect 5476 2804 5484 2873
rect 5456 2796 5484 2804
rect 5456 2787 5464 2796
rect 5436 2776 5453 2787
rect 5440 2773 5453 2776
rect 5496 2744 5504 2896
rect 5576 2887 5584 3013
rect 5476 2740 5504 2744
rect 5473 2736 5504 2740
rect 5473 2727 5487 2736
rect 5416 2716 5433 2727
rect 5420 2713 5433 2716
rect 5296 2367 5304 2413
rect 5316 2347 5324 2493
rect 5356 2407 5364 2493
rect 4976 2167 4984 2193
rect 5096 2147 5104 2193
rect 4776 1827 4784 2033
rect 4796 1996 4853 2004
rect 4796 1947 4804 1996
rect 4836 1887 4844 1913
rect 4876 1847 4884 1973
rect 4916 1967 4924 2133
rect 5136 2127 5144 2193
rect 4936 2007 4944 2093
rect 4956 1987 4964 2033
rect 4976 1967 4984 2113
rect 5016 2087 5024 2113
rect 5080 2064 5094 2067
rect 5076 2053 5094 2064
rect 5076 2007 5084 2053
rect 5176 2027 5184 2313
rect 5196 2267 5204 2293
rect 5196 2067 5204 2153
rect 5116 1987 5124 2013
rect 5216 1987 5224 2313
rect 5333 2304 5347 2313
rect 5316 2300 5347 2304
rect 5316 2296 5344 2300
rect 5236 2067 5244 2293
rect 5316 2224 5324 2296
rect 5356 2267 5364 2393
rect 5376 2307 5384 2573
rect 5356 2256 5373 2267
rect 5360 2253 5373 2256
rect 5296 2220 5324 2224
rect 5293 2216 5324 2220
rect 5293 2207 5307 2216
rect 5256 2107 5264 2193
rect 5336 2187 5344 2253
rect 5416 2224 5424 2593
rect 5436 2504 5444 2613
rect 5436 2500 5464 2504
rect 5436 2496 5467 2500
rect 5436 2387 5444 2496
rect 5453 2487 5467 2496
rect 5516 2487 5524 2533
rect 5496 2407 5504 2433
rect 5436 2327 5444 2373
rect 5416 2220 5444 2224
rect 5416 2216 5447 2220
rect 5433 2207 5447 2216
rect 5380 2204 5393 2207
rect 5376 2200 5393 2204
rect 5373 2193 5393 2200
rect 5373 2187 5387 2193
rect 5296 1987 5304 2013
rect 4976 1956 4993 1967
rect 4980 1953 4993 1956
rect 5120 1924 5133 1927
rect 5116 1913 5133 1924
rect 5116 1904 5124 1913
rect 5096 1896 5124 1904
rect 4936 1867 4944 1893
rect 4976 1847 4984 1893
rect 5096 1867 5104 1896
rect 5156 1887 5164 1973
rect 4836 1807 4844 1833
rect 5016 1807 5024 1833
rect 5196 1807 5204 1913
rect 4756 1796 4784 1804
rect 4756 1647 4764 1773
rect 4756 1467 4764 1493
rect 4447 1456 4464 1467
rect 4447 1453 4460 1456
rect 4700 1464 4713 1467
rect 4696 1453 4713 1464
rect 4376 1307 4384 1373
rect 4416 1347 4424 1393
rect 4533 1384 4547 1393
rect 4516 1380 4547 1384
rect 4516 1376 4544 1380
rect 4516 1347 4524 1376
rect 4596 1367 4604 1433
rect 4236 1204 4244 1233
rect 4256 1227 4264 1253
rect 4436 1247 4444 1313
rect 4476 1247 4484 1333
rect 4576 1227 4584 1333
rect 4333 1213 4334 1220
rect 4407 1216 4513 1224
rect 4576 1216 4593 1227
rect 4580 1213 4593 1216
rect 4333 1204 4347 1213
rect 4236 1200 4347 1204
rect 4236 1196 4344 1200
rect 4387 1176 4413 1184
rect 4216 1156 4233 1167
rect 4220 1153 4233 1156
rect 4276 1107 4284 1153
rect 4316 1127 4324 1173
rect 4136 947 4144 972
rect 4176 947 4184 1013
rect 4236 1007 4244 1093
rect 4256 947 4264 973
rect 4296 947 4304 1013
rect 4336 947 4344 1033
rect 3676 847 3684 873
rect 3796 847 3804 873
rect 3776 747 3784 773
rect 3626 696 3693 704
rect 3716 647 3724 733
rect 3776 647 3784 733
rect 3793 707 3807 713
rect 3793 700 3813 707
rect 3796 696 3813 700
rect 3800 693 3813 696
rect 3776 636 3793 647
rect 3780 633 3793 636
rect 3676 567 3684 633
rect 3576 436 3604 444
rect 3436 127 3444 213
rect 3476 187 3484 233
rect 3436 116 3453 127
rect 3440 113 3453 116
rect 3496 87 3504 113
rect 3536 27 3544 173
rect 3576 27 3584 436
rect 3636 427 3644 553
rect 3596 287 3604 413
rect 3716 367 3724 473
rect 3756 427 3764 593
rect 3796 427 3804 573
rect 3836 567 3844 633
rect 3876 547 3884 693
rect 3876 388 3884 533
rect 3916 507 3924 733
rect 3936 647 3944 773
rect 3976 747 3984 913
rect 4376 907 4384 1113
rect 4396 987 4404 1053
rect 4456 1047 4464 1153
rect 4496 1147 4504 1173
rect 4476 947 4484 993
rect 4407 936 4433 944
rect 4116 787 4124 853
rect 4156 847 4164 873
rect 4276 847 4284 873
rect 3953 707 3967 713
rect 3953 700 3973 707
rect 3956 696 3973 700
rect 3960 693 3973 696
rect 3936 636 3953 647
rect 3940 633 3953 636
rect 3996 587 4004 633
rect 4036 507 4044 693
rect 4076 507 4084 733
rect 4100 704 4113 707
rect 4096 693 4113 704
rect 4026 493 4044 507
rect 3956 444 3964 493
rect 3936 440 3964 444
rect 3933 436 3964 440
rect 3933 427 3947 436
rect 3987 424 4000 427
rect 4036 424 4044 493
rect 4096 487 4104 693
rect 4196 647 4204 693
rect 4187 636 4204 647
rect 4276 647 4284 773
rect 4336 747 4344 873
rect 4356 807 4364 833
rect 4336 647 4344 733
rect 4356 707 4364 793
rect 4276 636 4293 647
rect 4187 633 4200 636
rect 4280 633 4293 636
rect 4136 607 4144 633
rect 4176 567 4184 633
rect 4136 467 4144 493
rect 4196 487 4204 533
rect 4396 487 4404 873
rect 4416 767 4424 893
rect 4556 887 4564 1033
rect 4636 947 4644 973
rect 4556 884 4573 887
rect 4536 876 4573 884
rect 4516 707 4524 753
rect 4536 664 4544 876
rect 4560 873 4573 876
rect 4516 656 4544 664
rect 4516 647 4524 656
rect 4556 647 4564 813
rect 4576 704 4584 873
rect 4596 747 4604 933
rect 4676 927 4684 1433
rect 4696 1407 4704 1453
rect 4696 1347 4704 1393
rect 4716 1247 4724 1353
rect 4736 1287 4744 1373
rect 4776 1367 4784 1796
rect 4796 1747 4804 1793
rect 4976 1747 4984 1773
rect 4816 1567 4824 1673
rect 4856 1607 4864 1673
rect 4956 1647 4964 1673
rect 4996 1627 5004 1673
rect 4796 1307 4804 1493
rect 4816 1327 4824 1393
rect 4876 1347 4884 1453
rect 4896 1367 4904 1393
rect 4916 1347 4924 1453
rect 4700 1244 4713 1247
rect 4696 1233 4713 1244
rect 4696 1167 4704 1233
rect 4756 1107 4764 1233
rect 4767 1096 4784 1104
rect 4776 1047 4784 1096
rect 4716 887 4724 973
rect 4736 947 4744 993
rect 4776 947 4784 993
rect 4740 884 4753 887
rect 4736 880 4753 884
rect 4733 873 4753 880
rect 4733 867 4747 873
rect 4656 767 4664 853
rect 4676 787 4684 813
rect 4576 696 4613 704
rect 4636 647 4644 733
rect 4507 636 4524 647
rect 4507 633 4520 636
rect 4547 636 4564 647
rect 4547 633 4560 636
rect 4536 607 4544 633
rect 4676 607 4684 633
rect 4676 524 4684 553
rect 4716 547 4724 813
rect 4776 647 4784 793
rect 4796 707 4804 773
rect 4816 767 4824 1173
rect 4856 1167 4864 1313
rect 4876 1227 4884 1333
rect 4916 1184 4924 1273
rect 4956 1267 4964 1593
rect 5016 1447 5024 1733
rect 5056 1647 5064 1773
rect 5036 1467 5044 1553
rect 5096 1467 5104 1773
rect 5136 1747 5144 1793
rect 5116 1647 5124 1673
rect 5136 1567 5144 1633
rect 5156 1627 5164 1673
rect 5176 1647 5184 1733
rect 5196 1567 5204 1613
rect 5036 1456 5053 1467
rect 5040 1453 5053 1456
rect 4976 1367 4984 1433
rect 4976 1287 4984 1353
rect 4996 1227 5004 1273
rect 5016 1227 5024 1333
rect 5036 1307 5044 1393
rect 5096 1327 5104 1453
rect 5136 1267 5144 1553
rect 5216 1547 5224 1933
rect 5276 1887 5284 1913
rect 5236 1567 5244 1873
rect 5156 1407 5164 1493
rect 5176 1404 5184 1513
rect 5196 1467 5204 1493
rect 5216 1467 5224 1533
rect 5256 1507 5264 1853
rect 5316 1687 5324 1833
rect 5376 1827 5384 2093
rect 5436 2087 5444 2133
rect 5416 1987 5424 2053
rect 5456 2027 5464 2353
rect 5536 2267 5544 2393
rect 5496 2147 5504 2253
rect 5536 2168 5544 2253
rect 5467 2016 5484 2024
rect 5356 1687 5364 1793
rect 5416 1684 5424 1913
rect 5456 1887 5464 1973
rect 5456 1707 5464 1833
rect 5476 1787 5484 2016
rect 5516 1927 5524 2073
rect 5496 1747 5504 1793
rect 5536 1747 5544 2132
rect 5556 2067 5564 2773
rect 5576 2587 5584 2833
rect 5596 2787 5604 2853
rect 5636 2847 5644 3293
rect 5676 3267 5684 3413
rect 5656 2967 5664 3193
rect 5676 3027 5684 3153
rect 5716 3067 5724 3472
rect 5736 3207 5744 3333
rect 5776 3307 5784 3333
rect 5816 3247 5824 3473
rect 5876 3447 5884 3473
rect 5896 3408 5904 3533
rect 5807 3236 5824 3247
rect 5807 3233 5820 3236
rect 5756 3187 5764 3233
rect 5896 3184 5904 3372
rect 5936 3284 5944 3613
rect 5996 3587 6004 3813
rect 6016 3627 6024 3693
rect 6076 3667 6084 3753
rect 6016 3547 6024 3613
rect 6076 3587 6084 3653
rect 6016 3536 6033 3547
rect 6020 3533 6033 3536
rect 5996 3407 6004 3533
rect 6096 3487 6104 3813
rect 6116 3767 6124 3893
rect 6016 3447 6024 3473
rect 5956 3327 5964 3353
rect 6096 3347 6104 3473
rect 6116 3447 6124 3753
rect 6136 3424 6144 3953
rect 6236 3884 6244 4633
rect 6296 4567 6304 4613
rect 6416 4567 6424 4873
rect 6456 4864 6464 5193
rect 6436 4856 6464 4864
rect 6296 4287 6304 4393
rect 6316 4387 6324 4513
rect 6356 4407 6364 4553
rect 6436 4387 6444 4856
rect 6316 4347 6324 4373
rect 6316 4067 6324 4233
rect 6356 4227 6364 4293
rect 6316 4053 6333 4067
rect 6260 4004 6273 4007
rect 6216 3876 6244 3884
rect 6256 3993 6273 4004
rect 6216 3627 6224 3876
rect 6256 3867 6264 3993
rect 6256 3828 6264 3853
rect 6276 3767 6284 3853
rect 6296 3827 6304 4053
rect 6316 3867 6324 4053
rect 6376 3967 6384 4373
rect 6476 4347 6484 5173
rect 6396 3887 6404 4333
rect 6276 3756 6293 3767
rect 6280 3753 6293 3756
rect 6216 3547 6224 3573
rect 6160 3544 6173 3547
rect 6156 3533 6173 3544
rect 6156 3487 6164 3533
rect 6196 3447 6204 3473
rect 6116 3416 6144 3424
rect 6013 3327 6027 3333
rect 6007 3320 6027 3327
rect 6007 3316 6024 3320
rect 6007 3313 6020 3316
rect 6080 3304 6093 3307
rect 6076 3293 6093 3304
rect 5936 3276 5964 3284
rect 5956 3264 5964 3276
rect 5956 3256 6013 3264
rect 5936 3207 5944 3253
rect 6076 3227 6084 3293
rect 6116 3247 6124 3416
rect 6176 3307 6184 3353
rect 5896 3176 5924 3184
rect 5727 3024 5740 3027
rect 5727 3013 5744 3024
rect 5696 2927 5704 2953
rect 5736 2887 5744 3013
rect 5687 2776 5713 2784
rect 5616 2567 5624 2713
rect 5656 2667 5664 2713
rect 5636 2547 5644 2633
rect 5636 2487 5644 2533
rect 5616 2367 5624 2413
rect 5656 2347 5664 2413
rect 5716 2407 5724 2633
rect 5776 2607 5784 3113
rect 5816 3107 5824 3153
rect 5876 3067 5884 3113
rect 5876 3027 5884 3053
rect 5820 3024 5833 3027
rect 5816 3013 5833 3024
rect 5816 2967 5824 3013
rect 5836 2984 5844 3013
rect 5836 2976 5884 2984
rect 5856 2927 5864 2953
rect 5876 2944 5884 2976
rect 5916 2967 5924 3176
rect 5996 3067 6004 3153
rect 6016 3027 6024 3073
rect 6036 3027 6044 3113
rect 6076 3087 6084 3213
rect 6116 3184 6124 3233
rect 6156 3207 6164 3233
rect 6116 3176 6144 3184
rect 6036 3016 6053 3027
rect 6040 3013 6053 3016
rect 5876 2936 5933 2944
rect 5836 2787 5844 2833
rect 5876 2767 5884 2893
rect 5976 2887 5984 2953
rect 6036 2927 6044 2953
rect 5976 2787 5984 2833
rect 5876 2727 5884 2753
rect 5867 2716 5884 2727
rect 5936 2727 5944 2753
rect 5996 2727 6004 2853
rect 5936 2716 5953 2727
rect 5867 2713 5880 2716
rect 5940 2713 5953 2716
rect 5816 2687 5824 2713
rect 5733 2504 5747 2513
rect 5796 2507 5804 2533
rect 5856 2507 5864 2653
rect 5956 2627 5964 2713
rect 5996 2687 6004 2713
rect 5733 2500 5773 2504
rect 5736 2496 5773 2500
rect 5796 2496 5813 2507
rect 5800 2493 5813 2496
rect 5780 2444 5793 2447
rect 5776 2433 5793 2444
rect 5776 2407 5784 2433
rect 5856 2387 5864 2493
rect 5916 2447 5924 2533
rect 5976 2447 5984 2593
rect 6036 2547 6044 2773
rect 6096 2607 6104 3113
rect 6136 3104 6144 3176
rect 6116 3096 6144 3104
rect 6116 2967 6124 3096
rect 6216 3088 6224 3413
rect 6236 3127 6244 3573
rect 6276 3427 6284 3613
rect 6316 3547 6324 3814
rect 6436 3787 6444 3993
rect 6496 3964 6504 4913
rect 6476 3956 6504 3964
rect 6307 3476 6333 3484
rect 6216 3027 6224 3052
rect 6256 3027 6264 3333
rect 6276 3244 6284 3353
rect 6296 3347 6304 3473
rect 6336 3307 6344 3413
rect 6276 3236 6313 3244
rect 6356 3167 6364 3233
rect 6116 2724 6124 2953
rect 6136 2787 6144 2893
rect 6176 2807 6184 2893
rect 6196 2848 6204 2933
rect 6236 2927 6244 2953
rect 6276 2927 6284 2953
rect 6196 2727 6204 2812
rect 6116 2716 6153 2724
rect 6076 2507 6084 2573
rect 5596 2107 5604 2333
rect 5616 2087 5624 2253
rect 5676 2207 5684 2293
rect 5716 2207 5724 2313
rect 5756 2267 5764 2313
rect 5747 2256 5764 2267
rect 5747 2253 5760 2256
rect 5616 1987 5624 2073
rect 5576 1827 5584 1973
rect 5656 1927 5664 2013
rect 5596 1867 5604 1913
rect 5573 1764 5587 1773
rect 5573 1760 5613 1764
rect 5576 1756 5613 1760
rect 5396 1676 5424 1684
rect 5396 1627 5404 1676
rect 5216 1456 5233 1467
rect 5220 1453 5233 1456
rect 5316 1427 5324 1553
rect 5356 1467 5364 1513
rect 5416 1467 5424 1533
rect 5407 1456 5424 1467
rect 5407 1453 5420 1456
rect 5176 1396 5213 1404
rect 5156 1367 5164 1393
rect 5016 1216 5033 1227
rect 5020 1213 5033 1216
rect 4916 1176 4944 1184
rect 4896 1127 4904 1153
rect 4936 1007 4944 1176
rect 5076 1167 5084 1253
rect 5176 1227 5184 1293
rect 5067 1156 5084 1167
rect 5067 1153 5080 1156
rect 5016 1127 5024 1153
rect 5096 1027 5104 1213
rect 5236 1167 5244 1333
rect 5296 1327 5304 1393
rect 5167 1156 5193 1164
rect 5316 1127 5324 1373
rect 5356 1267 5364 1373
rect 5376 1367 5384 1393
rect 5496 1287 5504 1393
rect 5516 1367 5524 1673
rect 5536 1527 5544 1593
rect 5536 1467 5544 1513
rect 5576 1467 5584 1693
rect 5656 1627 5664 1753
rect 5696 1507 5704 2113
rect 5716 1547 5724 2053
rect 5736 1987 5744 2073
rect 5796 2067 5804 2373
rect 5836 2287 5844 2353
rect 5896 2327 5904 2433
rect 6036 2367 6044 2493
rect 5876 2267 5884 2293
rect 6036 2267 6044 2313
rect 5840 2204 5853 2207
rect 5836 2193 5853 2204
rect 5836 2064 5844 2193
rect 5896 2147 5904 2193
rect 6016 2147 6024 2193
rect 5836 2056 5853 2064
rect 5787 1984 5800 1987
rect 5787 1973 5804 1984
rect 5767 1924 5780 1927
rect 5767 1913 5784 1924
rect 5736 1787 5744 1873
rect 5756 1747 5764 1813
rect 5776 1687 5784 1913
rect 5796 1867 5804 1973
rect 5796 1807 5804 1853
rect 5376 1227 5384 1273
rect 5336 1167 5344 1213
rect 5336 1156 5353 1167
rect 5340 1153 5353 1156
rect 5356 1127 5364 1153
rect 4816 587 4824 633
rect 4836 607 4844 993
rect 4896 947 4904 973
rect 4936 947 4944 993
rect 4856 847 4864 873
rect 4916 847 4924 873
rect 4876 624 4884 753
rect 4916 747 4924 773
rect 4976 767 4984 873
rect 4916 647 4924 733
rect 4956 707 4964 733
rect 4916 636 4933 647
rect 4920 633 4933 636
rect 4876 616 4904 624
rect 4676 516 4704 524
rect 3987 413 4004 424
rect 4036 416 4073 424
rect 3996 387 4004 413
rect 4116 384 4124 413
rect 4067 376 4124 384
rect 3716 356 3733 367
rect 3720 353 3733 356
rect 3656 244 3664 353
rect 3736 267 3744 293
rect 3816 287 3824 373
rect 3967 364 3980 367
rect 3967 360 3984 364
rect 3967 353 3987 360
rect 3656 240 3684 244
rect 3656 236 3687 240
rect 3636 187 3644 233
rect 3673 227 3687 236
rect 3696 207 3704 253
rect 3816 187 3824 233
rect 3856 167 3864 333
rect 3676 127 3684 153
rect 3667 116 3684 127
rect 3667 113 3680 116
rect 3613 104 3627 113
rect 3613 100 3644 104
rect 3616 96 3644 100
rect 3636 64 3644 96
rect 3656 87 3664 113
rect 3716 87 3724 153
rect 3876 144 3884 353
rect 3973 347 3987 353
rect 3896 187 3904 253
rect 3996 247 4004 373
rect 4056 360 4093 364
rect 4053 356 4093 360
rect 4053 347 4067 356
rect 4136 284 4144 333
rect 4116 276 4144 284
rect 4096 187 4104 213
rect 4007 176 4033 184
rect 4087 176 4104 187
rect 4087 173 4100 176
rect 4116 144 4124 276
rect 3836 140 3884 144
rect 4096 140 4124 144
rect 3833 136 3884 140
rect 4093 136 4124 140
rect 3636 56 3664 64
rect 3176 -44 3224 -36
rect 3656 -36 3664 56
rect 3736 27 3744 133
rect 3833 127 3847 136
rect 4093 127 4107 136
rect 4156 127 4164 253
rect 4196 227 4204 433
rect 4256 407 4264 453
rect 4416 427 4424 453
rect 4336 364 4344 393
rect 4336 356 4384 364
rect 4236 340 4273 344
rect 4233 336 4273 340
rect 4233 327 4247 336
rect 4327 344 4340 347
rect 4327 340 4344 344
rect 4327 333 4347 340
rect 4333 327 4347 333
rect 4276 187 4284 293
rect 4376 287 4384 356
rect 4436 247 4444 333
rect 4456 287 4464 413
rect 4576 287 4584 393
rect 4616 367 4624 453
rect 4616 327 4624 353
rect 4676 307 4684 393
rect 4376 187 4384 213
rect 4456 187 4464 273
rect 4596 187 4604 233
rect 4587 176 4604 187
rect 4587 173 4600 176
rect 3987 124 4000 127
rect 3987 120 4004 124
rect 3987 113 4007 120
rect 4147 116 4164 127
rect 4147 113 4160 116
rect 3796 67 3804 113
rect 3836 87 3844 113
rect 3676 -24 3684 13
rect 3876 4 3884 93
rect 3936 67 3944 113
rect 3993 107 4007 113
rect 3856 -4 3884 4
rect 3856 -16 3864 -4
rect 3976 -16 3984 73
rect 4176 47 4184 173
rect 4327 116 4353 124
rect 4433 124 4447 133
rect 4407 120 4447 124
rect 4407 116 4444 120
rect 4656 124 4664 213
rect 4696 187 4704 516
rect 4756 427 4764 473
rect 4796 427 4804 453
rect 4756 187 4764 413
rect 4836 367 4844 393
rect 4827 356 4844 367
rect 4827 353 4840 356
rect 4656 116 4693 124
rect 4747 124 4760 127
rect 4747 120 4764 124
rect 4747 113 4767 120
rect 4596 87 4604 113
rect 4753 107 4767 113
rect 4816 107 4824 353
rect 4896 347 4904 616
rect 4976 607 4984 633
rect 5016 607 5024 1013
rect 5056 847 5064 933
rect 5076 887 5084 993
rect 5096 947 5104 973
rect 5136 947 5144 1053
rect 5176 787 5184 873
rect 5056 644 5064 733
rect 5076 704 5084 773
rect 5076 696 5113 704
rect 5056 636 5093 644
rect 5136 607 5144 633
rect 4936 347 4944 533
rect 5116 427 5124 453
rect 5056 347 5064 393
rect 4896 307 4904 333
rect 4836 247 4844 293
rect 4836 127 4844 233
rect 4936 204 4944 333
rect 5096 307 5104 353
rect 4916 196 4944 204
rect 4916 144 4924 196
rect 4896 140 4924 144
rect 4893 136 4924 140
rect 4893 127 4907 136
rect 4836 116 4853 127
rect 4840 113 4853 116
rect 4896 87 4904 113
rect 4956 27 4964 173
rect 5016 127 5024 233
rect 5136 227 5144 353
rect 5196 287 5204 1113
rect 5396 1087 5404 1153
rect 5476 1087 5484 1253
rect 5536 1227 5544 1333
rect 5516 1107 5524 1153
rect 5556 1127 5564 1153
rect 5316 947 5324 1073
rect 5307 936 5324 947
rect 5380 944 5393 947
rect 5307 933 5320 936
rect 5376 933 5393 944
rect 5256 647 5264 793
rect 5296 724 5304 773
rect 5296 716 5324 724
rect 5256 564 5264 633
rect 5276 607 5284 693
rect 5316 647 5324 716
rect 5356 707 5364 813
rect 5376 807 5384 933
rect 5416 807 5424 853
rect 5436 787 5444 933
rect 5456 767 5464 873
rect 5307 633 5324 647
rect 5287 596 5304 604
rect 5256 556 5284 564
rect 5236 444 5244 553
rect 5236 440 5264 444
rect 5236 436 5267 440
rect 5253 427 5267 436
rect 5276 367 5284 556
rect 5296 427 5304 596
rect 5316 587 5324 633
rect 5376 427 5384 573
rect 5396 467 5404 753
rect 5416 696 5453 704
rect 5416 607 5424 696
rect 5476 664 5484 1033
rect 5536 947 5544 973
rect 5596 884 5604 973
rect 5616 904 5624 1493
rect 5660 1464 5673 1467
rect 5656 1453 5673 1464
rect 5636 1404 5644 1453
rect 5656 1427 5664 1453
rect 5636 1396 5693 1404
rect 5816 1364 5824 2033
rect 5856 1987 5864 2053
rect 5896 1984 5904 2010
rect 5956 1927 5964 2133
rect 6056 2127 6064 2193
rect 6116 2024 6124 2390
rect 6136 1984 6144 2593
rect 6216 2507 6224 2553
rect 6236 2507 6244 2533
rect 6256 2524 6264 2893
rect 6296 2687 6304 2873
rect 6316 2867 6324 3053
rect 6356 2928 6364 3093
rect 6376 3067 6384 3773
rect 6396 3367 6404 3733
rect 6456 3667 6464 3953
rect 6476 3687 6484 3956
rect 6476 3307 6484 3673
rect 6467 3296 6484 3307
rect 6467 3293 6480 3296
rect 6416 3227 6424 3293
rect 6496 3284 6504 3653
rect 6516 3587 6524 5013
rect 6456 3276 6504 3284
rect 6416 3027 6424 3213
rect 6436 3064 6444 3253
rect 6456 3084 6464 3276
rect 6476 3107 6484 3213
rect 6516 3107 6524 3153
rect 6456 3076 6484 3084
rect 6436 3056 6464 3064
rect 6373 3004 6387 3013
rect 6373 3000 6424 3004
rect 6376 2996 6424 3000
rect 6396 2927 6404 2953
rect 6316 2727 6324 2813
rect 6336 2787 6344 2833
rect 6356 2827 6364 2892
rect 6396 2847 6404 2913
rect 6416 2887 6424 2996
rect 6436 2787 6444 2973
rect 6356 2687 6364 2713
rect 6256 2516 6284 2524
rect 6236 2496 6253 2507
rect 6240 2493 6253 2496
rect 6196 2404 6204 2430
rect 6216 2347 6224 2373
rect 6176 2267 6184 2293
rect 6216 2287 6224 2333
rect 6156 2167 6164 2193
rect 6176 2127 6184 2253
rect 6236 2204 6244 2313
rect 6276 2307 6284 2516
rect 6207 2196 6244 2204
rect 6296 2167 6304 2673
rect 6316 2327 6324 2493
rect 6416 2447 6424 2613
rect 6376 2267 6384 2293
rect 6356 2124 6364 2193
rect 6396 2167 6404 2193
rect 6356 2116 6384 2124
rect 6087 1976 6144 1984
rect 5887 1916 5953 1924
rect 5836 1587 5844 1733
rect 5916 1704 5924 1893
rect 6036 1867 6044 1973
rect 6096 1847 6104 1913
rect 6136 1887 6144 1976
rect 6196 1847 6204 2013
rect 6156 1747 6164 1813
rect 5987 1744 6000 1747
rect 5987 1733 6004 1744
rect 5916 1700 5964 1704
rect 5916 1696 5967 1700
rect 5953 1687 5967 1696
rect 5887 1676 5913 1684
rect 5996 1647 6004 1733
rect 6067 1676 6093 1684
rect 6136 1647 6144 1673
rect 5836 1447 5844 1473
rect 5973 1464 5987 1473
rect 5973 1460 6013 1464
rect 5976 1456 6013 1460
rect 5876 1367 5884 1393
rect 5796 1360 5824 1364
rect 5793 1356 5824 1360
rect 5793 1347 5807 1356
rect 5636 947 5644 1053
rect 5616 896 5644 904
rect 5596 876 5624 884
rect 5553 864 5567 873
rect 5536 860 5567 864
rect 5536 856 5564 860
rect 5536 807 5544 856
rect 5456 656 5484 664
rect 5436 427 5444 453
rect 5376 416 5393 427
rect 5380 413 5393 416
rect 5456 384 5464 656
rect 5516 647 5524 773
rect 5556 707 5564 773
rect 5476 587 5484 633
rect 5436 376 5464 384
rect 5156 144 5164 273
rect 5136 136 5164 144
rect 5056 87 5064 113
rect 5136 27 5144 136
rect 5216 127 5224 213
rect 5276 187 5284 353
rect 5316 267 5324 353
rect 5356 187 5364 213
rect 5396 144 5404 313
rect 5436 287 5444 376
rect 5496 367 5504 553
rect 5576 467 5584 833
rect 5616 824 5624 876
rect 5596 816 5624 824
rect 5596 787 5604 816
rect 5616 707 5624 753
rect 5636 664 5644 896
rect 5656 747 5664 1333
rect 5736 1227 5744 1293
rect 5756 1167 5764 1253
rect 5716 1107 5724 1153
rect 5676 964 5684 1053
rect 5816 987 5824 1213
rect 5836 1167 5844 1273
rect 5896 1167 5904 1313
rect 5936 1307 5944 1433
rect 5927 1224 5940 1227
rect 5927 1213 5944 1224
rect 5936 1167 5944 1213
rect 5976 1167 5984 1393
rect 6056 1367 6064 1453
rect 6036 1356 6053 1364
rect 5996 1267 6004 1313
rect 5996 1227 6004 1253
rect 5996 1216 6013 1227
rect 6000 1213 6013 1216
rect 6036 1204 6044 1356
rect 6016 1196 6044 1204
rect 5836 1156 5853 1167
rect 5840 1153 5853 1156
rect 5976 1156 5993 1167
rect 5980 1153 5993 1156
rect 5856 1127 5864 1153
rect 5896 1107 5904 1153
rect 5996 1067 6004 1153
rect 6016 1007 6024 1196
rect 6036 1127 6044 1153
rect 6096 1047 6104 1633
rect 6196 1607 6204 1833
rect 6236 1787 6244 2113
rect 6276 1987 6284 2013
rect 6316 1926 6324 2013
rect 6256 1887 6264 1912
rect 6316 1867 6324 1912
rect 6136 1327 6144 1453
rect 6156 1287 6164 1393
rect 6176 1347 6184 1453
rect 6216 1444 6224 1573
rect 6276 1547 6284 1673
rect 6296 1587 6304 1833
rect 6316 1687 6324 1773
rect 6356 1647 6364 2033
rect 6376 1927 6384 2116
rect 6416 2027 6424 2433
rect 6436 2307 6444 2773
rect 6436 2047 6444 2293
rect 6456 1987 6464 3056
rect 6416 1887 6424 1973
rect 6456 1848 6464 1973
rect 6476 1884 6484 3076
rect 6516 2647 6524 3013
rect 6476 1876 6493 1884
rect 6416 1747 6424 1773
rect 6456 1767 6464 1812
rect 6476 1704 6484 1793
rect 6456 1696 6484 1704
rect 6456 1687 6464 1696
rect 6447 1676 6464 1687
rect 6447 1673 6460 1676
rect 6196 1436 6224 1444
rect 6176 1307 6184 1333
rect 6196 1247 6204 1436
rect 6236 1307 6244 1533
rect 6256 1267 6264 1493
rect 6296 1407 6304 1513
rect 6316 1447 6324 1473
rect 6356 1467 6364 1593
rect 6396 1547 6404 1673
rect 6396 1447 6404 1493
rect 6416 1407 6424 1633
rect 6387 1376 6444 1384
rect 6336 1327 6344 1373
rect 6247 1224 6260 1227
rect 6300 1224 6313 1227
rect 6247 1213 6264 1224
rect 6160 1164 6173 1167
rect 6156 1153 6173 1164
rect 6156 1067 6164 1153
rect 6216 1107 6224 1153
rect 6256 1087 6264 1213
rect 6296 1213 6313 1224
rect 6296 1087 6304 1213
rect 6376 1167 6384 1333
rect 6336 1107 6344 1153
rect 5676 956 5724 964
rect 5716 947 5724 956
rect 5896 947 5904 973
rect 6056 947 6064 993
rect 6216 947 6224 973
rect 5716 936 5733 947
rect 5720 933 5733 936
rect 5760 944 5773 947
rect 5756 933 5773 944
rect 5827 936 5853 944
rect 6056 936 6073 947
rect 6060 933 6073 936
rect 6160 944 6173 947
rect 6156 933 6173 944
rect 5696 807 5704 933
rect 5756 807 5764 933
rect 5776 807 5784 873
rect 5636 656 5664 664
rect 5636 607 5644 633
rect 5596 547 5604 593
rect 5656 547 5664 656
rect 5676 587 5684 633
rect 5636 536 5653 544
rect 5587 424 5600 427
rect 5587 413 5604 424
rect 5467 356 5493 364
rect 5436 187 5444 273
rect 5436 176 5453 187
rect 5440 173 5453 176
rect 5376 140 5404 144
rect 5373 136 5404 140
rect 5373 127 5387 136
rect 5476 127 5484 253
rect 5516 204 5524 293
rect 5536 247 5544 413
rect 5596 367 5604 413
rect 5636 267 5644 536
rect 5736 487 5744 733
rect 5776 647 5784 753
rect 5816 747 5824 773
rect 5816 707 5824 733
rect 5836 647 5844 853
rect 5876 827 5884 873
rect 5976 827 5984 873
rect 5876 767 5884 813
rect 5776 636 5793 647
rect 5780 633 5793 636
rect 5876 587 5884 693
rect 5756 427 5764 453
rect 5716 307 5724 413
rect 5796 367 5804 493
rect 5876 427 5884 573
rect 5936 527 5944 693
rect 5976 567 5984 813
rect 6016 807 6024 873
rect 6036 827 6044 933
rect 6156 887 6164 933
rect 6256 887 6264 1033
rect 6296 944 6304 993
rect 6296 936 6333 944
rect 5996 796 6013 804
rect 5996 647 6004 796
rect 6056 747 6064 833
rect 6016 707 6024 733
rect 6116 707 6124 793
rect 6196 707 6204 873
rect 6036 607 6044 633
rect 6136 567 6144 633
rect 6176 607 6184 633
rect 5976 447 5984 553
rect 5933 427 5947 433
rect 5927 420 5947 427
rect 5927 416 5944 420
rect 5927 413 5940 416
rect 5733 344 5747 353
rect 5733 340 5764 344
rect 5736 336 5764 340
rect 5756 247 5764 336
rect 5496 196 5524 204
rect 5496 127 5504 196
rect 5536 187 5544 233
rect 5696 187 5704 213
rect 5836 187 5844 413
rect 5936 327 5944 353
rect 6036 347 6044 533
rect 6296 524 6304 936
rect 6387 944 6400 947
rect 6387 933 6404 944
rect 6356 847 6364 873
rect 6336 836 6353 844
rect 6336 707 6344 836
rect 6316 587 6324 633
rect 6356 607 6364 633
rect 6296 516 6324 524
rect 6196 427 6204 473
rect 6316 467 6324 516
rect 6116 420 6153 424
rect 6113 416 6153 420
rect 6113 407 6127 416
rect 5956 187 5964 233
rect 5976 227 5984 293
rect 5976 127 5984 213
rect 5496 116 5513 127
rect 5500 113 5513 116
rect 5727 116 5753 124
rect 5907 116 5933 124
rect 5176 67 5184 113
rect 5336 87 5344 113
rect 5676 87 5684 113
rect 6036 107 6044 333
rect 6076 287 6084 333
rect 6087 276 6104 284
rect 6096 187 6104 276
rect 6116 247 6124 353
rect 6136 247 6144 416
rect 6316 367 6324 453
rect 6356 427 6364 593
rect 6396 587 6404 933
rect 6416 747 6424 1293
rect 6436 1287 6444 1376
rect 6456 887 6464 1633
rect 6476 987 6484 1593
rect 6496 1527 6504 1873
rect 6516 1487 6524 2153
rect 6496 1327 6504 1393
rect 6396 187 6404 473
rect 6396 176 6413 187
rect 6400 173 6413 176
rect 6216 136 6304 144
rect 6100 124 6113 127
rect 6096 120 6113 124
rect 6093 113 6113 120
rect 6216 124 6224 136
rect 6296 127 6304 136
rect 6240 124 6253 127
rect 6167 116 6224 124
rect 6236 113 6253 124
rect 6307 116 6333 124
rect 6093 107 6107 113
rect 6236 104 6244 113
rect 6207 96 6244 104
rect 3836 -24 3864 -16
rect 3956 -24 3984 -16
rect 5176 -24 5184 13
rect 3836 -36 3844 -24
rect 3656 -44 3844 -36
use INVX1  _927_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493700
transform 1 0 5630 0 -1 5470
box -6 -8 66 272
use NOR2X1  _928_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727495070
transform -1 0 5690 0 1 4950
box -6 -8 86 272
use NAND2X1  _929_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494699
transform -1 0 5970 0 1 4950
box -6 -8 86 272
use INVX1  _930_
timestamp 1727493700
transform 1 0 6050 0 1 4950
box -6 -8 66 272
use INVX1  _931_
timestamp 1727493700
transform -1 0 5390 0 1 5470
box -6 -8 66 272
use INVX2  _932_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493898
transform -1 0 3490 0 -1 4950
box -6 -8 66 272
use NOR2X1  _933_
timestamp 1727495070
transform 1 0 5490 0 -1 5470
box -6 -8 86 272
use NAND2X1  _934_
timestamp 1727494699
transform 1 0 5450 0 1 5470
box -6 -8 86 272
use INVX1  _935_
timestamp 1727493700
transform 1 0 6010 0 1 5990
box -6 -8 66 272
use NOR2X1  _936_
timestamp 1727495070
transform -1 0 5450 0 -1 5990
box -6 -8 86 272
use AOI21X1  _937_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform 1 0 5610 0 1 5470
box -6 -8 106 272
use NOR2X1  _938_
timestamp 1727495070
transform -1 0 5990 0 -1 6510
box -6 -8 86 272
use OAI21X1  _939_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727498925
transform 1 0 6050 0 -1 6510
box -6 -8 106 272
use INVX1  _940_
timestamp 1727493700
transform 1 0 6270 0 1 5470
box -6 -8 66 272
use INVX4  _941_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494067
transform 1 0 3850 0 -1 4950
box -6 -8 86 272
use OAI21X1  _942_
timestamp 1727498925
transform 1 0 5750 0 -1 5470
box -6 -8 106 272
use INVX1  _943_
timestamp 1727493700
transform 1 0 6010 0 -1 5990
box -6 -8 66 272
use NOR2X1  _944_
timestamp 1727495070
transform 1 0 5750 0 1 4950
box -6 -8 86 272
use INVX1  _945_
timestamp 1727493700
transform 1 0 6290 0 -1 5470
box -6 -8 66 272
use INVX1  _946_
timestamp 1727493700
transform -1 0 5850 0 -1 6510
box -6 -8 66 272
use OAI21X1  _947_
timestamp 1727498925
transform 1 0 5770 0 1 5470
box -6 -8 106 272
use OAI21X1  _948_
timestamp 1727498925
transform -1 0 6050 0 1 5470
box -6 -8 106 272
use AOI22X1  _949_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487144
transform 1 0 5910 0 -1 5470
box -6 -8 126 272
use NAND2X1  _950_
timestamp 1727494699
transform -1 0 5730 0 -1 6510
box -6 -8 86 272
use OAI21X1  _951_
timestamp 1727498925
transform -1 0 6230 0 -1 5990
box -6 -8 106 272
use OAI21X1  _952_
timestamp 1727498925
transform -1 0 5790 0 -1 5990
box -6 -8 106 272
use NAND2X1  _953_
timestamp 1727494699
transform 1 0 5230 0 -1 5990
box -6 -8 86 272
use NOR2X1  _954_
timestamp 1727495070
transform 1 0 6290 0 -1 5990
box -6 -8 86 272
use NOR2X1  _955_
timestamp 1727495070
transform 1 0 6210 0 -1 6510
box -6 -8 86 272
use OAI22X1  _956_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727495774
transform -1 0 5950 0 1 5990
box -6 -8 126 272
use OR2X2  _957_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727496117
transform -1 0 5610 0 -1 5990
box -6 -8 106 272
use INVX1  _958_
timestamp 1727493700
transform 1 0 6310 0 1 5990
box -6 -8 66 272
use AOI22X1  _959_
timestamp 1727487144
transform -1 0 6250 0 1 5990
box -6 -8 126 272
use NAND3X1  _960_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494898
transform 1 0 6110 0 -1 5470
box -6 -8 106 272
use AND2X2  _961_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform -1 0 6210 0 1 5470
box -6 -8 106 273
use OAI21X1  _962_
timestamp 1727498925
transform 1 0 5850 0 -1 5990
box -6 -8 106 272
use INVX1  _963_
timestamp 1727493700
transform -1 0 5590 0 -1 6510
box -6 -8 66 272
use INVX1  _964_
timestamp 1727493700
transform -1 0 5410 0 -1 5470
box -6 -8 66 272
use NAND2X1  _965_
timestamp 1727494699
transform 1 0 4510 0 -1 5470
box -6 -8 86 272
use OAI21X1  _966_
timestamp 1727498925
transform -1 0 4750 0 -1 5470
box -6 -8 106 272
use INVX1  _967_
timestamp 1727493700
transform 1 0 4970 0 1 5470
box -6 -8 66 272
use NAND2X1  _968_
timestamp 1727494699
transform 1 0 5170 0 1 4950
box -6 -8 86 272
use OAI21X1  _969_
timestamp 1727498925
transform 1 0 5050 0 -1 5470
box -6 -8 106 272
use INVX1  _970_
timestamp 1727493700
transform 1 0 4090 0 -1 6510
box -6 -8 66 272
use NAND2X1  _971_
timestamp 1727494699
transform 1 0 4890 0 -1 6510
box -6 -8 86 272
use OAI21X1  _972_
timestamp 1727498925
transform 1 0 4710 0 -1 6510
box -6 -8 106 272
use INVX1  _973_
timestamp 1727493700
transform 1 0 4370 0 -1 5990
box -6 -8 66 272
use NAND2X1  _974_
timestamp 1727494699
transform 1 0 4390 0 1 3390
box -6 -8 86 272
use OAI21X1  _975_
timestamp 1727498925
transform 1 0 4470 0 -1 3910
box -6 -8 106 272
use INVX1  _976_
timestamp 1727493700
transform 1 0 3710 0 -1 4950
box -6 -8 66 272
use NAND2X1  _977_
timestamp 1727494699
transform 1 0 3990 0 1 3390
box -6 -8 86 272
use OAI21X1  _978_
timestamp 1727498925
transform 1 0 3770 0 1 3910
box -6 -8 106 272
use INVX1  _979_
timestamp 1727493700
transform 1 0 3190 0 1 3910
box -6 -8 66 272
use NAND2X1  _980_
timestamp 1727494699
transform 1 0 3330 0 -1 3910
box -6 -8 86 272
use OAI21X1  _981_
timestamp 1727498925
transform -1 0 3270 0 -1 3910
box -6 -8 106 272
use INVX1  _982_
timestamp 1727493700
transform 1 0 2110 0 -1 4430
box -6 -8 66 272
use NAND2X1  _983_
timestamp 1727494699
transform 1 0 2710 0 1 3910
box -6 -8 86 272
use OAI21X1  _984_
timestamp 1727498925
transform -1 0 2950 0 1 3910
box -6 -8 106 272
use INVX4  _985_
timestamp 1727494067
transform 1 0 3650 0 -1 3390
box -6 -8 86 272
use NAND2X1  _986_
timestamp 1727494699
transform 1 0 3950 0 1 3910
box -6 -8 86 272
use OAI21X1  _987_
timestamp 1727498925
transform -1 0 4190 0 1 3910
box -6 -8 106 272
use INVX1  _988_
timestamp 1727493700
transform -1 0 2390 0 1 4430
box -6 -8 66 272
use INVX1  _989_
timestamp 1727493700
transform 1 0 5270 0 1 1830
box -6 -8 66 272
use INVX2  _990_
timestamp 1727493898
transform -1 0 1850 0 -1 2350
box -6 -8 66 272
use NOR2X1  _991_
timestamp 1727495070
transform 1 0 5610 0 1 2350
box -6 -8 86 272
use AND2X2  _992_
timestamp 1727487319
transform 1 0 5450 0 1 2350
box -6 -8 106 273
use NAND2X1  _993_
timestamp 1727494699
transform 1 0 5770 0 1 2350
box -6 -8 86 272
use NAND2X1  _994_
timestamp 1727494699
transform -1 0 4390 0 -1 4430
box -6 -8 86 272
use NAND2X1  _995_
timestamp 1727494699
transform -1 0 4710 0 -1 3910
box -6 -8 86 272
use OR2X2  _996_
timestamp 1727496117
transform 1 0 6290 0 -1 4430
box -6 -8 106 272
use NAND2X1  _997_
timestamp 1727494699
transform 1 0 5510 0 1 4430
box -6 -8 86 272
use AND2X2  _998_
timestamp 1727487319
transform -1 0 6370 0 1 4430
box -6 -8 106 273
use OAI21X1  _999_
timestamp 1727498925
transform 1 0 6110 0 1 4430
box -6 -8 106 272
use NAND2X1  _1000_
timestamp 1727494699
transform -1 0 4990 0 1 3910
box -6 -8 86 272
use INVX1  _1001_
timestamp 1727493700
transform 1 0 5350 0 1 3910
box -6 -8 66 272
use NAND2X1  _1002_
timestamp 1727494699
transform 1 0 4690 0 1 3390
box -6 -8 86 272
use OR2X2  _1003_
timestamp 1727496117
transform 1 0 4770 0 -1 3910
box -6 -8 106 272
use AOI22X1  _1004_
timestamp 1727487144
transform 1 0 4710 0 1 3910
box -6 -8 126 272
use INVX1  _1005_
timestamp 1727493700
transform -1 0 5290 0 1 3910
box -6 -8 66 272
use NAND3X1  _1006_
timestamp 1727494898
transform 1 0 5630 0 1 3910
box -6 -8 106 272
use NOR2X1  _1007_
timestamp 1727495070
transform -1 0 5010 0 -1 3910
box -6 -8 86 272
use OAI21X1  _1008_
timestamp 1727498925
transform -1 0 5170 0 1 3910
box -6 -8 106 272
use NAND3X1  _1009_
timestamp 1727494898
transform 1 0 5950 0 1 3910
box -6 -8 106 272
use INVX1  _1010_
timestamp 1727493700
transform -1 0 5430 0 -1 4430
box -6 -8 66 272
use NAND2X1  _1011_
timestamp 1727494699
transform 1 0 4990 0 1 3390
box -6 -8 86 272
use INVX2  _1012_
timestamp 1727493898
transform -1 0 3550 0 1 2350
box -6 -8 66 272
use NAND2X1  _1013_
timestamp 1727494699
transform -1 0 4430 0 1 2350
box -6 -8 86 272
use OAI21X1  _1014_
timestamp 1727498925
transform 1 0 5290 0 1 2350
box -6 -8 106 272
use OAI21X1  _1015_
timestamp 1727498925
transform 1 0 5310 0 1 3390
box -6 -8 106 272
use AOI21X1  _1016_
timestamp 1727487319
transform -1 0 5890 0 1 3910
box -6 -8 106 272
use OAI21X1  _1017_
timestamp 1727498925
transform 1 0 5630 0 1 3390
box -6 -8 106 272
use OAI21X1  _1018_
timestamp 1727498925
transform 1 0 5070 0 -1 3910
box -6 -8 106 272
use AND2X2  _1019_
timestamp 1727487319
transform 1 0 4010 0 -1 2870
box -6 -8 106 273
use NAND3X1  _1020_
timestamp 1727494898
transform 1 0 4170 0 -1 2870
box -6 -8 106 272
use AOI22X1  _1021_
timestamp 1727487144
transform -1 0 4330 0 -1 3390
box -6 -8 126 272
use INVX1  _1022_
timestamp 1727493700
transform 1 0 4550 0 -1 3390
box -6 -8 66 272
use NAND2X1  _1023_
timestamp 1727494699
transform -1 0 4170 0 1 2870
box -6 -8 86 272
use INVX1  _1024_
timestamp 1727493700
transform -1 0 4890 0 -1 3390
box -6 -8 66 272
use NAND3X1  _1025_
timestamp 1727494898
transform 1 0 4670 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1026_
timestamp 1727494699
transform -1 0 4630 0 1 3390
box -6 -8 86 272
use NOR2X1  _1027_
timestamp 1727495070
transform 1 0 4830 0 1 3390
box -6 -8 86 272
use OAI21X1  _1028_
timestamp 1727498925
transform 1 0 4950 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1029_
timestamp 1727494898
transform 1 0 5270 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1030_
timestamp 1727487319
transform -1 0 5350 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1031_
timestamp 1727498925
transform -1 0 4810 0 1 2870
box -6 -8 106 272
use NAND3X1  _1032_
timestamp 1727494898
transform -1 0 4490 0 1 2870
box -6 -8 106 272
use NAND3X1  _1033_
timestamp 1727494898
transform 1 0 4870 0 1 2870
box -6 -8 106 272
use NAND2X1  _1034_
timestamp 1727494699
transform -1 0 4430 0 -1 2870
box -6 -8 86 272
use INVX1  _1035_
timestamp 1727493700
transform 1 0 4650 0 -1 2870
box -6 -8 66 272
use AND2X2  _1036_
timestamp 1727487319
transform 1 0 4490 0 -1 2870
box -6 -8 106 273
use NAND2X1  _1037_
timestamp 1727494699
transform -1 0 5230 0 1 2350
box -6 -8 86 272
use INVX1  _1038_
timestamp 1727493700
transform 1 0 4590 0 -1 1310
box -6 -8 66 272
use OAI21X1  _1039_
timestamp 1727498925
transform 1 0 4810 0 1 2350
box -6 -8 106 272
use NAND3X1  _1040_
timestamp 1727494898
transform 1 0 4770 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1041_
timestamp 1727498925
transform 1 0 4990 0 1 2350
box -6 -8 106 272
use INVX1  _1042_
timestamp 1727493700
transform 1 0 5530 0 -1 2350
box -6 -8 66 272
use OAI21X1  _1043_
timestamp 1727498925
transform -1 0 5170 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1044_
timestamp 1727494898
transform 1 0 4930 0 -1 2870
box -6 -8 106 272
use AND2X2  _1045_
timestamp 1727487319
transform 1 0 5270 0 -1 2870
box -6 -8 106 273
use NAND3X1  _1046_
timestamp 1727494898
transform 1 0 5670 0 1 2870
box -6 -8 106 272
use AOI21X1  _1047_
timestamp 1727487319
transform 1 0 5030 0 1 2870
box -6 -8 106 272
use AOI21X1  _1048_
timestamp 1727487319
transform 1 0 5110 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1049_
timestamp 1727494699
transform 1 0 5110 0 -1 2870
box -6 -8 86 272
use OAI21X1  _1050_
timestamp 1727498925
transform 1 0 5350 0 1 2870
box -6 -8 106 272
use NAND3X1  _1051_
timestamp 1727494898
transform 1 0 5830 0 1 2870
box -6 -8 106 272
use AOI21X1  _1052_
timestamp 1727487319
transform 1 0 6010 0 1 2870
box -6 -8 106 272
use OAI21X1  _1053_
timestamp 1727498925
transform 1 0 6390 0 1 5470
box -6 -8 106 272
use AOI21X1  _1054_
timestamp 1727487319
transform 1 0 5430 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1055_
timestamp 1727498925
transform -1 0 4330 0 1 2870
box -6 -8 106 272
use AND2X2  _1056_
timestamp 1727487319
transform -1 0 3030 0 1 1830
box -6 -8 106 273
use NAND2X1  _1057_
timestamp 1727494699
transform -1 0 4130 0 1 1830
box -6 -8 86 272
use INVX1  _1058_
timestamp 1727493700
transform -1 0 4290 0 1 2350
box -6 -8 66 272
use INVX2  _1059_
timestamp 1727493898
transform 1 0 3150 0 1 2870
box -6 -8 66 272
use NAND2X1  _1060_
timestamp 1727494699
transform 1 0 3930 0 1 2350
box -6 -8 86 272
use OAI21X1  _1061_
timestamp 1727498925
transform 1 0 4070 0 1 2350
box -6 -8 106 272
use NAND2X1  _1062_
timestamp 1727494699
transform 1 0 4330 0 -1 2350
box -6 -8 86 272
use INVX1  _1063_
timestamp 1727493700
transform -1 0 4390 0 1 1830
box -6 -8 66 272
use NAND3X1  _1064_
timestamp 1727494898
transform -1 0 4130 0 1 1310
box -6 -8 106 272
use NAND2X1  _1065_
timestamp 1727494699
transform -1 0 4010 0 -1 1830
box -6 -8 86 272
use NOR2X1  _1066_
timestamp 1727495070
transform -1 0 4270 0 1 1830
box -6 -8 86 272
use AOI22X1  _1067_
timestamp 1727487144
transform 1 0 4090 0 -1 1830
box -6 -8 126 272
use OAI21X1  _1068_
timestamp 1727498925
transform -1 0 4710 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1069_
timestamp 1727487319
transform -1 0 4450 0 1 1310
box -6 -8 106 272
use AOI21X1  _1070_
timestamp 1727487319
transform 1 0 4550 0 1 2870
box -6 -8 106 272
use OAI21X1  _1071_
timestamp 1727498925
transform 1 0 4790 0 -1 1830
box -6 -8 106 272
use NAND3X1  _1072_
timestamp 1727494898
transform 1 0 4450 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1073_
timestamp 1727487319
transform 1 0 5110 0 -1 1830
box -6 -8 106 272
use NAND2X1  _1074_
timestamp 1727494699
transform 1 0 4470 0 -1 2350
box -6 -8 86 272
use INVX1  _1075_
timestamp 1727493700
transform -1 0 4850 0 1 1830
box -6 -8 66 272
use AND2X2  _1076_
timestamp 1727487319
transform -1 0 4710 0 -1 2350
box -6 -8 106 273
use AND2X2  _1077_
timestamp 1727487319
transform 1 0 4490 0 1 2350
box -6 -8 106 273
use NAND2X1  _1078_
timestamp 1727494699
transform -1 0 4850 0 -1 2350
box -6 -8 86 272
use INVX2  _1079_
timestamp 1727493898
transform 1 0 3810 0 1 2870
box -6 -8 66 272
use NAND2X1  _1080_
timestamp 1727494699
transform -1 0 5310 0 -1 2350
box -6 -8 86 272
use OAI21X1  _1081_
timestamp 1727498925
transform -1 0 5010 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1082_
timestamp 1727494898
transform 1 0 5110 0 1 1830
box -6 -8 106 272
use OAI21X1  _1083_
timestamp 1727498925
transform 1 0 4450 0 1 1830
box -6 -8 106 272
use OAI21X1  _1084_
timestamp 1727498925
transform 1 0 4650 0 1 2350
box -6 -8 106 272
use NAND3X1  _1085_
timestamp 1727494898
transform 1 0 4610 0 1 1830
box -6 -8 106 272
use AND2X2  _1086_
timestamp 1727487319
transform 1 0 5450 0 -1 1830
box -6 -8 106 273
use OAI21X1  _1087_
timestamp 1727498925
transform 1 0 5170 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1088_
timestamp 1727494898
transform 1 0 4950 0 -1 1830
box -6 -8 106 272
use NAND3X1  _1089_
timestamp 1727494898
transform 1 0 4510 0 1 1310
box -6 -8 106 272
use NAND2X1  _1090_
timestamp 1727494699
transform -1 0 5370 0 -1 1830
box -6 -8 86 272
use NAND3X1  _1091_
timestamp 1727494898
transform 1 0 4850 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1092_
timestamp 1727494898
transform 1 0 5510 0 -1 1310
box -6 -8 106 272
use OAI21X1  _1093_
timestamp 1727498925
transform 1 0 5190 0 1 2870
box -6 -8 106 272
use NAND3X1  _1094_
timestamp 1727494898
transform 1 0 4870 0 1 1310
box -6 -8 106 272
use OAI21X1  _1095_
timestamp 1727498925
transform 1 0 5030 0 1 1310
box -6 -8 106 272
use NAND3X1  _1096_
timestamp 1727494898
transform 1 0 5350 0 1 1310
box -6 -8 106 272
use INVX4  _1097_
timestamp 1727494067
transform -1 0 1710 0 -1 3910
box -6 -8 86 272
use NOR2X1  _1098_
timestamp 1727495070
transform 1 0 5610 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1099_
timestamp 1727498925
transform 1 0 5370 0 -1 2350
box -6 -8 106 272
use NAND2X1  _1100_
timestamp 1727494699
transform -1 0 5590 0 1 1310
box -6 -8 86 272
use OR2X2  _1101_
timestamp 1727496117
transform 1 0 5670 0 1 1310
box -6 -8 106 272
use AND2X2  _1102_
timestamp 1727487319
transform 1 0 5830 0 1 1310
box -6 -8 106 273
use NAND3X1  _1103_
timestamp 1727494898
transform 1 0 6130 0 1 1310
box -6 -8 106 272
use AOI21X1  _1104_
timestamp 1727487319
transform 1 0 5190 0 1 1310
box -6 -8 106 272
use AOI21X1  _1105_
timestamp 1727487319
transform 1 0 5350 0 -1 1310
box -6 -8 106 272
use NAND2X1  _1106_
timestamp 1727494699
transform -1 0 6070 0 1 1310
box -6 -8 86 272
use OAI21X1  _1107_
timestamp 1727498925
transform -1 0 6250 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1108_
timestamp 1727494898
transform 1 0 6410 0 -1 5470
box -6 -8 106 272
use INVX1  _1109_
timestamp 1727493700
transform 1 0 6310 0 1 270
box -6 -8 66 272
use OAI21X1  _1110_
timestamp 1727498925
transform -1 0 5930 0 -1 1310
box -6 -8 106 272
use AOI21X1  _1111_
timestamp 1727487319
transform 1 0 5010 0 -1 1310
box -6 -8 106 272
use OAI21X1  _1112_
timestamp 1727498925
transform -1 0 4390 0 -1 1830
box -6 -8 106 272
use NAND3X1  _1113_
timestamp 1727494898
transform -1 0 3870 0 -1 1830
box -6 -8 106 272
use AOI22X1  _1114_
timestamp 1727487144
transform -1 0 3710 0 -1 1830
box -6 -8 126 272
use INVX1  _1115_
timestamp 1727493700
transform -1 0 3230 0 -1 1310
box -6 -8 66 272
use NAND2X1  _1116_
timestamp 1727494699
transform -1 0 3370 0 1 1830
box -6 -8 86 272
use INVX1  _1117_
timestamp 1727493700
transform -1 0 3530 0 -1 1310
box -6 -8 66 272
use NAND3X1  _1118_
timestamp 1727494898
transform 1 0 3770 0 1 790
box -6 -8 106 272
use NAND2X1  _1119_
timestamp 1727494699
transform -1 0 3850 0 1 2350
box -6 -8 86 272
use NOR2X1  _1120_
timestamp 1727495070
transform -1 0 3950 0 -1 2350
box -6 -8 86 272
use OAI21X1  _1121_
timestamp 1727498925
transform -1 0 3690 0 -1 1310
box -6 -8 106 272
use AOI21X1  _1122_
timestamp 1727487319
transform 1 0 4250 0 1 790
box -6 -8 106 272
use OAI21X1  _1123_
timestamp 1727498925
transform 1 0 3750 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1124_
timestamp 1727494898
transform -1 0 3410 0 -1 1310
box -6 -8 106 272
use AOI22X1  _1125_
timestamp 1727487144
transform -1 0 4510 0 -1 1310
box -6 -8 126 272
use NAND2X1  _1126_
timestamp 1727494699
transform -1 0 3510 0 1 1830
box -6 -8 86 272
use INVX1  _1127_
timestamp 1727493700
transform -1 0 3510 0 1 1310
box -6 -8 66 272
use AND2X2  _1128_
timestamp 1727487319
transform 1 0 3690 0 -1 2350
box -6 -8 106 273
use AND2X2  _1129_
timestamp 1727487319
transform 1 0 4010 0 -1 2350
box -6 -8 106 273
use NAND2X1  _1130_
timestamp 1727494699
transform 1 0 3910 0 1 1830
box -6 -8 86 272
use AOI22X1  _1131_
timestamp 1727487144
transform -1 0 3630 0 -1 2350
box -6 -8 126 272
use INVX1  _1132_
timestamp 1727493700
transform 1 0 3570 0 1 1310
box -6 -8 66 272
use NAND3X1  _1133_
timestamp 1727494898
transform 1 0 3690 0 1 1310
box -6 -8 106 272
use INVX1  _1134_
timestamp 1727493700
transform -1 0 3430 0 1 2350
box -6 -8 66 272
use OAI21X1  _1135_
timestamp 1727498925
transform 1 0 3590 0 1 1830
box -6 -8 106 272
use OAI21X1  _1136_
timestamp 1727498925
transform -1 0 4270 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1137_
timestamp 1727494898
transform 1 0 3750 0 1 1830
box -6 -8 106 272
use AND2X2  _1138_
timestamp 1727487319
transform 1 0 4070 0 -1 1310
box -6 -8 106 273
use OAI21X1  _1139_
timestamp 1727498925
transform 1 0 4610 0 -1 790
box -6 -8 106 272
use AOI21X1  _1140_
timestamp 1727487319
transform 1 0 4190 0 1 1310
box -6 -8 106 272
use NAND3X1  _1141_
timestamp 1727494898
transform 1 0 4230 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1142_
timestamp 1727494898
transform -1 0 4190 0 1 790
box -6 -8 106 272
use NAND2X1  _1143_
timestamp 1727494699
transform -1 0 3990 0 -1 1310
box -6 -8 86 272
use NAND3X1  _1144_
timestamp 1727494898
transform 1 0 4770 0 -1 790
box -6 -8 106 272
use NAND3X1  _1145_
timestamp 1727494898
transform 1 0 5090 0 -1 790
box -6 -8 106 272
use OAI21X1  _1146_
timestamp 1727498925
transform -1 0 4790 0 1 1310
box -6 -8 106 272
use NAND3X1  _1147_
timestamp 1727494898
transform 1 0 4730 0 1 790
box -6 -8 106 272
use OAI21X1  _1148_
timestamp 1727498925
transform 1 0 4570 0 1 790
box -6 -8 106 272
use NAND3X1  _1149_
timestamp 1727494898
transform 1 0 5050 0 1 790
box -6 -8 106 272
use NAND2X1  _1150_
timestamp 1727494699
transform -1 0 5310 0 1 790
box -6 -8 86 272
use INVX1  _1151_
timestamp 1727493700
transform -1 0 5850 0 -1 270
box -6 -8 66 272
use AOI22X1  _1152_
timestamp 1727487144
transform 1 0 4910 0 1 1830
box -6 -8 126 272
use INVX1  _1153_
timestamp 1727493700
transform 1 0 6410 0 -1 270
box -6 -8 66 272
use OAI21X1  _1154_
timestamp 1727498925
transform 1 0 6090 0 -1 270
box -6 -8 106 272
use NOR2X1  _1155_
timestamp 1727495070
transform -1 0 6090 0 1 270
box -6 -8 86 272
use NAND2X1  _1156_
timestamp 1727494699
transform 1 0 6150 0 1 270
box -6 -8 86 272
use NAND3X1  _1157_
timestamp 1727494898
transform 1 0 5930 0 -1 270
box -6 -8 106 272
use NAND2X1  _1158_
timestamp 1727494699
transform 1 0 6250 0 -1 270
box -6 -8 86 272
use OAI21X1  _1159_
timestamp 1727498925
transform 1 0 5450 0 -1 270
box -6 -8 106 272
use NAND3X1  _1160_
timestamp 1727494898
transform -1 0 5390 0 -1 270
box -6 -8 106 272
use NAND2X1  _1161_
timestamp 1727494699
transform -1 0 5230 0 -1 270
box -6 -8 86 272
use NAND3X1  _1162_
timestamp 1727494898
transform 1 0 5250 0 -1 790
box -6 -8 106 272
use AOI21X1  _1163_
timestamp 1727487319
transform 1 0 4890 0 1 790
box -6 -8 106 272
use AOI21X1  _1164_
timestamp 1727487319
transform 1 0 4930 0 -1 790
box -6 -8 106 272
use NAND3X1  _1165_
timestamp 1727494898
transform -1 0 5730 0 -1 270
box -6 -8 106 272
use NAND3X1  _1166_
timestamp 1727494898
transform -1 0 5770 0 1 270
box -6 -8 106 272
use NAND2X1  _1167_
timestamp 1727494699
transform 1 0 5530 0 1 270
box -6 -8 86 272
use OAI21X1  _1168_
timestamp 1727498925
transform 1 0 5610 0 -1 790
box -6 -8 106 272
use AOI21X1  _1169_
timestamp 1727487319
transform 1 0 5850 0 1 790
box -6 -8 106 272
use AOI21X1  _1170_
timestamp 1727487319
transform -1 0 5770 0 -1 1310
box -6 -8 106 272
use OAI21X1  _1171_
timestamp 1727498925
transform -1 0 5470 0 1 790
box -6 -8 106 272
use NAND3X1  _1172_
timestamp 1727494898
transform 1 0 5430 0 -1 790
box -6 -8 106 272
use AOI21X1  _1173_
timestamp 1727487319
transform 1 0 5690 0 1 790
box -6 -8 106 272
use OAI21X1  _1174_
timestamp 1727498925
transform 1 0 6110 0 -1 790
box -6 -8 106 272
use NAND3X1  _1175_
timestamp 1727494898
transform 1 0 5530 0 1 790
box -6 -8 106 272
use NAND3X1  _1176_
timestamp 1727494898
transform 1 0 5790 0 -1 790
box -6 -8 106 272
use NAND3X1  _1177_
timestamp 1727494898
transform 1 0 6330 0 1 790
box -6 -8 106 272
use AOI21X1  _1178_
timestamp 1727487319
transform 1 0 6390 0 -1 1830
box -6 -8 106 272
use INVX1  _1179_
timestamp 1727493700
transform 1 0 5750 0 -1 1830
box -6 -8 66 272
use INVX1  _1180_
timestamp 1727493700
transform 1 0 6450 0 -1 3390
box -6 -8 66 272
use NOR2X1  _1181_
timestamp 1727495070
transform 1 0 6150 0 -1 4430
box -6 -8 86 272
use INVX1  _1182_
timestamp 1727493700
transform -1 0 5890 0 1 4430
box -6 -8 66 272
use INVX1  _1183_
timestamp 1727493700
transform -1 0 4630 0 1 3910
box -6 -8 66 272
use OAI21X1  _1184_
timestamp 1727498925
transform 1 0 4450 0 -1 4430
box -6 -8 106 272
use AOI21X1  _1185_
timestamp 1727487319
transform 1 0 5990 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1186_
timestamp 1727498925
transform 1 0 5410 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1187_
timestamp 1727494898
transform 1 0 5590 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1188_
timestamp 1727487319
transform 1 0 5750 0 -1 3910
box -6 -8 106 272
use AND2X2  _1189_
timestamp 1727487319
transform -1 0 5690 0 -1 3390
box -6 -8 106 273
use NAND3X1  _1190_
timestamp 1727494898
transform 1 0 5910 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1191_
timestamp 1727487319
transform -1 0 5910 0 1 3390
box -6 -8 106 272
use OAI21X1  _1192_
timestamp 1727498925
transform 1 0 5510 0 1 2870
box -6 -8 106 272
use NAND3X1  _1193_
timestamp 1727494898
transform 1 0 5430 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1194_
timestamp 1727494898
transform 1 0 5750 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1195_
timestamp 1727494898
transform 1 0 6310 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1196_
timestamp 1727498925
transform 1 0 6310 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1197_
timestamp 1727494898
transform 1 0 5990 0 -1 1310
box -6 -8 106 272
use AOI22X1  _1198_
timestamp 1727487144
transform 1 0 6310 0 1 1310
box -6 -8 126 272
use NAND3X1  _1199_
timestamp 1727494898
transform -1 0 6370 0 -1 790
box -6 -8 106 272
use OAI21X1  _1200_
timestamp 1727498925
transform 1 0 6010 0 1 790
box -6 -8 106 272
use AOI21X1  _1201_
timestamp 1727487319
transform 1 0 6170 0 1 790
box -6 -8 106 272
use NAND3X1  _1202_
timestamp 1727494898
transform 1 0 5990 0 1 3390
box -6 -8 106 272
use NAND3X1  _1203_
timestamp 1727494898
transform -1 0 5930 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1204_
timestamp 1727494699
transform 1 0 5050 0 -1 4950
box -6 -8 86 272
use NAND2X1  _1205_
timestamp 1727494699
transform 1 0 5470 0 1 4950
box -6 -8 86 272
use AOI22X1  _1206_
timestamp 1727487144
transform -1 0 5330 0 -1 4950
box -6 -8 126 272
use OAI22X1  _1207_
timestamp 1727495774
transform 1 0 5650 0 1 4430
box -6 -8 126 272
use OAI21X1  _1208_
timestamp 1727498925
transform -1 0 6050 0 1 4430
box -6 -8 106 272
use NAND3X1  _1209_
timestamp 1727494898
transform -1 0 5590 0 -1 4430
box -6 -8 106 272
use AOI21X1  _1210_
timestamp 1727487319
transform -1 0 5770 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1211_
timestamp 1727498925
transform 1 0 5470 0 1 3910
box -6 -8 106 272
use OAI21X1  _1212_
timestamp 1727498925
transform -1 0 5570 0 1 3390
box -6 -8 106 272
use NAND3X1  _1213_
timestamp 1727494898
transform 1 0 6170 0 1 3390
box -6 -8 106 272
use INVX1  _1214_
timestamp 1727493700
transform 1 0 6330 0 1 3390
box -6 -8 66 272
use AOI22X1  _1215_
timestamp 1727487144
transform -1 0 6030 0 -1 3390
box -6 -8 126 272
use OAI21X1  _1216_
timestamp 1727498925
transform 1 0 6090 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1217_
timestamp 1727494898
transform -1 0 6370 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1218_
timestamp 1727487319
transform 1 0 6350 0 -1 6510
box -6 -8 106 272
use NOR3X1  _1219_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727495302
transform -1 0 6350 0 1 1830
box -6 -8 186 272
use INVX1  _1220_
timestamp 1727493700
transform -1 0 4830 0 -1 4430
box -6 -8 66 272
use NAND3X1  _1221_
timestamp 1727494898
transform -1 0 5010 0 -1 4430
box -6 -8 106 272
use INVX1  _1222_
timestamp 1727493700
transform 1 0 6310 0 1 4950
box -6 -8 66 272
use NOR2X1  _1223_
timestamp 1727495070
transform -1 0 6430 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1224_
timestamp 1727495070
transform 1 0 6210 0 -1 4950
box -6 -8 86 272
use NAND2X1  _1225_
timestamp 1727494699
transform -1 0 6250 0 1 4950
box -6 -8 86 272
use NAND2X1  _1226_
timestamp 1727494699
transform 1 0 4790 0 1 4430
box -6 -8 86 272
use NOR2X1  _1227_
timestamp 1727495070
transform -1 0 5630 0 -1 4950
box -6 -8 86 272
use OAI21X1  _1228_
timestamp 1727498925
transform -1 0 6130 0 -1 4950
box -6 -8 106 272
use NAND3X1  _1229_
timestamp 1727494898
transform 1 0 5850 0 -1 4950
box -6 -8 106 272
use INVX1  _1230_
timestamp 1727493700
transform 1 0 5370 0 1 4430
box -6 -8 66 272
use INVX1  _1231_
timestamp 1727493700
transform -1 0 5130 0 -1 4430
box -6 -8 66 272
use OAI21X1  _1232_
timestamp 1727498925
transform 1 0 5210 0 -1 4430
box -6 -8 106 272
use NAND3X1  _1233_
timestamp 1727494898
transform -1 0 5310 0 1 4430
box -6 -8 106 272
use AOI21X1  _1234_
timestamp 1727487319
transform 1 0 6070 0 -1 3910
box -6 -8 106 272
use NOR3X1  _1235_
timestamp 1727495302
transform 1 0 6230 0 -1 3910
box -6 -8 186 272
use OAI21X1  _1236_
timestamp 1727498925
transform 1 0 6130 0 -1 2870
box -6 -8 106 272
use NAND3X1  _1237_
timestamp 1727494898
transform -1 0 6430 0 1 2870
box -6 -8 106 272
use NAND3X1  _1238_
timestamp 1727494898
transform -1 0 6270 0 1 2870
box -6 -8 106 272
use NAND3X1  _1239_
timestamp 1727494898
transform 1 0 5950 0 -1 2870
box -6 -8 106 272
use INVX1  _1240_
timestamp 1727493700
transform 1 0 5910 0 1 2350
box -6 -8 66 272
use OAI21X1  _1241_
timestamp 1727498925
transform -1 0 6110 0 1 1830
box -6 -8 106 272
use AOI21X1  _1242_
timestamp 1727487319
transform 1 0 5850 0 1 1830
box -6 -8 106 272
use OAI21X1  _1243_
timestamp 1727498925
transform -1 0 5990 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1244_
timestamp 1727487319
transform -1 0 6050 0 -1 790
box -6 -8 106 272
use NAND2X1  _1245_
timestamp 1727494699
transform -1 0 5070 0 -1 270
box -6 -8 86 272
use OAI21X1  _1246_
timestamp 1727498925
transform -1 0 5470 0 1 270
box -6 -8 106 272
use NAND2X1  _1247_
timestamp 1727494699
transform 1 0 4430 0 1 790
box -6 -8 86 272
use INVX1  _1248_
timestamp 1727493700
transform -1 0 4290 0 -1 270
box -6 -8 66 272
use NOR2X1  _1249_
timestamp 1727495070
transform 1 0 4710 0 -1 1310
box -6 -8 86 272
use OAI21X1  _1250_
timestamp 1727498925
transform 1 0 3850 0 1 1310
box -6 -8 106 272
use NAND2X1  _1251_
timestamp 1727494699
transform 1 0 4850 0 -1 270
box -6 -8 86 272
use OR2X2  _1252_
timestamp 1727496117
transform -1 0 4610 0 -1 270
box -6 -8 106 272
use NAND3X1  _1253_
timestamp 1727494898
transform 1 0 4350 0 -1 270
box -6 -8 106 272
use AND2X2  _1254_
timestamp 1727487319
transform 1 0 5050 0 1 270
box -6 -8 106 273
use NOR2X1  _1255_
timestamp 1727495070
transform 1 0 4890 0 1 270
box -6 -8 86 272
use OAI21X1  _1256_
timestamp 1727498925
transform -1 0 4830 0 1 270
box -6 -8 106 272
use NAND2X1  _1257_
timestamp 1727494699
transform 1 0 4410 0 1 270
box -6 -8 86 272
use AOI21X1  _1258_
timestamp 1727487319
transform -1 0 4550 0 -1 790
box -6 -8 106 272
use NAND2X1  _1259_
timestamp 1727494699
transform 1 0 2610 0 1 2350
box -6 -8 86 272
use AND2X2  _1260_
timestamp 1727487319
transform -1 0 3310 0 1 2350
box -6 -8 106 273
use OAI21X1  _1261_
timestamp 1727498925
transform 1 0 3050 0 1 2350
box -6 -8 106 272
use AND2X2  _1262_
timestamp 1727487319
transform -1 0 3250 0 -1 2350
box -6 -8 106 273
use OAI21X1  _1263_
timestamp 1727498925
transform 1 0 2810 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1264_
timestamp 1727494898
transform 1 0 2890 0 1 2350
box -6 -8 106 272
use INVX1  _1265_
timestamp 1727493700
transform -1 0 2270 0 -1 2350
box -6 -8 66 272
use NAND2X1  _1266_
timestamp 1727494699
transform -1 0 3070 0 -1 2350
box -6 -8 86 272
use AOI22X1  _1267_
timestamp 1727487144
transform 1 0 3310 0 -1 2350
box -6 -8 126 272
use INVX1  _1268_
timestamp 1727493700
transform -1 0 2570 0 -1 2350
box -6 -8 66 272
use NAND3X1  _1269_
timestamp 1727494898
transform -1 0 2750 0 -1 2350
box -6 -8 106 272
use NAND2X1  _1270_
timestamp 1727494699
transform 1 0 2750 0 -1 1310
box -6 -8 86 272
use AOI21X1  _1271_
timestamp 1727487319
transform -1 0 3710 0 1 790
box -6 -8 106 272
use NAND2X1  _1272_
timestamp 1727494699
transform 1 0 2770 0 1 1830
box -6 -8 86 272
use INVX1  _1273_
timestamp 1727493700
transform -1 0 2890 0 1 1310
box -6 -8 66 272
use AOI22X1  _1274_
timestamp 1727487144
transform -1 0 3210 0 1 1830
box -6 -8 126 272
use AOI21X1  _1275_
timestamp 1727487319
transform 1 0 3090 0 1 1310
box -6 -8 106 272
use NAND2X1  _1276_
timestamp 1727494699
transform 1 0 3310 0 1 790
box -6 -8 86 272
use OAI21X1  _1277_
timestamp 1727498925
transform 1 0 3270 0 1 1310
box -6 -8 106 272
use INVX1  _1278_
timestamp 1727493700
transform 1 0 3310 0 -1 1830
box -6 -8 66 272
use OAI21X1  _1279_
timestamp 1727498925
transform -1 0 3530 0 -1 1830
box -6 -8 106 272
use NAND2X1  _1280_
timestamp 1727494699
transform -1 0 3110 0 -1 1310
box -6 -8 86 272
use NAND3X1  _1281_
timestamp 1727494898
transform 1 0 3150 0 1 790
box -6 -8 106 272
use AND2X2  _1282_
timestamp 1727487319
transform -1 0 3050 0 -1 790
box -6 -8 106 273
use NAND2X1  _1283_
timestamp 1727494699
transform 1 0 2890 0 -1 1310
box -6 -8 86 272
use NAND2X1  _1284_
timestamp 1727494699
transform 1 0 3470 0 1 790
box -6 -8 86 272
use NAND3X1  _1285_
timestamp 1727494898
transform 1 0 3470 0 -1 790
box -6 -8 106 272
use NAND3X1  _1286_
timestamp 1727494898
transform 1 0 3950 0 -1 790
box -6 -8 106 272
use OAI21X1  _1287_
timestamp 1727498925
transform -1 0 4370 0 -1 790
box -6 -8 106 272
use AOI22X1  _1288_
timestamp 1727487144
transform 1 0 3130 0 -1 790
box -6 -8 126 272
use AOI21X1  _1289_
timestamp 1727487319
transform -1 0 3070 0 1 790
box -6 -8 106 272
use OAI21X1  _1290_
timestamp 1727498925
transform 1 0 4110 0 -1 790
box -6 -8 106 272
use NAND3X1  _1291_
timestamp 1727494898
transform -1 0 3990 0 1 270
box -6 -8 106 272
use AND2X2  _1292_
timestamp 1727487319
transform 1 0 4570 0 1 270
box -6 -8 106 273
use NAND3X1  _1293_
timestamp 1727494898
transform 1 0 3790 0 -1 790
box -6 -8 106 272
use OAI21X1  _1294_
timestamp 1727498925
transform 1 0 3730 0 1 270
box -6 -8 106 272
use NAND3X1  _1295_
timestamp 1727494898
transform -1 0 3490 0 1 270
box -6 -8 106 272
use NAND3X1  _1296_
timestamp 1727494898
transform -1 0 3510 0 -1 270
box -6 -8 106 272
use AOI21X1  _1297_
timestamp 1727487319
transform -1 0 5310 0 1 270
box -6 -8 106 272
use AOI22X1  _1298_
timestamp 1727487144
transform -1 0 4350 0 1 270
box -6 -8 126 272
use AOI21X1  _1299_
timestamp 1727487319
transform 1 0 4070 0 1 270
box -6 -8 106 272
use OAI21X1  _1300_
timestamp 1727498925
transform -1 0 4010 0 -1 270
box -6 -8 106 272
use AOI21X1  _1301_
timestamp 1727487319
transform 1 0 2490 0 -1 270
box -6 -8 106 272
use INVX1  _1302_
timestamp 1727493700
transform -1 0 2710 0 -1 270
box -6 -8 66 272
use NAND3X1  _1303_
timestamp 1727494898
transform -1 0 3850 0 -1 270
box -6 -8 106 272
use OAI21X1  _1304_
timestamp 1727498925
transform 1 0 4070 0 -1 270
box -6 -8 106 272
use AOI21X1  _1305_
timestamp 1727487319
transform -1 0 2870 0 -1 270
box -6 -8 106 272
use OAI21X1  _1306_
timestamp 1727498925
transform 1 0 2630 0 1 270
box -6 -8 106 272
use OAI21X1  _1307_
timestamp 1727498925
transform -1 0 5950 0 1 270
box -6 -8 106 272
use NAND3X1  _1308_
timestamp 1727494898
transform 1 0 2930 0 -1 270
box -6 -8 106 272
use NAND3X1  _1309_
timestamp 1727494898
transform 1 0 2330 0 -1 270
box -6 -8 106 272
use NAND3X1  _1310_
timestamp 1727494898
transform -1 0 2910 0 1 270
box -6 -8 106 272
use AND2X2  _1311_
timestamp 1727487319
transform -1 0 2610 0 1 1310
box -6 -8 106 273
use NAND2X1  _1312_
timestamp 1727494699
transform -1 0 2470 0 -1 1830
box -6 -8 86 272
use NAND3X1  _1313_
timestamp 1727494898
transform -1 0 6330 0 -1 1830
box -6 -8 106 272
use INVX1  _1314_
timestamp 1727493700
transform -1 0 6430 0 1 2350
box -6 -8 66 272
use NAND2X1  _1315_
timestamp 1727494699
transform 1 0 6410 0 1 1830
box -6 -8 86 272
use NAND3X1  _1316_
timestamp 1727494898
transform -1 0 6410 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1317_
timestamp 1727494898
transform -1 0 6070 0 -1 2350
box -6 -8 106 272
use AOI21X1  _1318_
timestamp 1727487319
transform 1 0 6150 0 -1 2350
box -6 -8 106 272
use OAI21X1  _1319_
timestamp 1727498925
transform -1 0 5750 0 -1 2350
box -6 -8 106 272
use AOI21X1  _1320_
timestamp 1727487319
transform -1 0 5630 0 1 1830
box -6 -8 106 272
use NAND2X1  _1321_
timestamp 1727494699
transform 1 0 2610 0 -1 1310
box -6 -8 86 272
use NAND2X1  _1322_
timestamp 1727494699
transform 1 0 2890 0 -1 1830
box -6 -8 86 272
use AND2X2  _1323_
timestamp 1727487319
transform -1 0 2550 0 1 1830
box -6 -8 106 273
use NOR2X1  _1324_
timestamp 1727495070
transform -1 0 2890 0 1 4950
box -6 -8 86 272
use NOR2X1  _1325_
timestamp 1727495070
transform -1 0 3050 0 1 4950
box -6 -8 86 272
use OAI21X1  _1326_
timestamp 1727498925
transform 1 0 2770 0 -1 4950
box -6 -8 106 272
use AOI21X1  _1327_
timestamp 1727487319
transform -1 0 3650 0 -1 4950
box -6 -8 106 272
use OAI21X1  _1328_
timestamp 1727498925
transform 1 0 2870 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1329_
timestamp 1727498925
transform -1 0 3050 0 -1 4950
box -6 -8 106 272
use NAND2X1  _1330_
timestamp 1727494699
transform 1 0 2850 0 1 4430
box -6 -8 86 272
use OAI21X1  _1331_
timestamp 1727498925
transform 1 0 2690 0 1 4430
box -6 -8 106 272
use INVX1  _1332_
timestamp 1727493700
transform 1 0 2230 0 -1 4430
box -6 -8 66 272
use INVX1  _1333_
timestamp 1727493700
transform 1 0 2090 0 -1 3910
box -6 -8 66 272
use OAI21X1  _1334_
timestamp 1727498925
transform -1 0 2630 0 -1 3910
box -6 -8 106 272
use OAI21X1  _1335_
timestamp 1727498925
transform 1 0 2210 0 -1 3910
box -6 -8 106 272
use AOI21X1  _1336_
timestamp 1727487319
transform -1 0 3670 0 -1 270
box -6 -8 106 272
use OAI21X1  _1337_
timestamp 1727498925
transform 1 0 3110 0 -1 270
box -6 -8 106 272
use OAI21X1  _1338_
timestamp 1727498925
transform -1 0 4770 0 -1 270
box -6 -8 106 272
use AOI21X1  _1339_
timestamp 1727487319
transform -1 0 3730 0 -1 790
box -6 -8 106 272
use OAI21X1  _1340_
timestamp 1727498925
transform -1 0 3670 0 1 270
box -6 -8 106 272
use NAND2X1  _1341_
timestamp 1727494699
transform -1 0 2910 0 1 790
box -6 -8 86 272
use INVX1  _1342_
timestamp 1727493700
transform -1 0 2770 0 1 790
box -6 -8 66 272
use NOR2X1  _1343_
timestamp 1727495070
transform -1 0 3110 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1344_
timestamp 1727498925
transform -1 0 2450 0 -1 2350
box -6 -8 106 272
use NAND2X1  _1345_
timestamp 1727494699
transform -1 0 2450 0 1 1310
box -6 -8 86 272
use OR2X2  _1346_
timestamp 1727496117
transform 1 0 2270 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1347_
timestamp 1727494898
transform -1 0 2650 0 1 790
box -6 -8 106 272
use AND2X2  _1348_
timestamp 1727487319
transform -1 0 2070 0 -1 1310
box -6 -8 106 273
use NOR2X1  _1349_
timestamp 1727495070
transform -1 0 2210 0 -1 1310
box -6 -8 86 272
use OAI21X1  _1350_
timestamp 1727498925
transform 1 0 2230 0 1 790
box -6 -8 106 272
use NAND2X1  _1351_
timestamp 1727494699
transform 1 0 2090 0 1 790
box -6 -8 86 272
use NOR2X1  _1352_
timestamp 1727495070
transform 1 0 3330 0 -1 790
box -6 -8 86 272
use AOI21X1  _1353_
timestamp 1727487319
transform -1 0 2890 0 -1 790
box -6 -8 106 272
use NAND2X1  _1354_
timestamp 1727494699
transform -1 0 1610 0 1 2350
box -6 -8 86 272
use INVX1  _1355_
timestamp 1727493700
transform -1 0 1370 0 -1 2350
box -6 -8 66 272
use AND2X2  _1356_
timestamp 1727487319
transform 1 0 1850 0 1 2350
box -6 -8 106 273
use AND2X2  _1357_
timestamp 1727487319
transform -1 0 2250 0 1 2350
box -6 -8 106 273
use NAND2X1  _1358_
timestamp 1727494699
transform 1 0 2010 0 1 2350
box -6 -8 86 272
use AOI22X1  _1359_
timestamp 1727487144
transform 1 0 1350 0 1 2350
box -6 -8 126 272
use INVX1  _1360_
timestamp 1727493700
transform -1 0 1030 0 1 1830
box -6 -8 66 272
use AOI21X1  _1361_
timestamp 1727487319
transform 1 0 1250 0 1 1830
box -6 -8 106 272
use INVX2  _1362_
timestamp 1727493898
transform 1 0 1350 0 1 2870
box -6 -8 66 272
use OAI21X1  _1363_
timestamp 1727498925
transform 1 0 1690 0 1 2350
box -6 -8 106 272
use OAI21X1  _1364_
timestamp 1727498925
transform -1 0 2550 0 1 2350
box -6 -8 106 272
use AOI21X1  _1365_
timestamp 1727487319
transform -1 0 1530 0 -1 2350
box -6 -8 106 272
use OAI22X1  _1366_
timestamp 1727495774
transform -1 0 1510 0 -1 1830
box -6 -8 126 272
use NAND3X1  _1367_
timestamp 1727494898
transform 1 0 1610 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1368_
timestamp 1727494898
transform -1 0 1190 0 1 1830
box -6 -8 106 272
use NOR2X1  _1369_
timestamp 1727495070
transform 1 0 1590 0 1 1830
box -6 -8 86 272
use NAND3X1  _1370_
timestamp 1727494898
transform -1 0 1530 0 1 1830
box -6 -8 106 272
use NAND2X1  _1371_
timestamp 1727494699
transform -1 0 1550 0 1 790
box -6 -8 86 272
use NOR2X1  _1372_
timestamp 1727495070
transform 1 0 2190 0 -1 790
box -6 -8 86 272
use NOR2X1  _1373_
timestamp 1727495070
transform 1 0 2950 0 1 1310
box -6 -8 86 272
use OAI21X1  _1374_
timestamp 1727498925
transform 1 0 2450 0 -1 1310
box -6 -8 106 272
use AOI21X1  _1375_
timestamp 1727487319
transform 1 0 1790 0 -1 1310
box -6 -8 106 272
use OAI21X1  _1376_
timestamp 1727498925
transform 1 0 1870 0 -1 790
box -6 -8 106 272
use AND2X2  _1377_
timestamp 1727487319
transform -1 0 2030 0 1 790
box -6 -8 106 273
use NAND3X1  _1378_
timestamp 1727494898
transform 1 0 1630 0 -1 1310
box -6 -8 106 272
use NAND2X1  _1379_
timestamp 1727494699
transform 1 0 1610 0 1 790
box -6 -8 86 272
use NAND3X1  _1380_
timestamp 1727494898
transform -1 0 1590 0 1 270
box -6 -8 106 272
use NAND3X1  _1381_
timestamp 1727494898
transform -1 0 1010 0 -1 270
box -6 -8 106 272
use NOR3X1  _1382_
timestamp 1727495302
transform -1 0 3310 0 1 270
box -6 -8 186 272
use AOI21X1  _1383_
timestamp 1727487319
transform -1 0 3070 0 1 270
box -6 -8 106 272
use AOI21X1  _1384_
timestamp 1727487319
transform 1 0 1650 0 1 270
box -6 -8 106 272
use NAND3X1  _1385_
timestamp 1727494898
transform 1 0 1770 0 1 790
box -6 -8 106 272
use OAI21X1  _1386_
timestamp 1727498925
transform -1 0 2730 0 -1 790
box -6 -8 106 272
use AOI21X1  _1387_
timestamp 1727487319
transform 1 0 2030 0 -1 790
box -6 -8 106 272
use OAI21X1  _1388_
timestamp 1727498925
transform -1 0 1430 0 1 270
box -6 -8 106 272
use NAND3X1  _1389_
timestamp 1727494898
transform -1 0 1310 0 -1 270
box -6 -8 106 272
use INVX1  _1390_
timestamp 1727493700
transform -1 0 1130 0 -1 270
box -6 -8 66 272
use NAND3X1  _1391_
timestamp 1727494898
transform 1 0 1170 0 1 270
box -6 -8 106 272
use OAI21X1  _1392_
timestamp 1727498925
transform 1 0 1810 0 1 270
box -6 -8 106 272
use NAND3X1  _1393_
timestamp 1727494898
transform 1 0 1550 0 -1 270
box -6 -8 106 272
use AOI21X1  _1394_
timestamp 1727487319
transform 1 0 1890 0 -1 270
box -6 -8 106 272
use NAND3X1  _1395_
timestamp 1727494898
transform 1 0 1370 0 -1 270
box -6 -8 106 272
use NAND3X1  _1396_
timestamp 1727494898
transform 1 0 1990 0 1 270
box -6 -8 106 272
use AOI22X1  _1397_
timestamp 1727487144
transform -1 0 2430 0 1 270
box -6 -8 126 272
use NOR2X1  _1398_
timestamp 1727495070
transform 1 0 2490 0 1 270
box -6 -8 86 272
use AOI21X1  _1399_
timestamp 1727487319
transform 1 0 2530 0 -1 1830
box -6 -8 106 272
use OAI21X1  _1400_
timestamp 1727498925
transform -1 0 2810 0 -1 1830
box -6 -8 106 272
use INVX1  _1401_
timestamp 1727493700
transform -1 0 2110 0 -1 270
box -6 -8 66 272
use AOI21X1  _1402_
timestamp 1727487319
transform -1 0 2270 0 -1 270
box -6 -8 106 272
use NAND3X1  _1403_
timestamp 1727494898
transform 1 0 2150 0 1 270
box -6 -8 106 272
use NAND3X1  _1404_
timestamp 1727494898
transform 1 0 1730 0 -1 270
box -6 -8 106 272
use NAND2X1  _1405_
timestamp 1727494699
transform 1 0 2490 0 -1 790
box -6 -8 86 272
use OAI21X1  _1406_
timestamp 1727498925
transform -1 0 2710 0 1 1830
box -6 -8 106 272
use OAI21X1  _1407_
timestamp 1727498925
transform -1 0 2670 0 -1 2870
box -6 -8 106 272
use AND2X2  _1408_
timestamp 1727487319
transform -1 0 4990 0 -1 4950
box -6 -8 106 273
use NAND2X1  _1409_
timestamp 1727494699
transform 1 0 4350 0 1 4950
box -6 -8 86 272
use OAI21X1  _1410_
timestamp 1727498925
transform -1 0 4810 0 -1 4950
box -6 -8 106 272
use OAI21X1  _1411_
timestamp 1727498925
transform -1 0 4650 0 -1 4950
box -6 -8 106 272
use AOI21X1  _1412_
timestamp 1727487319
transform -1 0 3350 0 1 4430
box -6 -8 106 272
use AOI22X1  _1413_
timestamp 1727487144
transform 1 0 2590 0 -1 4430
box -6 -8 126 272
use OAI21X1  _1414_
timestamp 1727498925
transform -1 0 5410 0 1 4950
box -6 -8 106 272
use NAND3X1  _1415_
timestamp 1727494898
transform -1 0 2330 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1416_
timestamp 1727487319
transform -1 0 2430 0 -1 790
box -6 -8 106 272
use INVX1  _1417_
timestamp 1727493700
transform 1 0 1890 0 1 1310
box -6 -8 66 272
use OAI21X1  _1418_
timestamp 1727498925
transform 1 0 2390 0 1 790
box -6 -8 106 272
use INVX1  _1419_
timestamp 1727493700
transform -1 0 1410 0 1 790
box -6 -8 66 272
use AOI21X1  _1420_
timestamp 1727487319
transform -1 0 1630 0 -1 790
box -6 -8 106 272
use NAND2X1  _1421_
timestamp 1727494699
transform -1 0 1030 0 -1 1830
box -6 -8 86 272
use INVX1  _1422_
timestamp 1727493700
transform 1 0 1050 0 1 1310
box -6 -8 66 272
use NOR2X1  _1423_
timestamp 1727495070
transform -1 0 770 0 1 1830
box -6 -8 86 272
use OAI21X1  _1424_
timestamp 1727498925
transform -1 0 1230 0 -1 2350
box -6 -8 106 272
use NAND2X1  _1425_
timestamp 1727494699
transform -1 0 550 0 -1 1830
box -6 -8 86 272
use OR2X2  _1426_
timestamp 1727496117
transform 1 0 790 0 -1 1830
box -6 -8 106 272
use NAND3X1  _1427_
timestamp 1727494898
transform -1 0 990 0 1 1310
box -6 -8 106 272
use AND2X2  _1428_
timestamp 1727487319
transform 1 0 610 0 -1 1830
box -6 -8 106 273
use NOR2X1  _1429_
timestamp 1727495070
transform -1 0 410 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1430_
timestamp 1727498925
transform 1 0 730 0 1 1310
box -6 -8 106 272
use NAND2X1  _1431_
timestamp 1727494699
transform 1 0 870 0 1 790
box -6 -8 86 272
use NAND2X1  _1432_
timestamp 1727494699
transform 1 0 1590 0 1 1310
box -6 -8 86 272
use NAND2X1  _1433_
timestamp 1727494699
transform -1 0 910 0 1 1830
box -6 -8 86 272
use INVX1  _1434_
timestamp 1727493700
transform -1 0 450 0 1 1830
box -6 -8 66 272
use NAND2X1  _1435_
timestamp 1727494699
transform -1 0 1070 0 -1 2350
box -6 -8 86 272
use NAND2X1  _1436_
timestamp 1727494699
transform 1 0 1010 0 1 2350
box -6 -8 86 272
use NOR2X1  _1437_
timestamp 1727495070
transform 1 0 850 0 -1 2350
box -6 -8 86 272
use INVX1  _1438_
timestamp 1727493700
transform -1 0 290 0 -1 2350
box -6 -8 66 272
use AOI22X1  _1439_
timestamp 1727487144
transform 1 0 1150 0 1 2350
box -6 -8 126 272
use INVX1  _1440_
timestamp 1727493700
transform -1 0 130 0 1 1830
box -6 -8 66 272
use NAND3X1  _1441_
timestamp 1727494898
transform -1 0 310 0 1 1830
box -6 -8 106 272
use OAI21X1  _1442_
timestamp 1727498925
transform -1 0 610 0 1 1830
box -6 -8 106 272
use NAND2X1  _1443_
timestamp 1727494699
transform -1 0 470 0 1 790
box -6 -8 86 272
use AOI21X1  _1444_
timestamp 1727487319
transform -1 0 630 0 1 790
box -6 -8 106 272
use NAND3X1  _1445_
timestamp 1727494898
transform -1 0 810 0 1 790
box -6 -8 106 272
use INVX1  _1446_
timestamp 1727493700
transform -1 0 130 0 -1 790
box -6 -8 66 272
use OAI21X1  _1447_
timestamp 1727498925
transform 1 0 350 0 -1 790
box -6 -8 106 272
use AND2X2  _1448_
timestamp 1727487319
transform -1 0 790 0 -1 1310
box -6 -8 106 273
use NAND2X1  _1449_
timestamp 1727494699
transform 1 0 1030 0 1 790
box -6 -8 86 272
use NAND3X1  _1450_
timestamp 1727494898
transform -1 0 330 0 1 790
box -6 -8 106 272
use NAND3X1  _1451_
timestamp 1727494898
transform 1 0 510 0 -1 790
box -6 -8 106 272
use NAND3X1  _1452_
timestamp 1727494898
transform 1 0 850 0 -1 790
box -6 -8 106 272
use OAI21X1  _1453_
timestamp 1727498925
transform -1 0 1810 0 -1 790
box -6 -8 106 272
use AOI22X1  _1454_
timestamp 1727487144
transform -1 0 790 0 -1 790
box -6 -8 126 272
use OR2X2  _1455_
timestamp 1727496117
transform 1 0 230 0 1 270
box -6 -8 106 272
use NAND2X1  _1456_
timestamp 1727494699
transform -1 0 170 0 1 270
box -6 -8 86 272
use AOI21X1  _1457_
timestamp 1727487319
transform 1 0 390 0 1 270
box -6 -8 106 272
use OAI21X1  _1458_
timestamp 1727498925
transform 1 0 710 0 1 270
box -6 -8 106 272
use NAND3X1  _1459_
timestamp 1727494898
transform -1 0 650 0 1 270
box -6 -8 106 272
use NAND3X1  _1460_
timestamp 1727494898
transform 1 0 1210 0 -1 790
box -6 -8 106 272
use OAI21X1  _1461_
timestamp 1727498925
transform 1 0 870 0 1 270
box -6 -8 106 272
use NAND3X1  _1462_
timestamp 1727494898
transform -1 0 1470 0 -1 790
box -6 -8 106 272
use NAND2X1  _1463_
timestamp 1727494699
transform -1 0 150 0 -1 270
box -6 -8 86 272
use NAND3X1  _1464_
timestamp 1727494898
transform -1 0 330 0 -1 270
box -6 -8 106 272
use AOI21X1  _1465_
timestamp 1727487319
transform -1 0 830 0 -1 270
box -6 -8 106 272
use OAI21X1  _1466_
timestamp 1727498925
transform -1 0 670 0 -1 270
box -6 -8 106 272
use NAND3X1  _1467_
timestamp 1727494898
transform 1 0 410 0 -1 270
box -6 -8 106 272
use NAND2X1  _1468_
timestamp 1727494699
transform -1 0 1110 0 1 270
box -6 -8 86 272
use AOI21X1  _1469_
timestamp 1727487319
transform -1 0 1670 0 -1 1830
box -6 -8 106 272
use NAND2X1  _1470_
timestamp 1727494699
transform -1 0 2150 0 -1 1830
box -6 -8 86 272
use OAI21X1  _1471_
timestamp 1727498925
transform -1 0 2010 0 -1 1830
box -6 -8 106 272
use INVX1  _1472_
timestamp 1727493700
transform -1 0 1150 0 -1 1830
box -6 -8 66 272
use NOR2X1  _1473_
timestamp 1727495070
transform 1 0 2150 0 1 1830
box -6 -8 86 272
use OAI21X1  _1474_
timestamp 1727498925
transform 1 0 2290 0 1 1830
box -6 -8 106 272
use NOR2X1  _1475_
timestamp 1727495070
transform -1 0 2710 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1476_
timestamp 1727495070
transform 1 0 3110 0 -1 4950
box -6 -8 86 272
use AOI21X1  _1477_
timestamp 1727487319
transform -1 0 5790 0 -1 4950
box -6 -8 106 272
use OAI21X1  _1478_
timestamp 1727498925
transform -1 0 5490 0 -1 4950
box -6 -8 106 272
use NOR2X1  _1479_
timestamp 1727495070
transform -1 0 2310 0 -1 6510
box -6 -8 86 272
use NOR2X1  _1480_
timestamp 1727495070
transform 1 0 3230 0 -1 5470
box -6 -8 86 272
use AOI22X1  _1481_
timestamp 1727487144
transform -1 0 3370 0 -1 4950
box -6 -8 126 272
use OAI21X1  _1482_
timestamp 1727498925
transform 1 0 4130 0 -1 4950
box -6 -8 106 272
use INVX1  _1483_
timestamp 1727493700
transform 1 0 3570 0 -1 2870
box -6 -8 66 272
use INVX1  _1484_
timestamp 1727493700
transform 1 0 1210 0 1 3910
box -6 -8 66 272
use OAI21X1  _1485_
timestamp 1727498925
transform 1 0 2370 0 -1 3910
box -6 -8 106 272
use INVX1  _1486_
timestamp 1727493700
transform 1 0 1470 0 1 1310
box -6 -8 66 272
use OAI21X1  _1487_
timestamp 1727498925
transform -1 0 650 0 1 1310
box -6 -8 106 272
use INVX1  _1488_
timestamp 1727493700
transform 1 0 570 0 -1 1310
box -6 -8 66 272
use AOI21X1  _1489_
timestamp 1727487319
transform -1 0 170 0 1 790
box -6 -8 106 272
use NAND2X1  _1490_
timestamp 1727494699
transform -1 0 1590 0 -1 2870
box -6 -8 86 272
use INVX1  _1491_
timestamp 1727493700
transform 1 0 950 0 -1 2870
box -6 -8 66 272
use NOR2X1  _1492_
timestamp 1727495070
transform -1 0 950 0 1 2350
box -6 -8 86 272
use OAI22X1  _1493_
timestamp 1727495774
transform -1 0 790 0 -1 2350
box -6 -8 126 272
use NAND2X1  _1494_
timestamp 1727494699
transform -1 0 610 0 -1 2350
box -6 -8 86 272
use OR2X2  _1495_
timestamp 1727496117
transform -1 0 450 0 -1 2350
box -6 -8 106 272
use NAND3X1  _1496_
timestamp 1727494898
transform -1 0 510 0 1 2350
box -6 -8 106 272
use INVX2  _1497_
timestamp 1727493898
transform 1 0 1150 0 -1 3390
box -6 -8 66 272
use NAND2X1  _1498_
timestamp 1727494699
transform -1 0 650 0 1 2350
box -6 -8 86 272
use OAI21X1  _1499_
timestamp 1727498925
transform 1 0 710 0 1 2350
box -6 -8 106 272
use NAND2X1  _1500_
timestamp 1727494699
transform 1 0 1190 0 -1 3910
box -6 -8 86 272
use NAND2X1  _1501_
timestamp 1727494699
transform 1 0 1350 0 -1 3910
box -6 -8 86 272
use NOR2X1  _1502_
timestamp 1727495070
transform -1 0 1150 0 1 3910
box -6 -8 86 272
use INVX1  _1503_
timestamp 1727493700
transform -1 0 710 0 1 3910
box -6 -8 66 272
use INVX1  _1504_
timestamp 1727493700
transform 1 0 930 0 1 2870
box -6 -8 66 272
use OAI21X1  _1505_
timestamp 1727498925
transform -1 0 870 0 1 2870
box -6 -8 106 272
use AND2X2  _1506_
timestamp 1727487319
transform -1 0 690 0 1 2870
box -6 -8 106 273
use AOI21X1  _1507_
timestamp 1727487319
transform -1 0 350 0 1 2350
box -6 -8 106 272
use INVX1  _1508_
timestamp 1727493700
transform -1 0 130 0 -1 1830
box -6 -8 66 272
use NAND3X1  _1509_
timestamp 1727494898
transform -1 0 190 0 1 2350
box -6 -8 106 272
use NAND3X1  _1510_
timestamp 1727494898
transform 1 0 70 0 1 1310
box -6 -8 106 272
use OAI21X1  _1511_
timestamp 1727498925
transform -1 0 290 0 -1 790
box -6 -8 106 272
use INVX1  _1512_
timestamp 1727493700
transform -1 0 150 0 -1 2350
box -6 -8 66 272
use OAI21X1  _1513_
timestamp 1727498925
transform 1 0 250 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1514_
timestamp 1727494898
transform -1 0 510 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1515_
timestamp 1727494898
transform 1 0 230 0 1 1310
box -6 -8 106 272
use OAI21X1  _1516_
timestamp 1727498925
transform -1 0 190 0 -1 1310
box -6 -8 106 272
use NAND3X1  _1517_
timestamp 1727494898
transform -1 0 490 0 1 1310
box -6 -8 106 272
use NAND2X1  _1518_
timestamp 1727494699
transform -1 0 930 0 -1 1310
box -6 -8 86 272
use NAND3X1  _1519_
timestamp 1727494898
transform -1 0 1250 0 -1 1310
box -6 -8 106 272
use AOI21X1  _1520_
timestamp 1727487319
transform 1 0 1030 0 -1 790
box -6 -8 106 272
use OAI21X1  _1521_
timestamp 1727498925
transform 1 0 1170 0 1 790
box -6 -8 106 272
use NAND3X1  _1522_
timestamp 1727494898
transform 1 0 990 0 -1 1310
box -6 -8 106 272
use NAND2X1  _1523_
timestamp 1727494699
transform -1 0 1390 0 1 1310
box -6 -8 86 272
use NOR3X1  _1524_
timestamp 1727495302
transform 1 0 1750 0 1 1830
box -6 -8 186 272
use AOI21X1  _1525_
timestamp 1727487319
transform 1 0 1990 0 1 1830
box -6 -8 106 272
use INVX1  _1526_
timestamp 1727493700
transform -1 0 1970 0 -1 2350
box -6 -8 66 272
use OAI21X1  _1527_
timestamp 1727498925
transform 1 0 2050 0 -1 2350
box -6 -8 106 272
use OAI21X1  _1528_
timestamp 1727498925
transform 1 0 2730 0 -1 2870
box -6 -8 106 272
use NAND2X1  _1529_
timestamp 1727494699
transform -1 0 5150 0 1 4430
box -6 -8 86 272
use NAND2X1  _1530_
timestamp 1727494699
transform -1 0 5010 0 1 4430
box -6 -8 86 272
use NAND2X1  _1531_
timestamp 1727494699
transform -1 0 4710 0 -1 4430
box -6 -8 86 272
use NAND2X1  _1532_
timestamp 1727494699
transform 1 0 3110 0 1 4950
box -6 -8 86 272
use OAI21X1  _1533_
timestamp 1727498925
transform -1 0 3430 0 -1 4430
box -6 -8 106 272
use AOI21X1  _1534_
timestamp 1727487319
transform 1 0 3490 0 -1 3390
box -6 -8 106 272
use AOI22X1  _1535_
timestamp 1727487144
transform -1 0 3270 0 -1 2870
box -6 -8 126 272
use INVX1  _1536_
timestamp 1727493700
transform 1 0 3510 0 1 2870
box -6 -8 66 272
use NAND2X1  _1537_
timestamp 1727494699
transform -1 0 270 0 -1 1830
box -6 -8 86 272
use INVX1  _1538_
timestamp 1727493700
transform 1 0 1210 0 -1 2870
box -6 -8 66 272
use OAI21X1  _1539_
timestamp 1727498925
transform -1 0 890 0 -1 2870
box -6 -8 106 272
use INVX1  _1540_
timestamp 1727493700
transform -1 0 710 0 -1 2870
box -6 -8 66 272
use INVX1  _1541_
timestamp 1727493700
transform 1 0 1010 0 -1 3390
box -6 -8 66 272
use NOR2X1  _1542_
timestamp 1727495070
transform 1 0 1050 0 -1 3910
box -6 -8 86 272
use NOR2X1  _1543_
timestamp 1727495070
transform 1 0 870 0 -1 3390
box -6 -8 86 272
use NOR2X1  _1544_
timestamp 1727495070
transform 1 0 930 0 1 3910
box -6 -8 86 272
use AOI21X1  _1545_
timestamp 1727487319
transform -1 0 870 0 1 3910
box -6 -8 106 272
use NAND2X1  _1546_
timestamp 1727494699
transform 1 0 510 0 1 3910
box -6 -8 86 272
use NOR2X1  _1547_
timestamp 1727495070
transform -1 0 790 0 -1 3910
box -6 -8 86 272
use OAI22X1  _1548_
timestamp 1727495774
transform -1 0 970 0 -1 3910
box -6 -8 126 272
use NAND2X1  _1549_
timestamp 1727494699
transform 1 0 350 0 1 3910
box -6 -8 86 272
use OAI21X1  _1550_
timestamp 1727498925
transform -1 0 810 0 -1 3390
box -6 -8 106 272
use INVX1  _1551_
timestamp 1727493700
transform -1 0 130 0 1 3910
box -6 -8 66 272
use NAND3X1  _1552_
timestamp 1727494898
transform 1 0 190 0 1 3910
box -6 -8 106 272
use NAND2X1  _1553_
timestamp 1727494699
transform 1 0 90 0 -1 3390
box -6 -8 86 272
use NOR2X1  _1554_
timestamp 1727495070
transform -1 0 150 0 -1 2870
box -6 -8 86 272
use AOI21X1  _1555_
timestamp 1727487319
transform 1 0 230 0 -1 3390
box -6 -8 106 272
use OAI21X1  _1556_
timestamp 1727498925
transform 1 0 330 0 -1 2870
box -6 -8 106 272
use OR2X2  _1557_
timestamp 1727496117
transform 1 0 90 0 1 2870
box -6 -8 106 272
use INVX1  _1558_
timestamp 1727493700
transform -1 0 270 0 -1 2870
box -6 -8 66 272
use NAND3X1  _1559_
timestamp 1727494898
transform -1 0 590 0 -1 2870
box -6 -8 106 272
use NAND2X1  _1560_
timestamp 1727494699
transform 1 0 1070 0 -1 2870
box -6 -8 86 272
use NAND2X1  _1561_
timestamp 1727494699
transform 1 0 1350 0 -1 2870
box -6 -8 86 272
use NAND3X1  _1562_
timestamp 1727494898
transform 1 0 1050 0 1 2870
box -6 -8 106 272
use NAND2X1  _1563_
timestamp 1727494699
transform -1 0 1550 0 1 2870
box -6 -8 86 272
use NOR2X1  _1564_
timestamp 1727495070
transform 1 0 2670 0 1 1310
box -6 -8 86 272
use NOR2X1  _1565_
timestamp 1727495070
transform -1 0 1550 0 -1 1310
box -6 -8 86 272
use NAND3X1  _1566_
timestamp 1727494898
transform 1 0 2210 0 1 1310
box -6 -8 106 272
use NAND2X1  _1567_
timestamp 1727494699
transform 1 0 1310 0 -1 1310
box -6 -8 86 272
use AOI22X1  _1568_
timestamp 1727487144
transform 1 0 2030 0 1 1310
box -6 -8 126 272
use AOI21X1  _1569_
timestamp 1727487319
transform 1 0 2290 0 -1 2870
box -6 -8 106 272
use INVX1  _1570_
timestamp 1727493700
transform 1 0 2450 0 -1 2870
box -6 -8 66 272
use NAND2X1  _1571_
timestamp 1727494699
transform -1 0 1250 0 1 1310
box -6 -8 86 272
use OAI21X1  _1572_
timestamp 1727498925
transform -1 0 1330 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1573_
timestamp 1727487319
transform -1 0 1830 0 1 1310
box -6 -8 106 272
use OAI21X1  _1574_
timestamp 1727498925
transform -1 0 1830 0 -1 1830
box -6 -8 106 272
use AOI21X1  _1575_
timestamp 1727487319
transform 1 0 2130 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1576_
timestamp 1727498925
transform 1 0 2410 0 1 2870
box -6 -8 106 272
use OR2X2  _1577_
timestamp 1727496117
transform -1 0 1870 0 -1 3910
box -6 -8 106 272
use NAND3X1  _1578_
timestamp 1727494898
transform 1 0 2550 0 1 3390
box -6 -8 106 272
use INVX1  _1579_
timestamp 1727493700
transform 1 0 6430 0 1 3910
box -6 -8 66 272
use OAI21X1  _1580_
timestamp 1727498925
transform 1 0 6270 0 1 3910
box -6 -8 106 272
use NAND2X1  _1581_
timestamp 1727494699
transform 1 0 6110 0 1 3910
box -6 -8 86 272
use NAND2X1  _1582_
timestamp 1727494699
transform 1 0 2990 0 1 4430
box -6 -8 86 272
use OAI21X1  _1583_
timestamp 1727498925
transform -1 0 3130 0 1 3910
box -6 -8 106 272
use AOI21X1  _1584_
timestamp 1727487319
transform 1 0 3250 0 1 3390
box -6 -8 106 272
use AOI22X1  _1585_
timestamp 1727487144
transform -1 0 3430 0 -1 3390
box -6 -8 126 272
use INVX1  _1586_
timestamp 1727493700
transform 1 0 2910 0 1 2870
box -6 -8 66 272
use AOI21X1  _1587_
timestamp 1727487319
transform -1 0 650 0 -1 3910
box -6 -8 106 272
use NOR2X1  _1588_
timestamp 1727495070
transform 1 0 1030 0 1 3390
box -6 -8 86 272
use NAND2X1  _1589_
timestamp 1727494699
transform 1 0 890 0 1 3390
box -6 -8 86 272
use OAI22X1  _1590_
timestamp 1727495774
transform 1 0 710 0 1 3390
box -6 -8 126 272
use NAND2X1  _1591_
timestamp 1727494699
transform -1 0 650 0 1 3390
box -6 -8 86 272
use OR2X2  _1592_
timestamp 1727496117
transform 1 0 70 0 1 3390
box -6 -8 106 272
use OAI21X1  _1593_
timestamp 1727498925
transform -1 0 170 0 -1 3910
box -6 -8 106 272
use NAND2X1  _1594_
timestamp 1727494699
transform 1 0 230 0 -1 3910
box -6 -8 86 272
use NAND2X1  _1595_
timestamp 1727494699
transform -1 0 330 0 1 3390
box -6 -8 86 272
use OR2X2  _1596_
timestamp 1727496117
transform 1 0 390 0 1 3390
box -6 -8 106 272
use NAND2X1  _1597_
timestamp 1727494699
transform 1 0 390 0 -1 3390
box -6 -8 86 272
use NAND3X1  _1598_
timestamp 1727494898
transform -1 0 530 0 1 2870
box -6 -8 106 272
use OAI21X1  _1599_
timestamp 1727498925
transform -1 0 350 0 1 2870
box -6 -8 106 272
use NAND3X1  _1600_
timestamp 1727494898
transform 1 0 530 0 -1 3390
box -6 -8 106 272
use NAND2X1  _1601_
timestamp 1727494699
transform 1 0 1210 0 1 2870
box -6 -8 86 272
use NOR2X1  _1602_
timestamp 1727495070
transform -1 0 1750 0 -1 2870
box -6 -8 86 272
use NAND3X1  _1603_
timestamp 1727494898
transform 1 0 1810 0 -1 2870
box -6 -8 106 272
use NAND3X1  _1604_
timestamp 1727494898
transform -1 0 2070 0 -1 2870
box -6 -8 106 272
use NAND3X1  _1605_
timestamp 1727494898
transform 1 0 1610 0 1 2870
box -6 -8 106 272
use INVX1  _1606_
timestamp 1727493700
transform 1 0 2290 0 1 3390
box -6 -8 66 272
use OR2X2  _1607_
timestamp 1727496117
transform 1 0 1450 0 -1 3390
box -6 -8 106 272
use AND2X2  _1608_
timestamp 1727487319
transform 1 0 1610 0 -1 3390
box -6 -8 106 273
use NAND3X1  _1609_
timestamp 1727494898
transform 1 0 1770 0 1 2870
box -6 -8 106 272
use AOI21X1  _1610_
timestamp 1727487319
transform -1 0 5870 0 -1 2870
box -6 -8 106 272
use OAI21X1  _1611_
timestamp 1727498925
transform -1 0 5690 0 -1 2870
box -6 -8 106 272
use INVX1  _1612_
timestamp 1727493700
transform 1 0 810 0 -1 4430
box -6 -8 66 272
use AOI21X1  _1613_
timestamp 1727487319
transform 1 0 2550 0 1 3910
box -6 -8 106 272
use AOI21X1  _1614_
timestamp 1727487319
transform -1 0 2670 0 1 2870
box -6 -8 106 272
use AOI22X1  _1615_
timestamp 1727487144
transform -1 0 2850 0 1 2870
box -6 -8 126 272
use INVX1  _1616_
timestamp 1727493700
transform -1 0 3090 0 1 2870
box -6 -8 66 272
use OAI21X1  _1617_
timestamp 1727498925
transform -1 0 1390 0 -1 3390
box -6 -8 106 272
use INVX1  _1618_
timestamp 1727493700
transform -1 0 1830 0 -1 3390
box -6 -8 66 272
use OAI21X1  _1619_
timestamp 1727498925
transform 1 0 370 0 -1 3910
box -6 -8 106 272
use INVX1  _1620_
timestamp 1727493700
transform 1 0 1490 0 -1 3910
box -6 -8 66 272
use OAI21X1  _1621_
timestamp 1727498925
transform -1 0 1290 0 1 3390
box -6 -8 106 272
use OR2X2  _1622_
timestamp 1727496117
transform 1 0 1650 0 1 3390
box -6 -8 106 272
use NAND2X1  _1623_
timestamp 1727494699
transform -1 0 1590 0 1 3390
box -6 -8 86 272
use NAND2X1  _1624_
timestamp 1727494699
transform 1 0 1830 0 1 3390
box -6 -8 86 272
use NAND3X1  _1625_
timestamp 1727494898
transform 1 0 2070 0 -1 3390
box -6 -8 106 272
use OR2X2  _1626_
timestamp 1727496117
transform 1 0 2070 0 1 2870
box -6 -8 106 272
use AOI21X1  _1627_
timestamp 1727487319
transform -1 0 2330 0 1 2870
box -6 -8 106 272
use INVX1  _1628_
timestamp 1727493700
transform 1 0 2150 0 1 3390
box -6 -8 66 272
use OAI21X1  _1629_
timestamp 1727498925
transform 1 0 2230 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1630_
timestamp 1727494898
transform 1 0 2390 0 -1 3390
box -6 -8 106 272
use NAND3X1  _1631_
timestamp 1727494898
transform -1 0 5910 0 -1 2350
box -6 -8 106 272
use OAI21X1  _1632_
timestamp 1727498925
transform 1 0 6190 0 1 2350
box -6 -8 106 272
use NAND2X1  _1633_
timestamp 1727494699
transform 1 0 6030 0 1 2350
box -6 -8 86 272
use NAND2X1  _1634_
timestamp 1727494699
transform 1 0 2390 0 1 3910
box -6 -8 86 272
use OAI21X1  _1635_
timestamp 1727498925
transform -1 0 3690 0 1 3390
box -6 -8 106 272
use AOI21X1  _1636_
timestamp 1727487319
transform -1 0 3530 0 1 3390
box -6 -8 106 272
use AOI22X1  _1637_
timestamp 1727487144
transform -1 0 3010 0 -1 3390
box -6 -8 126 272
use INVX1  _1638_
timestamp 1727493700
transform 1 0 2890 0 1 3390
box -6 -8 66 272
use AOI21X1  _1639_
timestamp 1727487319
transform 1 0 1910 0 -1 3390
box -6 -8 106 272
use OAI21X1  _1640_
timestamp 1727498925
transform -1 0 1450 0 1 3390
box -6 -8 106 272
use OAI21X1  _1641_
timestamp 1727498925
transform 1 0 1970 0 1 3390
box -6 -8 106 272
use NAND3X1  _1642_
timestamp 1727494898
transform -1 0 5790 0 1 1830
box -6 -8 106 272
use OAI21X1  _1643_
timestamp 1727498925
transform -1 0 6170 0 -1 1830
box -6 -8 106 272
use NAND2X1  _1644_
timestamp 1727494699
transform -1 0 5470 0 1 1830
box -6 -8 86 272
use NAND2X1  _1645_
timestamp 1727494699
transform 1 0 2410 0 1 3390
box -6 -8 86 272
use OAI21X1  _1646_
timestamp 1727498925
transform -1 0 2650 0 -1 3390
box -6 -8 106 272
use AOI21X1  _1647_
timestamp 1727487319
transform 1 0 2730 0 -1 3390
box -6 -8 106 272
use AOI22X1  _1648_
timestamp 1727487144
transform -1 0 2830 0 1 3390
box -6 -8 126 272
use NAND2X1  _1649_
timestamp 1727494699
transform -1 0 4730 0 1 5470
box -6 -8 86 272
use OAI21X1  _1650_
timestamp 1727498925
transform -1 0 4890 0 1 5470
box -6 -8 106 272
use NAND2X1  _1651_
timestamp 1727494699
transform 1 0 4650 0 -1 5990
box -6 -8 86 272
use OAI21X1  _1652_
timestamp 1727498925
transform -1 0 4590 0 1 5470
box -6 -8 106 272
use NAND2X1  _1653_
timestamp 1727494699
transform 1 0 4710 0 1 5990
box -6 -8 86 272
use OAI21X1  _1654_
timestamp 1727498925
transform 1 0 4550 0 1 5990
box -6 -8 106 272
use NAND2X1  _1655_
timestamp 1727494699
transform 1 0 4510 0 1 4430
box -6 -8 86 272
use OAI21X1  _1656_
timestamp 1727498925
transform 1 0 4350 0 1 4430
box -6 -8 106 272
use NAND2X1  _1657_
timestamp 1727494699
transform 1 0 3970 0 1 4430
box -6 -8 86 272
use OAI21X1  _1658_
timestamp 1727498925
transform -1 0 3770 0 1 4430
box -6 -8 106 272
use NAND2X1  _1659_
timestamp 1727494699
transform -1 0 3550 0 1 3910
box -6 -8 86 272
use OAI21X1  _1660_
timestamp 1727498925
transform 1 0 3310 0 1 3910
box -6 -8 106 272
use NAND2X1  _1661_
timestamp 1727494699
transform 1 0 3190 0 -1 4430
box -6 -8 86 272
use OAI21X1  _1662_
timestamp 1727498925
transform 1 0 3030 0 -1 4430
box -6 -8 106 272
use NAND2X1  _1663_
timestamp 1727494699
transform -1 0 3910 0 1 4430
box -6 -8 86 272
use OAI21X1  _1664_
timestamp 1727498925
transform 1 0 3730 0 -1 4430
box -6 -8 106 272
use DFFPOSX1  _1665_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727503886
transform -1 0 4990 0 -1 5470
box -6 -8 246 272
use DFFPOSX1  _1666_
timestamp 1727503886
transform -1 0 5110 0 1 4950
box -6 -8 246 272
use DFFPOSX1  _1667_
timestamp 1727503886
transform -1 0 4650 0 -1 6510
box -6 -8 246 272
use DFFPOSX1  _1668_
timestamp 1727503886
transform -1 0 3890 0 -1 3910
box -6 -8 246 272
use DFFPOSX1  _1669_
timestamp 1727503886
transform -1 0 3930 0 1 3390
box -6 -8 246 272
use DFFPOSX1  _1670_
timestamp 1727503886
transform -1 0 3110 0 -1 3910
box -6 -8 246 272
use DFFPOSX1  _1671_
timestamp 1727503886
transform -1 0 2870 0 -1 3910
box -6 -8 246 272
use DFFPOSX1  _1672_
timestamp 1727503886
transform -1 0 4130 0 -1 3910
box -6 -8 246 272
use DFFPOSX1  _1673_
timestamp 1727503886
transform -1 0 2630 0 1 4430
box -6 -8 246 272
use DFFPOSX1  _1674_
timestamp 1727503886
transform -1 0 2530 0 -1 4430
box -6 -8 246 272
use DFFPOSX1  _1675_
timestamp 1727503886
transform 1 0 4230 0 -1 4950
box -6 -8 246 272
use DFFPOSX1  _1676_
timestamp 1727503886
transform 1 0 3270 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1677_
timestamp 1727503886
transform 1 0 3210 0 1 2870
box -6 -8 246 272
use DFFPOSX1  _1678_
timestamp 1727503886
transform -1 0 3070 0 -1 2870
box -6 -8 246 272
use DFFPOSX1  _1679_
timestamp 1727503886
transform -1 0 3250 0 -1 3390
box -6 -8 246 272
use DFFPOSX1  _1680_
timestamp 1727503886
transform -1 0 3190 0 1 3390
box -6 -8 246 272
use DFFPOSX1  _1681_
timestamp 1727503886
transform 1 0 5030 0 1 5470
box -6 -8 246 272
use DFFPOSX1  _1682_
timestamp 1727503886
transform -1 0 4430 0 1 5470
box -6 -8 246 272
use DFFPOSX1  _1683_
timestamp 1727503886
transform -1 0 4470 0 1 5990
box -6 -8 246 272
use DFFPOSX1  _1684_
timestamp 1727503886
transform -1 0 4290 0 1 4430
box -6 -8 246 272
use DFFPOSX1  _1685_
timestamp 1727503886
transform -1 0 3590 0 1 4430
box -6 -8 246 272
use DFFPOSX1  _1686_
timestamp 1727503886
transform 1 0 3410 0 -1 3910
box -6 -8 246 272
use DFFPOSX1  _1687_
timestamp 1727503886
transform -1 0 2950 0 -1 4430
box -6 -8 246 272
use DFFPOSX1  _1688_
timestamp 1727503886
transform -1 0 3670 0 -1 4430
box -6 -8 246 272
use DFFSR  _1689_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727492080
transform -1 0 5450 0 -1 6510
box -6 -8 486 273
use DFFSR  _1690_
timestamp 1727492080
transform -1 0 5270 0 1 5990
box -6 -8 486 273
use DFFSR  _1691_
timestamp 1727492080
transform 1 0 5270 0 1 5990
box -6 -8 486 273
use INVX1  _1692_
timestamp 1727493700
transform -1 0 3730 0 1 5990
box -6 -8 66 272
use INVX4  _1693_
timestamp 1727494067
transform -1 0 4030 0 -1 6510
box -6 -8 86 272
use OAI21X1  _1694_
timestamp 1727498925
transform -1 0 3610 0 1 5990
box -6 -8 106 272
use NOR2X1  _1695_
timestamp 1727495070
transform 1 0 3330 0 -1 6510
box -6 -8 86 272
use INVX1  _1696_
timestamp 1727493700
transform -1 0 3070 0 -1 6510
box -6 -8 66 272
use INVX2  _1697_
timestamp 1727493898
transform -1 0 3850 0 1 5470
box -6 -8 66 272
use NAND2X1  _1698_
timestamp 1727494699
transform 1 0 4210 0 1 4950
box -6 -8 86 272
use INVX2  _1699_
timestamp 1727493898
transform 1 0 3530 0 -1 5470
box -6 -8 66 272
use NAND2X1  _1700_
timestamp 1727494699
transform 1 0 3850 0 -1 5470
box -6 -8 86 272
use NAND2X1  _1701_
timestamp 1727494699
transform 1 0 3650 0 1 5470
box -6 -8 86 272
use AOI22X1  _1702_
timestamp 1727487144
transform 1 0 3650 0 -1 5470
box -6 -8 126 272
use INVX2  _1703_
timestamp 1727493898
transform 1 0 3130 0 1 4430
box -6 -8 66 272
use INVX1  _1704_
timestamp 1727493700
transform 1 0 4510 0 -1 5990
box -6 -8 66 272
use INVX1  _1705_
timestamp 1727493700
transform -1 0 3590 0 1 5470
box -6 -8 66 272
use OAI21X1  _1706_
timestamp 1727498925
transform -1 0 4010 0 1 5470
box -6 -8 106 272
use NAND2X1  _1707_
timestamp 1727494699
transform 1 0 3750 0 -1 5990
box -6 -8 86 272
use NAND2X1  _1708_
timestamp 1727494699
transform -1 0 3530 0 -1 5990
box -6 -8 86 272
use OAI21X1  _1709_
timestamp 1727498925
transform -1 0 3690 0 -1 5990
box -6 -8 106 272
use OAI21X1  _1710_
timestamp 1727498925
transform -1 0 4070 0 1 5990
box -6 -8 106 272
use AOI21X1  _1711_
timestamp 1727487319
transform -1 0 3910 0 1 5990
box -6 -8 106 272
use NOR2X1  _1712_
timestamp 1727495070
transform 1 0 2050 0 1 5470
box -6 -8 86 272
use OAI21X1  _1713_
timestamp 1727498925
transform 1 0 2510 0 -1 6510
box -6 -8 106 272
use OAI21X1  _1714_
timestamp 1727498925
transform -1 0 2850 0 1 5990
box -6 -8 106 272
use OR2X2  _1715_
timestamp 1727496117
transform 1 0 3050 0 1 5990
box -6 -8 106 272
use OAI21X1  _1716_
timestamp 1727498925
transform -1 0 3450 0 1 5990
box -6 -8 106 272
use NAND2X1  _1717_
timestamp 1727494699
transform -1 0 3290 0 1 5990
box -6 -8 86 272
use INVX1  _1718_
timestamp 1727493700
transform -1 0 2970 0 1 5990
box -6 -8 66 272
use NOR2X1  _1719_
timestamp 1727495070
transform 1 0 2850 0 -1 6510
box -6 -8 86 272
use OAI21X1  _1720_
timestamp 1727498925
transform -1 0 2770 0 -1 6510
box -6 -8 106 272
use NAND2X1  _1721_
timestamp 1727494699
transform 1 0 2790 0 1 5470
box -6 -8 86 272
use NAND3X1  _1722_
timestamp 1727494898
transform -1 0 3470 0 -1 5470
box -6 -8 106 272
use AOI22X1  _1723_
timestamp 1727487144
transform 1 0 3050 0 -1 5470
box -6 -8 126 272
use INVX1  _1724_
timestamp 1727493700
transform -1 0 3330 0 1 5470
box -6 -8 66 272
use NOR2X1  _1725_
timestamp 1727495070
transform -1 0 3470 0 1 5470
box -6 -8 86 272
use OAI21X1  _1726_
timestamp 1727498925
transform -1 0 3210 0 1 5470
box -6 -8 106 272
use OAI21X1  _1727_
timestamp 1727498925
transform -1 0 3030 0 1 5470
box -6 -8 106 272
use OAI21X1  _1728_
timestamp 1727498925
transform -1 0 2730 0 1 5470
box -6 -8 106 272
use AOI21X1  _1729_
timestamp 1727487319
transform -1 0 2570 0 1 5470
box -6 -8 106 272
use INVX1  _1730_
timestamp 1727493700
transform 1 0 2290 0 1 5990
box -6 -8 66 272
use OAI21X1  _1731_
timestamp 1727498925
transform -1 0 2690 0 1 5990
box -6 -8 106 272
use MUX2X1  _1732_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727494482
transform 1 0 2410 0 1 5990
box -6 -8 126 272
use NAND2X1  _1733_
timestamp 1727494699
transform -1 0 2450 0 -1 6510
box -6 -8 86 272
use INVX1  _1734_
timestamp 1727493700
transform 1 0 3810 0 -1 6510
box -6 -8 66 272
use OAI21X1  _1735_
timestamp 1727498925
transform -1 0 3730 0 -1 6510
box -6 -8 106 272
use MUX2X1  _1736_
timestamp 1727494482
transform -1 0 4190 0 1 5470
box -6 -8 126 272
use OAI21X1  _1737_
timestamp 1727498925
transform 1 0 4210 0 -1 5990
box -6 -8 106 272
use NAND2X1  _1738_
timestamp 1727494699
transform -1 0 4130 0 -1 5990
box -6 -8 86 272
use NAND3X1  _1739_
timestamp 1727494898
transform 1 0 3890 0 -1 5990
box -6 -8 106 272
use NAND3X1  _1740_
timestamp 1727494898
transform -1 0 3570 0 -1 6510
box -6 -8 106 272
use AOI22X1  _1741_
timestamp 1727487144
transform 1 0 3150 0 -1 6510
box -6 -8 126 272
use OAI21X1  _1742_
timestamp 1727498925
transform 1 0 2510 0 -1 5990
box -6 -8 106 272
use OAI21X1  _1743_
timestamp 1727498925
transform -1 0 2070 0 1 5990
box -6 -8 106 272
use NAND2X1  _1744_
timestamp 1727494699
transform 1 0 1950 0 -1 6510
box -6 -8 86 272
use NAND2X1  _1745_
timestamp 1727494699
transform -1 0 1890 0 -1 6510
box -6 -8 86 272
use INVX1  _1746_
timestamp 1727493700
transform 1 0 3990 0 -1 5470
box -6 -8 66 272
use NOR2X1  _1747_
timestamp 1727495070
transform 1 0 2130 0 1 5990
box -6 -8 86 272
use OAI21X1  _1748_
timestamp 1727498925
transform -1 0 1910 0 1 5990
box -6 -8 106 272
use NAND2X1  _1749_
timestamp 1727494699
transform -1 0 3350 0 1 4950
box -6 -8 86 272
use INVX1  _1750_
timestamp 1727493700
transform -1 0 4050 0 -1 4950
box -6 -8 66 272
use NOR2X1  _1751_
timestamp 1727495070
transform 1 0 4070 0 1 4950
box -6 -8 86 272
use NAND2X1  _1752_
timestamp 1727494699
transform 1 0 3930 0 1 4950
box -6 -8 86 272
use AOI22X1  _1753_
timestamp 1727487144
transform 1 0 3570 0 1 4950
box -6 -8 126 272
use OAI21X1  _1754_
timestamp 1727498925
transform -1 0 3850 0 1 4950
box -6 -8 106 272
use OAI21X1  _1755_
timestamp 1727498925
transform -1 0 3510 0 1 4950
box -6 -8 106 272
use OAI21X1  _1756_
timestamp 1727498925
transform -1 0 3070 0 -1 5990
box -6 -8 106 272
use AOI21X1  _1757_
timestamp 1727487319
transform -1 0 2890 0 -1 5990
box -6 -8 106 272
use INVX1  _1758_
timestamp 1727493700
transform -1 0 2730 0 -1 5990
box -6 -8 66 272
use OAI21X1  _1759_
timestamp 1727498925
transform 1 0 2350 0 -1 5990
box -6 -8 106 272
use MUX2X1  _1760_
timestamp 1727494482
transform -1 0 2290 0 -1 5990
box -6 -8 126 272
use NAND2X1  _1761_
timestamp 1727494699
transform 1 0 1510 0 1 5990
box -6 -8 86 272
use OAI21X1  _1762_
timestamp 1727498925
transform -1 0 1390 0 -1 6510
box -6 -8 106 272
use OAI21X1  _1763_
timestamp 1727498925
transform -1 0 1550 0 -1 6510
box -6 -8 106 272
use NAND3X1  _1764_
timestamp 1727494898
transform -1 0 1730 0 -1 6510
box -6 -8 106 272
use NAND2X1  _1765_
timestamp 1727494699
transform 1 0 1150 0 -1 6510
box -6 -8 86 272
use INVX1  _1766_
timestamp 1727493700
transform 1 0 2090 0 -1 6510
box -6 -8 66 272
use INVX1  _1767_
timestamp 1727493700
transform -1 0 150 0 -1 6510
box -6 -8 66 272
use AND2X2  _1768_
timestamp 1727487319
transform -1 0 1450 0 1 5990
box -6 -8 106 273
use NAND2X1  _1769_
timestamp 1727494699
transform -1 0 1890 0 -1 4950
box -6 -8 86 272
use AND2X2  _1770_
timestamp 1727487319
transform -1 0 2750 0 1 4950
box -6 -8 106 273
use NAND2X1  _1771_
timestamp 1727494699
transform -1 0 2590 0 1 4950
box -6 -8 86 272
use AOI22X1  _1772_
timestamp 1727487144
transform 1 0 2110 0 -1 5470
box -6 -8 126 272
use OAI21X1  _1773_
timestamp 1727498925
transform 1 0 2590 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1774_
timestamp 1727498925
transform -1 0 2050 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1775_
timestamp 1727498925
transform 1 0 1830 0 -1 5990
box -6 -8 106 272
use AOI21X1  _1776_
timestamp 1727487319
transform -1 0 1750 0 -1 5990
box -6 -8 106 272
use OAI21X1  _1777_
timestamp 1727498925
transform -1 0 1590 0 -1 5990
box -6 -8 106 272
use OAI21X1  _1778_
timestamp 1727498925
transform -1 0 1430 0 -1 5990
box -6 -8 106 272
use INVX1  _1779_
timestamp 1727493700
transform -1 0 390 0 1 5990
box -6 -8 66 272
use OAI21X1  _1780_
timestamp 1727498925
transform 1 0 210 0 -1 6510
box -6 -8 106 272
use NAND3X1  _1781_
timestamp 1727494898
transform 1 0 370 0 -1 6510
box -6 -8 106 272
use NAND2X1  _1782_
timestamp 1727494699
transform -1 0 630 0 -1 6510
box -6 -8 86 272
use INVX1  _1783_
timestamp 1727493700
transform 1 0 2750 0 -1 5470
box -6 -8 66 272
use INVX1  _1784_
timestamp 1727493700
transform 1 0 1030 0 -1 6510
box -6 -8 66 272
use AOI21X1  _1785_
timestamp 1727487319
transform -1 0 970 0 -1 6510
box -6 -8 106 272
use NAND3X1  _1786_
timestamp 1727494898
transform 1 0 710 0 -1 6510
box -6 -8 106 272
use NAND2X1  _1787_
timestamp 1727494699
transform -1 0 530 0 1 5990
box -6 -8 86 272
use INVX1  _1788_
timestamp 1727493700
transform -1 0 1270 0 -1 5990
box -6 -8 66 272
use AOI21X1  _1789_
timestamp 1727487319
transform 1 0 590 0 1 5990
box -6 -8 106 272
use NAND2X1  _1790_
timestamp 1727494699
transform 1 0 1650 0 1 3910
box -6 -8 86 272
use AND2X2  _1791_
timestamp 1727487319
transform -1 0 2190 0 1 3910
box -6 -8 106 273
use NAND2X1  _1792_
timestamp 1727494699
transform -1 0 2030 0 1 3910
box -6 -8 86 272
use AOI22X1  _1793_
timestamp 1727487144
transform 1 0 1910 0 -1 4430
box -6 -8 126 272
use OAI21X1  _1794_
timestamp 1727498925
transform -1 0 1850 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1795_
timestamp 1727498925
transform -1 0 1670 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1796_
timestamp 1727498925
transform -1 0 1990 0 1 5470
box -6 -8 106 272
use AOI21X1  _1797_
timestamp 1727487319
transform -1 0 1830 0 1 5470
box -6 -8 106 272
use OAI21X1  _1798_
timestamp 1727498925
transform -1 0 1650 0 1 5470
box -6 -8 106 272
use OAI21X1  _1799_
timestamp 1727498925
transform -1 0 1490 0 1 5470
box -6 -8 106 272
use AOI21X1  _1800_
timestamp 1727487319
transform 1 0 910 0 -1 5990
box -6 -8 106 272
use NOR2X1  _1801_
timestamp 1727495070
transform 1 0 1670 0 1 5990
box -6 -8 86 272
use OAI21X1  _1802_
timestamp 1727498925
transform -1 0 1290 0 1 5990
box -6 -8 106 272
use NAND2X1  _1803_
timestamp 1727494699
transform 1 0 1050 0 1 5990
box -6 -8 86 272
use OAI21X1  _1804_
timestamp 1727498925
transform -1 0 990 0 1 5990
box -6 -8 106 272
use INVX1  _1805_
timestamp 1727493700
transform -1 0 850 0 -1 5990
box -6 -8 66 272
use NOR2X1  _1806_
timestamp 1727495070
transform -1 0 830 0 1 5990
box -6 -8 86 272
use NOR2X1  _1807_
timestamp 1727495070
transform -1 0 1150 0 -1 5990
box -6 -8 86 272
use INVX1  _1808_
timestamp 1727493700
transform -1 0 1330 0 1 5470
box -6 -8 66 272
use NAND2X1  _1809_
timestamp 1727494699
transform -1 0 1150 0 -1 4430
box -6 -8 86 272
use AND2X2  _1810_
timestamp 1727487319
transform -1 0 1890 0 1 3910
box -6 -8 106 273
use NAND2X1  _1811_
timestamp 1727494699
transform 1 0 1490 0 1 3910
box -6 -8 86 272
use AOI22X1  _1812_
timestamp 1727487144
transform 1 0 1390 0 -1 4430
box -6 -8 126 272
use OAI21X1  _1813_
timestamp 1727498925
transform -1 0 1430 0 1 3910
box -6 -8 106 272
use OAI21X1  _1814_
timestamp 1727498925
transform -1 0 1310 0 -1 4430
box -6 -8 106 272
use OAI21X1  _1815_
timestamp 1727498925
transform 1 0 1790 0 -1 5470
box -6 -8 106 272
use AOI21X1  _1816_
timestamp 1727487319
transform -1 0 1730 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1817_
timestamp 1727498925
transform -1 0 1550 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1818_
timestamp 1727498925
transform -1 0 1390 0 -1 5470
box -6 -8 106 272
use OAI21X1  _1819_
timestamp 1727498925
transform 1 0 1110 0 1 5470
box -6 -8 106 272
use AOI21X1  _1820_
timestamp 1727487319
transform -1 0 710 0 -1 5990
box -6 -8 106 272
use INVX1  _1821_
timestamp 1727493700
transform 1 0 830 0 1 5470
box -6 -8 66 272
use NAND2X1  _1822_
timestamp 1727494699
transform -1 0 770 0 1 5470
box -6 -8 86 272
use NAND2X1  _1823_
timestamp 1727494699
transform -1 0 910 0 -1 5470
box -6 -8 86 272
use OAI21X1  _1824_
timestamp 1727498925
transform -1 0 630 0 1 5470
box -6 -8 106 272
use INVX1  _1825_
timestamp 1727493700
transform 1 0 930 0 -1 4430
box -6 -8 66 272
use AND2X2  _1826_
timestamp 1727487319
transform -1 0 1790 0 1 4430
box -6 -8 106 273
use NAND2X1  _1827_
timestamp 1727494699
transform 1 0 1550 0 1 4430
box -6 -8 86 272
use AOI22X1  _1828_
timestamp 1727487144
transform 1 0 1350 0 1 4430
box -6 -8 126 272
use OAI21X1  _1829_
timestamp 1727498925
transform -1 0 1290 0 1 4430
box -6 -8 106 272
use OAI22X1  _1830_
timestamp 1727495774
transform -1 0 1130 0 1 4430
box -6 -8 126 272
use OAI21X1  _1831_
timestamp 1727498925
transform 1 0 2010 0 1 4950
box -6 -8 106 272
use AOI21X1  _1832_
timestamp 1727487319
transform -1 0 1930 0 1 4950
box -6 -8 106 272
use OAI21X1  _1833_
timestamp 1727498925
transform -1 0 1430 0 1 4950
box -6 -8 106 272
use OAI21X1  _1834_
timestamp 1727498925
transform -1 0 1270 0 1 4950
box -6 -8 106 272
use NAND2X1  _1835_
timestamp 1727494699
transform -1 0 1070 0 -1 5470
box -6 -8 86 272
use OAI21X1  _1836_
timestamp 1727498925
transform -1 0 1050 0 1 5470
box -6 -8 106 272
use INVX1  _1837_
timestamp 1727493700
transform -1 0 410 0 -1 5470
box -6 -8 66 272
use NAND3X1  _1838_
timestamp 1727494898
transform 1 0 650 0 -1 5470
box -6 -8 106 272
use NAND2X1  _1839_
timestamp 1727494699
transform 1 0 1030 0 1 4950
box -6 -8 86 272
use INVX1  _1840_
timestamp 1727493700
transform 1 0 530 0 -1 4950
box -6 -8 66 272
use AOI21X1  _1841_
timestamp 1727487319
transform 1 0 470 0 -1 5470
box -6 -8 106 272
use NAND2X1  _1842_
timestamp 1727494699
transform 1 0 2310 0 -1 4950
box -6 -8 86 272
use AND2X2  _1843_
timestamp 1727487319
transform 1 0 1850 0 1 4430
box -6 -8 106 273
use NAND2X1  _1844_
timestamp 1727494699
transform -1 0 2090 0 1 4430
box -6 -8 86 272
use AOI22X1  _1845_
timestamp 1727487144
transform -1 0 2270 0 1 4430
box -6 -8 126 272
use OAI21X1  _1846_
timestamp 1727498925
transform 1 0 1970 0 -1 4950
box -6 -8 106 272
use OAI21X1  _1847_
timestamp 1727498925
transform 1 0 2130 0 -1 4950
box -6 -8 106 272
use OAI21X1  _1848_
timestamp 1727498925
transform 1 0 2330 0 1 4950
box -6 -8 106 272
use AOI21X1  _1849_
timestamp 1727487319
transform -1 0 2270 0 1 4950
box -6 -8 106 272
use OAI21X1  _1850_
timestamp 1727498925
transform -1 0 1770 0 1 4950
box -6 -8 106 272
use OAI21X1  _1851_
timestamp 1727498925
transform -1 0 1590 0 1 4950
box -6 -8 106 272
use OAI21X1  _1852_
timestamp 1727498925
transform 1 0 570 0 1 4950
box -6 -8 106 272
use NAND2X1  _1853_
timestamp 1727494699
transform -1 0 170 0 -1 5470
box -6 -8 86 272
use INVX1  _1854_
timestamp 1727493700
transform -1 0 290 0 -1 5470
box -6 -8 66 272
use NAND3X1  _1855_
timestamp 1727494898
transform 1 0 230 0 1 4950
box -6 -8 106 272
use NAND2X1  _1856_
timestamp 1727494699
transform 1 0 650 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1857_
timestamp 1727495070
transform -1 0 2090 0 -1 5990
box -6 -8 86 272
use NAND2X1  _1858_
timestamp 1727494699
transform -1 0 2270 0 1 5470
box -6 -8 86 272
use NOR2X1  _1859_
timestamp 1727495070
transform 1 0 2450 0 -1 5470
box -6 -8 86 272
use INVX1  _1860_
timestamp 1727493700
transform 1 0 730 0 1 4950
box -6 -8 66 272
use NAND3X1  _1861_
timestamp 1727494898
transform -1 0 970 0 1 4950
box -6 -8 106 272
use NOR2X1  _1862_
timestamp 1727495070
transform 1 0 1670 0 -1 4950
box -6 -8 86 272
use AND2X2  _1863_
timestamp 1727487319
transform 1 0 2450 0 -1 4950
box -6 -8 106 273
use NAND3X1  _1864_
timestamp 1727494898
transform -1 0 170 0 1 4950
box -6 -8 106 272
use OAI21X1  _1865_
timestamp 1727498925
transform -1 0 510 0 1 4950
box -6 -8 106 272
use NAND2X1  _1866_
timestamp 1727494699
transform 1 0 70 0 1 4430
box -6 -8 86 272
use OAI21X1  _1867_
timestamp 1727498925
transform -1 0 750 0 -1 4430
box -6 -8 106 272
use NOR2X1  _1868_
timestamp 1727495070
transform -1 0 3370 0 -1 5990
box -6 -8 86 272
use OAI21X1  _1869_
timestamp 1727498925
transform 1 0 1130 0 -1 5470
box -6 -8 106 272
use INVX1  _1870_
timestamp 1727493700
transform -1 0 130 0 1 5990
box -6 -8 66 272
use NAND3X1  _1871_
timestamp 1727494898
transform -1 0 170 0 1 5470
box -6 -8 106 272
use NAND3X1  _1872_
timestamp 1727494898
transform -1 0 190 0 -1 5990
box -6 -8 106 272
use INVX1  _1873_
timestamp 1727493700
transform -1 0 250 0 1 5990
box -6 -8 66 272
use NAND2X1  _1874_
timestamp 1727494699
transform -1 0 310 0 1 5470
box -6 -8 86 272
use AOI21X1  _1875_
timestamp 1727487319
transform -1 0 470 0 1 5470
box -6 -8 106 272
use OAI21X1  _1876_
timestamp 1727498925
transform -1 0 370 0 -1 5990
box -6 -8 106 272
use AND2X2  _1877_
timestamp 1727487319
transform 1 0 430 0 -1 5990
box -6 -8 106 273
use OAI21X1  _1878_
timestamp 1727498925
transform 1 0 350 0 -1 4430
box -6 -8 106 272
use NAND3X1  _1879_
timestamp 1727494898
transform -1 0 790 0 1 4430
box -6 -8 106 272
use INVX1  _1880_
timestamp 1727493700
transform -1 0 1470 0 -1 4950
box -6 -8 66 272
use NAND2X1  _1881_
timestamp 1727494699
transform 1 0 1530 0 -1 4950
box -6 -8 86 272
use AOI21X1  _1882_
timestamp 1727487319
transform -1 0 1170 0 -1 4950
box -6 -8 106 272
use NAND2X1  _1883_
timestamp 1727494699
transform 1 0 1250 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1884_
timestamp 1727495070
transform 1 0 930 0 -1 4950
box -6 -8 86 272
use NOR2X1  _1885_
timestamp 1727495070
transform -1 0 870 0 -1 4950
box -6 -8 86 272
use NAND3X1  _1886_
timestamp 1727494898
transform -1 0 470 0 -1 4950
box -6 -8 106 272
use INVX1  _1887_
timestamp 1727493700
transform -1 0 310 0 -1 4950
box -6 -8 66 272
use NAND3X1  _1888_
timestamp 1727494898
transform 1 0 70 0 -1 4950
box -6 -8 106 272
use NAND2X1  _1889_
timestamp 1727494699
transform 1 0 390 0 1 4430
box -6 -8 86 272
use NAND3X1  _1890_
timestamp 1727494898
transform 1 0 530 0 1 4430
box -6 -8 106 272
use AND2X2  _1891_
timestamp 1727487319
transform -1 0 330 0 1 4430
box -6 -8 106 273
use NAND2X1  _1892_
timestamp 1727494699
transform -1 0 290 0 -1 4430
box -6 -8 86 272
use NAND2X1  _1893_
timestamp 1727494699
transform 1 0 510 0 -1 4430
box -6 -8 86 272
use BUFX2  _1894_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727487319
transform -1 0 950 0 1 4430
box -6 -8 86 272
use BUFX2  _1895_
timestamp 1727487319
transform -1 0 150 0 -1 4430
box -6 -8 86 272
use BUFX2  _1896_
timestamp 1727487319
transform -1 0 4570 0 1 4950
box -6 -8 86 272
use BUFX2  _1897_
timestamp 1727487319
transform 1 0 3930 0 1 790
box -6 -8 86 272
use BUFX2  _1898_
timestamp 1727487319
transform 1 0 3650 0 1 2870
box -6 -8 86 272
use BUFX2  _1899_
timestamp 1727487319
transform 1 0 3270 0 -1 270
box -6 -8 86 272
use BUFX2  _1900_
timestamp 1727487319
transform 1 0 3170 0 -1 1830
box -6 -8 86 272
use BUFX2  _1901_
timestamp 1727487319
transform -1 0 2830 0 1 2350
box -6 -8 86 272
use BUFX2  _1902_
timestamp 1727487319
transform -1 0 5230 0 1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert0
timestamp 1727487319
transform -1 0 2390 0 1 2350
box -6 -8 86 272
use BUFX2  BUFX2_insert1
timestamp 1727487319
transform -1 0 2330 0 1 3910
box -6 -8 86 272
use BUFX2  BUFX2_insert2
timestamp 1727487319
transform 1 0 3930 0 1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert3
timestamp 1727487319
transform 1 0 3630 0 1 2350
box -6 -8 86 272
use BUFX2  BUFX2_insert4
timestamp 1727487319
transform -1 0 4870 0 1 4950
box -6 -8 86 272
use BUFX2  BUFX2_insert5
timestamp 1727487319
transform -1 0 4150 0 -1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert6
timestamp 1727487319
transform 1 0 4410 0 -1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert7
timestamp 1727487319
transform -1 0 4190 0 -1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert8
timestamp 1727487319
transform -1 0 4250 0 -1 4430
box -6 -8 86 272
use BUFX2  BUFX2_insert9
timestamp 1727487319
transform -1 0 4730 0 1 4430
box -6 -8 86 272
use BUFX2  BUFX2_insert10
timestamp 1727487319
transform 1 0 5090 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert11
timestamp 1727487319
transform 1 0 4790 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert17
timestamp 1727487319
transform -1 0 3690 0 1 3910
box -6 -8 86 272
use BUFX2  BUFX2_insert18
timestamp 1727487319
transform 1 0 4270 0 1 3910
box -6 -8 86 272
use BUFX2  BUFX2_insert19
timestamp 1727487319
transform -1 0 5290 0 -1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert20
timestamp 1727487319
transform -1 0 5010 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert21
timestamp 1727487319
transform 1 0 3850 0 -1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert22
timestamp 1727487319
transform -1 0 3770 0 -1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert23
timestamp 1727487319
transform -1 0 2010 0 1 2870
box -6 -8 86 272
use BUFX2  BUFX2_insert24
timestamp 1727487319
transform -1 0 2010 0 -1 3910
box -6 -8 86 272
use BUFX2  BUFX2_insert25
timestamp 1727487319
transform -1 0 4730 0 1 4950
box -6 -8 86 272
use BUFX2  BUFX2_insert26
timestamp 1727487319
transform 1 0 3930 0 -1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert27
timestamp 1727487319
transform 1 0 4410 0 1 3910
box -6 -8 86 272
use BUFX2  BUFX2_insert28
timestamp 1727487319
transform -1 0 3870 0 -1 3390
box -6 -8 86 272
use BUFX2  BUFX2_insert29
timestamp 1727487319
transform -1 0 2390 0 -1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert30
timestamp 1727487319
transform 1 0 2330 0 1 5470
box -6 -8 86 272
use BUFX2  BUFX2_insert31
timestamp 1727487319
transform 1 0 3130 0 -1 5990
box -6 -8 86 272
use BUFX2  BUFX2_insert32
timestamp 1727487319
transform -1 0 4230 0 1 5990
box -6 -8 86 272
use CLKBUF1  CLKBUF1_insert12 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727490190
transform 1 0 4250 0 -1 5470
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert13
timestamp 1727490190
transform -1 0 4330 0 1 3390
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert14
timestamp 1727490190
transform -1 0 4110 0 -1 4430
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert15
timestamp 1727490190
transform -1 0 4390 0 -1 3910
box -6 -8 206 272
use CLKBUF1  CLKBUF1_insert16
timestamp 1727490190
transform 1 0 4210 0 -1 6510
box -6 -8 206 272
use FILL  FILL95550x4050 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727493435
transform 1 0 6370 0 1 270
box -6 -8 26 272
use FILL  FILL95550x7950
timestamp 1727493435
transform -1 0 6390 0 -1 790
box -6 -8 26 272
use FILL  FILL95550x66450
timestamp 1727493435
transform 1 0 6370 0 1 4430
box -6 -8 26 272
use FILL  FILL95550x74250
timestamp 1727493435
transform 1 0 6370 0 1 4950
box -6 -8 26 272
use FILL  FILL95550x85950
timestamp 1727493435
transform -1 0 6390 0 -1 5990
box -6 -8 26 272
use FILL  FILL95550x89850
timestamp 1727493435
transform 1 0 6370 0 1 5990
box -6 -8 26 272
use FILL  FILL95850x4050
timestamp 1727493435
transform 1 0 6390 0 1 270
box -6 -8 26 272
use FILL  FILL95850x7950
timestamp 1727493435
transform -1 0 6410 0 -1 790
box -6 -8 26 272
use FILL  FILL95850x50850
timestamp 1727493435
transform 1 0 6390 0 1 3390
box -6 -8 26 272
use FILL  FILL95850x62550
timestamp 1727493435
transform -1 0 6410 0 -1 4430
box -6 -8 26 272
use FILL  FILL95850x66450
timestamp 1727493435
transform 1 0 6390 0 1 4430
box -6 -8 26 272
use FILL  FILL95850x74250
timestamp 1727493435
transform 1 0 6390 0 1 4950
box -6 -8 26 272
use FILL  FILL95850x85950
timestamp 1727493435
transform -1 0 6410 0 -1 5990
box -6 -8 26 272
use FILL  FILL95850x89850
timestamp 1727493435
transform 1 0 6390 0 1 5990
box -6 -8 26 272
use FILL  FILL96150x4050
timestamp 1727493435
transform 1 0 6410 0 1 270
box -6 -8 26 272
use FILL  FILL96150x7950
timestamp 1727493435
transform -1 0 6430 0 -1 790
box -6 -8 26 272
use FILL  FILL96150x15750
timestamp 1727493435
transform -1 0 6430 0 -1 1310
box -6 -8 26 272
use FILL  FILL96150x31350
timestamp 1727493435
transform -1 0 6430 0 -1 2350
box -6 -8 26 272
use FILL  FILL96150x39150
timestamp 1727493435
transform -1 0 6430 0 -1 2870
box -6 -8 26 272
use FILL  FILL96150x50850
timestamp 1727493435
transform 1 0 6410 0 1 3390
box -6 -8 26 272
use FILL  FILL96150x54750
timestamp 1727493435
transform -1 0 6430 0 -1 3910
box -6 -8 26 272
use FILL  FILL96150x62550
timestamp 1727493435
transform -1 0 6430 0 -1 4430
box -6 -8 26 272
use FILL  FILL96150x66450
timestamp 1727493435
transform 1 0 6410 0 1 4430
box -6 -8 26 272
use FILL  FILL96150x74250
timestamp 1727493435
transform 1 0 6410 0 1 4950
box -6 -8 26 272
use FILL  FILL96150x85950
timestamp 1727493435
transform -1 0 6430 0 -1 5990
box -6 -8 26 272
use FILL  FILL96150x89850
timestamp 1727493435
transform 1 0 6410 0 1 5990
box -6 -8 26 272
use FILL  FILL96450x4050
timestamp 1727493435
transform 1 0 6430 0 1 270
box -6 -8 26 272
use FILL  FILL96450x7950
timestamp 1727493435
transform -1 0 6450 0 -1 790
box -6 -8 26 272
use FILL  FILL96450x11850
timestamp 1727493435
transform 1 0 6430 0 1 790
box -6 -8 26 272
use FILL  FILL96450x15750
timestamp 1727493435
transform -1 0 6450 0 -1 1310
box -6 -8 26 272
use FILL  FILL96450x19650
timestamp 1727493435
transform 1 0 6430 0 1 1310
box -6 -8 26 272
use FILL  FILL96450x31350
timestamp 1727493435
transform -1 0 6450 0 -1 2350
box -6 -8 26 272
use FILL  FILL96450x35250
timestamp 1727493435
transform 1 0 6430 0 1 2350
box -6 -8 26 272
use FILL  FILL96450x39150
timestamp 1727493435
transform -1 0 6450 0 -1 2870
box -6 -8 26 272
use FILL  FILL96450x43050
timestamp 1727493435
transform 1 0 6430 0 1 2870
box -6 -8 26 272
use FILL  FILL96450x50850
timestamp 1727493435
transform 1 0 6430 0 1 3390
box -6 -8 26 272
use FILL  FILL96450x54750
timestamp 1727493435
transform -1 0 6450 0 -1 3910
box -6 -8 26 272
use FILL  FILL96450x62550
timestamp 1727493435
transform -1 0 6450 0 -1 4430
box -6 -8 26 272
use FILL  FILL96450x66450
timestamp 1727493435
transform 1 0 6430 0 1 4430
box -6 -8 26 272
use FILL  FILL96450x70350
timestamp 1727493435
transform -1 0 6450 0 -1 4950
box -6 -8 26 272
use FILL  FILL96450x74250
timestamp 1727493435
transform 1 0 6430 0 1 4950
box -6 -8 26 272
use FILL  FILL96450x85950
timestamp 1727493435
transform -1 0 6450 0 -1 5990
box -6 -8 26 272
use FILL  FILL96450x89850
timestamp 1727493435
transform 1 0 6430 0 1 5990
box -6 -8 26 272
use FILL  FILL96750x4050
timestamp 1727493435
transform 1 0 6450 0 1 270
box -6 -8 26 272
use FILL  FILL96750x7950
timestamp 1727493435
transform -1 0 6470 0 -1 790
box -6 -8 26 272
use FILL  FILL96750x11850
timestamp 1727493435
transform 1 0 6450 0 1 790
box -6 -8 26 272
use FILL  FILL96750x15750
timestamp 1727493435
transform -1 0 6470 0 -1 1310
box -6 -8 26 272
use FILL  FILL96750x19650
timestamp 1727493435
transform 1 0 6450 0 1 1310
box -6 -8 26 272
use FILL  FILL96750x31350
timestamp 1727493435
transform -1 0 6470 0 -1 2350
box -6 -8 26 272
use FILL  FILL96750x35250
timestamp 1727493435
transform 1 0 6450 0 1 2350
box -6 -8 26 272
use FILL  FILL96750x39150
timestamp 1727493435
transform -1 0 6470 0 -1 2870
box -6 -8 26 272
use FILL  FILL96750x43050
timestamp 1727493435
transform 1 0 6450 0 1 2870
box -6 -8 26 272
use FILL  FILL96750x50850
timestamp 1727493435
transform 1 0 6450 0 1 3390
box -6 -8 26 272
use FILL  FILL96750x54750
timestamp 1727493435
transform -1 0 6470 0 -1 3910
box -6 -8 26 272
use FILL  FILL96750x62550
timestamp 1727493435
transform -1 0 6470 0 -1 4430
box -6 -8 26 272
use FILL  FILL96750x66450
timestamp 1727493435
transform 1 0 6450 0 1 4430
box -6 -8 26 272
use FILL  FILL96750x70350
timestamp 1727493435
transform -1 0 6470 0 -1 4950
box -6 -8 26 272
use FILL  FILL96750x74250
timestamp 1727493435
transform 1 0 6450 0 1 4950
box -6 -8 26 272
use FILL  FILL96750x85950
timestamp 1727493435
transform -1 0 6470 0 -1 5990
box -6 -8 26 272
use FILL  FILL96750x89850
timestamp 1727493435
transform 1 0 6450 0 1 5990
box -6 -8 26 272
use FILL  FILL96750x93750
timestamp 1727493435
transform -1 0 6470 0 -1 6510
box -6 -8 26 272
use FILL  FILL97050x150
timestamp 1727493435
transform -1 0 6490 0 -1 270
box -6 -8 26 272
use FILL  FILL97050x4050
timestamp 1727493435
transform 1 0 6470 0 1 270
box -6 -8 26 272
use FILL  FILL97050x7950
timestamp 1727493435
transform -1 0 6490 0 -1 790
box -6 -8 26 272
use FILL  FILL97050x11850
timestamp 1727493435
transform 1 0 6470 0 1 790
box -6 -8 26 272
use FILL  FILL97050x15750
timestamp 1727493435
transform -1 0 6490 0 -1 1310
box -6 -8 26 272
use FILL  FILL97050x19650
timestamp 1727493435
transform 1 0 6470 0 1 1310
box -6 -8 26 272
use FILL  FILL97050x31350
timestamp 1727493435
transform -1 0 6490 0 -1 2350
box -6 -8 26 272
use FILL  FILL97050x35250
timestamp 1727493435
transform 1 0 6470 0 1 2350
box -6 -8 26 272
use FILL  FILL97050x39150
timestamp 1727493435
transform -1 0 6490 0 -1 2870
box -6 -8 26 272
use FILL  FILL97050x43050
timestamp 1727493435
transform 1 0 6470 0 1 2870
box -6 -8 26 272
use FILL  FILL97050x50850
timestamp 1727493435
transform 1 0 6470 0 1 3390
box -6 -8 26 272
use FILL  FILL97050x54750
timestamp 1727493435
transform -1 0 6490 0 -1 3910
box -6 -8 26 272
use FILL  FILL97050x62550
timestamp 1727493435
transform -1 0 6490 0 -1 4430
box -6 -8 26 272
use FILL  FILL97050x66450
timestamp 1727493435
transform 1 0 6470 0 1 4430
box -6 -8 26 272
use FILL  FILL97050x70350
timestamp 1727493435
transform -1 0 6490 0 -1 4950
box -6 -8 26 272
use FILL  FILL97050x74250
timestamp 1727493435
transform 1 0 6470 0 1 4950
box -6 -8 26 272
use FILL  FILL97050x85950
timestamp 1727493435
transform -1 0 6490 0 -1 5990
box -6 -8 26 272
use FILL  FILL97050x89850
timestamp 1727493435
transform 1 0 6470 0 1 5990
box -6 -8 26 272
use FILL  FILL97050x93750
timestamp 1727493435
transform -1 0 6490 0 -1 6510
box -6 -8 26 272
use FILL  FILL97350x150
timestamp 1727493435
transform -1 0 6510 0 -1 270
box -6 -8 26 272
use FILL  FILL97350x4050
timestamp 1727493435
transform 1 0 6490 0 1 270
box -6 -8 26 272
use FILL  FILL97350x7950
timestamp 1727493435
transform -1 0 6510 0 -1 790
box -6 -8 26 272
use FILL  FILL97350x11850
timestamp 1727493435
transform 1 0 6490 0 1 790
box -6 -8 26 272
use FILL  FILL97350x15750
timestamp 1727493435
transform -1 0 6510 0 -1 1310
box -6 -8 26 272
use FILL  FILL97350x19650
timestamp 1727493435
transform 1 0 6490 0 1 1310
box -6 -8 26 272
use FILL  FILL97350x23550
timestamp 1727493435
transform -1 0 6510 0 -1 1830
box -6 -8 26 272
use FILL  FILL97350x27450
timestamp 1727493435
transform 1 0 6490 0 1 1830
box -6 -8 26 272
use FILL  FILL97350x31350
timestamp 1727493435
transform -1 0 6510 0 -1 2350
box -6 -8 26 272
use FILL  FILL97350x35250
timestamp 1727493435
transform 1 0 6490 0 1 2350
box -6 -8 26 272
use FILL  FILL97350x39150
timestamp 1727493435
transform -1 0 6510 0 -1 2870
box -6 -8 26 272
use FILL  FILL97350x43050
timestamp 1727493435
transform 1 0 6490 0 1 2870
box -6 -8 26 272
use FILL  FILL97350x50850
timestamp 1727493435
transform 1 0 6490 0 1 3390
box -6 -8 26 272
use FILL  FILL97350x54750
timestamp 1727493435
transform -1 0 6510 0 -1 3910
box -6 -8 26 272
use FILL  FILL97350x58650
timestamp 1727493435
transform 1 0 6490 0 1 3910
box -6 -8 26 272
use FILL  FILL97350x62550
timestamp 1727493435
transform -1 0 6510 0 -1 4430
box -6 -8 26 272
use FILL  FILL97350x66450
timestamp 1727493435
transform 1 0 6490 0 1 4430
box -6 -8 26 272
use FILL  FILL97350x70350
timestamp 1727493435
transform -1 0 6510 0 -1 4950
box -6 -8 26 272
use FILL  FILL97350x74250
timestamp 1727493435
transform 1 0 6490 0 1 4950
box -6 -8 26 272
use FILL  FILL97350x82050
timestamp 1727493435
transform 1 0 6490 0 1 5470
box -6 -8 26 272
use FILL  FILL97350x85950
timestamp 1727493435
transform -1 0 6510 0 -1 5990
box -6 -8 26 272
use FILL  FILL97350x89850
timestamp 1727493435
transform 1 0 6490 0 1 5990
box -6 -8 26 272
use FILL  FILL97350x93750
timestamp 1727493435
transform -1 0 6510 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__927_
timestamp 1727493435
transform 1 0 5570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__928_
timestamp 1727493435
transform -1 0 5570 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__929_
timestamp 1727493435
transform -1 0 5850 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__930_
timestamp 1727493435
transform 1 0 5970 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__931_
timestamp 1727493435
transform -1 0 5290 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__932_
timestamp 1727493435
transform -1 0 3390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__933_
timestamp 1727493435
transform 1 0 5410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__934_
timestamp 1727493435
transform 1 0 5390 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__935_
timestamp 1727493435
transform 1 0 5950 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__936_
timestamp 1727493435
transform -1 0 5330 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__937_
timestamp 1727493435
transform 1 0 5530 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__938_
timestamp 1727493435
transform -1 0 5870 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__939_
timestamp 1727493435
transform 1 0 5990 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__940_
timestamp 1727493435
transform 1 0 6210 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__941_
timestamp 1727493435
transform 1 0 3770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__942_
timestamp 1727493435
transform 1 0 5690 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__943_
timestamp 1727493435
transform 1 0 5950 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__944_
timestamp 1727493435
transform 1 0 5690 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__945_
timestamp 1727493435
transform 1 0 6210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__946_
timestamp 1727493435
transform -1 0 5750 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__947_
timestamp 1727493435
transform 1 0 5710 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__948_
timestamp 1727493435
transform -1 0 5890 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__949_
timestamp 1727493435
transform 1 0 5850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__950_
timestamp 1727493435
transform -1 0 5610 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__951_
timestamp 1727493435
transform -1 0 6090 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__952_
timestamp 1727493435
transform -1 0 5630 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__953_
timestamp 1727493435
transform 1 0 5170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__954_
timestamp 1727493435
transform 1 0 6230 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__955_
timestamp 1727493435
transform 1 0 6150 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__956_
timestamp 1727493435
transform -1 0 5770 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__957_
timestamp 1727493435
transform -1 0 5470 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__958_
timestamp 1727493435
transform 1 0 6250 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__959_
timestamp 1727493435
transform -1 0 6090 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__960_
timestamp 1727493435
transform 1 0 6030 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__961_
timestamp 1727493435
transform -1 0 6070 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__962_
timestamp 1727493435
transform 1 0 5790 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__963_
timestamp 1727493435
transform -1 0 5470 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__964_
timestamp 1727493435
transform -1 0 5310 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__965_
timestamp 1727493435
transform 1 0 4450 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__966_
timestamp 1727493435
transform -1 0 4610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__967_
timestamp 1727493435
transform 1 0 4890 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__968_
timestamp 1727493435
transform 1 0 5110 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__969_
timestamp 1727493435
transform 1 0 4990 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__970_
timestamp 1727493435
transform 1 0 4030 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__971_
timestamp 1727493435
transform 1 0 4810 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__972_
timestamp 1727493435
transform 1 0 4650 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__973_
timestamp 1727493435
transform 1 0 4310 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__974_
timestamp 1727493435
transform 1 0 4330 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__975_
timestamp 1727493435
transform 1 0 4390 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__976_
timestamp 1727493435
transform 1 0 3650 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__977_
timestamp 1727493435
transform 1 0 3930 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__978_
timestamp 1727493435
transform 1 0 3690 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__979_
timestamp 1727493435
transform 1 0 3130 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__980_
timestamp 1727493435
transform 1 0 3270 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__981_
timestamp 1727493435
transform -1 0 3130 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__982_
timestamp 1727493435
transform 1 0 2030 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__983_
timestamp 1727493435
transform 1 0 2650 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__984_
timestamp 1727493435
transform -1 0 2810 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__985_
timestamp 1727493435
transform 1 0 3590 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__986_
timestamp 1727493435
transform 1 0 3870 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__987_
timestamp 1727493435
transform -1 0 4050 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__988_
timestamp 1727493435
transform -1 0 2290 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__989_
timestamp 1727493435
transform 1 0 5210 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__990_
timestamp 1727493435
transform -1 0 1730 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__991_
timestamp 1727493435
transform 1 0 5550 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__992_
timestamp 1727493435
transform 1 0 5390 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__993_
timestamp 1727493435
transform 1 0 5690 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__994_
timestamp 1727493435
transform -1 0 4270 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__995_
timestamp 1727493435
transform -1 0 4590 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__996_
timestamp 1727493435
transform 1 0 6230 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__997_
timestamp 1727493435
transform 1 0 5430 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__998_
timestamp 1727493435
transform -1 0 6230 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__999_
timestamp 1727493435
transform 1 0 6050 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1000_
timestamp 1727493435
transform -1 0 4850 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1001_
timestamp 1727493435
transform 1 0 5290 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1002_
timestamp 1727493435
transform 1 0 4630 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1003_
timestamp 1727493435
transform 1 0 4710 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1004_
timestamp 1727493435
transform 1 0 4630 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1005_
timestamp 1727493435
transform -1 0 5190 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1006_
timestamp 1727493435
transform 1 0 5570 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1007_
timestamp 1727493435
transform -1 0 4890 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1008_
timestamp 1727493435
transform -1 0 5010 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1009_
timestamp 1727493435
transform 1 0 5890 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1010_
timestamp 1727493435
transform -1 0 5330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1011_
timestamp 1727493435
transform 1 0 4910 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1012_
timestamp 1727493435
transform -1 0 3450 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1013_
timestamp 1727493435
transform -1 0 4310 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1014_
timestamp 1727493435
transform 1 0 5230 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1015_
timestamp 1727493435
transform 1 0 5230 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1016_
timestamp 1727493435
transform -1 0 5750 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1017_
timestamp 1727493435
transform 1 0 5570 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1018_
timestamp 1727493435
transform 1 0 5010 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1019_
timestamp 1727493435
transform 1 0 3930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1020_
timestamp 1727493435
transform 1 0 4110 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1021_
timestamp 1727493435
transform -1 0 4170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1022_
timestamp 1727493435
transform 1 0 4490 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1023_
timestamp 1727493435
transform -1 0 4030 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1024_
timestamp 1727493435
transform -1 0 4790 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1025_
timestamp 1727493435
transform 1 0 4610 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1026_
timestamp 1727493435
transform -1 0 4490 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1027_
timestamp 1727493435
transform 1 0 4770 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1028_
timestamp 1727493435
transform 1 0 4890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1029_
timestamp 1727493435
transform 1 0 5210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1030_
timestamp 1727493435
transform -1 0 5190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1031_
timestamp 1727493435
transform -1 0 4670 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1032_
timestamp 1727493435
transform -1 0 4350 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1033_
timestamp 1727493435
transform 1 0 4810 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1034_
timestamp 1727493435
transform -1 0 4290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1035_
timestamp 1727493435
transform 1 0 4590 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1036_
timestamp 1727493435
transform 1 0 4430 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1037_
timestamp 1727493435
transform -1 0 5110 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1038_
timestamp 1727493435
transform 1 0 4510 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1039_
timestamp 1727493435
transform 1 0 4750 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1040_
timestamp 1727493435
transform 1 0 4710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1041_
timestamp 1727493435
transform 1 0 4910 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1042_
timestamp 1727493435
transform 1 0 5470 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1043_
timestamp 1727493435
transform -1 0 5030 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1044_
timestamp 1727493435
transform 1 0 4870 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1045_
timestamp 1727493435
transform 1 0 5190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1046_
timestamp 1727493435
transform 1 0 5610 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1047_
timestamp 1727493435
transform 1 0 4970 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1048_
timestamp 1727493435
transform 1 0 5050 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1049_
timestamp 1727493435
transform 1 0 5030 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1050_
timestamp 1727493435
transform 1 0 5290 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1051_
timestamp 1727493435
transform 1 0 5770 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1052_
timestamp 1727493435
transform 1 0 5930 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1053_
timestamp 1727493435
transform 1 0 6330 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1054_
timestamp 1727493435
transform 1 0 5370 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1055_
timestamp 1727493435
transform -1 0 4190 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1056_
timestamp 1727493435
transform -1 0 2870 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1057_
timestamp 1727493435
transform -1 0 4010 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1058_
timestamp 1727493435
transform -1 0 4190 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1059_
timestamp 1727493435
transform 1 0 3090 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1060_
timestamp 1727493435
transform 1 0 3850 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1061_
timestamp 1727493435
transform 1 0 4010 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1062_
timestamp 1727493435
transform 1 0 4270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1063_
timestamp 1727493435
transform -1 0 4290 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1064_
timestamp 1727493435
transform -1 0 3970 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1065_
timestamp 1727493435
transform -1 0 3890 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1066_
timestamp 1727493435
transform -1 0 4150 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1067_
timestamp 1727493435
transform 1 0 4010 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1068_
timestamp 1727493435
transform -1 0 4570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1069_
timestamp 1727493435
transform -1 0 4310 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1070_
timestamp 1727493435
transform 1 0 4490 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1071_
timestamp 1727493435
transform 1 0 4710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1072_
timestamp 1727493435
transform 1 0 4390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1073_
timestamp 1727493435
transform 1 0 5050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1074_
timestamp 1727493435
transform 1 0 4410 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1075_
timestamp 1727493435
transform -1 0 4730 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1076_
timestamp 1727493435
transform -1 0 4570 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1077_
timestamp 1727493435
transform 1 0 4430 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1078_
timestamp 1727493435
transform -1 0 4730 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1079_
timestamp 1727493435
transform 1 0 3730 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1080_
timestamp 1727493435
transform -1 0 5190 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1081_
timestamp 1727493435
transform -1 0 4870 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1082_
timestamp 1727493435
transform 1 0 5030 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1083_
timestamp 1727493435
transform 1 0 4390 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1084_
timestamp 1727493435
transform 1 0 4590 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1085_
timestamp 1727493435
transform 1 0 4550 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1086_
timestamp 1727493435
transform 1 0 5370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1087_
timestamp 1727493435
transform 1 0 5110 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1088_
timestamp 1727493435
transform 1 0 4890 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1089_
timestamp 1727493435
transform 1 0 4450 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1090_
timestamp 1727493435
transform -1 0 5230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1091_
timestamp 1727493435
transform 1 0 4790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1092_
timestamp 1727493435
transform 1 0 5450 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1093_
timestamp 1727493435
transform 1 0 5130 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1094_
timestamp 1727493435
transform 1 0 4790 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1095_
timestamp 1727493435
transform 1 0 4970 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1096_
timestamp 1727493435
transform 1 0 5290 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1097_
timestamp 1727493435
transform -1 0 1570 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1098_
timestamp 1727493435
transform 1 0 5550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1099_
timestamp 1727493435
transform 1 0 5310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1100_
timestamp 1727493435
transform -1 0 5470 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1101_
timestamp 1727493435
transform 1 0 5590 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1102_
timestamp 1727493435
transform 1 0 5770 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1103_
timestamp 1727493435
transform 1 0 6070 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1104_
timestamp 1727493435
transform 1 0 5130 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1105_
timestamp 1727493435
transform 1 0 5270 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1106_
timestamp 1727493435
transform -1 0 5950 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1107_
timestamp 1727493435
transform -1 0 6110 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1108_
timestamp 1727493435
transform 1 0 6350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1109_
timestamp 1727493435
transform 1 0 6230 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1110_
timestamp 1727493435
transform -1 0 5790 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1111_
timestamp 1727493435
transform 1 0 4950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1112_
timestamp 1727493435
transform -1 0 4230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1113_
timestamp 1727493435
transform -1 0 3730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1114_
timestamp 1727493435
transform -1 0 3550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1115_
timestamp 1727493435
transform -1 0 3130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1116_
timestamp 1727493435
transform -1 0 3230 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1117_
timestamp 1727493435
transform -1 0 3430 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1118_
timestamp 1727493435
transform 1 0 3710 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1119_
timestamp 1727493435
transform -1 0 3730 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1120_
timestamp 1727493435
transform -1 0 3810 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1121_
timestamp 1727493435
transform -1 0 3550 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1122_
timestamp 1727493435
transform 1 0 4190 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1123_
timestamp 1727493435
transform 1 0 3690 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1124_
timestamp 1727493435
transform -1 0 3250 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1125_
timestamp 1727493435
transform -1 0 4350 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1126_
timestamp 1727493435
transform -1 0 3390 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1127_
timestamp 1727493435
transform -1 0 3390 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1128_
timestamp 1727493435
transform 1 0 3630 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1129_
timestamp 1727493435
transform 1 0 3950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1130_
timestamp 1727493435
transform 1 0 3850 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1131_
timestamp 1727493435
transform -1 0 3450 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1132_
timestamp 1727493435
transform 1 0 3510 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1133_
timestamp 1727493435
transform 1 0 3630 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1134_
timestamp 1727493435
transform -1 0 3330 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1135_
timestamp 1727493435
transform 1 0 3510 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1136_
timestamp 1727493435
transform -1 0 4130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1137_
timestamp 1727493435
transform 1 0 3690 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1138_
timestamp 1727493435
transform 1 0 3990 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1139_
timestamp 1727493435
transform 1 0 4550 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1140_
timestamp 1727493435
transform 1 0 4130 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1141_
timestamp 1727493435
transform 1 0 4170 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1142_
timestamp 1727493435
transform -1 0 4030 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1143_
timestamp 1727493435
transform -1 0 3870 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1144_
timestamp 1727493435
transform 1 0 4710 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1145_
timestamp 1727493435
transform 1 0 5030 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1146_
timestamp 1727493435
transform -1 0 4630 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1147_
timestamp 1727493435
transform 1 0 4670 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1148_
timestamp 1727493435
transform 1 0 4510 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1149_
timestamp 1727493435
transform 1 0 4990 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1150_
timestamp 1727493435
transform -1 0 5170 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1151_
timestamp 1727493435
transform -1 0 5750 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1152_
timestamp 1727493435
transform 1 0 4850 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1153_
timestamp 1727493435
transform 1 0 6330 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1154_
timestamp 1727493435
transform 1 0 6030 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1155_
timestamp 1727493435
transform -1 0 5970 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1156_
timestamp 1727493435
transform 1 0 6090 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1157_
timestamp 1727493435
transform 1 0 5850 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1158_
timestamp 1727493435
transform 1 0 6190 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1159_
timestamp 1727493435
transform 1 0 5390 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1160_
timestamp 1727493435
transform -1 0 5250 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1161_
timestamp 1727493435
transform -1 0 5090 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1162_
timestamp 1727493435
transform 1 0 5190 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1163_
timestamp 1727493435
transform 1 0 4830 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1164_
timestamp 1727493435
transform 1 0 4870 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1165_
timestamp 1727493435
transform -1 0 5570 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1166_
timestamp 1727493435
transform -1 0 5630 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1167_
timestamp 1727493435
transform 1 0 5470 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1168_
timestamp 1727493435
transform 1 0 5530 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1169_
timestamp 1727493435
transform 1 0 5790 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1170_
timestamp 1727493435
transform -1 0 5630 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1171_
timestamp 1727493435
transform -1 0 5330 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1172_
timestamp 1727493435
transform 1 0 5350 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1173_
timestamp 1727493435
transform 1 0 5630 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1174_
timestamp 1727493435
transform 1 0 6050 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1175_
timestamp 1727493435
transform 1 0 5470 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1176_
timestamp 1727493435
transform 1 0 5710 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1177_
timestamp 1727493435
transform 1 0 6270 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1178_
timestamp 1727493435
transform 1 0 6330 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1179_
timestamp 1727493435
transform 1 0 5690 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1180_
timestamp 1727493435
transform 1 0 6370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1181_
timestamp 1727493435
transform 1 0 6090 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1182_
timestamp 1727493435
transform -1 0 5790 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1183_
timestamp 1727493435
transform -1 0 4510 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1184_
timestamp 1727493435
transform 1 0 4390 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1185_
timestamp 1727493435
transform 1 0 5930 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1186_
timestamp 1727493435
transform 1 0 5350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1187_
timestamp 1727493435
transform 1 0 5510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1188_
timestamp 1727493435
transform 1 0 5690 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1189_
timestamp 1727493435
transform -1 0 5550 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1190_
timestamp 1727493435
transform 1 0 5850 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1191_
timestamp 1727493435
transform -1 0 5750 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1192_
timestamp 1727493435
transform 1 0 5450 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1193_
timestamp 1727493435
transform 1 0 5370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1194_
timestamp 1727493435
transform 1 0 5690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1195_
timestamp 1727493435
transform 1 0 6230 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1196_
timestamp 1727493435
transform 1 0 6250 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1197_
timestamp 1727493435
transform 1 0 5930 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1198_
timestamp 1727493435
transform 1 0 6230 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1199_
timestamp 1727493435
transform -1 0 6230 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1200_
timestamp 1727493435
transform 1 0 5950 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1201_
timestamp 1727493435
transform 1 0 6110 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1202_
timestamp 1727493435
transform 1 0 5910 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1203_
timestamp 1727493435
transform -1 0 5790 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1204_
timestamp 1727493435
transform 1 0 4990 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1205_
timestamp 1727493435
transform 1 0 5410 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1206_
timestamp 1727493435
transform -1 0 5150 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1207_
timestamp 1727493435
transform 1 0 5590 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1208_
timestamp 1727493435
transform -1 0 5910 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1209_
timestamp 1727493435
transform -1 0 5450 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1210_
timestamp 1727493435
transform -1 0 5610 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1211_
timestamp 1727493435
transform 1 0 5410 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1212_
timestamp 1727493435
transform -1 0 5430 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1213_
timestamp 1727493435
transform 1 0 6090 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1214_
timestamp 1727493435
transform 1 0 6270 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1215_
timestamp 1727493435
transform -1 0 5870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1216_
timestamp 1727493435
transform 1 0 6030 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1217_
timestamp 1727493435
transform -1 0 6210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1218_
timestamp 1727493435
transform 1 0 6290 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1219_
timestamp 1727493435
transform -1 0 6130 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1220_
timestamp 1727493435
transform -1 0 4730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1221_
timestamp 1727493435
transform -1 0 4850 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1222_
timestamp 1727493435
transform 1 0 6250 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1223_
timestamp 1727493435
transform -1 0 6310 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1224_
timestamp 1727493435
transform 1 0 6130 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1225_
timestamp 1727493435
transform -1 0 6130 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1226_
timestamp 1727493435
transform 1 0 4730 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1227_
timestamp 1727493435
transform -1 0 5510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1228_
timestamp 1727493435
transform -1 0 5970 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1229_
timestamp 1727493435
transform 1 0 5790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1230_
timestamp 1727493435
transform 1 0 5310 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1231_
timestamp 1727493435
transform -1 0 5030 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1232_
timestamp 1727493435
transform 1 0 5130 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1233_
timestamp 1727493435
transform -1 0 5170 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1234_
timestamp 1727493435
transform 1 0 6010 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1235_
timestamp 1727493435
transform 1 0 6170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1236_
timestamp 1727493435
transform 1 0 6050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1237_
timestamp 1727493435
transform -1 0 6290 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1238_
timestamp 1727493435
transform -1 0 6130 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1239_
timestamp 1727493435
transform 1 0 5870 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1240_
timestamp 1727493435
transform 1 0 5850 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1241_
timestamp 1727493435
transform -1 0 5970 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1242_
timestamp 1727493435
transform 1 0 5790 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1243_
timestamp 1727493435
transform -1 0 5830 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1244_
timestamp 1727493435
transform -1 0 5910 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1245_
timestamp 1727493435
transform -1 0 4950 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1246_
timestamp 1727493435
transform -1 0 5330 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1247_
timestamp 1727493435
transform 1 0 4350 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1248_
timestamp 1727493435
transform -1 0 4190 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1249_
timestamp 1727493435
transform 1 0 4650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1250_
timestamp 1727493435
transform 1 0 3790 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1251_
timestamp 1727493435
transform 1 0 4770 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1252_
timestamp 1727493435
transform -1 0 4470 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1253_
timestamp 1727493435
transform 1 0 4290 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1254_
timestamp 1727493435
transform 1 0 4970 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1255_
timestamp 1727493435
transform 1 0 4830 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1256_
timestamp 1727493435
transform -1 0 4690 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1257_
timestamp 1727493435
transform 1 0 4350 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1258_
timestamp 1727493435
transform -1 0 4390 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1259_
timestamp 1727493435
transform 1 0 2550 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1260_
timestamp 1727493435
transform -1 0 3170 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1261_
timestamp 1727493435
transform 1 0 2990 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1262_
timestamp 1727493435
transform -1 0 3090 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1263_
timestamp 1727493435
transform 1 0 2750 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1264_
timestamp 1727493435
transform 1 0 2830 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1265_
timestamp 1727493435
transform -1 0 2170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1266_
timestamp 1727493435
transform -1 0 2930 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1267_
timestamp 1727493435
transform 1 0 3250 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1268_
timestamp 1727493435
transform -1 0 2470 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1269_
timestamp 1727493435
transform -1 0 2590 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1270_
timestamp 1727493435
transform 1 0 2690 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1271_
timestamp 1727493435
transform -1 0 3570 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1272_
timestamp 1727493435
transform 1 0 2710 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1273_
timestamp 1727493435
transform -1 0 2770 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1274_
timestamp 1727493435
transform -1 0 3050 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1275_
timestamp 1727493435
transform 1 0 3030 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1276_
timestamp 1727493435
transform 1 0 3250 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1277_
timestamp 1727493435
transform 1 0 3190 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1278_
timestamp 1727493435
transform 1 0 3250 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1279_
timestamp 1727493435
transform -1 0 3390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1280_
timestamp 1727493435
transform -1 0 2990 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1281_
timestamp 1727493435
transform 1 0 3070 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1282_
timestamp 1727493435
transform -1 0 2910 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1283_
timestamp 1727493435
transform 1 0 2830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1284_
timestamp 1727493435
transform 1 0 3390 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1285_
timestamp 1727493435
transform 1 0 3410 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1286_
timestamp 1727493435
transform 1 0 3890 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1287_
timestamp 1727493435
transform -1 0 4230 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1288_
timestamp 1727493435
transform 1 0 3050 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1289_
timestamp 1727493435
transform -1 0 2930 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1290_
timestamp 1727493435
transform 1 0 4050 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1291_
timestamp 1727493435
transform -1 0 3850 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1292_
timestamp 1727493435
transform 1 0 4490 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1293_
timestamp 1727493435
transform 1 0 3730 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1294_
timestamp 1727493435
transform 1 0 3670 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1295_
timestamp 1727493435
transform -1 0 3330 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1296_
timestamp 1727493435
transform -1 0 3370 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1297_
timestamp 1727493435
transform -1 0 5170 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1298_
timestamp 1727493435
transform -1 0 4190 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1299_
timestamp 1727493435
transform 1 0 3990 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1300_
timestamp 1727493435
transform -1 0 3870 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1301_
timestamp 1727493435
transform 1 0 2430 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1302_
timestamp 1727493435
transform -1 0 2610 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1303_
timestamp 1727493435
transform -1 0 3690 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1304_
timestamp 1727493435
transform 1 0 4010 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1305_
timestamp 1727493435
transform -1 0 2730 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1306_
timestamp 1727493435
transform 1 0 2570 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1307_
timestamp 1727493435
transform -1 0 5790 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1308_
timestamp 1727493435
transform 1 0 2870 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1309_
timestamp 1727493435
transform 1 0 2270 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1310_
timestamp 1727493435
transform -1 0 2750 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1311_
timestamp 1727493435
transform -1 0 2470 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1312_
timestamp 1727493435
transform -1 0 2350 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1313_
timestamp 1727493435
transform -1 0 6190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1314_
timestamp 1727493435
transform -1 0 6310 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1315_
timestamp 1727493435
transform 1 0 6350 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1316_
timestamp 1727493435
transform -1 0 6270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1317_
timestamp 1727493435
transform -1 0 5930 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1318_
timestamp 1727493435
transform 1 0 6070 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1319_
timestamp 1727493435
transform -1 0 5610 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1320_
timestamp 1727493435
transform -1 0 5490 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1321_
timestamp 1727493435
transform 1 0 2550 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1322_
timestamp 1727493435
transform 1 0 2810 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1323_
timestamp 1727493435
transform -1 0 2410 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1324_
timestamp 1727493435
transform -1 0 2770 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1325_
timestamp 1727493435
transform -1 0 2910 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1326_
timestamp 1727493435
transform 1 0 2710 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1327_
timestamp 1727493435
transform -1 0 3510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1328_
timestamp 1727493435
transform 1 0 2810 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1329_
timestamp 1727493435
transform -1 0 2890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1330_
timestamp 1727493435
transform 1 0 2790 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1331_
timestamp 1727493435
transform 1 0 2630 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1332_
timestamp 1727493435
transform 1 0 2170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1333_
timestamp 1727493435
transform 1 0 2010 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1334_
timestamp 1727493435
transform -1 0 2490 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1335_
timestamp 1727493435
transform 1 0 2150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1336_
timestamp 1727493435
transform -1 0 3530 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1337_
timestamp 1727493435
transform 1 0 3030 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1338_
timestamp 1727493435
transform -1 0 4630 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1339_
timestamp 1727493435
transform -1 0 3590 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1340_
timestamp 1727493435
transform -1 0 3510 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1341_
timestamp 1727493435
transform -1 0 2790 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1342_
timestamp 1727493435
transform -1 0 2670 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1343_
timestamp 1727493435
transform -1 0 2990 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1344_
timestamp 1727493435
transform -1 0 2290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1345_
timestamp 1727493435
transform -1 0 2330 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1346_
timestamp 1727493435
transform 1 0 2210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1347_
timestamp 1727493435
transform -1 0 2510 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1348_
timestamp 1727493435
transform -1 0 1910 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1349_
timestamp 1727493435
transform -1 0 2090 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1350_
timestamp 1727493435
transform 1 0 2170 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1351_
timestamp 1727493435
transform 1 0 2030 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1352_
timestamp 1727493435
transform 1 0 3250 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1353_
timestamp 1727493435
transform -1 0 2750 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1354_
timestamp 1727493435
transform -1 0 1490 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1355_
timestamp 1727493435
transform -1 0 1250 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1356_
timestamp 1727493435
transform 1 0 1790 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1357_
timestamp 1727493435
transform -1 0 2110 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1358_
timestamp 1727493435
transform 1 0 1950 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1359_
timestamp 1727493435
transform 1 0 1270 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1360_
timestamp 1727493435
transform -1 0 930 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1361_
timestamp 1727493435
transform 1 0 1190 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1362_
timestamp 1727493435
transform 1 0 1290 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1363_
timestamp 1727493435
transform 1 0 1610 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1364_
timestamp 1727493435
transform -1 0 2410 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1365_
timestamp 1727493435
transform -1 0 1390 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1366_
timestamp 1727493435
transform -1 0 1350 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1367_
timestamp 1727493435
transform 1 0 1530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1368_
timestamp 1727493435
transform -1 0 1050 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1369_
timestamp 1727493435
transform 1 0 1530 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1370_
timestamp 1727493435
transform -1 0 1370 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1371_
timestamp 1727493435
transform -1 0 1430 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1372_
timestamp 1727493435
transform 1 0 2130 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1373_
timestamp 1727493435
transform 1 0 2890 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1374_
timestamp 1727493435
transform 1 0 2370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1375_
timestamp 1727493435
transform 1 0 1730 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1376_
timestamp 1727493435
transform 1 0 1810 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1377_
timestamp 1727493435
transform -1 0 1890 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1378_
timestamp 1727493435
transform 1 0 1550 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1379_
timestamp 1727493435
transform 1 0 1550 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1380_
timestamp 1727493435
transform -1 0 1450 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1381_
timestamp 1727493435
transform -1 0 850 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1382_
timestamp 1727493435
transform -1 0 3090 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1383_
timestamp 1727493435
transform -1 0 2930 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1384_
timestamp 1727493435
transform 1 0 1590 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1385_
timestamp 1727493435
transform 1 0 1690 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1386_
timestamp 1727493435
transform -1 0 2590 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1387_
timestamp 1727493435
transform 1 0 1970 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1388_
timestamp 1727493435
transform -1 0 1290 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1389_
timestamp 1727493435
transform -1 0 1150 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1390_
timestamp 1727493435
transform -1 0 1030 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1391_
timestamp 1727493435
transform 1 0 1110 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1392_
timestamp 1727493435
transform 1 0 1750 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1393_
timestamp 1727493435
transform 1 0 1470 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1394_
timestamp 1727493435
transform 1 0 1830 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1395_
timestamp 1727493435
transform 1 0 1310 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1396_
timestamp 1727493435
transform 1 0 1910 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1397_
timestamp 1727493435
transform -1 0 2270 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1398_
timestamp 1727493435
transform 1 0 2430 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1399_
timestamp 1727493435
transform 1 0 2470 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1400_
timestamp 1727493435
transform -1 0 2650 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1401_
timestamp 1727493435
transform -1 0 2010 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1402_
timestamp 1727493435
transform -1 0 2130 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1403_
timestamp 1727493435
transform 1 0 2090 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1404_
timestamp 1727493435
transform 1 0 1650 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1405_
timestamp 1727493435
transform 1 0 2430 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1406_
timestamp 1727493435
transform -1 0 2570 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1407_
timestamp 1727493435
transform -1 0 2530 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1408_
timestamp 1727493435
transform -1 0 4830 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1409_
timestamp 1727493435
transform 1 0 4290 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1410_
timestamp 1727493435
transform -1 0 4670 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1411_
timestamp 1727493435
transform -1 0 4490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1412_
timestamp 1727493435
transform -1 0 3210 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1413_
timestamp 1727493435
transform 1 0 2530 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1414_
timestamp 1727493435
transform -1 0 5270 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1415_
timestamp 1727493435
transform -1 0 2170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1416_
timestamp 1727493435
transform -1 0 2290 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1417_
timestamp 1727493435
transform 1 0 1830 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1418_
timestamp 1727493435
transform 1 0 2330 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1419_
timestamp 1727493435
transform -1 0 1290 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1420_
timestamp 1727493435
transform -1 0 1490 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1421_
timestamp 1727493435
transform -1 0 910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1422_
timestamp 1727493435
transform 1 0 990 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1423_
timestamp 1727493435
transform -1 0 630 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1424_
timestamp 1727493435
transform -1 0 1090 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1425_
timestamp 1727493435
transform -1 0 430 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1426_
timestamp 1727493435
transform 1 0 710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1427_
timestamp 1727493435
transform -1 0 850 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1428_
timestamp 1727493435
transform 1 0 550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1429_
timestamp 1727493435
transform -1 0 290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1430_
timestamp 1727493435
transform 1 0 650 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1431_
timestamp 1727493435
transform 1 0 810 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1432_
timestamp 1727493435
transform 1 0 1530 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1433_
timestamp 1727493435
transform -1 0 790 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1434_
timestamp 1727493435
transform -1 0 330 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1435_
timestamp 1727493435
transform -1 0 950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1436_
timestamp 1727493435
transform 1 0 950 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1437_
timestamp 1727493435
transform 1 0 790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1438_
timestamp 1727493435
transform -1 0 170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1439_
timestamp 1727493435
transform 1 0 1090 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1440_
timestamp 1727493435
transform -1 0 30 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1441_
timestamp 1727493435
transform -1 0 150 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1442_
timestamp 1727493435
transform -1 0 470 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1443_
timestamp 1727493435
transform -1 0 350 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1444_
timestamp 1727493435
transform -1 0 490 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1445_
timestamp 1727493435
transform -1 0 650 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1446_
timestamp 1727493435
transform -1 0 30 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1447_
timestamp 1727493435
transform 1 0 290 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1448_
timestamp 1727493435
transform -1 0 650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1449_
timestamp 1727493435
transform 1 0 950 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1450_
timestamp 1727493435
transform -1 0 190 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1451_
timestamp 1727493435
transform 1 0 450 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1452_
timestamp 1727493435
transform 1 0 790 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1453_
timestamp 1727493435
transform -1 0 1650 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1454_
timestamp 1727493435
transform -1 0 630 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1455_
timestamp 1727493435
transform 1 0 170 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1456_
timestamp 1727493435
transform -1 0 30 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1457_
timestamp 1727493435
transform 1 0 330 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1458_
timestamp 1727493435
transform 1 0 650 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1459_
timestamp 1727493435
transform -1 0 510 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1460_
timestamp 1727493435
transform 1 0 1130 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1461_
timestamp 1727493435
transform 1 0 810 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1462_
timestamp 1727493435
transform -1 0 1330 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1463_
timestamp 1727493435
transform -1 0 30 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1464_
timestamp 1727493435
transform -1 0 170 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1465_
timestamp 1727493435
transform -1 0 690 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1466_
timestamp 1727493435
transform -1 0 530 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1467_
timestamp 1727493435
transform 1 0 330 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1468_
timestamp 1727493435
transform -1 0 990 0 1 270
box -6 -8 26 272
use FILL  FILL_0__1469_
timestamp 1727493435
transform -1 0 1530 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1470_
timestamp 1727493435
transform -1 0 2030 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1471_
timestamp 1727493435
transform -1 0 1850 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1472_
timestamp 1727493435
transform -1 0 1050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1473_
timestamp 1727493435
transform 1 0 2090 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1474_
timestamp 1727493435
transform 1 0 2230 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1475_
timestamp 1727493435
transform -1 0 2570 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1476_
timestamp 1727493435
transform 1 0 3050 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1477_
timestamp 1727493435
transform -1 0 5650 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1478_
timestamp 1727493435
transform -1 0 5350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1479_
timestamp 1727493435
transform -1 0 2170 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1480_
timestamp 1727493435
transform 1 0 3170 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1481_
timestamp 1727493435
transform -1 0 3210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1482_
timestamp 1727493435
transform 1 0 4050 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1483_
timestamp 1727493435
transform 1 0 3510 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1484_
timestamp 1727493435
transform 1 0 1150 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1485_
timestamp 1727493435
transform 1 0 2310 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1486_
timestamp 1727493435
transform 1 0 1390 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1487_
timestamp 1727493435
transform -1 0 510 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1488_
timestamp 1727493435
transform 1 0 510 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1489_
timestamp 1727493435
transform -1 0 30 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1490_
timestamp 1727493435
transform -1 0 1450 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1491_
timestamp 1727493435
transform 1 0 890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1492_
timestamp 1727493435
transform -1 0 830 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1493_
timestamp 1727493435
transform -1 0 630 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1494_
timestamp 1727493435
transform -1 0 470 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1495_
timestamp 1727493435
transform -1 0 310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1496_
timestamp 1727493435
transform -1 0 370 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1497_
timestamp 1727493435
transform 1 0 1070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1498_
timestamp 1727493435
transform -1 0 530 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1499_
timestamp 1727493435
transform 1 0 650 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1500_
timestamp 1727493435
transform 1 0 1130 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1501_
timestamp 1727493435
transform 1 0 1270 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1502_
timestamp 1727493435
transform -1 0 1030 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1503_
timestamp 1727493435
transform -1 0 610 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1504_
timestamp 1727493435
transform 1 0 870 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1505_
timestamp 1727493435
transform -1 0 710 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1506_
timestamp 1727493435
transform -1 0 550 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1507_
timestamp 1727493435
transform -1 0 210 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1508_
timestamp 1727493435
transform -1 0 30 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1509_
timestamp 1727493435
transform -1 0 30 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1510_
timestamp 1727493435
transform 1 0 10 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1511_
timestamp 1727493435
transform -1 0 150 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1512_
timestamp 1727493435
transform -1 0 30 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1513_
timestamp 1727493435
transform 1 0 190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1514_
timestamp 1727493435
transform -1 0 370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1515_
timestamp 1727493435
transform 1 0 170 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1516_
timestamp 1727493435
transform -1 0 30 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1517_
timestamp 1727493435
transform -1 0 350 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1518_
timestamp 1727493435
transform -1 0 810 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1519_
timestamp 1727493435
transform -1 0 1110 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1520_
timestamp 1727493435
transform 1 0 950 0 -1 790
box -6 -8 26 272
use FILL  FILL_0__1521_
timestamp 1727493435
transform 1 0 1110 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1522_
timestamp 1727493435
transform 1 0 930 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1523_
timestamp 1727493435
transform -1 0 1270 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1524_
timestamp 1727493435
transform 1 0 1670 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1525_
timestamp 1727493435
transform 1 0 1930 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1526_
timestamp 1727493435
transform -1 0 1870 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1527_
timestamp 1727493435
transform 1 0 1970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1528_
timestamp 1727493435
transform 1 0 2670 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1529_
timestamp 1727493435
transform -1 0 5030 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1530_
timestamp 1727493435
transform -1 0 4890 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1531_
timestamp 1727493435
transform -1 0 4570 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1532_
timestamp 1727493435
transform 1 0 3050 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1533_
timestamp 1727493435
transform -1 0 3290 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1534_
timestamp 1727493435
transform 1 0 3430 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1535_
timestamp 1727493435
transform -1 0 3090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1536_
timestamp 1727493435
transform 1 0 3450 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1537_
timestamp 1727493435
transform -1 0 150 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1538_
timestamp 1727493435
transform 1 0 1150 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1539_
timestamp 1727493435
transform -1 0 730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1540_
timestamp 1727493435
transform -1 0 610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1541_
timestamp 1727493435
transform 1 0 950 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1542_
timestamp 1727493435
transform 1 0 970 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1543_
timestamp 1727493435
transform 1 0 810 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1544_
timestamp 1727493435
transform 1 0 870 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1545_
timestamp 1727493435
transform -1 0 730 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1546_
timestamp 1727493435
transform 1 0 430 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1547_
timestamp 1727493435
transform -1 0 670 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1548_
timestamp 1727493435
transform -1 0 810 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1549_
timestamp 1727493435
transform 1 0 290 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1550_
timestamp 1727493435
transform -1 0 650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1551_
timestamp 1727493435
transform -1 0 30 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1552_
timestamp 1727493435
transform 1 0 130 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1553_
timestamp 1727493435
transform 1 0 10 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1554_
timestamp 1727493435
transform -1 0 30 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1555_
timestamp 1727493435
transform 1 0 170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1556_
timestamp 1727493435
transform 1 0 270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1557_
timestamp 1727493435
transform 1 0 10 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1558_
timestamp 1727493435
transform -1 0 170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1559_
timestamp 1727493435
transform -1 0 450 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1560_
timestamp 1727493435
transform 1 0 1010 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1561_
timestamp 1727493435
transform 1 0 1270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1562_
timestamp 1727493435
transform 1 0 990 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1563_
timestamp 1727493435
transform -1 0 1430 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1564_
timestamp 1727493435
transform 1 0 2610 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1565_
timestamp 1727493435
transform -1 0 1410 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1566_
timestamp 1727493435
transform 1 0 2150 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1567_
timestamp 1727493435
transform 1 0 1250 0 -1 1310
box -6 -8 26 272
use FILL  FILL_0__1568_
timestamp 1727493435
transform 1 0 1950 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1569_
timestamp 1727493435
transform 1 0 2230 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1570_
timestamp 1727493435
transform 1 0 2390 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1571_
timestamp 1727493435
transform -1 0 1130 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1572_
timestamp 1727493435
transform -1 0 1170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1573_
timestamp 1727493435
transform -1 0 1690 0 1 1310
box -6 -8 26 272
use FILL  FILL_0__1574_
timestamp 1727493435
transform -1 0 1690 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1575_
timestamp 1727493435
transform 1 0 2070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1576_
timestamp 1727493435
transform 1 0 2330 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1577_
timestamp 1727493435
transform -1 0 1730 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1578_
timestamp 1727493435
transform 1 0 2490 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1579_
timestamp 1727493435
transform 1 0 6370 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1580_
timestamp 1727493435
transform 1 0 6190 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1581_
timestamp 1727493435
transform 1 0 6050 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1582_
timestamp 1727493435
transform 1 0 2930 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1583_
timestamp 1727493435
transform -1 0 2970 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1584_
timestamp 1727493435
transform 1 0 3190 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1585_
timestamp 1727493435
transform -1 0 3270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1586_
timestamp 1727493435
transform 1 0 2850 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1587_
timestamp 1727493435
transform -1 0 490 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1588_
timestamp 1727493435
transform 1 0 970 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1589_
timestamp 1727493435
transform 1 0 830 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1590_
timestamp 1727493435
transform 1 0 650 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1591_
timestamp 1727493435
transform -1 0 510 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1592_
timestamp 1727493435
transform 1 0 10 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1593_
timestamp 1727493435
transform -1 0 30 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1594_
timestamp 1727493435
transform 1 0 170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1595_
timestamp 1727493435
transform -1 0 190 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1596_
timestamp 1727493435
transform 1 0 330 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1597_
timestamp 1727493435
transform 1 0 330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1598_
timestamp 1727493435
transform -1 0 370 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1599_
timestamp 1727493435
transform -1 0 210 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1600_
timestamp 1727493435
transform 1 0 470 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1601_
timestamp 1727493435
transform 1 0 1150 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1602_
timestamp 1727493435
transform -1 0 1610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1603_
timestamp 1727493435
transform 1 0 1750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1604_
timestamp 1727493435
transform -1 0 1930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1605_
timestamp 1727493435
transform 1 0 1550 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1606_
timestamp 1727493435
transform 1 0 2210 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1607_
timestamp 1727493435
transform 1 0 1390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1608_
timestamp 1727493435
transform 1 0 1550 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1609_
timestamp 1727493435
transform 1 0 1710 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1610_
timestamp 1727493435
transform -1 0 5710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1611_
timestamp 1727493435
transform -1 0 5550 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0__1612_
timestamp 1727493435
transform 1 0 750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1613_
timestamp 1727493435
transform 1 0 2470 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1614_
timestamp 1727493435
transform -1 0 2530 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1615_
timestamp 1727493435
transform -1 0 2690 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1616_
timestamp 1727493435
transform -1 0 2990 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1617_
timestamp 1727493435
transform -1 0 1230 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1618_
timestamp 1727493435
transform -1 0 1730 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1619_
timestamp 1727493435
transform 1 0 310 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1620_
timestamp 1727493435
transform 1 0 1430 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0__1621_
timestamp 1727493435
transform -1 0 1130 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1622_
timestamp 1727493435
transform 1 0 1590 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1623_
timestamp 1727493435
transform -1 0 1470 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1624_
timestamp 1727493435
transform 1 0 1750 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1625_
timestamp 1727493435
transform 1 0 2010 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1626_
timestamp 1727493435
transform 1 0 2010 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1627_
timestamp 1727493435
transform -1 0 2190 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1628_
timestamp 1727493435
transform 1 0 2070 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1629_
timestamp 1727493435
transform 1 0 2170 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1630_
timestamp 1727493435
transform 1 0 2330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1631_
timestamp 1727493435
transform -1 0 5770 0 -1 2350
box -6 -8 26 272
use FILL  FILL_0__1632_
timestamp 1727493435
transform 1 0 6110 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1633_
timestamp 1727493435
transform 1 0 5970 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1634_
timestamp 1727493435
transform 1 0 2330 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1635_
timestamp 1727493435
transform -1 0 3550 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1636_
timestamp 1727493435
transform -1 0 3370 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1637_
timestamp 1727493435
transform -1 0 2850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1638_
timestamp 1727493435
transform 1 0 2830 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1639_
timestamp 1727493435
transform 1 0 1830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1640_
timestamp 1727493435
transform -1 0 1310 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1641_
timestamp 1727493435
transform 1 0 1910 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1642_
timestamp 1727493435
transform -1 0 5650 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1643_
timestamp 1727493435
transform -1 0 6010 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1644_
timestamp 1727493435
transform -1 0 5350 0 1 1830
box -6 -8 26 272
use FILL  FILL_0__1645_
timestamp 1727493435
transform 1 0 2350 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1646_
timestamp 1727493435
transform -1 0 2510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1647_
timestamp 1727493435
transform 1 0 2650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0__1648_
timestamp 1727493435
transform -1 0 2670 0 1 3390
box -6 -8 26 272
use FILL  FILL_0__1649_
timestamp 1727493435
transform -1 0 4610 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1650_
timestamp 1727493435
transform -1 0 4750 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1651_
timestamp 1727493435
transform 1 0 4570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1652_
timestamp 1727493435
transform -1 0 4450 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1653_
timestamp 1727493435
transform 1 0 4650 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1654_
timestamp 1727493435
transform 1 0 4470 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1655_
timestamp 1727493435
transform 1 0 4450 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1656_
timestamp 1727493435
transform 1 0 4290 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1657_
timestamp 1727493435
transform 1 0 3910 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1658_
timestamp 1727493435
transform -1 0 3610 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1659_
timestamp 1727493435
transform -1 0 3430 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1660_
timestamp 1727493435
transform 1 0 3250 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1661_
timestamp 1727493435
transform 1 0 3130 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1662_
timestamp 1727493435
transform 1 0 2950 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1663_
timestamp 1727493435
transform -1 0 3790 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1664_
timestamp 1727493435
transform 1 0 3670 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1692_
timestamp 1727493435
transform -1 0 3630 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1693_
timestamp 1727493435
transform -1 0 3890 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1694_
timestamp 1727493435
transform -1 0 3470 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1695_
timestamp 1727493435
transform 1 0 3270 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1696_
timestamp 1727493435
transform -1 0 2950 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1697_
timestamp 1727493435
transform -1 0 3750 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1698_
timestamp 1727493435
transform 1 0 4150 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1699_
timestamp 1727493435
transform 1 0 3470 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1700_
timestamp 1727493435
transform 1 0 3770 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1701_
timestamp 1727493435
transform 1 0 3590 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1702_
timestamp 1727493435
transform 1 0 3590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1703_
timestamp 1727493435
transform 1 0 3070 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1704_
timestamp 1727493435
transform 1 0 4430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1705_
timestamp 1727493435
transform -1 0 3490 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1706_
timestamp 1727493435
transform -1 0 3870 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1707_
timestamp 1727493435
transform 1 0 3690 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1708_
timestamp 1727493435
transform -1 0 3390 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1709_
timestamp 1727493435
transform -1 0 3550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1710_
timestamp 1727493435
transform -1 0 3930 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1711_
timestamp 1727493435
transform -1 0 3750 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1712_
timestamp 1727493435
transform 1 0 1990 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1713_
timestamp 1727493435
transform 1 0 2450 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1714_
timestamp 1727493435
transform -1 0 2710 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1715_
timestamp 1727493435
transform 1 0 2970 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1716_
timestamp 1727493435
transform -1 0 3310 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1717_
timestamp 1727493435
transform -1 0 3170 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1718_
timestamp 1727493435
transform -1 0 2870 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1719_
timestamp 1727493435
transform 1 0 2770 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1720_
timestamp 1727493435
transform -1 0 2630 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1721_
timestamp 1727493435
transform 1 0 2730 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1722_
timestamp 1727493435
transform -1 0 3330 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1723_
timestamp 1727493435
transform 1 0 2970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1724_
timestamp 1727493435
transform -1 0 3230 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1725_
timestamp 1727493435
transform -1 0 3350 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1726_
timestamp 1727493435
transform -1 0 3050 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1727_
timestamp 1727493435
transform -1 0 2890 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1728_
timestamp 1727493435
transform -1 0 2590 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1729_
timestamp 1727493435
transform -1 0 2430 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1730_
timestamp 1727493435
transform 1 0 2210 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1731_
timestamp 1727493435
transform -1 0 2550 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1732_
timestamp 1727493435
transform 1 0 2350 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1733_
timestamp 1727493435
transform -1 0 2330 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1734_
timestamp 1727493435
transform 1 0 3730 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1735_
timestamp 1727493435
transform -1 0 3590 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1736_
timestamp 1727493435
transform -1 0 4030 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1737_
timestamp 1727493435
transform 1 0 4130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1738_
timestamp 1727493435
transform -1 0 4010 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1739_
timestamp 1727493435
transform 1 0 3830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1740_
timestamp 1727493435
transform -1 0 3430 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1741_
timestamp 1727493435
transform 1 0 3070 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1742_
timestamp 1727493435
transform 1 0 2450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1743_
timestamp 1727493435
transform -1 0 1930 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1744_
timestamp 1727493435
transform 1 0 1890 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1745_
timestamp 1727493435
transform -1 0 1750 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1746_
timestamp 1727493435
transform 1 0 3930 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1747_
timestamp 1727493435
transform 1 0 2070 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1748_
timestamp 1727493435
transform -1 0 1770 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1749_
timestamp 1727493435
transform -1 0 3210 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1750_
timestamp 1727493435
transform -1 0 3950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1751_
timestamp 1727493435
transform 1 0 4010 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1752_
timestamp 1727493435
transform 1 0 3850 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1753_
timestamp 1727493435
transform 1 0 3510 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1754_
timestamp 1727493435
transform -1 0 3710 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1755_
timestamp 1727493435
transform -1 0 3370 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1756_
timestamp 1727493435
transform -1 0 2910 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1757_
timestamp 1727493435
transform -1 0 2750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1758_
timestamp 1727493435
transform -1 0 2630 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1759_
timestamp 1727493435
transform 1 0 2290 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1760_
timestamp 1727493435
transform -1 0 2110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1761_
timestamp 1727493435
transform 1 0 1450 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1762_
timestamp 1727493435
transform -1 0 1250 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1763_
timestamp 1727493435
transform -1 0 1410 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1764_
timestamp 1727493435
transform -1 0 1570 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1765_
timestamp 1727493435
transform 1 0 1090 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1766_
timestamp 1727493435
transform 1 0 2030 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1767_
timestamp 1727493435
transform -1 0 30 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1768_
timestamp 1727493435
transform -1 0 1310 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1769_
timestamp 1727493435
transform -1 0 1770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1770_
timestamp 1727493435
transform -1 0 2610 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1771_
timestamp 1727493435
transform -1 0 2450 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1772_
timestamp 1727493435
transform 1 0 2050 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1773_
timestamp 1727493435
transform 1 0 2530 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1774_
timestamp 1727493435
transform -1 0 1910 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1775_
timestamp 1727493435
transform 1 0 1750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1776_
timestamp 1727493435
transform -1 0 1610 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1777_
timestamp 1727493435
transform -1 0 1450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1778_
timestamp 1727493435
transform -1 0 1290 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1779_
timestamp 1727493435
transform -1 0 270 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1780_
timestamp 1727493435
transform 1 0 150 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1781_
timestamp 1727493435
transform 1 0 310 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1782_
timestamp 1727493435
transform -1 0 490 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1783_
timestamp 1727493435
transform 1 0 2690 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1784_
timestamp 1727493435
transform 1 0 970 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1785_
timestamp 1727493435
transform -1 0 830 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1786_
timestamp 1727493435
transform 1 0 630 0 -1 6510
box -6 -8 26 272
use FILL  FILL_0__1787_
timestamp 1727493435
transform -1 0 410 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1788_
timestamp 1727493435
transform -1 0 1170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1789_
timestamp 1727493435
transform 1 0 530 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1790_
timestamp 1727493435
transform 1 0 1570 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1791_
timestamp 1727493435
transform -1 0 2050 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1792_
timestamp 1727493435
transform -1 0 1910 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1793_
timestamp 1727493435
transform 1 0 1850 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1794_
timestamp 1727493435
transform -1 0 1690 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1795_
timestamp 1727493435
transform -1 0 1530 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1796_
timestamp 1727493435
transform -1 0 1850 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1797_
timestamp 1727493435
transform -1 0 1670 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1798_
timestamp 1727493435
transform -1 0 1510 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1799_
timestamp 1727493435
transform -1 0 1350 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1800_
timestamp 1727493435
transform 1 0 850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1801_
timestamp 1727493435
transform 1 0 1590 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1802_
timestamp 1727493435
transform -1 0 1150 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1803_
timestamp 1727493435
transform 1 0 990 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1804_
timestamp 1727493435
transform -1 0 850 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1805_
timestamp 1727493435
transform -1 0 730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1806_
timestamp 1727493435
transform -1 0 710 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1807_
timestamp 1727493435
transform -1 0 1030 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1808_
timestamp 1727493435
transform -1 0 1230 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1809_
timestamp 1727493435
transform -1 0 1010 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1810_
timestamp 1727493435
transform -1 0 1750 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1811_
timestamp 1727493435
transform 1 0 1430 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1812_
timestamp 1727493435
transform 1 0 1310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1813_
timestamp 1727493435
transform -1 0 1290 0 1 3910
box -6 -8 26 272
use FILL  FILL_0__1814_
timestamp 1727493435
transform -1 0 1170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1815_
timestamp 1727493435
transform 1 0 1730 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1816_
timestamp 1727493435
transform -1 0 1570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1817_
timestamp 1727493435
transform -1 0 1410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1818_
timestamp 1727493435
transform -1 0 1250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1819_
timestamp 1727493435
transform 1 0 1050 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1820_
timestamp 1727493435
transform -1 0 550 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1821_
timestamp 1727493435
transform 1 0 770 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1822_
timestamp 1727493435
transform -1 0 650 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1823_
timestamp 1727493435
transform -1 0 770 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1824_
timestamp 1727493435
transform -1 0 490 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1825_
timestamp 1727493435
transform 1 0 870 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1826_
timestamp 1727493435
transform -1 0 1650 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1827_
timestamp 1727493435
transform 1 0 1470 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1828_
timestamp 1727493435
transform 1 0 1290 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1829_
timestamp 1727493435
transform -1 0 1150 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1830_
timestamp 1727493435
transform -1 0 970 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1831_
timestamp 1727493435
transform 1 0 1930 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1832_
timestamp 1727493435
transform -1 0 1790 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1833_
timestamp 1727493435
transform -1 0 1290 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1834_
timestamp 1727493435
transform -1 0 1130 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1835_
timestamp 1727493435
transform -1 0 930 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1836_
timestamp 1727493435
transform -1 0 910 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1837_
timestamp 1727493435
transform -1 0 310 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1838_
timestamp 1727493435
transform 1 0 570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1839_
timestamp 1727493435
transform 1 0 970 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1840_
timestamp 1727493435
transform 1 0 470 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1841_
timestamp 1727493435
transform 1 0 410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1842_
timestamp 1727493435
transform 1 0 2230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1843_
timestamp 1727493435
transform 1 0 1790 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1844_
timestamp 1727493435
transform -1 0 1970 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1845_
timestamp 1727493435
transform -1 0 2110 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1846_
timestamp 1727493435
transform 1 0 1890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1847_
timestamp 1727493435
transform 1 0 2070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1848_
timestamp 1727493435
transform 1 0 2270 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1849_
timestamp 1727493435
transform -1 0 2130 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1850_
timestamp 1727493435
transform -1 0 1610 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1851_
timestamp 1727493435
transform -1 0 1450 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1852_
timestamp 1727493435
transform 1 0 510 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1853_
timestamp 1727493435
transform -1 0 30 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1854_
timestamp 1727493435
transform -1 0 190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1855_
timestamp 1727493435
transform 1 0 170 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1856_
timestamp 1727493435
transform 1 0 590 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1857_
timestamp 1727493435
transform -1 0 1950 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1858_
timestamp 1727493435
transform -1 0 2150 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1859_
timestamp 1727493435
transform 1 0 2390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1860_
timestamp 1727493435
transform 1 0 670 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1861_
timestamp 1727493435
transform -1 0 810 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1862_
timestamp 1727493435
transform 1 0 1610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1863_
timestamp 1727493435
transform 1 0 2390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1864_
timestamp 1727493435
transform -1 0 30 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1865_
timestamp 1727493435
transform -1 0 350 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1866_
timestamp 1727493435
transform 1 0 10 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1867_
timestamp 1727493435
transform -1 0 610 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1868_
timestamp 1727493435
transform -1 0 3230 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1869_
timestamp 1727493435
transform 1 0 1070 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0__1870_
timestamp 1727493435
transform -1 0 30 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1871_
timestamp 1727493435
transform -1 0 30 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1872_
timestamp 1727493435
transform -1 0 30 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1873_
timestamp 1727493435
transform -1 0 150 0 1 5990
box -6 -8 26 272
use FILL  FILL_0__1874_
timestamp 1727493435
transform -1 0 190 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1875_
timestamp 1727493435
transform -1 0 330 0 1 5470
box -6 -8 26 272
use FILL  FILL_0__1876_
timestamp 1727493435
transform -1 0 210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1877_
timestamp 1727493435
transform 1 0 370 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0__1878_
timestamp 1727493435
transform 1 0 290 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1879_
timestamp 1727493435
transform -1 0 650 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1880_
timestamp 1727493435
transform -1 0 1350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1881_
timestamp 1727493435
transform 1 0 1470 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1882_
timestamp 1727493435
transform -1 0 1030 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1883_
timestamp 1727493435
transform 1 0 1170 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1884_
timestamp 1727493435
transform 1 0 870 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1885_
timestamp 1727493435
transform -1 0 750 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1886_
timestamp 1727493435
transform -1 0 330 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1887_
timestamp 1727493435
transform -1 0 190 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1888_
timestamp 1727493435
transform 1 0 10 0 -1 4950
box -6 -8 26 272
use FILL  FILL_0__1889_
timestamp 1727493435
transform 1 0 330 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1890_
timestamp 1727493435
transform 1 0 470 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1891_
timestamp 1727493435
transform -1 0 170 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1892_
timestamp 1727493435
transform -1 0 170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1893_
timestamp 1727493435
transform 1 0 450 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1894_
timestamp 1727493435
transform -1 0 810 0 1 4430
box -6 -8 26 272
use FILL  FILL_0__1895_
timestamp 1727493435
transform -1 0 30 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0__1896_
timestamp 1727493435
transform -1 0 4450 0 1 4950
box -6 -8 26 272
use FILL  FILL_0__1897_
timestamp 1727493435
transform 1 0 3870 0 1 790
box -6 -8 26 272
use FILL  FILL_0__1898_
timestamp 1727493435
transform 1 0 3570 0 1 2870
box -6 -8 26 272
use FILL  FILL_0__1899_
timestamp 1727493435
transform 1 0 3210 0 -1 270
box -6 -8 26 272
use FILL  FILL_0__1900_
timestamp 1727493435
transform 1 0 3110 0 -1 1830
box -6 -8 26 272
use FILL  FILL_0__1901_
timestamp 1727493435
transform -1 0 2710 0 1 2350
box -6 -8 26 272
use FILL  FILL_0__1902_
timestamp 1727493435
transform -1 0 5090 0 1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1727493435
transform -1 0 2270 0 1 2350
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1727493435
transform -1 0 2210 0 1 3910
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1727493435
transform 1 0 3870 0 1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1727493435
transform 1 0 3550 0 1 2350
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1727493435
transform -1 0 4750 0 1 4950
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1727493435
transform -1 0 4030 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1727493435
transform 1 0 4330 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1727493435
transform -1 0 4070 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert8
timestamp 1727493435
transform -1 0 4130 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert9
timestamp 1727493435
transform -1 0 4610 0 1 4430
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert10
timestamp 1727493435
transform 1 0 5010 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert11
timestamp 1727493435
transform 1 0 4730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1727493435
transform -1 0 3570 0 1 3910
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1727493435
transform 1 0 4190 0 1 3910
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1727493435
transform -1 0 5170 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1727493435
transform -1 0 4890 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1727493435
transform 1 0 3770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1727493435
transform -1 0 3650 0 -1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1727493435
transform -1 0 1890 0 1 2870
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1727493435
transform -1 0 1890 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1727493435
transform -1 0 4590 0 1 4950
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1727493435
transform 1 0 3870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1727493435
transform 1 0 4350 0 1 3910
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1727493435
transform -1 0 3750 0 -1 3390
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1727493435
transform -1 0 2250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1727493435
transform 1 0 2270 0 1 5470
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1727493435
transform 1 0 3070 0 -1 5990
box -6 -8 26 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1727493435
transform -1 0 4090 0 1 5990
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1727493435
transform 1 0 4190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert13
timestamp 1727493435
transform -1 0 4090 0 1 3390
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 3850 0 -1 4430
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 4150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_0_CLKBUF1_insert16
timestamp 1727493435
transform 1 0 4150 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__927_
timestamp 1727493435
transform 1 0 5590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__928_
timestamp 1727493435
transform -1 0 5590 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__929_
timestamp 1727493435
transform -1 0 5870 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__930_
timestamp 1727493435
transform 1 0 5990 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__931_
timestamp 1727493435
transform -1 0 5310 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__932_
timestamp 1727493435
transform -1 0 3410 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__933_
timestamp 1727493435
transform 1 0 5430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__934_
timestamp 1727493435
transform 1 0 5410 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__935_
timestamp 1727493435
transform 1 0 5970 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__936_
timestamp 1727493435
transform -1 0 5350 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__937_
timestamp 1727493435
transform 1 0 5550 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__938_
timestamp 1727493435
transform -1 0 5890 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__939_
timestamp 1727493435
transform 1 0 6010 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__940_
timestamp 1727493435
transform 1 0 6230 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__941_
timestamp 1727493435
transform 1 0 3790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__942_
timestamp 1727493435
transform 1 0 5710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__943_
timestamp 1727493435
transform 1 0 5970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__944_
timestamp 1727493435
transform 1 0 5710 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__945_
timestamp 1727493435
transform 1 0 6230 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__946_
timestamp 1727493435
transform -1 0 5770 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__947_
timestamp 1727493435
transform 1 0 5730 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__948_
timestamp 1727493435
transform -1 0 5910 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__949_
timestamp 1727493435
transform 1 0 5870 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__950_
timestamp 1727493435
transform -1 0 5630 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__951_
timestamp 1727493435
transform -1 0 6110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__952_
timestamp 1727493435
transform -1 0 5650 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__953_
timestamp 1727493435
transform 1 0 5190 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__954_
timestamp 1727493435
transform 1 0 6250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__955_
timestamp 1727493435
transform 1 0 6170 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__956_
timestamp 1727493435
transform -1 0 5790 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__957_
timestamp 1727493435
transform -1 0 5490 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__958_
timestamp 1727493435
transform 1 0 6270 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__959_
timestamp 1727493435
transform -1 0 6110 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__960_
timestamp 1727493435
transform 1 0 6050 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__961_
timestamp 1727493435
transform -1 0 6090 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__962_
timestamp 1727493435
transform 1 0 5810 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__963_
timestamp 1727493435
transform -1 0 5490 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__964_
timestamp 1727493435
transform -1 0 5330 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__965_
timestamp 1727493435
transform 1 0 4470 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__966_
timestamp 1727493435
transform -1 0 4630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__967_
timestamp 1727493435
transform 1 0 4910 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__968_
timestamp 1727493435
transform 1 0 5130 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__969_
timestamp 1727493435
transform 1 0 5010 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__970_
timestamp 1727493435
transform 1 0 4050 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__971_
timestamp 1727493435
transform 1 0 4830 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__972_
timestamp 1727493435
transform 1 0 4670 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__973_
timestamp 1727493435
transform 1 0 4330 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__974_
timestamp 1727493435
transform 1 0 4350 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__975_
timestamp 1727493435
transform 1 0 4410 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__976_
timestamp 1727493435
transform 1 0 3670 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__977_
timestamp 1727493435
transform 1 0 3950 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__978_
timestamp 1727493435
transform 1 0 3710 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__979_
timestamp 1727493435
transform 1 0 3150 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__980_
timestamp 1727493435
transform 1 0 3290 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__981_
timestamp 1727493435
transform -1 0 3150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__982_
timestamp 1727493435
transform 1 0 2050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__983_
timestamp 1727493435
transform 1 0 2670 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__984_
timestamp 1727493435
transform -1 0 2830 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__985_
timestamp 1727493435
transform 1 0 3610 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__986_
timestamp 1727493435
transform 1 0 3890 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__987_
timestamp 1727493435
transform -1 0 4070 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__988_
timestamp 1727493435
transform -1 0 2310 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__989_
timestamp 1727493435
transform 1 0 5230 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__990_
timestamp 1727493435
transform -1 0 1750 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__991_
timestamp 1727493435
transform 1 0 5570 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__992_
timestamp 1727493435
transform 1 0 5410 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__993_
timestamp 1727493435
transform 1 0 5710 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__994_
timestamp 1727493435
transform -1 0 4290 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__995_
timestamp 1727493435
transform -1 0 4610 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__996_
timestamp 1727493435
transform 1 0 6250 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__997_
timestamp 1727493435
transform 1 0 5450 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__998_
timestamp 1727493435
transform -1 0 6250 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__999_
timestamp 1727493435
transform 1 0 6070 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1000_
timestamp 1727493435
transform -1 0 4870 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1001_
timestamp 1727493435
transform 1 0 5310 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1002_
timestamp 1727493435
transform 1 0 4650 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1003_
timestamp 1727493435
transform 1 0 4730 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1004_
timestamp 1727493435
transform 1 0 4650 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1005_
timestamp 1727493435
transform -1 0 5210 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1006_
timestamp 1727493435
transform 1 0 5590 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1007_
timestamp 1727493435
transform -1 0 4910 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1008_
timestamp 1727493435
transform -1 0 5030 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1009_
timestamp 1727493435
transform 1 0 5910 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1010_
timestamp 1727493435
transform -1 0 5350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1011_
timestamp 1727493435
transform 1 0 4930 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1012_
timestamp 1727493435
transform -1 0 3470 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1013_
timestamp 1727493435
transform -1 0 4330 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1014_
timestamp 1727493435
transform 1 0 5250 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1015_
timestamp 1727493435
transform 1 0 5250 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1016_
timestamp 1727493435
transform -1 0 5770 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1017_
timestamp 1727493435
transform 1 0 5590 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1018_
timestamp 1727493435
transform 1 0 5030 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1019_
timestamp 1727493435
transform 1 0 3950 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1020_
timestamp 1727493435
transform 1 0 4130 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1021_
timestamp 1727493435
transform -1 0 4190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1022_
timestamp 1727493435
transform 1 0 4510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1023_
timestamp 1727493435
transform -1 0 4050 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1024_
timestamp 1727493435
transform -1 0 4810 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1025_
timestamp 1727493435
transform 1 0 4630 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1026_
timestamp 1727493435
transform -1 0 4510 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1027_
timestamp 1727493435
transform 1 0 4790 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1028_
timestamp 1727493435
transform 1 0 4910 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1029_
timestamp 1727493435
transform 1 0 5230 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1030_
timestamp 1727493435
transform -1 0 5210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1031_
timestamp 1727493435
transform -1 0 4690 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1032_
timestamp 1727493435
transform -1 0 4370 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1033_
timestamp 1727493435
transform 1 0 4830 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1034_
timestamp 1727493435
transform -1 0 4310 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1035_
timestamp 1727493435
transform 1 0 4610 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1036_
timestamp 1727493435
transform 1 0 4450 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1037_
timestamp 1727493435
transform -1 0 5130 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1038_
timestamp 1727493435
transform 1 0 4530 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1039_
timestamp 1727493435
transform 1 0 4770 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1040_
timestamp 1727493435
transform 1 0 4730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1041_
timestamp 1727493435
transform 1 0 4930 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1042_
timestamp 1727493435
transform 1 0 5490 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1043_
timestamp 1727493435
transform -1 0 5050 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1044_
timestamp 1727493435
transform 1 0 4890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1045_
timestamp 1727493435
transform 1 0 5210 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1046_
timestamp 1727493435
transform 1 0 5630 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1047_
timestamp 1727493435
transform 1 0 4990 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1048_
timestamp 1727493435
transform 1 0 5070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1049_
timestamp 1727493435
transform 1 0 5050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1050_
timestamp 1727493435
transform 1 0 5310 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1051_
timestamp 1727493435
transform 1 0 5790 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1052_
timestamp 1727493435
transform 1 0 5950 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1053_
timestamp 1727493435
transform 1 0 6350 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1054_
timestamp 1727493435
transform 1 0 5390 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1055_
timestamp 1727493435
transform -1 0 4210 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1056_
timestamp 1727493435
transform -1 0 2890 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1057_
timestamp 1727493435
transform -1 0 4030 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1058_
timestamp 1727493435
transform -1 0 4210 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1059_
timestamp 1727493435
transform 1 0 3110 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1060_
timestamp 1727493435
transform 1 0 3870 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1061_
timestamp 1727493435
transform 1 0 4030 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1062_
timestamp 1727493435
transform 1 0 4290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1063_
timestamp 1727493435
transform -1 0 4310 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1064_
timestamp 1727493435
transform -1 0 3990 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1065_
timestamp 1727493435
transform -1 0 3910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1066_
timestamp 1727493435
transform -1 0 4170 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1067_
timestamp 1727493435
transform 1 0 4030 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1068_
timestamp 1727493435
transform -1 0 4590 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1069_
timestamp 1727493435
transform -1 0 4330 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1070_
timestamp 1727493435
transform 1 0 4510 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1071_
timestamp 1727493435
transform 1 0 4730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1072_
timestamp 1727493435
transform 1 0 4410 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1073_
timestamp 1727493435
transform 1 0 5070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1074_
timestamp 1727493435
transform 1 0 4430 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1075_
timestamp 1727493435
transform -1 0 4750 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1076_
timestamp 1727493435
transform -1 0 4590 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1077_
timestamp 1727493435
transform 1 0 4450 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1078_
timestamp 1727493435
transform -1 0 4750 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1079_
timestamp 1727493435
transform 1 0 3750 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1080_
timestamp 1727493435
transform -1 0 5210 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1081_
timestamp 1727493435
transform -1 0 4890 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1082_
timestamp 1727493435
transform 1 0 5050 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1083_
timestamp 1727493435
transform 1 0 4410 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1084_
timestamp 1727493435
transform 1 0 4610 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1085_
timestamp 1727493435
transform 1 0 4570 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1086_
timestamp 1727493435
transform 1 0 5390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1087_
timestamp 1727493435
transform 1 0 5130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1088_
timestamp 1727493435
transform 1 0 4910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1089_
timestamp 1727493435
transform 1 0 4470 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1090_
timestamp 1727493435
transform -1 0 5250 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1091_
timestamp 1727493435
transform 1 0 4810 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1092_
timestamp 1727493435
transform 1 0 5470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1093_
timestamp 1727493435
transform 1 0 5150 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1094_
timestamp 1727493435
transform 1 0 4810 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1095_
timestamp 1727493435
transform 1 0 4990 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1096_
timestamp 1727493435
transform 1 0 5310 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1097_
timestamp 1727493435
transform -1 0 1590 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1098_
timestamp 1727493435
transform 1 0 5570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1099_
timestamp 1727493435
transform 1 0 5330 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1100_
timestamp 1727493435
transform -1 0 5490 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1101_
timestamp 1727493435
transform 1 0 5610 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1102_
timestamp 1727493435
transform 1 0 5790 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1103_
timestamp 1727493435
transform 1 0 6090 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1104_
timestamp 1727493435
transform 1 0 5150 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1105_
timestamp 1727493435
transform 1 0 5290 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1106_
timestamp 1727493435
transform -1 0 5970 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1107_
timestamp 1727493435
transform -1 0 6130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1108_
timestamp 1727493435
transform 1 0 6370 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1109_
timestamp 1727493435
transform 1 0 6250 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1110_
timestamp 1727493435
transform -1 0 5810 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1111_
timestamp 1727493435
transform 1 0 4970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1112_
timestamp 1727493435
transform -1 0 4250 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1113_
timestamp 1727493435
transform -1 0 3750 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1114_
timestamp 1727493435
transform -1 0 3570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1115_
timestamp 1727493435
transform -1 0 3150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1116_
timestamp 1727493435
transform -1 0 3250 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1117_
timestamp 1727493435
transform -1 0 3450 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1118_
timestamp 1727493435
transform 1 0 3730 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1119_
timestamp 1727493435
transform -1 0 3750 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1120_
timestamp 1727493435
transform -1 0 3830 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1121_
timestamp 1727493435
transform -1 0 3570 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1122_
timestamp 1727493435
transform 1 0 4210 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1123_
timestamp 1727493435
transform 1 0 3710 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1124_
timestamp 1727493435
transform -1 0 3270 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1125_
timestamp 1727493435
transform -1 0 4370 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1126_
timestamp 1727493435
transform -1 0 3410 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1127_
timestamp 1727493435
transform -1 0 3410 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1128_
timestamp 1727493435
transform 1 0 3650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1129_
timestamp 1727493435
transform 1 0 3970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1130_
timestamp 1727493435
transform 1 0 3870 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1131_
timestamp 1727493435
transform -1 0 3470 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1132_
timestamp 1727493435
transform 1 0 3530 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1133_
timestamp 1727493435
transform 1 0 3650 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1134_
timestamp 1727493435
transform -1 0 3350 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1135_
timestamp 1727493435
transform 1 0 3530 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1136_
timestamp 1727493435
transform -1 0 4150 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1137_
timestamp 1727493435
transform 1 0 3710 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1138_
timestamp 1727493435
transform 1 0 4010 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1139_
timestamp 1727493435
transform 1 0 4570 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1140_
timestamp 1727493435
transform 1 0 4150 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1141_
timestamp 1727493435
transform 1 0 4190 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1142_
timestamp 1727493435
transform -1 0 4050 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1143_
timestamp 1727493435
transform -1 0 3890 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1144_
timestamp 1727493435
transform 1 0 4730 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1145_
timestamp 1727493435
transform 1 0 5050 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1146_
timestamp 1727493435
transform -1 0 4650 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1147_
timestamp 1727493435
transform 1 0 4690 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1148_
timestamp 1727493435
transform 1 0 4530 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1149_
timestamp 1727493435
transform 1 0 5010 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1150_
timestamp 1727493435
transform -1 0 5190 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1151_
timestamp 1727493435
transform -1 0 5770 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1152_
timestamp 1727493435
transform 1 0 4870 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1153_
timestamp 1727493435
transform 1 0 6350 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1154_
timestamp 1727493435
transform 1 0 6050 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1155_
timestamp 1727493435
transform -1 0 5990 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1156_
timestamp 1727493435
transform 1 0 6110 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1157_
timestamp 1727493435
transform 1 0 5870 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1158_
timestamp 1727493435
transform 1 0 6210 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1159_
timestamp 1727493435
transform 1 0 5410 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1160_
timestamp 1727493435
transform -1 0 5270 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1161_
timestamp 1727493435
transform -1 0 5110 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1162_
timestamp 1727493435
transform 1 0 5210 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1163_
timestamp 1727493435
transform 1 0 4850 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1164_
timestamp 1727493435
transform 1 0 4890 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1165_
timestamp 1727493435
transform -1 0 5590 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1166_
timestamp 1727493435
transform -1 0 5650 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1167_
timestamp 1727493435
transform 1 0 5490 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1168_
timestamp 1727493435
transform 1 0 5550 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1169_
timestamp 1727493435
transform 1 0 5810 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1170_
timestamp 1727493435
transform -1 0 5650 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1171_
timestamp 1727493435
transform -1 0 5350 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1172_
timestamp 1727493435
transform 1 0 5370 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1173_
timestamp 1727493435
transform 1 0 5650 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1174_
timestamp 1727493435
transform 1 0 6070 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1175_
timestamp 1727493435
transform 1 0 5490 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1176_
timestamp 1727493435
transform 1 0 5730 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1177_
timestamp 1727493435
transform 1 0 6290 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1178_
timestamp 1727493435
transform 1 0 6350 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1179_
timestamp 1727493435
transform 1 0 5710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1180_
timestamp 1727493435
transform 1 0 6390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1181_
timestamp 1727493435
transform 1 0 6110 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1182_
timestamp 1727493435
transform -1 0 5810 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1183_
timestamp 1727493435
transform -1 0 4530 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1184_
timestamp 1727493435
transform 1 0 4410 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1185_
timestamp 1727493435
transform 1 0 5950 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1186_
timestamp 1727493435
transform 1 0 5370 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1187_
timestamp 1727493435
transform 1 0 5530 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1188_
timestamp 1727493435
transform 1 0 5710 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1189_
timestamp 1727493435
transform -1 0 5570 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1190_
timestamp 1727493435
transform 1 0 5870 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1191_
timestamp 1727493435
transform -1 0 5770 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1192_
timestamp 1727493435
transform 1 0 5470 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1193_
timestamp 1727493435
transform 1 0 5390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1194_
timestamp 1727493435
transform 1 0 5710 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1195_
timestamp 1727493435
transform 1 0 6250 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1196_
timestamp 1727493435
transform 1 0 6270 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1197_
timestamp 1727493435
transform 1 0 5950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1198_
timestamp 1727493435
transform 1 0 6250 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1199_
timestamp 1727493435
transform -1 0 6250 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1200_
timestamp 1727493435
transform 1 0 5970 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1201_
timestamp 1727493435
transform 1 0 6130 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1202_
timestamp 1727493435
transform 1 0 5930 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1203_
timestamp 1727493435
transform -1 0 5810 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1204_
timestamp 1727493435
transform 1 0 5010 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1205_
timestamp 1727493435
transform 1 0 5430 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1206_
timestamp 1727493435
transform -1 0 5170 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1207_
timestamp 1727493435
transform 1 0 5610 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1208_
timestamp 1727493435
transform -1 0 5930 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1209_
timestamp 1727493435
transform -1 0 5470 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1210_
timestamp 1727493435
transform -1 0 5630 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1211_
timestamp 1727493435
transform 1 0 5430 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1212_
timestamp 1727493435
transform -1 0 5450 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1213_
timestamp 1727493435
transform 1 0 6110 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1214_
timestamp 1727493435
transform 1 0 6290 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1215_
timestamp 1727493435
transform -1 0 5890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1216_
timestamp 1727493435
transform 1 0 6050 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1217_
timestamp 1727493435
transform -1 0 6230 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1218_
timestamp 1727493435
transform 1 0 6310 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1219_
timestamp 1727493435
transform -1 0 6150 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1220_
timestamp 1727493435
transform -1 0 4750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1221_
timestamp 1727493435
transform -1 0 4870 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1222_
timestamp 1727493435
transform 1 0 6270 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1223_
timestamp 1727493435
transform -1 0 6330 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1224_
timestamp 1727493435
transform 1 0 6150 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1225_
timestamp 1727493435
transform -1 0 6150 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1226_
timestamp 1727493435
transform 1 0 4750 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1227_
timestamp 1727493435
transform -1 0 5530 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1228_
timestamp 1727493435
transform -1 0 5990 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1229_
timestamp 1727493435
transform 1 0 5810 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1230_
timestamp 1727493435
transform 1 0 5330 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1231_
timestamp 1727493435
transform -1 0 5050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1232_
timestamp 1727493435
transform 1 0 5150 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1233_
timestamp 1727493435
transform -1 0 5190 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1234_
timestamp 1727493435
transform 1 0 6030 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1235_
timestamp 1727493435
transform 1 0 6190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1236_
timestamp 1727493435
transform 1 0 6070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1237_
timestamp 1727493435
transform -1 0 6310 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1238_
timestamp 1727493435
transform -1 0 6150 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1239_
timestamp 1727493435
transform 1 0 5890 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1240_
timestamp 1727493435
transform 1 0 5870 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1241_
timestamp 1727493435
transform -1 0 5990 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1242_
timestamp 1727493435
transform 1 0 5810 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1243_
timestamp 1727493435
transform -1 0 5850 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1244_
timestamp 1727493435
transform -1 0 5930 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1245_
timestamp 1727493435
transform -1 0 4970 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1246_
timestamp 1727493435
transform -1 0 5350 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1247_
timestamp 1727493435
transform 1 0 4370 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1248_
timestamp 1727493435
transform -1 0 4210 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1249_
timestamp 1727493435
transform 1 0 4670 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1250_
timestamp 1727493435
transform 1 0 3810 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1251_
timestamp 1727493435
transform 1 0 4790 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1252_
timestamp 1727493435
transform -1 0 4490 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1253_
timestamp 1727493435
transform 1 0 4310 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1254_
timestamp 1727493435
transform 1 0 4990 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1255_
timestamp 1727493435
transform 1 0 4850 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1256_
timestamp 1727493435
transform -1 0 4710 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1257_
timestamp 1727493435
transform 1 0 4370 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1258_
timestamp 1727493435
transform -1 0 4410 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1259_
timestamp 1727493435
transform 1 0 2570 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1260_
timestamp 1727493435
transform -1 0 3190 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1261_
timestamp 1727493435
transform 1 0 3010 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1262_
timestamp 1727493435
transform -1 0 3110 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1263_
timestamp 1727493435
transform 1 0 2770 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1264_
timestamp 1727493435
transform 1 0 2850 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1265_
timestamp 1727493435
transform -1 0 2190 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1266_
timestamp 1727493435
transform -1 0 2950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1267_
timestamp 1727493435
transform 1 0 3270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1268_
timestamp 1727493435
transform -1 0 2490 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1269_
timestamp 1727493435
transform -1 0 2610 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1270_
timestamp 1727493435
transform 1 0 2710 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1271_
timestamp 1727493435
transform -1 0 3590 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1272_
timestamp 1727493435
transform 1 0 2730 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1273_
timestamp 1727493435
transform -1 0 2790 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1274_
timestamp 1727493435
transform -1 0 3070 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1275_
timestamp 1727493435
transform 1 0 3050 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1276_
timestamp 1727493435
transform 1 0 3270 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1277_
timestamp 1727493435
transform 1 0 3210 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1278_
timestamp 1727493435
transform 1 0 3270 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1279_
timestamp 1727493435
transform -1 0 3410 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1280_
timestamp 1727493435
transform -1 0 3010 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1281_
timestamp 1727493435
transform 1 0 3090 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1282_
timestamp 1727493435
transform -1 0 2930 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1283_
timestamp 1727493435
transform 1 0 2850 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1284_
timestamp 1727493435
transform 1 0 3410 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1285_
timestamp 1727493435
transform 1 0 3430 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1286_
timestamp 1727493435
transform 1 0 3910 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1287_
timestamp 1727493435
transform -1 0 4250 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1288_
timestamp 1727493435
transform 1 0 3070 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1289_
timestamp 1727493435
transform -1 0 2950 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1290_
timestamp 1727493435
transform 1 0 4070 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1291_
timestamp 1727493435
transform -1 0 3870 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1292_
timestamp 1727493435
transform 1 0 4510 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1293_
timestamp 1727493435
transform 1 0 3750 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1294_
timestamp 1727493435
transform 1 0 3690 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1295_
timestamp 1727493435
transform -1 0 3350 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1296_
timestamp 1727493435
transform -1 0 3390 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1297_
timestamp 1727493435
transform -1 0 5190 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1298_
timestamp 1727493435
transform -1 0 4210 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1299_
timestamp 1727493435
transform 1 0 4010 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1300_
timestamp 1727493435
transform -1 0 3890 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1301_
timestamp 1727493435
transform 1 0 2450 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1302_
timestamp 1727493435
transform -1 0 2630 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1303_
timestamp 1727493435
transform -1 0 3710 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1304_
timestamp 1727493435
transform 1 0 4030 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1305_
timestamp 1727493435
transform -1 0 2750 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1306_
timestamp 1727493435
transform 1 0 2590 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1307_
timestamp 1727493435
transform -1 0 5810 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1308_
timestamp 1727493435
transform 1 0 2890 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1309_
timestamp 1727493435
transform 1 0 2290 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1310_
timestamp 1727493435
transform -1 0 2770 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1311_
timestamp 1727493435
transform -1 0 2490 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1312_
timestamp 1727493435
transform -1 0 2370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1313_
timestamp 1727493435
transform -1 0 6210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1314_
timestamp 1727493435
transform -1 0 6330 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1315_
timestamp 1727493435
transform 1 0 6370 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1316_
timestamp 1727493435
transform -1 0 6290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1317_
timestamp 1727493435
transform -1 0 5950 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1318_
timestamp 1727493435
transform 1 0 6090 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1319_
timestamp 1727493435
transform -1 0 5630 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1320_
timestamp 1727493435
transform -1 0 5510 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1321_
timestamp 1727493435
transform 1 0 2570 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1322_
timestamp 1727493435
transform 1 0 2830 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1323_
timestamp 1727493435
transform -1 0 2430 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1324_
timestamp 1727493435
transform -1 0 2790 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1325_
timestamp 1727493435
transform -1 0 2930 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1326_
timestamp 1727493435
transform 1 0 2730 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1327_
timestamp 1727493435
transform -1 0 3530 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1328_
timestamp 1727493435
transform 1 0 2830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1329_
timestamp 1727493435
transform -1 0 2910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1330_
timestamp 1727493435
transform 1 0 2810 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1331_
timestamp 1727493435
transform 1 0 2650 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1332_
timestamp 1727493435
transform 1 0 2190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1333_
timestamp 1727493435
transform 1 0 2030 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1334_
timestamp 1727493435
transform -1 0 2510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1335_
timestamp 1727493435
transform 1 0 2170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1336_
timestamp 1727493435
transform -1 0 3550 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1337_
timestamp 1727493435
transform 1 0 3050 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1338_
timestamp 1727493435
transform -1 0 4650 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1339_
timestamp 1727493435
transform -1 0 3610 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1340_
timestamp 1727493435
transform -1 0 3530 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1341_
timestamp 1727493435
transform -1 0 2810 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1342_
timestamp 1727493435
transform -1 0 2690 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1343_
timestamp 1727493435
transform -1 0 3010 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1344_
timestamp 1727493435
transform -1 0 2310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1345_
timestamp 1727493435
transform -1 0 2350 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1346_
timestamp 1727493435
transform 1 0 2230 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1347_
timestamp 1727493435
transform -1 0 2530 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1348_
timestamp 1727493435
transform -1 0 1930 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1349_
timestamp 1727493435
transform -1 0 2110 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1350_
timestamp 1727493435
transform 1 0 2190 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1351_
timestamp 1727493435
transform 1 0 2050 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1352_
timestamp 1727493435
transform 1 0 3270 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1353_
timestamp 1727493435
transform -1 0 2770 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1354_
timestamp 1727493435
transform -1 0 1510 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1355_
timestamp 1727493435
transform -1 0 1270 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1356_
timestamp 1727493435
transform 1 0 1810 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1357_
timestamp 1727493435
transform -1 0 2130 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1358_
timestamp 1727493435
transform 1 0 1970 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1359_
timestamp 1727493435
transform 1 0 1290 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1360_
timestamp 1727493435
transform -1 0 950 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1361_
timestamp 1727493435
transform 1 0 1210 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1362_
timestamp 1727493435
transform 1 0 1310 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1363_
timestamp 1727493435
transform 1 0 1630 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1364_
timestamp 1727493435
transform -1 0 2430 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1365_
timestamp 1727493435
transform -1 0 1410 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1366_
timestamp 1727493435
transform -1 0 1370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1367_
timestamp 1727493435
transform 1 0 1550 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1368_
timestamp 1727493435
transform -1 0 1070 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1369_
timestamp 1727493435
transform 1 0 1550 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1370_
timestamp 1727493435
transform -1 0 1390 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1371_
timestamp 1727493435
transform -1 0 1450 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1372_
timestamp 1727493435
transform 1 0 2150 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1373_
timestamp 1727493435
transform 1 0 2910 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1374_
timestamp 1727493435
transform 1 0 2390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1375_
timestamp 1727493435
transform 1 0 1750 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1376_
timestamp 1727493435
transform 1 0 1830 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1377_
timestamp 1727493435
transform -1 0 1910 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1378_
timestamp 1727493435
transform 1 0 1570 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1379_
timestamp 1727493435
transform 1 0 1570 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1380_
timestamp 1727493435
transform -1 0 1470 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1381_
timestamp 1727493435
transform -1 0 870 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1382_
timestamp 1727493435
transform -1 0 3110 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1383_
timestamp 1727493435
transform -1 0 2950 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1384_
timestamp 1727493435
transform 1 0 1610 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1385_
timestamp 1727493435
transform 1 0 1710 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1386_
timestamp 1727493435
transform -1 0 2610 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1387_
timestamp 1727493435
transform 1 0 1990 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1388_
timestamp 1727493435
transform -1 0 1310 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1389_
timestamp 1727493435
transform -1 0 1170 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1390_
timestamp 1727493435
transform -1 0 1050 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1391_
timestamp 1727493435
transform 1 0 1130 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1392_
timestamp 1727493435
transform 1 0 1770 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1393_
timestamp 1727493435
transform 1 0 1490 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1394_
timestamp 1727493435
transform 1 0 1850 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1395_
timestamp 1727493435
transform 1 0 1330 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1396_
timestamp 1727493435
transform 1 0 1930 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1397_
timestamp 1727493435
transform -1 0 2290 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1398_
timestamp 1727493435
transform 1 0 2450 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1399_
timestamp 1727493435
transform 1 0 2490 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1400_
timestamp 1727493435
transform -1 0 2670 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1401_
timestamp 1727493435
transform -1 0 2030 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1402_
timestamp 1727493435
transform -1 0 2150 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1403_
timestamp 1727493435
transform 1 0 2110 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1404_
timestamp 1727493435
transform 1 0 1670 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1405_
timestamp 1727493435
transform 1 0 2450 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1406_
timestamp 1727493435
transform -1 0 2590 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1407_
timestamp 1727493435
transform -1 0 2550 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1408_
timestamp 1727493435
transform -1 0 4850 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1409_
timestamp 1727493435
transform 1 0 4310 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1410_
timestamp 1727493435
transform -1 0 4690 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1411_
timestamp 1727493435
transform -1 0 4510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1412_
timestamp 1727493435
transform -1 0 3230 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1413_
timestamp 1727493435
transform 1 0 2550 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1414_
timestamp 1727493435
transform -1 0 5290 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1415_
timestamp 1727493435
transform -1 0 2190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1416_
timestamp 1727493435
transform -1 0 2310 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1417_
timestamp 1727493435
transform 1 0 1850 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1418_
timestamp 1727493435
transform 1 0 2350 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1419_
timestamp 1727493435
transform -1 0 1310 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1420_
timestamp 1727493435
transform -1 0 1510 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1421_
timestamp 1727493435
transform -1 0 930 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1422_
timestamp 1727493435
transform 1 0 1010 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1423_
timestamp 1727493435
transform -1 0 650 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1424_
timestamp 1727493435
transform -1 0 1110 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1425_
timestamp 1727493435
transform -1 0 450 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1426_
timestamp 1727493435
transform 1 0 730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1427_
timestamp 1727493435
transform -1 0 870 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1428_
timestamp 1727493435
transform 1 0 570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1429_
timestamp 1727493435
transform -1 0 310 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1430_
timestamp 1727493435
transform 1 0 670 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1431_
timestamp 1727493435
transform 1 0 830 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1432_
timestamp 1727493435
transform 1 0 1550 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1433_
timestamp 1727493435
transform -1 0 810 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1434_
timestamp 1727493435
transform -1 0 350 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1435_
timestamp 1727493435
transform -1 0 970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1436_
timestamp 1727493435
transform 1 0 970 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1437_
timestamp 1727493435
transform 1 0 810 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1438_
timestamp 1727493435
transform -1 0 190 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1439_
timestamp 1727493435
transform 1 0 1110 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1440_
timestamp 1727493435
transform -1 0 50 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1441_
timestamp 1727493435
transform -1 0 170 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1442_
timestamp 1727493435
transform -1 0 490 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1443_
timestamp 1727493435
transform -1 0 370 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1444_
timestamp 1727493435
transform -1 0 510 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1445_
timestamp 1727493435
transform -1 0 670 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1446_
timestamp 1727493435
transform -1 0 50 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1447_
timestamp 1727493435
transform 1 0 310 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1448_
timestamp 1727493435
transform -1 0 670 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1449_
timestamp 1727493435
transform 1 0 970 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1450_
timestamp 1727493435
transform -1 0 210 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1451_
timestamp 1727493435
transform 1 0 470 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1452_
timestamp 1727493435
transform 1 0 810 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1453_
timestamp 1727493435
transform -1 0 1670 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1454_
timestamp 1727493435
transform -1 0 650 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1455_
timestamp 1727493435
transform 1 0 190 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1456_
timestamp 1727493435
transform -1 0 50 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1457_
timestamp 1727493435
transform 1 0 350 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1458_
timestamp 1727493435
transform 1 0 670 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1459_
timestamp 1727493435
transform -1 0 530 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1460_
timestamp 1727493435
transform 1 0 1150 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1461_
timestamp 1727493435
transform 1 0 830 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1462_
timestamp 1727493435
transform -1 0 1350 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1463_
timestamp 1727493435
transform -1 0 50 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1464_
timestamp 1727493435
transform -1 0 190 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1465_
timestamp 1727493435
transform -1 0 710 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1466_
timestamp 1727493435
transform -1 0 550 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1467_
timestamp 1727493435
transform 1 0 350 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1468_
timestamp 1727493435
transform -1 0 1010 0 1 270
box -6 -8 26 272
use FILL  FILL_1__1469_
timestamp 1727493435
transform -1 0 1550 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1470_
timestamp 1727493435
transform -1 0 2050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1471_
timestamp 1727493435
transform -1 0 1870 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1472_
timestamp 1727493435
transform -1 0 1070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1473_
timestamp 1727493435
transform 1 0 2110 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1474_
timestamp 1727493435
transform 1 0 2250 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1475_
timestamp 1727493435
transform -1 0 2590 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1476_
timestamp 1727493435
transform 1 0 3070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1477_
timestamp 1727493435
transform -1 0 5670 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1478_
timestamp 1727493435
transform -1 0 5370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1479_
timestamp 1727493435
transform -1 0 2190 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1480_
timestamp 1727493435
transform 1 0 3190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1481_
timestamp 1727493435
transform -1 0 3230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1482_
timestamp 1727493435
transform 1 0 4070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1483_
timestamp 1727493435
transform 1 0 3530 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1484_
timestamp 1727493435
transform 1 0 1170 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1485_
timestamp 1727493435
transform 1 0 2330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1486_
timestamp 1727493435
transform 1 0 1410 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1487_
timestamp 1727493435
transform -1 0 530 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1488_
timestamp 1727493435
transform 1 0 530 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1489_
timestamp 1727493435
transform -1 0 50 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1490_
timestamp 1727493435
transform -1 0 1470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1491_
timestamp 1727493435
transform 1 0 910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1492_
timestamp 1727493435
transform -1 0 850 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1493_
timestamp 1727493435
transform -1 0 650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1494_
timestamp 1727493435
transform -1 0 490 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1495_
timestamp 1727493435
transform -1 0 330 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1496_
timestamp 1727493435
transform -1 0 390 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1497_
timestamp 1727493435
transform 1 0 1090 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1498_
timestamp 1727493435
transform -1 0 550 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1499_
timestamp 1727493435
transform 1 0 670 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1500_
timestamp 1727493435
transform 1 0 1150 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1501_
timestamp 1727493435
transform 1 0 1290 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1502_
timestamp 1727493435
transform -1 0 1050 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1503_
timestamp 1727493435
transform -1 0 630 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1504_
timestamp 1727493435
transform 1 0 890 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1505_
timestamp 1727493435
transform -1 0 730 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1506_
timestamp 1727493435
transform -1 0 570 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1507_
timestamp 1727493435
transform -1 0 230 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1508_
timestamp 1727493435
transform -1 0 50 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1509_
timestamp 1727493435
transform -1 0 50 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1510_
timestamp 1727493435
transform 1 0 30 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1511_
timestamp 1727493435
transform -1 0 170 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1512_
timestamp 1727493435
transform -1 0 50 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1513_
timestamp 1727493435
transform 1 0 210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1514_
timestamp 1727493435
transform -1 0 390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1515_
timestamp 1727493435
transform 1 0 190 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1516_
timestamp 1727493435
transform -1 0 50 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1517_
timestamp 1727493435
transform -1 0 370 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1518_
timestamp 1727493435
transform -1 0 830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1519_
timestamp 1727493435
transform -1 0 1130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1520_
timestamp 1727493435
transform 1 0 970 0 -1 790
box -6 -8 26 272
use FILL  FILL_1__1521_
timestamp 1727493435
transform 1 0 1130 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1522_
timestamp 1727493435
transform 1 0 950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1523_
timestamp 1727493435
transform -1 0 1290 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1524_
timestamp 1727493435
transform 1 0 1690 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1525_
timestamp 1727493435
transform 1 0 1950 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1526_
timestamp 1727493435
transform -1 0 1890 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1527_
timestamp 1727493435
transform 1 0 1990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1528_
timestamp 1727493435
transform 1 0 2690 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1529_
timestamp 1727493435
transform -1 0 5050 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1530_
timestamp 1727493435
transform -1 0 4910 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1531_
timestamp 1727493435
transform -1 0 4590 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1532_
timestamp 1727493435
transform 1 0 3070 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1533_
timestamp 1727493435
transform -1 0 3310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1534_
timestamp 1727493435
transform 1 0 3450 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1535_
timestamp 1727493435
transform -1 0 3110 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1536_
timestamp 1727493435
transform 1 0 3470 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1537_
timestamp 1727493435
transform -1 0 170 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1538_
timestamp 1727493435
transform 1 0 1170 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1539_
timestamp 1727493435
transform -1 0 750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1540_
timestamp 1727493435
transform -1 0 630 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1541_
timestamp 1727493435
transform 1 0 970 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1542_
timestamp 1727493435
transform 1 0 990 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1543_
timestamp 1727493435
transform 1 0 830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1544_
timestamp 1727493435
transform 1 0 890 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1545_
timestamp 1727493435
transform -1 0 750 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1546_
timestamp 1727493435
transform 1 0 450 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1547_
timestamp 1727493435
transform -1 0 690 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1548_
timestamp 1727493435
transform -1 0 830 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1549_
timestamp 1727493435
transform 1 0 310 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1550_
timestamp 1727493435
transform -1 0 670 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1551_
timestamp 1727493435
transform -1 0 50 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1552_
timestamp 1727493435
transform 1 0 150 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1553_
timestamp 1727493435
transform 1 0 30 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1554_
timestamp 1727493435
transform -1 0 50 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1555_
timestamp 1727493435
transform 1 0 190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1556_
timestamp 1727493435
transform 1 0 290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1557_
timestamp 1727493435
transform 1 0 30 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1558_
timestamp 1727493435
transform -1 0 190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1559_
timestamp 1727493435
transform -1 0 470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1560_
timestamp 1727493435
transform 1 0 1030 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1561_
timestamp 1727493435
transform 1 0 1290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1562_
timestamp 1727493435
transform 1 0 1010 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1563_
timestamp 1727493435
transform -1 0 1450 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1564_
timestamp 1727493435
transform 1 0 2630 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1565_
timestamp 1727493435
transform -1 0 1430 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1566_
timestamp 1727493435
transform 1 0 2170 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1567_
timestamp 1727493435
transform 1 0 1270 0 -1 1310
box -6 -8 26 272
use FILL  FILL_1__1568_
timestamp 1727493435
transform 1 0 1970 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1569_
timestamp 1727493435
transform 1 0 2250 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1570_
timestamp 1727493435
transform 1 0 2410 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1571_
timestamp 1727493435
transform -1 0 1150 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1572_
timestamp 1727493435
transform -1 0 1190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1573_
timestamp 1727493435
transform -1 0 1710 0 1 1310
box -6 -8 26 272
use FILL  FILL_1__1574_
timestamp 1727493435
transform -1 0 1710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1575_
timestamp 1727493435
transform 1 0 2090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1576_
timestamp 1727493435
transform 1 0 2350 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1577_
timestamp 1727493435
transform -1 0 1750 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1578_
timestamp 1727493435
transform 1 0 2510 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1579_
timestamp 1727493435
transform 1 0 6390 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1580_
timestamp 1727493435
transform 1 0 6210 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1581_
timestamp 1727493435
transform 1 0 6070 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1582_
timestamp 1727493435
transform 1 0 2950 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1583_
timestamp 1727493435
transform -1 0 2990 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1584_
timestamp 1727493435
transform 1 0 3210 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1585_
timestamp 1727493435
transform -1 0 3290 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1586_
timestamp 1727493435
transform 1 0 2870 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1587_
timestamp 1727493435
transform -1 0 510 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1588_
timestamp 1727493435
transform 1 0 990 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1589_
timestamp 1727493435
transform 1 0 850 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1590_
timestamp 1727493435
transform 1 0 670 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1591_
timestamp 1727493435
transform -1 0 530 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1592_
timestamp 1727493435
transform 1 0 30 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1593_
timestamp 1727493435
transform -1 0 50 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1594_
timestamp 1727493435
transform 1 0 190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1595_
timestamp 1727493435
transform -1 0 210 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1596_
timestamp 1727493435
transform 1 0 350 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1597_
timestamp 1727493435
transform 1 0 350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1598_
timestamp 1727493435
transform -1 0 390 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1599_
timestamp 1727493435
transform -1 0 230 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1600_
timestamp 1727493435
transform 1 0 490 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1601_
timestamp 1727493435
transform 1 0 1170 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1602_
timestamp 1727493435
transform -1 0 1630 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1603_
timestamp 1727493435
transform 1 0 1770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1604_
timestamp 1727493435
transform -1 0 1950 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1605_
timestamp 1727493435
transform 1 0 1570 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1606_
timestamp 1727493435
transform 1 0 2230 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1607_
timestamp 1727493435
transform 1 0 1410 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1608_
timestamp 1727493435
transform 1 0 1570 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1609_
timestamp 1727493435
transform 1 0 1730 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1610_
timestamp 1727493435
transform -1 0 5730 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1611_
timestamp 1727493435
transform -1 0 5570 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1__1612_
timestamp 1727493435
transform 1 0 770 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1613_
timestamp 1727493435
transform 1 0 2490 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1614_
timestamp 1727493435
transform -1 0 2550 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1615_
timestamp 1727493435
transform -1 0 2710 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1616_
timestamp 1727493435
transform -1 0 3010 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1617_
timestamp 1727493435
transform -1 0 1250 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1618_
timestamp 1727493435
transform -1 0 1750 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1619_
timestamp 1727493435
transform 1 0 330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1620_
timestamp 1727493435
transform 1 0 1450 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1__1621_
timestamp 1727493435
transform -1 0 1150 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1622_
timestamp 1727493435
transform 1 0 1610 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1623_
timestamp 1727493435
transform -1 0 1490 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1624_
timestamp 1727493435
transform 1 0 1770 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1625_
timestamp 1727493435
transform 1 0 2030 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1626_
timestamp 1727493435
transform 1 0 2030 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1627_
timestamp 1727493435
transform -1 0 2210 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1628_
timestamp 1727493435
transform 1 0 2090 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1629_
timestamp 1727493435
transform 1 0 2190 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1630_
timestamp 1727493435
transform 1 0 2350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1631_
timestamp 1727493435
transform -1 0 5790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_1__1632_
timestamp 1727493435
transform 1 0 6130 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1633_
timestamp 1727493435
transform 1 0 5990 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1634_
timestamp 1727493435
transform 1 0 2350 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1635_
timestamp 1727493435
transform -1 0 3570 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1636_
timestamp 1727493435
transform -1 0 3390 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1637_
timestamp 1727493435
transform -1 0 2870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1638_
timestamp 1727493435
transform 1 0 2850 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1639_
timestamp 1727493435
transform 1 0 1850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1640_
timestamp 1727493435
transform -1 0 1330 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1641_
timestamp 1727493435
transform 1 0 1930 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1642_
timestamp 1727493435
transform -1 0 5670 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1643_
timestamp 1727493435
transform -1 0 6030 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1644_
timestamp 1727493435
transform -1 0 5370 0 1 1830
box -6 -8 26 272
use FILL  FILL_1__1645_
timestamp 1727493435
transform 1 0 2370 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1646_
timestamp 1727493435
transform -1 0 2530 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1647_
timestamp 1727493435
transform 1 0 2670 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1__1648_
timestamp 1727493435
transform -1 0 2690 0 1 3390
box -6 -8 26 272
use FILL  FILL_1__1649_
timestamp 1727493435
transform -1 0 4630 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1650_
timestamp 1727493435
transform -1 0 4770 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1651_
timestamp 1727493435
transform 1 0 4590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1652_
timestamp 1727493435
transform -1 0 4470 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1653_
timestamp 1727493435
transform 1 0 4670 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1654_
timestamp 1727493435
transform 1 0 4490 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1655_
timestamp 1727493435
transform 1 0 4470 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1656_
timestamp 1727493435
transform 1 0 4310 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1657_
timestamp 1727493435
transform 1 0 3930 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1658_
timestamp 1727493435
transform -1 0 3630 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1659_
timestamp 1727493435
transform -1 0 3450 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1660_
timestamp 1727493435
transform 1 0 3270 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1661_
timestamp 1727493435
transform 1 0 3150 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1662_
timestamp 1727493435
transform 1 0 2970 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1663_
timestamp 1727493435
transform -1 0 3810 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1664_
timestamp 1727493435
transform 1 0 3690 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1692_
timestamp 1727493435
transform -1 0 3650 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1693_
timestamp 1727493435
transform -1 0 3910 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1694_
timestamp 1727493435
transform -1 0 3490 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1695_
timestamp 1727493435
transform 1 0 3290 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1696_
timestamp 1727493435
transform -1 0 2970 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1697_
timestamp 1727493435
transform -1 0 3770 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1698_
timestamp 1727493435
transform 1 0 4170 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1699_
timestamp 1727493435
transform 1 0 3490 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1700_
timestamp 1727493435
transform 1 0 3790 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1701_
timestamp 1727493435
transform 1 0 3610 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1702_
timestamp 1727493435
transform 1 0 3610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1703_
timestamp 1727493435
transform 1 0 3090 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1704_
timestamp 1727493435
transform 1 0 4450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1705_
timestamp 1727493435
transform -1 0 3510 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1706_
timestamp 1727493435
transform -1 0 3890 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1707_
timestamp 1727493435
transform 1 0 3710 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1708_
timestamp 1727493435
transform -1 0 3410 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1709_
timestamp 1727493435
transform -1 0 3570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1710_
timestamp 1727493435
transform -1 0 3950 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1711_
timestamp 1727493435
transform -1 0 3770 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1712_
timestamp 1727493435
transform 1 0 2010 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1713_
timestamp 1727493435
transform 1 0 2470 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1714_
timestamp 1727493435
transform -1 0 2730 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1715_
timestamp 1727493435
transform 1 0 2990 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1716_
timestamp 1727493435
transform -1 0 3330 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1717_
timestamp 1727493435
transform -1 0 3190 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1718_
timestamp 1727493435
transform -1 0 2890 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1719_
timestamp 1727493435
transform 1 0 2790 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1720_
timestamp 1727493435
transform -1 0 2650 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1721_
timestamp 1727493435
transform 1 0 2750 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1722_
timestamp 1727493435
transform -1 0 3350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1723_
timestamp 1727493435
transform 1 0 2990 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1724_
timestamp 1727493435
transform -1 0 3250 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1725_
timestamp 1727493435
transform -1 0 3370 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1726_
timestamp 1727493435
transform -1 0 3070 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1727_
timestamp 1727493435
transform -1 0 2910 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1728_
timestamp 1727493435
transform -1 0 2610 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1729_
timestamp 1727493435
transform -1 0 2450 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1730_
timestamp 1727493435
transform 1 0 2230 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1731_
timestamp 1727493435
transform -1 0 2570 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1732_
timestamp 1727493435
transform 1 0 2370 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1733_
timestamp 1727493435
transform -1 0 2350 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1734_
timestamp 1727493435
transform 1 0 3750 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1735_
timestamp 1727493435
transform -1 0 3610 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1736_
timestamp 1727493435
transform -1 0 4050 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1737_
timestamp 1727493435
transform 1 0 4150 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1738_
timestamp 1727493435
transform -1 0 4030 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1739_
timestamp 1727493435
transform 1 0 3850 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1740_
timestamp 1727493435
transform -1 0 3450 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1741_
timestamp 1727493435
transform 1 0 3090 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1742_
timestamp 1727493435
transform 1 0 2470 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1743_
timestamp 1727493435
transform -1 0 1950 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1744_
timestamp 1727493435
transform 1 0 1910 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1745_
timestamp 1727493435
transform -1 0 1770 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1746_
timestamp 1727493435
transform 1 0 3950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1747_
timestamp 1727493435
transform 1 0 2090 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1748_
timestamp 1727493435
transform -1 0 1790 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1749_
timestamp 1727493435
transform -1 0 3230 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1750_
timestamp 1727493435
transform -1 0 3970 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1751_
timestamp 1727493435
transform 1 0 4030 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1752_
timestamp 1727493435
transform 1 0 3870 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1753_
timestamp 1727493435
transform 1 0 3530 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1754_
timestamp 1727493435
transform -1 0 3730 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1755_
timestamp 1727493435
transform -1 0 3390 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1756_
timestamp 1727493435
transform -1 0 2930 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1757_
timestamp 1727493435
transform -1 0 2770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1758_
timestamp 1727493435
transform -1 0 2650 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1759_
timestamp 1727493435
transform 1 0 2310 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1760_
timestamp 1727493435
transform -1 0 2130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1761_
timestamp 1727493435
transform 1 0 1470 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1762_
timestamp 1727493435
transform -1 0 1270 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1763_
timestamp 1727493435
transform -1 0 1430 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1764_
timestamp 1727493435
transform -1 0 1590 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1765_
timestamp 1727493435
transform 1 0 1110 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1766_
timestamp 1727493435
transform 1 0 2050 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1767_
timestamp 1727493435
transform -1 0 50 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1768_
timestamp 1727493435
transform -1 0 1330 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1769_
timestamp 1727493435
transform -1 0 1790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1770_
timestamp 1727493435
transform -1 0 2630 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1771_
timestamp 1727493435
transform -1 0 2470 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1772_
timestamp 1727493435
transform 1 0 2070 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1773_
timestamp 1727493435
transform 1 0 2550 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1774_
timestamp 1727493435
transform -1 0 1930 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1775_
timestamp 1727493435
transform 1 0 1770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1776_
timestamp 1727493435
transform -1 0 1630 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1777_
timestamp 1727493435
transform -1 0 1470 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1778_
timestamp 1727493435
transform -1 0 1310 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1779_
timestamp 1727493435
transform -1 0 290 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1780_
timestamp 1727493435
transform 1 0 170 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1781_
timestamp 1727493435
transform 1 0 330 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1782_
timestamp 1727493435
transform -1 0 510 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1783_
timestamp 1727493435
transform 1 0 2710 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1784_
timestamp 1727493435
transform 1 0 990 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1785_
timestamp 1727493435
transform -1 0 850 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1786_
timestamp 1727493435
transform 1 0 650 0 -1 6510
box -6 -8 26 272
use FILL  FILL_1__1787_
timestamp 1727493435
transform -1 0 430 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1788_
timestamp 1727493435
transform -1 0 1190 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1789_
timestamp 1727493435
transform 1 0 550 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1790_
timestamp 1727493435
transform 1 0 1590 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1791_
timestamp 1727493435
transform -1 0 2070 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1792_
timestamp 1727493435
transform -1 0 1930 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1793_
timestamp 1727493435
transform 1 0 1870 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1794_
timestamp 1727493435
transform -1 0 1710 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1795_
timestamp 1727493435
transform -1 0 1550 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1796_
timestamp 1727493435
transform -1 0 1870 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1797_
timestamp 1727493435
transform -1 0 1690 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1798_
timestamp 1727493435
transform -1 0 1530 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1799_
timestamp 1727493435
transform -1 0 1370 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1800_
timestamp 1727493435
transform 1 0 870 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1801_
timestamp 1727493435
transform 1 0 1610 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1802_
timestamp 1727493435
transform -1 0 1170 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1803_
timestamp 1727493435
transform 1 0 1010 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1804_
timestamp 1727493435
transform -1 0 870 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1805_
timestamp 1727493435
transform -1 0 750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1806_
timestamp 1727493435
transform -1 0 730 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1807_
timestamp 1727493435
transform -1 0 1050 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1808_
timestamp 1727493435
transform -1 0 1250 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1809_
timestamp 1727493435
transform -1 0 1030 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1810_
timestamp 1727493435
transform -1 0 1770 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1811_
timestamp 1727493435
transform 1 0 1450 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1812_
timestamp 1727493435
transform 1 0 1330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1813_
timestamp 1727493435
transform -1 0 1310 0 1 3910
box -6 -8 26 272
use FILL  FILL_1__1814_
timestamp 1727493435
transform -1 0 1190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1815_
timestamp 1727493435
transform 1 0 1750 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1816_
timestamp 1727493435
transform -1 0 1590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1817_
timestamp 1727493435
transform -1 0 1430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1818_
timestamp 1727493435
transform -1 0 1270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1819_
timestamp 1727493435
transform 1 0 1070 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1820_
timestamp 1727493435
transform -1 0 570 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1821_
timestamp 1727493435
transform 1 0 790 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1822_
timestamp 1727493435
transform -1 0 670 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1823_
timestamp 1727493435
transform -1 0 790 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1824_
timestamp 1727493435
transform -1 0 510 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1825_
timestamp 1727493435
transform 1 0 890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1826_
timestamp 1727493435
transform -1 0 1670 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1827_
timestamp 1727493435
transform 1 0 1490 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1828_
timestamp 1727493435
transform 1 0 1310 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1829_
timestamp 1727493435
transform -1 0 1170 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1830_
timestamp 1727493435
transform -1 0 990 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1831_
timestamp 1727493435
transform 1 0 1950 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1832_
timestamp 1727493435
transform -1 0 1810 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1833_
timestamp 1727493435
transform -1 0 1310 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1834_
timestamp 1727493435
transform -1 0 1150 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1835_
timestamp 1727493435
transform -1 0 950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1836_
timestamp 1727493435
transform -1 0 930 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1837_
timestamp 1727493435
transform -1 0 330 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1838_
timestamp 1727493435
transform 1 0 590 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1839_
timestamp 1727493435
transform 1 0 990 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1840_
timestamp 1727493435
transform 1 0 490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1841_
timestamp 1727493435
transform 1 0 430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1842_
timestamp 1727493435
transform 1 0 2250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1843_
timestamp 1727493435
transform 1 0 1810 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1844_
timestamp 1727493435
transform -1 0 1990 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1845_
timestamp 1727493435
transform -1 0 2130 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1846_
timestamp 1727493435
transform 1 0 1910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1847_
timestamp 1727493435
transform 1 0 2090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1848_
timestamp 1727493435
transform 1 0 2290 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1849_
timestamp 1727493435
transform -1 0 2150 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1850_
timestamp 1727493435
transform -1 0 1630 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1851_
timestamp 1727493435
transform -1 0 1470 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1852_
timestamp 1727493435
transform 1 0 530 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1853_
timestamp 1727493435
transform -1 0 50 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1854_
timestamp 1727493435
transform -1 0 210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1855_
timestamp 1727493435
transform 1 0 190 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1856_
timestamp 1727493435
transform 1 0 610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1857_
timestamp 1727493435
transform -1 0 1970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1858_
timestamp 1727493435
transform -1 0 2170 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1859_
timestamp 1727493435
transform 1 0 2410 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1860_
timestamp 1727493435
transform 1 0 690 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1861_
timestamp 1727493435
transform -1 0 830 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1862_
timestamp 1727493435
transform 1 0 1630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1863_
timestamp 1727493435
transform 1 0 2410 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1864_
timestamp 1727493435
transform -1 0 50 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1865_
timestamp 1727493435
transform -1 0 370 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1866_
timestamp 1727493435
transform 1 0 30 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1867_
timestamp 1727493435
transform -1 0 630 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1868_
timestamp 1727493435
transform -1 0 3250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1869_
timestamp 1727493435
transform 1 0 1090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1__1870_
timestamp 1727493435
transform -1 0 50 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1871_
timestamp 1727493435
transform -1 0 50 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1872_
timestamp 1727493435
transform -1 0 50 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1873_
timestamp 1727493435
transform -1 0 170 0 1 5990
box -6 -8 26 272
use FILL  FILL_1__1874_
timestamp 1727493435
transform -1 0 210 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1875_
timestamp 1727493435
transform -1 0 350 0 1 5470
box -6 -8 26 272
use FILL  FILL_1__1876_
timestamp 1727493435
transform -1 0 230 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1877_
timestamp 1727493435
transform 1 0 390 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1__1878_
timestamp 1727493435
transform 1 0 310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1879_
timestamp 1727493435
transform -1 0 670 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1880_
timestamp 1727493435
transform -1 0 1370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1881_
timestamp 1727493435
transform 1 0 1490 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1882_
timestamp 1727493435
transform -1 0 1050 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1883_
timestamp 1727493435
transform 1 0 1190 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1884_
timestamp 1727493435
transform 1 0 890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1885_
timestamp 1727493435
transform -1 0 770 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1886_
timestamp 1727493435
transform -1 0 350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1887_
timestamp 1727493435
transform -1 0 210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1888_
timestamp 1727493435
transform 1 0 30 0 -1 4950
box -6 -8 26 272
use FILL  FILL_1__1889_
timestamp 1727493435
transform 1 0 350 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1890_
timestamp 1727493435
transform 1 0 490 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1891_
timestamp 1727493435
transform -1 0 190 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1892_
timestamp 1727493435
transform -1 0 190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1893_
timestamp 1727493435
transform 1 0 470 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1894_
timestamp 1727493435
transform -1 0 830 0 1 4430
box -6 -8 26 272
use FILL  FILL_1__1895_
timestamp 1727493435
transform -1 0 50 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1__1896_
timestamp 1727493435
transform -1 0 4470 0 1 4950
box -6 -8 26 272
use FILL  FILL_1__1897_
timestamp 1727493435
transform 1 0 3890 0 1 790
box -6 -8 26 272
use FILL  FILL_1__1898_
timestamp 1727493435
transform 1 0 3590 0 1 2870
box -6 -8 26 272
use FILL  FILL_1__1899_
timestamp 1727493435
transform 1 0 3230 0 -1 270
box -6 -8 26 272
use FILL  FILL_1__1900_
timestamp 1727493435
transform 1 0 3130 0 -1 1830
box -6 -8 26 272
use FILL  FILL_1__1901_
timestamp 1727493435
transform -1 0 2730 0 1 2350
box -6 -8 26 272
use FILL  FILL_1__1902_
timestamp 1727493435
transform -1 0 5110 0 1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1727493435
transform -1 0 2290 0 1 2350
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1727493435
transform -1 0 2230 0 1 3910
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1727493435
transform 1 0 3890 0 1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1727493435
transform 1 0 3570 0 1 2350
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1727493435
transform -1 0 4770 0 1 4950
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1727493435
transform -1 0 4050 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1727493435
transform 1 0 4350 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1727493435
transform -1 0 4090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert8
timestamp 1727493435
transform -1 0 4150 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert9
timestamp 1727493435
transform -1 0 4630 0 1 4430
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert10
timestamp 1727493435
transform 1 0 5030 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert11
timestamp 1727493435
transform 1 0 4750 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1727493435
transform -1 0 3590 0 1 3910
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1727493435
transform 1 0 4210 0 1 3910
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1727493435
transform -1 0 5190 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1727493435
transform -1 0 4910 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1727493435
transform 1 0 3790 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1727493435
transform -1 0 3670 0 -1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1727493435
transform -1 0 1910 0 1 2870
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1727493435
transform -1 0 1910 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1727493435
transform -1 0 4610 0 1 4950
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1727493435
transform 1 0 3890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1727493435
transform 1 0 4370 0 1 3910
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1727493435
transform -1 0 3770 0 -1 3390
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1727493435
transform -1 0 2270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1727493435
transform 1 0 2290 0 1 5470
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1727493435
transform 1 0 3090 0 -1 5990
box -6 -8 26 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1727493435
transform -1 0 4110 0 1 5990
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1727493435
transform 1 0 4210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert13
timestamp 1727493435
transform -1 0 4110 0 1 3390
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 3870 0 -1 4430
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 4170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_1_CLKBUF1_insert16
timestamp 1727493435
transform 1 0 4170 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__927_
timestamp 1727493435
transform 1 0 5610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__928_
timestamp 1727493435
transform -1 0 5610 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__929_
timestamp 1727493435
transform -1 0 5890 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__930_
timestamp 1727493435
transform 1 0 6010 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__931_
timestamp 1727493435
transform -1 0 5330 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__932_
timestamp 1727493435
transform -1 0 3430 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__933_
timestamp 1727493435
transform 1 0 5450 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__934_
timestamp 1727493435
transform 1 0 5430 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__935_
timestamp 1727493435
transform 1 0 5990 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__936_
timestamp 1727493435
transform -1 0 5370 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__937_
timestamp 1727493435
transform 1 0 5570 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__938_
timestamp 1727493435
transform -1 0 5910 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__939_
timestamp 1727493435
transform 1 0 6030 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__940_
timestamp 1727493435
transform 1 0 6250 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__941_
timestamp 1727493435
transform 1 0 3810 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__942_
timestamp 1727493435
transform 1 0 5730 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__943_
timestamp 1727493435
transform 1 0 5990 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__944_
timestamp 1727493435
transform 1 0 5730 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__945_
timestamp 1727493435
transform 1 0 6250 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__946_
timestamp 1727493435
transform -1 0 5790 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__947_
timestamp 1727493435
transform 1 0 5750 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__948_
timestamp 1727493435
transform -1 0 5930 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__949_
timestamp 1727493435
transform 1 0 5890 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__950_
timestamp 1727493435
transform -1 0 5650 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__951_
timestamp 1727493435
transform -1 0 6130 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__952_
timestamp 1727493435
transform -1 0 5670 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__953_
timestamp 1727493435
transform 1 0 5210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__954_
timestamp 1727493435
transform 1 0 6270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__955_
timestamp 1727493435
transform 1 0 6190 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__956_
timestamp 1727493435
transform -1 0 5810 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__957_
timestamp 1727493435
transform -1 0 5510 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__958_
timestamp 1727493435
transform 1 0 6290 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__959_
timestamp 1727493435
transform -1 0 6130 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__960_
timestamp 1727493435
transform 1 0 6070 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__961_
timestamp 1727493435
transform -1 0 6110 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__962_
timestamp 1727493435
transform 1 0 5830 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__963_
timestamp 1727493435
transform -1 0 5510 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__964_
timestamp 1727493435
transform -1 0 5350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__965_
timestamp 1727493435
transform 1 0 4490 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__966_
timestamp 1727493435
transform -1 0 4650 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__967_
timestamp 1727493435
transform 1 0 4930 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__968_
timestamp 1727493435
transform 1 0 5150 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__969_
timestamp 1727493435
transform 1 0 5030 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__970_
timestamp 1727493435
transform 1 0 4070 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__971_
timestamp 1727493435
transform 1 0 4850 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__972_
timestamp 1727493435
transform 1 0 4690 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__973_
timestamp 1727493435
transform 1 0 4350 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__974_
timestamp 1727493435
transform 1 0 4370 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__975_
timestamp 1727493435
transform 1 0 4430 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__976_
timestamp 1727493435
transform 1 0 3690 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__977_
timestamp 1727493435
transform 1 0 3970 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__978_
timestamp 1727493435
transform 1 0 3730 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__979_
timestamp 1727493435
transform 1 0 3170 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__980_
timestamp 1727493435
transform 1 0 3310 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__981_
timestamp 1727493435
transform -1 0 3170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__982_
timestamp 1727493435
transform 1 0 2070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__983_
timestamp 1727493435
transform 1 0 2690 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__984_
timestamp 1727493435
transform -1 0 2850 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__985_
timestamp 1727493435
transform 1 0 3630 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__986_
timestamp 1727493435
transform 1 0 3910 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__987_
timestamp 1727493435
transform -1 0 4090 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__988_
timestamp 1727493435
transform -1 0 2330 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__989_
timestamp 1727493435
transform 1 0 5250 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__990_
timestamp 1727493435
transform -1 0 1770 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__991_
timestamp 1727493435
transform 1 0 5590 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__992_
timestamp 1727493435
transform 1 0 5430 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__993_
timestamp 1727493435
transform 1 0 5730 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__994_
timestamp 1727493435
transform -1 0 4310 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__995_
timestamp 1727493435
transform -1 0 4630 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__996_
timestamp 1727493435
transform 1 0 6270 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__997_
timestamp 1727493435
transform 1 0 5470 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__998_
timestamp 1727493435
transform -1 0 6270 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__999_
timestamp 1727493435
transform 1 0 6090 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1000_
timestamp 1727493435
transform -1 0 4890 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1001_
timestamp 1727493435
transform 1 0 5330 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1002_
timestamp 1727493435
transform 1 0 4670 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1003_
timestamp 1727493435
transform 1 0 4750 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1004_
timestamp 1727493435
transform 1 0 4670 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1005_
timestamp 1727493435
transform -1 0 5230 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1006_
timestamp 1727493435
transform 1 0 5610 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1007_
timestamp 1727493435
transform -1 0 4930 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1008_
timestamp 1727493435
transform -1 0 5050 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1009_
timestamp 1727493435
transform 1 0 5930 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1010_
timestamp 1727493435
transform -1 0 5370 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1011_
timestamp 1727493435
transform 1 0 4950 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1012_
timestamp 1727493435
transform -1 0 3490 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1013_
timestamp 1727493435
transform -1 0 4350 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1014_
timestamp 1727493435
transform 1 0 5270 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1015_
timestamp 1727493435
transform 1 0 5270 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1016_
timestamp 1727493435
transform -1 0 5790 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1017_
timestamp 1727493435
transform 1 0 5610 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1018_
timestamp 1727493435
transform 1 0 5050 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1019_
timestamp 1727493435
transform 1 0 3970 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1020_
timestamp 1727493435
transform 1 0 4150 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1021_
timestamp 1727493435
transform -1 0 4210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1022_
timestamp 1727493435
transform 1 0 4530 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1023_
timestamp 1727493435
transform -1 0 4070 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1024_
timestamp 1727493435
transform -1 0 4830 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1025_
timestamp 1727493435
transform 1 0 4650 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1026_
timestamp 1727493435
transform -1 0 4530 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1027_
timestamp 1727493435
transform 1 0 4810 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1028_
timestamp 1727493435
transform 1 0 4930 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1029_
timestamp 1727493435
transform 1 0 5250 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1030_
timestamp 1727493435
transform -1 0 5230 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1031_
timestamp 1727493435
transform -1 0 4710 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1032_
timestamp 1727493435
transform -1 0 4390 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1033_
timestamp 1727493435
transform 1 0 4850 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1034_
timestamp 1727493435
transform -1 0 4330 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1035_
timestamp 1727493435
transform 1 0 4630 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1036_
timestamp 1727493435
transform 1 0 4470 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1037_
timestamp 1727493435
transform -1 0 5150 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1038_
timestamp 1727493435
transform 1 0 4550 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1039_
timestamp 1727493435
transform 1 0 4790 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1040_
timestamp 1727493435
transform 1 0 4750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1041_
timestamp 1727493435
transform 1 0 4950 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1042_
timestamp 1727493435
transform 1 0 5510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1043_
timestamp 1727493435
transform -1 0 5070 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1044_
timestamp 1727493435
transform 1 0 4910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1045_
timestamp 1727493435
transform 1 0 5230 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1046_
timestamp 1727493435
transform 1 0 5650 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1047_
timestamp 1727493435
transform 1 0 5010 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1048_
timestamp 1727493435
transform 1 0 5090 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1049_
timestamp 1727493435
transform 1 0 5070 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1050_
timestamp 1727493435
transform 1 0 5330 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1051_
timestamp 1727493435
transform 1 0 5810 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1052_
timestamp 1727493435
transform 1 0 5970 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1053_
timestamp 1727493435
transform 1 0 6370 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1054_
timestamp 1727493435
transform 1 0 5410 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1055_
timestamp 1727493435
transform -1 0 4230 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1056_
timestamp 1727493435
transform -1 0 2910 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1057_
timestamp 1727493435
transform -1 0 4050 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1058_
timestamp 1727493435
transform -1 0 4230 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1059_
timestamp 1727493435
transform 1 0 3130 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1060_
timestamp 1727493435
transform 1 0 3890 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1061_
timestamp 1727493435
transform 1 0 4050 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1062_
timestamp 1727493435
transform 1 0 4310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1063_
timestamp 1727493435
transform -1 0 4330 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1064_
timestamp 1727493435
transform -1 0 4010 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1065_
timestamp 1727493435
transform -1 0 3930 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1066_
timestamp 1727493435
transform -1 0 4190 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1067_
timestamp 1727493435
transform 1 0 4050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1068_
timestamp 1727493435
transform -1 0 4610 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1069_
timestamp 1727493435
transform -1 0 4350 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1070_
timestamp 1727493435
transform 1 0 4530 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1071_
timestamp 1727493435
transform 1 0 4750 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1072_
timestamp 1727493435
transform 1 0 4430 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1073_
timestamp 1727493435
transform 1 0 5090 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1074_
timestamp 1727493435
transform 1 0 4450 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1075_
timestamp 1727493435
transform -1 0 4770 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1076_
timestamp 1727493435
transform -1 0 4610 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1077_
timestamp 1727493435
transform 1 0 4470 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1078_
timestamp 1727493435
transform -1 0 4770 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1079_
timestamp 1727493435
transform 1 0 3770 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1080_
timestamp 1727493435
transform -1 0 5230 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1081_
timestamp 1727493435
transform -1 0 4910 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1082_
timestamp 1727493435
transform 1 0 5070 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1083_
timestamp 1727493435
transform 1 0 4430 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1084_
timestamp 1727493435
transform 1 0 4630 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1085_
timestamp 1727493435
transform 1 0 4590 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1086_
timestamp 1727493435
transform 1 0 5410 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1087_
timestamp 1727493435
transform 1 0 5150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1088_
timestamp 1727493435
transform 1 0 4930 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1089_
timestamp 1727493435
transform 1 0 4490 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1090_
timestamp 1727493435
transform -1 0 5270 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1091_
timestamp 1727493435
transform 1 0 4830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1092_
timestamp 1727493435
transform 1 0 5490 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1093_
timestamp 1727493435
transform 1 0 5170 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1094_
timestamp 1727493435
transform 1 0 4830 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1095_
timestamp 1727493435
transform 1 0 5010 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1096_
timestamp 1727493435
transform 1 0 5330 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1097_
timestamp 1727493435
transform -1 0 1610 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1098_
timestamp 1727493435
transform 1 0 5590 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1099_
timestamp 1727493435
transform 1 0 5350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1100_
timestamp 1727493435
transform -1 0 5510 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1101_
timestamp 1727493435
transform 1 0 5630 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1102_
timestamp 1727493435
transform 1 0 5810 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1103_
timestamp 1727493435
transform 1 0 6110 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1104_
timestamp 1727493435
transform 1 0 5170 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1105_
timestamp 1727493435
transform 1 0 5310 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1106_
timestamp 1727493435
transform -1 0 5990 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1107_
timestamp 1727493435
transform -1 0 6150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1108_
timestamp 1727493435
transform 1 0 6390 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1109_
timestamp 1727493435
transform 1 0 6270 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1110_
timestamp 1727493435
transform -1 0 5830 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1111_
timestamp 1727493435
transform 1 0 4990 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1112_
timestamp 1727493435
transform -1 0 4270 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1113_
timestamp 1727493435
transform -1 0 3770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1114_
timestamp 1727493435
transform -1 0 3590 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1115_
timestamp 1727493435
transform -1 0 3170 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1116_
timestamp 1727493435
transform -1 0 3270 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1117_
timestamp 1727493435
transform -1 0 3470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1118_
timestamp 1727493435
transform 1 0 3750 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1119_
timestamp 1727493435
transform -1 0 3770 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1120_
timestamp 1727493435
transform -1 0 3850 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1121_
timestamp 1727493435
transform -1 0 3590 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1122_
timestamp 1727493435
transform 1 0 4230 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1123_
timestamp 1727493435
transform 1 0 3730 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1124_
timestamp 1727493435
transform -1 0 3290 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1125_
timestamp 1727493435
transform -1 0 4390 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1126_
timestamp 1727493435
transform -1 0 3430 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1127_
timestamp 1727493435
transform -1 0 3430 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1128_
timestamp 1727493435
transform 1 0 3670 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1129_
timestamp 1727493435
transform 1 0 3990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1130_
timestamp 1727493435
transform 1 0 3890 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1131_
timestamp 1727493435
transform -1 0 3490 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1132_
timestamp 1727493435
transform 1 0 3550 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1133_
timestamp 1727493435
transform 1 0 3670 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1134_
timestamp 1727493435
transform -1 0 3370 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1135_
timestamp 1727493435
transform 1 0 3550 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1136_
timestamp 1727493435
transform -1 0 4170 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1137_
timestamp 1727493435
transform 1 0 3730 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1138_
timestamp 1727493435
transform 1 0 4030 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1139_
timestamp 1727493435
transform 1 0 4590 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1140_
timestamp 1727493435
transform 1 0 4170 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1141_
timestamp 1727493435
transform 1 0 4210 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1142_
timestamp 1727493435
transform -1 0 4070 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1143_
timestamp 1727493435
transform -1 0 3910 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1144_
timestamp 1727493435
transform 1 0 4750 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1145_
timestamp 1727493435
transform 1 0 5070 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1146_
timestamp 1727493435
transform -1 0 4670 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1147_
timestamp 1727493435
transform 1 0 4710 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1148_
timestamp 1727493435
transform 1 0 4550 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1149_
timestamp 1727493435
transform 1 0 5030 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1150_
timestamp 1727493435
transform -1 0 5210 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1151_
timestamp 1727493435
transform -1 0 5790 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1152_
timestamp 1727493435
transform 1 0 4890 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1153_
timestamp 1727493435
transform 1 0 6370 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1154_
timestamp 1727493435
transform 1 0 6070 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1155_
timestamp 1727493435
transform -1 0 6010 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1156_
timestamp 1727493435
transform 1 0 6130 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1157_
timestamp 1727493435
transform 1 0 5890 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1158_
timestamp 1727493435
transform 1 0 6230 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1159_
timestamp 1727493435
transform 1 0 5430 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1160_
timestamp 1727493435
transform -1 0 5290 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1161_
timestamp 1727493435
transform -1 0 5130 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1162_
timestamp 1727493435
transform 1 0 5230 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1163_
timestamp 1727493435
transform 1 0 4870 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1164_
timestamp 1727493435
transform 1 0 4910 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1165_
timestamp 1727493435
transform -1 0 5610 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1166_
timestamp 1727493435
transform -1 0 5670 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1167_
timestamp 1727493435
transform 1 0 5510 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1168_
timestamp 1727493435
transform 1 0 5570 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1169_
timestamp 1727493435
transform 1 0 5830 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1170_
timestamp 1727493435
transform -1 0 5670 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1171_
timestamp 1727493435
transform -1 0 5370 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1172_
timestamp 1727493435
transform 1 0 5390 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1173_
timestamp 1727493435
transform 1 0 5670 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1174_
timestamp 1727493435
transform 1 0 6090 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1175_
timestamp 1727493435
transform 1 0 5510 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1176_
timestamp 1727493435
transform 1 0 5750 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1177_
timestamp 1727493435
transform 1 0 6310 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1178_
timestamp 1727493435
transform 1 0 6370 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1179_
timestamp 1727493435
transform 1 0 5730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1180_
timestamp 1727493435
transform 1 0 6410 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1181_
timestamp 1727493435
transform 1 0 6130 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1182_
timestamp 1727493435
transform -1 0 5830 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1183_
timestamp 1727493435
transform -1 0 4550 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1184_
timestamp 1727493435
transform 1 0 4430 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1185_
timestamp 1727493435
transform 1 0 5970 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1186_
timestamp 1727493435
transform 1 0 5390 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1187_
timestamp 1727493435
transform 1 0 5550 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1188_
timestamp 1727493435
transform 1 0 5730 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1189_
timestamp 1727493435
transform -1 0 5590 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1190_
timestamp 1727493435
transform 1 0 5890 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1191_
timestamp 1727493435
transform -1 0 5790 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1192_
timestamp 1727493435
transform 1 0 5490 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1193_
timestamp 1727493435
transform 1 0 5410 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1194_
timestamp 1727493435
transform 1 0 5730 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1195_
timestamp 1727493435
transform 1 0 6270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1196_
timestamp 1727493435
transform 1 0 6290 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1197_
timestamp 1727493435
transform 1 0 5970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1198_
timestamp 1727493435
transform 1 0 6270 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1199_
timestamp 1727493435
transform -1 0 6270 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1200_
timestamp 1727493435
transform 1 0 5990 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1201_
timestamp 1727493435
transform 1 0 6150 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1202_
timestamp 1727493435
transform 1 0 5950 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1203_
timestamp 1727493435
transform -1 0 5830 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1204_
timestamp 1727493435
transform 1 0 5030 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1205_
timestamp 1727493435
transform 1 0 5450 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1206_
timestamp 1727493435
transform -1 0 5190 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1207_
timestamp 1727493435
transform 1 0 5630 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1208_
timestamp 1727493435
transform -1 0 5950 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1209_
timestamp 1727493435
transform -1 0 5490 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1210_
timestamp 1727493435
transform -1 0 5650 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1211_
timestamp 1727493435
transform 1 0 5450 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1212_
timestamp 1727493435
transform -1 0 5470 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1213_
timestamp 1727493435
transform 1 0 6130 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1214_
timestamp 1727493435
transform 1 0 6310 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1215_
timestamp 1727493435
transform -1 0 5910 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1216_
timestamp 1727493435
transform 1 0 6070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1217_
timestamp 1727493435
transform -1 0 6250 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1218_
timestamp 1727493435
transform 1 0 6330 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1219_
timestamp 1727493435
transform -1 0 6170 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1220_
timestamp 1727493435
transform -1 0 4770 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1221_
timestamp 1727493435
transform -1 0 4890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1222_
timestamp 1727493435
transform 1 0 6290 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1223_
timestamp 1727493435
transform -1 0 6350 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1224_
timestamp 1727493435
transform 1 0 6170 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1225_
timestamp 1727493435
transform -1 0 6170 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1226_
timestamp 1727493435
transform 1 0 4770 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1227_
timestamp 1727493435
transform -1 0 5550 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1228_
timestamp 1727493435
transform -1 0 6010 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1229_
timestamp 1727493435
transform 1 0 5830 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1230_
timestamp 1727493435
transform 1 0 5350 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1231_
timestamp 1727493435
transform -1 0 5070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1232_
timestamp 1727493435
transform 1 0 5170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1233_
timestamp 1727493435
transform -1 0 5210 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1234_
timestamp 1727493435
transform 1 0 6050 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1235_
timestamp 1727493435
transform 1 0 6210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1236_
timestamp 1727493435
transform 1 0 6090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1237_
timestamp 1727493435
transform -1 0 6330 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1238_
timestamp 1727493435
transform -1 0 6170 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1239_
timestamp 1727493435
transform 1 0 5910 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1240_
timestamp 1727493435
transform 1 0 5890 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1241_
timestamp 1727493435
transform -1 0 6010 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1242_
timestamp 1727493435
transform 1 0 5830 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1243_
timestamp 1727493435
transform -1 0 5870 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1244_
timestamp 1727493435
transform -1 0 5950 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1245_
timestamp 1727493435
transform -1 0 4990 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1246_
timestamp 1727493435
transform -1 0 5370 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1247_
timestamp 1727493435
transform 1 0 4390 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1248_
timestamp 1727493435
transform -1 0 4230 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1249_
timestamp 1727493435
transform 1 0 4690 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1250_
timestamp 1727493435
transform 1 0 3830 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1251_
timestamp 1727493435
transform 1 0 4810 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1252_
timestamp 1727493435
transform -1 0 4510 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1253_
timestamp 1727493435
transform 1 0 4330 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1254_
timestamp 1727493435
transform 1 0 5010 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1255_
timestamp 1727493435
transform 1 0 4870 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1256_
timestamp 1727493435
transform -1 0 4730 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1257_
timestamp 1727493435
transform 1 0 4390 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1258_
timestamp 1727493435
transform -1 0 4430 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1259_
timestamp 1727493435
transform 1 0 2590 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1260_
timestamp 1727493435
transform -1 0 3210 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1261_
timestamp 1727493435
transform 1 0 3030 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1262_
timestamp 1727493435
transform -1 0 3130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1263_
timestamp 1727493435
transform 1 0 2790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1264_
timestamp 1727493435
transform 1 0 2870 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1265_
timestamp 1727493435
transform -1 0 2210 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1266_
timestamp 1727493435
transform -1 0 2970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1267_
timestamp 1727493435
transform 1 0 3290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1268_
timestamp 1727493435
transform -1 0 2510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1269_
timestamp 1727493435
transform -1 0 2630 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1270_
timestamp 1727493435
transform 1 0 2730 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1271_
timestamp 1727493435
transform -1 0 3610 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1272_
timestamp 1727493435
transform 1 0 2750 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1273_
timestamp 1727493435
transform -1 0 2810 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1274_
timestamp 1727493435
transform -1 0 3090 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1275_
timestamp 1727493435
transform 1 0 3070 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1276_
timestamp 1727493435
transform 1 0 3290 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1277_
timestamp 1727493435
transform 1 0 3230 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1278_
timestamp 1727493435
transform 1 0 3290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1279_
timestamp 1727493435
transform -1 0 3430 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1280_
timestamp 1727493435
transform -1 0 3030 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1281_
timestamp 1727493435
transform 1 0 3110 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1282_
timestamp 1727493435
transform -1 0 2950 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1283_
timestamp 1727493435
transform 1 0 2870 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1284_
timestamp 1727493435
transform 1 0 3430 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1285_
timestamp 1727493435
transform 1 0 3450 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1286_
timestamp 1727493435
transform 1 0 3930 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1287_
timestamp 1727493435
transform -1 0 4270 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1288_
timestamp 1727493435
transform 1 0 3090 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1289_
timestamp 1727493435
transform -1 0 2970 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1290_
timestamp 1727493435
transform 1 0 4090 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1291_
timestamp 1727493435
transform -1 0 3890 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1292_
timestamp 1727493435
transform 1 0 4530 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1293_
timestamp 1727493435
transform 1 0 3770 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1294_
timestamp 1727493435
transform 1 0 3710 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1295_
timestamp 1727493435
transform -1 0 3370 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1296_
timestamp 1727493435
transform -1 0 3410 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1297_
timestamp 1727493435
transform -1 0 5210 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1298_
timestamp 1727493435
transform -1 0 4230 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1299_
timestamp 1727493435
transform 1 0 4030 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1300_
timestamp 1727493435
transform -1 0 3910 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1301_
timestamp 1727493435
transform 1 0 2470 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1302_
timestamp 1727493435
transform -1 0 2650 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1303_
timestamp 1727493435
transform -1 0 3730 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1304_
timestamp 1727493435
transform 1 0 4050 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1305_
timestamp 1727493435
transform -1 0 2770 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1306_
timestamp 1727493435
transform 1 0 2610 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1307_
timestamp 1727493435
transform -1 0 5830 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1308_
timestamp 1727493435
transform 1 0 2910 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1309_
timestamp 1727493435
transform 1 0 2310 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1310_
timestamp 1727493435
transform -1 0 2790 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1311_
timestamp 1727493435
transform -1 0 2510 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1312_
timestamp 1727493435
transform -1 0 2390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1313_
timestamp 1727493435
transform -1 0 6230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1314_
timestamp 1727493435
transform -1 0 6350 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1315_
timestamp 1727493435
transform 1 0 6390 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1316_
timestamp 1727493435
transform -1 0 6310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1317_
timestamp 1727493435
transform -1 0 5970 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1318_
timestamp 1727493435
transform 1 0 6110 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1319_
timestamp 1727493435
transform -1 0 5650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1320_
timestamp 1727493435
transform -1 0 5530 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1321_
timestamp 1727493435
transform 1 0 2590 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1322_
timestamp 1727493435
transform 1 0 2850 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1323_
timestamp 1727493435
transform -1 0 2450 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1324_
timestamp 1727493435
transform -1 0 2810 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1325_
timestamp 1727493435
transform -1 0 2950 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1326_
timestamp 1727493435
transform 1 0 2750 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1327_
timestamp 1727493435
transform -1 0 3550 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1328_
timestamp 1727493435
transform 1 0 2850 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1329_
timestamp 1727493435
transform -1 0 2930 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1330_
timestamp 1727493435
transform 1 0 2830 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1331_
timestamp 1727493435
transform 1 0 2670 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1332_
timestamp 1727493435
transform 1 0 2210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1333_
timestamp 1727493435
transform 1 0 2050 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1334_
timestamp 1727493435
transform -1 0 2530 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1335_
timestamp 1727493435
transform 1 0 2190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1336_
timestamp 1727493435
transform -1 0 3570 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1337_
timestamp 1727493435
transform 1 0 3070 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1338_
timestamp 1727493435
transform -1 0 4670 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1339_
timestamp 1727493435
transform -1 0 3630 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1340_
timestamp 1727493435
transform -1 0 3550 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1341_
timestamp 1727493435
transform -1 0 2830 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1342_
timestamp 1727493435
transform -1 0 2710 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1343_
timestamp 1727493435
transform -1 0 3030 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1344_
timestamp 1727493435
transform -1 0 2330 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1345_
timestamp 1727493435
transform -1 0 2370 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1346_
timestamp 1727493435
transform 1 0 2250 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1347_
timestamp 1727493435
transform -1 0 2550 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1348_
timestamp 1727493435
transform -1 0 1950 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1349_
timestamp 1727493435
transform -1 0 2130 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1350_
timestamp 1727493435
transform 1 0 2210 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1351_
timestamp 1727493435
transform 1 0 2070 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1352_
timestamp 1727493435
transform 1 0 3290 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1353_
timestamp 1727493435
transform -1 0 2790 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1354_
timestamp 1727493435
transform -1 0 1530 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1355_
timestamp 1727493435
transform -1 0 1290 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1356_
timestamp 1727493435
transform 1 0 1830 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1357_
timestamp 1727493435
transform -1 0 2150 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1358_
timestamp 1727493435
transform 1 0 1990 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1359_
timestamp 1727493435
transform 1 0 1310 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1360_
timestamp 1727493435
transform -1 0 970 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1361_
timestamp 1727493435
transform 1 0 1230 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1362_
timestamp 1727493435
transform 1 0 1330 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1363_
timestamp 1727493435
transform 1 0 1650 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1364_
timestamp 1727493435
transform -1 0 2450 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1365_
timestamp 1727493435
transform -1 0 1430 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1366_
timestamp 1727493435
transform -1 0 1390 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1367_
timestamp 1727493435
transform 1 0 1570 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1368_
timestamp 1727493435
transform -1 0 1090 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1369_
timestamp 1727493435
transform 1 0 1570 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1370_
timestamp 1727493435
transform -1 0 1410 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1371_
timestamp 1727493435
transform -1 0 1470 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1372_
timestamp 1727493435
transform 1 0 2170 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1373_
timestamp 1727493435
transform 1 0 2930 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1374_
timestamp 1727493435
transform 1 0 2410 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1375_
timestamp 1727493435
transform 1 0 1770 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1376_
timestamp 1727493435
transform 1 0 1850 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1377_
timestamp 1727493435
transform -1 0 1930 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1378_
timestamp 1727493435
transform 1 0 1590 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1379_
timestamp 1727493435
transform 1 0 1590 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1380_
timestamp 1727493435
transform -1 0 1490 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1381_
timestamp 1727493435
transform -1 0 890 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1382_
timestamp 1727493435
transform -1 0 3130 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1383_
timestamp 1727493435
transform -1 0 2970 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1384_
timestamp 1727493435
transform 1 0 1630 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1385_
timestamp 1727493435
transform 1 0 1730 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1386_
timestamp 1727493435
transform -1 0 2630 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1387_
timestamp 1727493435
transform 1 0 2010 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1388_
timestamp 1727493435
transform -1 0 1330 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1389_
timestamp 1727493435
transform -1 0 1190 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1390_
timestamp 1727493435
transform -1 0 1070 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1391_
timestamp 1727493435
transform 1 0 1150 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1392_
timestamp 1727493435
transform 1 0 1790 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1393_
timestamp 1727493435
transform 1 0 1510 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1394_
timestamp 1727493435
transform 1 0 1870 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1395_
timestamp 1727493435
transform 1 0 1350 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1396_
timestamp 1727493435
transform 1 0 1950 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1397_
timestamp 1727493435
transform -1 0 2310 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1398_
timestamp 1727493435
transform 1 0 2470 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1399_
timestamp 1727493435
transform 1 0 2510 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1400_
timestamp 1727493435
transform -1 0 2690 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1401_
timestamp 1727493435
transform -1 0 2050 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1402_
timestamp 1727493435
transform -1 0 2170 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1403_
timestamp 1727493435
transform 1 0 2130 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1404_
timestamp 1727493435
transform 1 0 1690 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1405_
timestamp 1727493435
transform 1 0 2470 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1406_
timestamp 1727493435
transform -1 0 2610 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1407_
timestamp 1727493435
transform -1 0 2570 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1408_
timestamp 1727493435
transform -1 0 4870 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1409_
timestamp 1727493435
transform 1 0 4330 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1410_
timestamp 1727493435
transform -1 0 4710 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1411_
timestamp 1727493435
transform -1 0 4530 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1412_
timestamp 1727493435
transform -1 0 3250 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1413_
timestamp 1727493435
transform 1 0 2570 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1414_
timestamp 1727493435
transform -1 0 5310 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1415_
timestamp 1727493435
transform -1 0 2210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1416_
timestamp 1727493435
transform -1 0 2330 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1417_
timestamp 1727493435
transform 1 0 1870 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1418_
timestamp 1727493435
transform 1 0 2370 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1419_
timestamp 1727493435
transform -1 0 1330 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1420_
timestamp 1727493435
transform -1 0 1530 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1421_
timestamp 1727493435
transform -1 0 950 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1422_
timestamp 1727493435
transform 1 0 1030 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1423_
timestamp 1727493435
transform -1 0 670 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1424_
timestamp 1727493435
transform -1 0 1130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1425_
timestamp 1727493435
transform -1 0 470 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1426_
timestamp 1727493435
transform 1 0 750 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1427_
timestamp 1727493435
transform -1 0 890 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1428_
timestamp 1727493435
transform 1 0 590 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1429_
timestamp 1727493435
transform -1 0 330 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1430_
timestamp 1727493435
transform 1 0 690 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1431_
timestamp 1727493435
transform 1 0 850 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1432_
timestamp 1727493435
transform 1 0 1570 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1433_
timestamp 1727493435
transform -1 0 830 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1434_
timestamp 1727493435
transform -1 0 370 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1435_
timestamp 1727493435
transform -1 0 990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1436_
timestamp 1727493435
transform 1 0 990 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1437_
timestamp 1727493435
transform 1 0 830 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1438_
timestamp 1727493435
transform -1 0 210 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1439_
timestamp 1727493435
transform 1 0 1130 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1440_
timestamp 1727493435
transform -1 0 70 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1441_
timestamp 1727493435
transform -1 0 190 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1442_
timestamp 1727493435
transform -1 0 510 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1443_
timestamp 1727493435
transform -1 0 390 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1444_
timestamp 1727493435
transform -1 0 530 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1445_
timestamp 1727493435
transform -1 0 690 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1446_
timestamp 1727493435
transform -1 0 70 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1447_
timestamp 1727493435
transform 1 0 330 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1448_
timestamp 1727493435
transform -1 0 690 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1449_
timestamp 1727493435
transform 1 0 990 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1450_
timestamp 1727493435
transform -1 0 230 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1451_
timestamp 1727493435
transform 1 0 490 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1452_
timestamp 1727493435
transform 1 0 830 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1453_
timestamp 1727493435
transform -1 0 1690 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1454_
timestamp 1727493435
transform -1 0 670 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1455_
timestamp 1727493435
transform 1 0 210 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1456_
timestamp 1727493435
transform -1 0 70 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1457_
timestamp 1727493435
transform 1 0 370 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1458_
timestamp 1727493435
transform 1 0 690 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1459_
timestamp 1727493435
transform -1 0 550 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1460_
timestamp 1727493435
transform 1 0 1170 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1461_
timestamp 1727493435
transform 1 0 850 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1462_
timestamp 1727493435
transform -1 0 1370 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1463_
timestamp 1727493435
transform -1 0 70 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1464_
timestamp 1727493435
transform -1 0 210 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1465_
timestamp 1727493435
transform -1 0 730 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1466_
timestamp 1727493435
transform -1 0 570 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1467_
timestamp 1727493435
transform 1 0 370 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1468_
timestamp 1727493435
transform -1 0 1030 0 1 270
box -6 -8 26 272
use FILL  FILL_2__1469_
timestamp 1727493435
transform -1 0 1570 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1470_
timestamp 1727493435
transform -1 0 2070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1471_
timestamp 1727493435
transform -1 0 1890 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1472_
timestamp 1727493435
transform -1 0 1090 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1473_
timestamp 1727493435
transform 1 0 2130 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1474_
timestamp 1727493435
transform 1 0 2270 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1475_
timestamp 1727493435
transform -1 0 2610 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1476_
timestamp 1727493435
transform 1 0 3090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1477_
timestamp 1727493435
transform -1 0 5690 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1478_
timestamp 1727493435
transform -1 0 5390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1479_
timestamp 1727493435
transform -1 0 2210 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1480_
timestamp 1727493435
transform 1 0 3210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1481_
timestamp 1727493435
transform -1 0 3250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1482_
timestamp 1727493435
transform 1 0 4090 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1483_
timestamp 1727493435
transform 1 0 3550 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1484_
timestamp 1727493435
transform 1 0 1190 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1485_
timestamp 1727493435
transform 1 0 2350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1486_
timestamp 1727493435
transform 1 0 1430 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1487_
timestamp 1727493435
transform -1 0 550 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1488_
timestamp 1727493435
transform 1 0 550 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1489_
timestamp 1727493435
transform -1 0 70 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1490_
timestamp 1727493435
transform -1 0 1490 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1491_
timestamp 1727493435
transform 1 0 930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1492_
timestamp 1727493435
transform -1 0 870 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1493_
timestamp 1727493435
transform -1 0 670 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1494_
timestamp 1727493435
transform -1 0 510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1495_
timestamp 1727493435
transform -1 0 350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1496_
timestamp 1727493435
transform -1 0 410 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1497_
timestamp 1727493435
transform 1 0 1110 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1498_
timestamp 1727493435
transform -1 0 570 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1499_
timestamp 1727493435
transform 1 0 690 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1500_
timestamp 1727493435
transform 1 0 1170 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1501_
timestamp 1727493435
transform 1 0 1310 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1502_
timestamp 1727493435
transform -1 0 1070 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1503_
timestamp 1727493435
transform -1 0 650 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1504_
timestamp 1727493435
transform 1 0 910 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1505_
timestamp 1727493435
transform -1 0 750 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1506_
timestamp 1727493435
transform -1 0 590 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1507_
timestamp 1727493435
transform -1 0 250 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1508_
timestamp 1727493435
transform -1 0 70 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1509_
timestamp 1727493435
transform -1 0 70 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1510_
timestamp 1727493435
transform 1 0 50 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1511_
timestamp 1727493435
transform -1 0 190 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1512_
timestamp 1727493435
transform -1 0 70 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1513_
timestamp 1727493435
transform 1 0 230 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1514_
timestamp 1727493435
transform -1 0 410 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1515_
timestamp 1727493435
transform 1 0 210 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1516_
timestamp 1727493435
transform -1 0 70 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1517_
timestamp 1727493435
transform -1 0 390 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1518_
timestamp 1727493435
transform -1 0 850 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1519_
timestamp 1727493435
transform -1 0 1150 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1520_
timestamp 1727493435
transform 1 0 990 0 -1 790
box -6 -8 26 272
use FILL  FILL_2__1521_
timestamp 1727493435
transform 1 0 1150 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1522_
timestamp 1727493435
transform 1 0 970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1523_
timestamp 1727493435
transform -1 0 1310 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1524_
timestamp 1727493435
transform 1 0 1710 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1525_
timestamp 1727493435
transform 1 0 1970 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1526_
timestamp 1727493435
transform -1 0 1910 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1527_
timestamp 1727493435
transform 1 0 2010 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1528_
timestamp 1727493435
transform 1 0 2710 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1529_
timestamp 1727493435
transform -1 0 5070 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1530_
timestamp 1727493435
transform -1 0 4930 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1531_
timestamp 1727493435
transform -1 0 4610 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1532_
timestamp 1727493435
transform 1 0 3090 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1533_
timestamp 1727493435
transform -1 0 3330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1534_
timestamp 1727493435
transform 1 0 3470 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1535_
timestamp 1727493435
transform -1 0 3130 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1536_
timestamp 1727493435
transform 1 0 3490 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1537_
timestamp 1727493435
transform -1 0 190 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1538_
timestamp 1727493435
transform 1 0 1190 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1539_
timestamp 1727493435
transform -1 0 770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1540_
timestamp 1727493435
transform -1 0 650 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1541_
timestamp 1727493435
transform 1 0 990 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1542_
timestamp 1727493435
transform 1 0 1010 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1543_
timestamp 1727493435
transform 1 0 850 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1544_
timestamp 1727493435
transform 1 0 910 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1545_
timestamp 1727493435
transform -1 0 770 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1546_
timestamp 1727493435
transform 1 0 470 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1547_
timestamp 1727493435
transform -1 0 710 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1548_
timestamp 1727493435
transform -1 0 850 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1549_
timestamp 1727493435
transform 1 0 330 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1550_
timestamp 1727493435
transform -1 0 690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1551_
timestamp 1727493435
transform -1 0 70 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1552_
timestamp 1727493435
transform 1 0 170 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1553_
timestamp 1727493435
transform 1 0 50 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1554_
timestamp 1727493435
transform -1 0 70 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1555_
timestamp 1727493435
transform 1 0 210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1556_
timestamp 1727493435
transform 1 0 310 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1557_
timestamp 1727493435
transform 1 0 50 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1558_
timestamp 1727493435
transform -1 0 210 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1559_
timestamp 1727493435
transform -1 0 490 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1560_
timestamp 1727493435
transform 1 0 1050 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1561_
timestamp 1727493435
transform 1 0 1310 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1562_
timestamp 1727493435
transform 1 0 1030 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1563_
timestamp 1727493435
transform -1 0 1470 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1564_
timestamp 1727493435
transform 1 0 2650 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1565_
timestamp 1727493435
transform -1 0 1450 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1566_
timestamp 1727493435
transform 1 0 2190 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1567_
timestamp 1727493435
transform 1 0 1290 0 -1 1310
box -6 -8 26 272
use FILL  FILL_2__1568_
timestamp 1727493435
transform 1 0 1990 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1569_
timestamp 1727493435
transform 1 0 2270 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1570_
timestamp 1727493435
transform 1 0 2430 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1571_
timestamp 1727493435
transform -1 0 1170 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1572_
timestamp 1727493435
transform -1 0 1210 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1573_
timestamp 1727493435
transform -1 0 1730 0 1 1310
box -6 -8 26 272
use FILL  FILL_2__1574_
timestamp 1727493435
transform -1 0 1730 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1575_
timestamp 1727493435
transform 1 0 2110 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1576_
timestamp 1727493435
transform 1 0 2370 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1577_
timestamp 1727493435
transform -1 0 1770 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1578_
timestamp 1727493435
transform 1 0 2530 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1579_
timestamp 1727493435
transform 1 0 6410 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1580_
timestamp 1727493435
transform 1 0 6230 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1581_
timestamp 1727493435
transform 1 0 6090 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1582_
timestamp 1727493435
transform 1 0 2970 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1583_
timestamp 1727493435
transform -1 0 3010 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1584_
timestamp 1727493435
transform 1 0 3230 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1585_
timestamp 1727493435
transform -1 0 3310 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1586_
timestamp 1727493435
transform 1 0 2890 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1587_
timestamp 1727493435
transform -1 0 530 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1588_
timestamp 1727493435
transform 1 0 1010 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1589_
timestamp 1727493435
transform 1 0 870 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1590_
timestamp 1727493435
transform 1 0 690 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1591_
timestamp 1727493435
transform -1 0 550 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1592_
timestamp 1727493435
transform 1 0 50 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1593_
timestamp 1727493435
transform -1 0 70 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1594_
timestamp 1727493435
transform 1 0 210 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1595_
timestamp 1727493435
transform -1 0 230 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1596_
timestamp 1727493435
transform 1 0 370 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1597_
timestamp 1727493435
transform 1 0 370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1598_
timestamp 1727493435
transform -1 0 410 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1599_
timestamp 1727493435
transform -1 0 250 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1600_
timestamp 1727493435
transform 1 0 510 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1601_
timestamp 1727493435
transform 1 0 1190 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1602_
timestamp 1727493435
transform -1 0 1650 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1603_
timestamp 1727493435
transform 1 0 1790 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1604_
timestamp 1727493435
transform -1 0 1970 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1605_
timestamp 1727493435
transform 1 0 1590 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1606_
timestamp 1727493435
transform 1 0 2250 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1607_
timestamp 1727493435
transform 1 0 1430 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1608_
timestamp 1727493435
transform 1 0 1590 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1609_
timestamp 1727493435
transform 1 0 1750 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1610_
timestamp 1727493435
transform -1 0 5750 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1611_
timestamp 1727493435
transform -1 0 5590 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2__1612_
timestamp 1727493435
transform 1 0 790 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1613_
timestamp 1727493435
transform 1 0 2510 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1614_
timestamp 1727493435
transform -1 0 2570 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1615_
timestamp 1727493435
transform -1 0 2730 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1616_
timestamp 1727493435
transform -1 0 3030 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1617_
timestamp 1727493435
transform -1 0 1270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1618_
timestamp 1727493435
transform -1 0 1770 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1619_
timestamp 1727493435
transform 1 0 350 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1620_
timestamp 1727493435
transform 1 0 1470 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2__1621_
timestamp 1727493435
transform -1 0 1170 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1622_
timestamp 1727493435
transform 1 0 1630 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1623_
timestamp 1727493435
transform -1 0 1510 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1624_
timestamp 1727493435
transform 1 0 1790 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1625_
timestamp 1727493435
transform 1 0 2050 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1626_
timestamp 1727493435
transform 1 0 2050 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1627_
timestamp 1727493435
transform -1 0 2230 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1628_
timestamp 1727493435
transform 1 0 2110 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1629_
timestamp 1727493435
transform 1 0 2210 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1630_
timestamp 1727493435
transform 1 0 2370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1631_
timestamp 1727493435
transform -1 0 5810 0 -1 2350
box -6 -8 26 272
use FILL  FILL_2__1632_
timestamp 1727493435
transform 1 0 6150 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1633_
timestamp 1727493435
transform 1 0 6010 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1634_
timestamp 1727493435
transform 1 0 2370 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1635_
timestamp 1727493435
transform -1 0 3590 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1636_
timestamp 1727493435
transform -1 0 3410 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1637_
timestamp 1727493435
transform -1 0 2890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1638_
timestamp 1727493435
transform 1 0 2870 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1639_
timestamp 1727493435
transform 1 0 1870 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1640_
timestamp 1727493435
transform -1 0 1350 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1641_
timestamp 1727493435
transform 1 0 1950 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1642_
timestamp 1727493435
transform -1 0 5690 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1643_
timestamp 1727493435
transform -1 0 6050 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1644_
timestamp 1727493435
transform -1 0 5390 0 1 1830
box -6 -8 26 272
use FILL  FILL_2__1645_
timestamp 1727493435
transform 1 0 2390 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1646_
timestamp 1727493435
transform -1 0 2550 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1647_
timestamp 1727493435
transform 1 0 2690 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2__1648_
timestamp 1727493435
transform -1 0 2710 0 1 3390
box -6 -8 26 272
use FILL  FILL_2__1649_
timestamp 1727493435
transform -1 0 4650 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1650_
timestamp 1727493435
transform -1 0 4790 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1651_
timestamp 1727493435
transform 1 0 4610 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1652_
timestamp 1727493435
transform -1 0 4490 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1653_
timestamp 1727493435
transform 1 0 4690 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1654_
timestamp 1727493435
transform 1 0 4510 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1655_
timestamp 1727493435
transform 1 0 4490 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1656_
timestamp 1727493435
transform 1 0 4330 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1657_
timestamp 1727493435
transform 1 0 3950 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1658_
timestamp 1727493435
transform -1 0 3650 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1659_
timestamp 1727493435
transform -1 0 3470 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1660_
timestamp 1727493435
transform 1 0 3290 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1661_
timestamp 1727493435
transform 1 0 3170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1662_
timestamp 1727493435
transform 1 0 2990 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1663_
timestamp 1727493435
transform -1 0 3830 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1664_
timestamp 1727493435
transform 1 0 3710 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1692_
timestamp 1727493435
transform -1 0 3670 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1693_
timestamp 1727493435
transform -1 0 3930 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1694_
timestamp 1727493435
transform -1 0 3510 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1695_
timestamp 1727493435
transform 1 0 3310 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1696_
timestamp 1727493435
transform -1 0 2990 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1697_
timestamp 1727493435
transform -1 0 3790 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1698_
timestamp 1727493435
transform 1 0 4190 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1699_
timestamp 1727493435
transform 1 0 3510 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1700_
timestamp 1727493435
transform 1 0 3810 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1701_
timestamp 1727493435
transform 1 0 3630 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1702_
timestamp 1727493435
transform 1 0 3630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1703_
timestamp 1727493435
transform 1 0 3110 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1704_
timestamp 1727493435
transform 1 0 4470 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1705_
timestamp 1727493435
transform -1 0 3530 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1706_
timestamp 1727493435
transform -1 0 3910 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1707_
timestamp 1727493435
transform 1 0 3730 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1708_
timestamp 1727493435
transform -1 0 3430 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1709_
timestamp 1727493435
transform -1 0 3590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1710_
timestamp 1727493435
transform -1 0 3970 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1711_
timestamp 1727493435
transform -1 0 3790 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1712_
timestamp 1727493435
transform 1 0 2030 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1713_
timestamp 1727493435
transform 1 0 2490 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1714_
timestamp 1727493435
transform -1 0 2750 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1715_
timestamp 1727493435
transform 1 0 3010 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1716_
timestamp 1727493435
transform -1 0 3350 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1717_
timestamp 1727493435
transform -1 0 3210 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1718_
timestamp 1727493435
transform -1 0 2910 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1719_
timestamp 1727493435
transform 1 0 2810 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1720_
timestamp 1727493435
transform -1 0 2670 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1721_
timestamp 1727493435
transform 1 0 2770 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1722_
timestamp 1727493435
transform -1 0 3370 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1723_
timestamp 1727493435
transform 1 0 3010 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1724_
timestamp 1727493435
transform -1 0 3270 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1725_
timestamp 1727493435
transform -1 0 3390 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1726_
timestamp 1727493435
transform -1 0 3090 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1727_
timestamp 1727493435
transform -1 0 2930 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1728_
timestamp 1727493435
transform -1 0 2630 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1729_
timestamp 1727493435
transform -1 0 2470 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1730_
timestamp 1727493435
transform 1 0 2250 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1731_
timestamp 1727493435
transform -1 0 2590 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1732_
timestamp 1727493435
transform 1 0 2390 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1733_
timestamp 1727493435
transform -1 0 2370 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1734_
timestamp 1727493435
transform 1 0 3770 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1735_
timestamp 1727493435
transform -1 0 3630 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1736_
timestamp 1727493435
transform -1 0 4070 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1737_
timestamp 1727493435
transform 1 0 4170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1738_
timestamp 1727493435
transform -1 0 4050 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1739_
timestamp 1727493435
transform 1 0 3870 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1740_
timestamp 1727493435
transform -1 0 3470 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1741_
timestamp 1727493435
transform 1 0 3110 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1742_
timestamp 1727493435
transform 1 0 2490 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1743_
timestamp 1727493435
transform -1 0 1970 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1744_
timestamp 1727493435
transform 1 0 1930 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1745_
timestamp 1727493435
transform -1 0 1790 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1746_
timestamp 1727493435
transform 1 0 3970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1747_
timestamp 1727493435
transform 1 0 2110 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1748_
timestamp 1727493435
transform -1 0 1810 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1749_
timestamp 1727493435
transform -1 0 3250 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1750_
timestamp 1727493435
transform -1 0 3990 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1751_
timestamp 1727493435
transform 1 0 4050 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1752_
timestamp 1727493435
transform 1 0 3890 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1753_
timestamp 1727493435
transform 1 0 3550 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1754_
timestamp 1727493435
transform -1 0 3750 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1755_
timestamp 1727493435
transform -1 0 3410 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1756_
timestamp 1727493435
transform -1 0 2950 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1757_
timestamp 1727493435
transform -1 0 2790 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1758_
timestamp 1727493435
transform -1 0 2670 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1759_
timestamp 1727493435
transform 1 0 2330 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1760_
timestamp 1727493435
transform -1 0 2150 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1761_
timestamp 1727493435
transform 1 0 1490 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1762_
timestamp 1727493435
transform -1 0 1290 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1763_
timestamp 1727493435
transform -1 0 1450 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1764_
timestamp 1727493435
transform -1 0 1610 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1765_
timestamp 1727493435
transform 1 0 1130 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1766_
timestamp 1727493435
transform 1 0 2070 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1767_
timestamp 1727493435
transform -1 0 70 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1768_
timestamp 1727493435
transform -1 0 1350 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1769_
timestamp 1727493435
transform -1 0 1810 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1770_
timestamp 1727493435
transform -1 0 2650 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1771_
timestamp 1727493435
transform -1 0 2490 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1772_
timestamp 1727493435
transform 1 0 2090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1773_
timestamp 1727493435
transform 1 0 2570 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1774_
timestamp 1727493435
transform -1 0 1950 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1775_
timestamp 1727493435
transform 1 0 1790 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1776_
timestamp 1727493435
transform -1 0 1650 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1777_
timestamp 1727493435
transform -1 0 1490 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1778_
timestamp 1727493435
transform -1 0 1330 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1779_
timestamp 1727493435
transform -1 0 310 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1780_
timestamp 1727493435
transform 1 0 190 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1781_
timestamp 1727493435
transform 1 0 350 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1782_
timestamp 1727493435
transform -1 0 530 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1783_
timestamp 1727493435
transform 1 0 2730 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1784_
timestamp 1727493435
transform 1 0 1010 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1785_
timestamp 1727493435
transform -1 0 870 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1786_
timestamp 1727493435
transform 1 0 670 0 -1 6510
box -6 -8 26 272
use FILL  FILL_2__1787_
timestamp 1727493435
transform -1 0 450 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1788_
timestamp 1727493435
transform -1 0 1210 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1789_
timestamp 1727493435
transform 1 0 570 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1790_
timestamp 1727493435
transform 1 0 1610 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1791_
timestamp 1727493435
transform -1 0 2090 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1792_
timestamp 1727493435
transform -1 0 1950 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1793_
timestamp 1727493435
transform 1 0 1890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1794_
timestamp 1727493435
transform -1 0 1730 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1795_
timestamp 1727493435
transform -1 0 1570 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1796_
timestamp 1727493435
transform -1 0 1890 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1797_
timestamp 1727493435
transform -1 0 1710 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1798_
timestamp 1727493435
transform -1 0 1550 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1799_
timestamp 1727493435
transform -1 0 1390 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1800_
timestamp 1727493435
transform 1 0 890 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1801_
timestamp 1727493435
transform 1 0 1630 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1802_
timestamp 1727493435
transform -1 0 1190 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1803_
timestamp 1727493435
transform 1 0 1030 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1804_
timestamp 1727493435
transform -1 0 890 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1805_
timestamp 1727493435
transform -1 0 770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1806_
timestamp 1727493435
transform -1 0 750 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1807_
timestamp 1727493435
transform -1 0 1070 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1808_
timestamp 1727493435
transform -1 0 1270 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1809_
timestamp 1727493435
transform -1 0 1050 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1810_
timestamp 1727493435
transform -1 0 1790 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1811_
timestamp 1727493435
transform 1 0 1470 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1812_
timestamp 1727493435
transform 1 0 1350 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1813_
timestamp 1727493435
transform -1 0 1330 0 1 3910
box -6 -8 26 272
use FILL  FILL_2__1814_
timestamp 1727493435
transform -1 0 1210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1815_
timestamp 1727493435
transform 1 0 1770 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1816_
timestamp 1727493435
transform -1 0 1610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1817_
timestamp 1727493435
transform -1 0 1450 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1818_
timestamp 1727493435
transform -1 0 1290 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1819_
timestamp 1727493435
transform 1 0 1090 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1820_
timestamp 1727493435
transform -1 0 590 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1821_
timestamp 1727493435
transform 1 0 810 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1822_
timestamp 1727493435
transform -1 0 690 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1823_
timestamp 1727493435
transform -1 0 810 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1824_
timestamp 1727493435
transform -1 0 530 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1825_
timestamp 1727493435
transform 1 0 910 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1826_
timestamp 1727493435
transform -1 0 1690 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1827_
timestamp 1727493435
transform 1 0 1510 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1828_
timestamp 1727493435
transform 1 0 1330 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1829_
timestamp 1727493435
transform -1 0 1190 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1830_
timestamp 1727493435
transform -1 0 1010 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1831_
timestamp 1727493435
transform 1 0 1970 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1832_
timestamp 1727493435
transform -1 0 1830 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1833_
timestamp 1727493435
transform -1 0 1330 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1834_
timestamp 1727493435
transform -1 0 1170 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1835_
timestamp 1727493435
transform -1 0 970 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1836_
timestamp 1727493435
transform -1 0 950 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1837_
timestamp 1727493435
transform -1 0 350 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1838_
timestamp 1727493435
transform 1 0 610 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1839_
timestamp 1727493435
transform 1 0 1010 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1840_
timestamp 1727493435
transform 1 0 510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1841_
timestamp 1727493435
transform 1 0 450 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1842_
timestamp 1727493435
transform 1 0 2270 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1843_
timestamp 1727493435
transform 1 0 1830 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1844_
timestamp 1727493435
transform -1 0 2010 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1845_
timestamp 1727493435
transform -1 0 2150 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1846_
timestamp 1727493435
transform 1 0 1930 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1847_
timestamp 1727493435
transform 1 0 2110 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1848_
timestamp 1727493435
transform 1 0 2310 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1849_
timestamp 1727493435
transform -1 0 2170 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1850_
timestamp 1727493435
transform -1 0 1650 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1851_
timestamp 1727493435
transform -1 0 1490 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1852_
timestamp 1727493435
transform 1 0 550 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1853_
timestamp 1727493435
transform -1 0 70 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1854_
timestamp 1727493435
transform -1 0 230 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1855_
timestamp 1727493435
transform 1 0 210 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1856_
timestamp 1727493435
transform 1 0 630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1857_
timestamp 1727493435
transform -1 0 1990 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1858_
timestamp 1727493435
transform -1 0 2190 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1859_
timestamp 1727493435
transform 1 0 2430 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1860_
timestamp 1727493435
transform 1 0 710 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1861_
timestamp 1727493435
transform -1 0 850 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1862_
timestamp 1727493435
transform 1 0 1650 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1863_
timestamp 1727493435
transform 1 0 2430 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1864_
timestamp 1727493435
transform -1 0 70 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1865_
timestamp 1727493435
transform -1 0 390 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1866_
timestamp 1727493435
transform 1 0 50 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1867_
timestamp 1727493435
transform -1 0 650 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1868_
timestamp 1727493435
transform -1 0 3270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1869_
timestamp 1727493435
transform 1 0 1110 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2__1870_
timestamp 1727493435
transform -1 0 70 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1871_
timestamp 1727493435
transform -1 0 70 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1872_
timestamp 1727493435
transform -1 0 70 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1873_
timestamp 1727493435
transform -1 0 190 0 1 5990
box -6 -8 26 272
use FILL  FILL_2__1874_
timestamp 1727493435
transform -1 0 230 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1875_
timestamp 1727493435
transform -1 0 370 0 1 5470
box -6 -8 26 272
use FILL  FILL_2__1876_
timestamp 1727493435
transform -1 0 250 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1877_
timestamp 1727493435
transform 1 0 410 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2__1878_
timestamp 1727493435
transform 1 0 330 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1879_
timestamp 1727493435
transform -1 0 690 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1880_
timestamp 1727493435
transform -1 0 1390 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1881_
timestamp 1727493435
transform 1 0 1510 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1882_
timestamp 1727493435
transform -1 0 1070 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1883_
timestamp 1727493435
transform 1 0 1210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1884_
timestamp 1727493435
transform 1 0 910 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1885_
timestamp 1727493435
transform -1 0 790 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1886_
timestamp 1727493435
transform -1 0 370 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1887_
timestamp 1727493435
transform -1 0 230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1888_
timestamp 1727493435
transform 1 0 50 0 -1 4950
box -6 -8 26 272
use FILL  FILL_2__1889_
timestamp 1727493435
transform 1 0 370 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1890_
timestamp 1727493435
transform 1 0 510 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1891_
timestamp 1727493435
transform -1 0 210 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1892_
timestamp 1727493435
transform -1 0 210 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1893_
timestamp 1727493435
transform 1 0 490 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1894_
timestamp 1727493435
transform -1 0 850 0 1 4430
box -6 -8 26 272
use FILL  FILL_2__1895_
timestamp 1727493435
transform -1 0 70 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2__1896_
timestamp 1727493435
transform -1 0 4490 0 1 4950
box -6 -8 26 272
use FILL  FILL_2__1897_
timestamp 1727493435
transform 1 0 3910 0 1 790
box -6 -8 26 272
use FILL  FILL_2__1898_
timestamp 1727493435
transform 1 0 3610 0 1 2870
box -6 -8 26 272
use FILL  FILL_2__1899_
timestamp 1727493435
transform 1 0 3250 0 -1 270
box -6 -8 26 272
use FILL  FILL_2__1900_
timestamp 1727493435
transform 1 0 3150 0 -1 1830
box -6 -8 26 272
use FILL  FILL_2__1901_
timestamp 1727493435
transform -1 0 2750 0 1 2350
box -6 -8 26 272
use FILL  FILL_2__1902_
timestamp 1727493435
transform -1 0 5130 0 1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1727493435
transform -1 0 2310 0 1 2350
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1727493435
transform -1 0 2250 0 1 3910
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1727493435
transform 1 0 3910 0 1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1727493435
transform 1 0 3590 0 1 2350
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1727493435
transform -1 0 4790 0 1 4950
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert5
timestamp 1727493435
transform -1 0 4070 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1727493435
transform 1 0 4370 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert7
timestamp 1727493435
transform -1 0 4110 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert8
timestamp 1727493435
transform -1 0 4170 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert9
timestamp 1727493435
transform -1 0 4650 0 1 4430
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert10
timestamp 1727493435
transform 1 0 5050 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert11
timestamp 1727493435
transform 1 0 4770 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1727493435
transform -1 0 3610 0 1 3910
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1727493435
transform 1 0 4230 0 1 3910
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1727493435
transform -1 0 5210 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1727493435
transform -1 0 4930 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1727493435
transform 1 0 3810 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1727493435
transform -1 0 3690 0 -1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1727493435
transform -1 0 1930 0 1 2870
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1727493435
transform -1 0 1930 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1727493435
transform -1 0 4630 0 1 4950
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1727493435
transform 1 0 3910 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert27
timestamp 1727493435
transform 1 0 4390 0 1 3910
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1727493435
transform -1 0 3790 0 -1 3390
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1727493435
transform -1 0 2290 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert30
timestamp 1727493435
transform 1 0 2310 0 1 5470
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1727493435
transform 1 0 3110 0 -1 5990
box -6 -8 26 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1727493435
transform -1 0 4130 0 1 5990
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1727493435
transform 1 0 4230 0 -1 5470
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert13
timestamp 1727493435
transform -1 0 4130 0 1 3390
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 3890 0 -1 4430
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert15
timestamp 1727493435
transform -1 0 4190 0 -1 3910
box -6 -8 26 272
use FILL  FILL_2_CLKBUF1_insert16
timestamp 1727493435
transform 1 0 4190 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__930_
timestamp 1727493435
transform 1 0 6030 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__933_
timestamp 1727493435
transform 1 0 5470 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__937_
timestamp 1727493435
transform 1 0 5590 0 1 5470
box -6 -8 26 272
use FILL  FILL_3__941_
timestamp 1727493435
transform 1 0 3830 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__945_
timestamp 1727493435
transform 1 0 6270 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__948_
timestamp 1727493435
transform -1 0 5950 0 1 5470
box -6 -8 26 272
use FILL  FILL_3__952_
timestamp 1727493435
transform -1 0 5690 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__956_
timestamp 1727493435
transform -1 0 5830 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__960_
timestamp 1727493435
transform 1 0 6090 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__963_
timestamp 1727493435
transform -1 0 5530 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__967_
timestamp 1727493435
transform 1 0 4950 0 1 5470
box -6 -8 26 272
use FILL  FILL_3__971_
timestamp 1727493435
transform 1 0 4870 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__975_
timestamp 1727493435
transform 1 0 4450 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__978_
timestamp 1727493435
transform 1 0 3750 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__982_
timestamp 1727493435
transform 1 0 2090 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__986_
timestamp 1727493435
transform 1 0 3930 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__990_
timestamp 1727493435
transform -1 0 1790 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__993_
timestamp 1727493435
transform 1 0 5750 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__997_
timestamp 1727493435
transform 1 0 5490 0 1 4430
box -6 -8 26 272
use FILL  FILL_3__1000_
timestamp 1727493435
transform -1 0 4910 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1004_
timestamp 1727493435
transform 1 0 4690 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1008_
timestamp 1727493435
transform -1 0 5070 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1011_
timestamp 1727493435
transform 1 0 4970 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1015_
timestamp 1727493435
transform 1 0 5290 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1019_
timestamp 1727493435
transform 1 0 3990 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1023_
timestamp 1727493435
transform -1 0 4090 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1026_
timestamp 1727493435
transform -1 0 4550 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1030_
timestamp 1727493435
transform -1 0 5250 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1034_
timestamp 1727493435
transform -1 0 4350 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1038_
timestamp 1727493435
transform 1 0 4570 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1041_
timestamp 1727493435
transform 1 0 4970 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1045_
timestamp 1727493435
transform 1 0 5250 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1049_
timestamp 1727493435
transform 1 0 5090 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1052_
timestamp 1727493435
transform 1 0 5990 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1056_
timestamp 1727493435
transform -1 0 2930 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1060_
timestamp 1727493435
transform 1 0 3910 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1064_
timestamp 1727493435
transform -1 0 4030 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1067_
timestamp 1727493435
transform 1 0 4070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1071_
timestamp 1727493435
transform 1 0 4770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1075_
timestamp 1727493435
transform -1 0 4790 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1079_
timestamp 1727493435
transform 1 0 3790 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1082_
timestamp 1727493435
transform 1 0 5090 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1086_
timestamp 1727493435
transform 1 0 5430 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1090_
timestamp 1727493435
transform -1 0 5290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1094_
timestamp 1727493435
transform 1 0 4850 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1097_
timestamp 1727493435
transform -1 0 1630 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1101_
timestamp 1727493435
transform 1 0 5650 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1105_
timestamp 1727493435
transform 1 0 5330 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1109_
timestamp 1727493435
transform 1 0 6290 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1112_
timestamp 1727493435
transform -1 0 4290 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1116_
timestamp 1727493435
transform -1 0 3290 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1120_
timestamp 1727493435
transform -1 0 3870 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1124_
timestamp 1727493435
transform -1 0 3310 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1127_
timestamp 1727493435
transform -1 0 3450 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1131_
timestamp 1727493435
transform -1 0 3510 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1135_
timestamp 1727493435
transform 1 0 3570 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1138_
timestamp 1727493435
transform 1 0 4050 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1142_
timestamp 1727493435
transform -1 0 4090 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1146_
timestamp 1727493435
transform -1 0 4690 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1150_
timestamp 1727493435
transform -1 0 5230 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1153_
timestamp 1727493435
transform 1 0 6390 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1157_
timestamp 1727493435
transform 1 0 5910 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1161_
timestamp 1727493435
transform -1 0 5150 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1165_
timestamp 1727493435
transform -1 0 5630 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1168_
timestamp 1727493435
transform 1 0 5590 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1172_
timestamp 1727493435
transform 1 0 5410 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1176_
timestamp 1727493435
transform 1 0 5770 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1180_
timestamp 1727493435
transform 1 0 6430 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1183_
timestamp 1727493435
transform -1 0 4570 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1187_
timestamp 1727493435
transform 1 0 5570 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1191_
timestamp 1727493435
transform -1 0 5810 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1195_
timestamp 1727493435
transform 1 0 6290 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1198_
timestamp 1727493435
transform 1 0 6290 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1202_
timestamp 1727493435
transform 1 0 5970 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1206_
timestamp 1727493435
transform -1 0 5210 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1210_
timestamp 1727493435
transform -1 0 5670 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1213_
timestamp 1727493435
transform 1 0 6150 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1217_
timestamp 1727493435
transform -1 0 6270 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1221_
timestamp 1727493435
transform -1 0 4910 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1224_
timestamp 1727493435
transform 1 0 6190 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1228_
timestamp 1727493435
transform -1 0 6030 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1232_
timestamp 1727493435
transform 1 0 5190 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1236_
timestamp 1727493435
transform 1 0 6110 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1239_
timestamp 1727493435
transform 1 0 5930 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1243_
timestamp 1727493435
transform -1 0 5890 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1247_
timestamp 1727493435
transform 1 0 4410 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1251_
timestamp 1727493435
transform 1 0 4830 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1254_
timestamp 1727493435
transform 1 0 5030 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1258_
timestamp 1727493435
transform -1 0 4450 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1262_
timestamp 1727493435
transform -1 0 3150 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1266_
timestamp 1727493435
transform -1 0 2990 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1269_
timestamp 1727493435
transform -1 0 2650 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1273_
timestamp 1727493435
transform -1 0 2830 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1277_
timestamp 1727493435
transform 1 0 3250 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1281_
timestamp 1727493435
transform 1 0 3130 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1284_
timestamp 1727493435
transform 1 0 3450 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1288_
timestamp 1727493435
transform 1 0 3110 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1292_
timestamp 1727493435
transform 1 0 4550 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1295_
timestamp 1727493435
transform -1 0 3390 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1299_
timestamp 1727493435
transform 1 0 4050 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1303_
timestamp 1727493435
transform -1 0 3750 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1307_
timestamp 1727493435
transform -1 0 5850 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1310_
timestamp 1727493435
transform -1 0 2810 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1314_
timestamp 1727493435
transform -1 0 6370 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1318_
timestamp 1727493435
transform 1 0 6130 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1322_
timestamp 1727493435
transform 1 0 2870 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1325_
timestamp 1727493435
transform -1 0 2970 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1329_
timestamp 1727493435
transform -1 0 2950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1333_
timestamp 1727493435
transform 1 0 2070 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1337_
timestamp 1727493435
transform 1 0 3090 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1340_
timestamp 1727493435
transform -1 0 3570 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1344_
timestamp 1727493435
transform -1 0 2350 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1348_
timestamp 1727493435
transform -1 0 1970 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1352_
timestamp 1727493435
transform 1 0 3310 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1355_
timestamp 1727493435
transform -1 0 1310 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1359_
timestamp 1727493435
transform 1 0 1330 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1363_
timestamp 1727493435
transform 1 0 1670 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1367_
timestamp 1727493435
transform 1 0 1590 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1370_
timestamp 1727493435
transform -1 0 1430 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1374_
timestamp 1727493435
transform 1 0 2430 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1378_
timestamp 1727493435
transform 1 0 1610 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1381_
timestamp 1727493435
transform -1 0 910 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1385_
timestamp 1727493435
transform 1 0 1750 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1389_
timestamp 1727493435
transform -1 0 1210 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1393_
timestamp 1727493435
transform 1 0 1530 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1396_
timestamp 1727493435
transform 1 0 1970 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1400_
timestamp 1727493435
transform -1 0 2710 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1404_
timestamp 1727493435
transform 1 0 1710 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1408_
timestamp 1727493435
transform -1 0 4890 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1411_
timestamp 1727493435
transform -1 0 4550 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1415_
timestamp 1727493435
transform -1 0 2230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1419_
timestamp 1727493435
transform -1 0 1350 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1423_
timestamp 1727493435
transform -1 0 690 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1426_
timestamp 1727493435
transform 1 0 770 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1430_
timestamp 1727493435
transform 1 0 710 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1434_
timestamp 1727493435
transform -1 0 390 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1438_
timestamp 1727493435
transform -1 0 230 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1441_
timestamp 1727493435
transform -1 0 210 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1445_
timestamp 1727493435
transform -1 0 710 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1449_
timestamp 1727493435
transform 1 0 1010 0 1 790
box -6 -8 26 272
use FILL  FILL_3__1453_
timestamp 1727493435
transform -1 0 1710 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1456_
timestamp 1727493435
transform -1 0 90 0 1 270
box -6 -8 26 272
use FILL  FILL_3__1460_
timestamp 1727493435
transform 1 0 1190 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1464_
timestamp 1727493435
transform -1 0 230 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1467_
timestamp 1727493435
transform 1 0 390 0 -1 270
box -6 -8 26 272
use FILL  FILL_3__1471_
timestamp 1727493435
transform -1 0 1910 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1475_
timestamp 1727493435
transform -1 0 2630 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1479_
timestamp 1727493435
transform -1 0 2230 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1482_
timestamp 1727493435
transform 1 0 4110 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1486_
timestamp 1727493435
transform 1 0 1450 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1490_
timestamp 1727493435
transform -1 0 1510 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1494_
timestamp 1727493435
transform -1 0 530 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1497_
timestamp 1727493435
transform 1 0 1130 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1501_
timestamp 1727493435
transform 1 0 1330 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1505_
timestamp 1727493435
transform -1 0 770 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1509_
timestamp 1727493435
transform -1 0 90 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1512_
timestamp 1727493435
transform -1 0 90 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1516_
timestamp 1727493435
transform -1 0 90 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1520_
timestamp 1727493435
transform 1 0 1010 0 -1 790
box -6 -8 26 272
use FILL  FILL_3__1524_
timestamp 1727493435
transform 1 0 1730 0 1 1830
box -6 -8 26 272
use FILL  FILL_3__1527_
timestamp 1727493435
transform 1 0 2030 0 -1 2350
box -6 -8 26 272
use FILL  FILL_3__1531_
timestamp 1727493435
transform -1 0 4630 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1535_
timestamp 1727493435
transform -1 0 3150 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1539_
timestamp 1727493435
transform -1 0 790 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1542_
timestamp 1727493435
transform 1 0 1030 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1546_
timestamp 1727493435
transform 1 0 490 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1550_
timestamp 1727493435
transform -1 0 710 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1553_
timestamp 1727493435
transform 1 0 70 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1557_
timestamp 1727493435
transform 1 0 70 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1561_
timestamp 1727493435
transform 1 0 1330 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1565_
timestamp 1727493435
transform -1 0 1470 0 -1 1310
box -6 -8 26 272
use FILL  FILL_3__1568_
timestamp 1727493435
transform 1 0 2010 0 1 1310
box -6 -8 26 272
use FILL  FILL_3__1572_
timestamp 1727493435
transform -1 0 1230 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1576_
timestamp 1727493435
transform 1 0 2390 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1580_
timestamp 1727493435
transform 1 0 6250 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1583_
timestamp 1727493435
transform -1 0 3030 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1587_
timestamp 1727493435
transform -1 0 550 0 -1 3910
box -6 -8 26 272
use FILL  FILL_3__1591_
timestamp 1727493435
transform -1 0 570 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1595_
timestamp 1727493435
transform -1 0 250 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1598_
timestamp 1727493435
transform -1 0 430 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1602_
timestamp 1727493435
transform -1 0 1670 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1606_
timestamp 1727493435
transform 1 0 2270 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1610_
timestamp 1727493435
transform -1 0 5770 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3__1613_
timestamp 1727493435
transform 1 0 2530 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1617_
timestamp 1727493435
transform -1 0 1290 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1621_
timestamp 1727493435
transform -1 0 1190 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1624_
timestamp 1727493435
transform 1 0 1810 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1628_
timestamp 1727493435
transform 1 0 2130 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1632_
timestamp 1727493435
transform 1 0 6170 0 1 2350
box -6 -8 26 272
use FILL  FILL_3__1636_
timestamp 1727493435
transform -1 0 3430 0 1 3390
box -6 -8 26 272
use FILL  FILL_3__1639_
timestamp 1727493435
transform 1 0 1890 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1643_
timestamp 1727493435
transform -1 0 6070 0 -1 1830
box -6 -8 26 272
use FILL  FILL_3__1647_
timestamp 1727493435
transform 1 0 2710 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3__1651_
timestamp 1727493435
transform 1 0 4630 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1654_
timestamp 1727493435
transform 1 0 4530 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1658_
timestamp 1727493435
transform -1 0 3670 0 1 4430
box -6 -8 26 272
use FILL  FILL_3__1662_
timestamp 1727493435
transform 1 0 3010 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1693_
timestamp 1727493435
transform -1 0 3950 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1696_
timestamp 1727493435
transform -1 0 3010 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1700_
timestamp 1727493435
transform 1 0 3830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1704_
timestamp 1727493435
transform 1 0 4490 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1708_
timestamp 1727493435
transform -1 0 3450 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1711_
timestamp 1727493435
transform -1 0 3810 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1715_
timestamp 1727493435
transform 1 0 3030 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1719_
timestamp 1727493435
transform 1 0 2830 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1723_
timestamp 1727493435
transform 1 0 3030 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1726_
timestamp 1727493435
transform -1 0 3110 0 1 5470
box -6 -8 26 272
use FILL  FILL_3__1730_
timestamp 1727493435
transform 1 0 2270 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1734_
timestamp 1727493435
transform 1 0 3790 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1737_
timestamp 1727493435
transform 1 0 4190 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1741_
timestamp 1727493435
transform 1 0 3130 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1745_
timestamp 1727493435
transform -1 0 1810 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1749_
timestamp 1727493435
transform -1 0 3270 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1752_
timestamp 1727493435
transform 1 0 3910 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1756_
timestamp 1727493435
transform -1 0 2970 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1760_
timestamp 1727493435
transform -1 0 2170 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1764_
timestamp 1727493435
transform -1 0 1630 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1767_
timestamp 1727493435
transform -1 0 90 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1771_
timestamp 1727493435
transform -1 0 2510 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1775_
timestamp 1727493435
transform 1 0 1810 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1779_
timestamp 1727493435
transform -1 0 330 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1782_
timestamp 1727493435
transform -1 0 550 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1786_
timestamp 1727493435
transform 1 0 690 0 -1 6510
box -6 -8 26 272
use FILL  FILL_3__1790_
timestamp 1727493435
transform 1 0 1630 0 1 3910
box -6 -8 26 272
use FILL  FILL_3__1794_
timestamp 1727493435
transform -1 0 1750 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1797_
timestamp 1727493435
transform -1 0 1730 0 1 5470
box -6 -8 26 272
use FILL  FILL_3__1801_
timestamp 1727493435
transform 1 0 1650 0 1 5990
box -6 -8 26 272
use FILL  FILL_3__1805_
timestamp 1727493435
transform -1 0 790 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1809_
timestamp 1727493435
transform -1 0 1070 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1812_
timestamp 1727493435
transform 1 0 1370 0 -1 4430
box -6 -8 26 272
use FILL  FILL_3__1816_
timestamp 1727493435
transform -1 0 1630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1820_
timestamp 1727493435
transform -1 0 610 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1823_
timestamp 1727493435
transform -1 0 830 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1827_
timestamp 1727493435
transform 1 0 1530 0 1 4430
box -6 -8 26 272
use FILL  FILL_3__1831_
timestamp 1727493435
transform 1 0 1990 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1835_
timestamp 1727493435
transform -1 0 990 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1838_
timestamp 1727493435
transform 1 0 630 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1842_
timestamp 1727493435
transform 1 0 2290 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1846_
timestamp 1727493435
transform 1 0 1950 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1850_
timestamp 1727493435
transform -1 0 1670 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1853_
timestamp 1727493435
transform -1 0 90 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3__1857_
timestamp 1727493435
transform -1 0 2010 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1861_
timestamp 1727493435
transform -1 0 870 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1865_
timestamp 1727493435
transform -1 0 410 0 1 4950
box -6 -8 26 272
use FILL  FILL_3__1868_
timestamp 1727493435
transform -1 0 3290 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1872_
timestamp 1727493435
transform -1 0 90 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1876_
timestamp 1727493435
transform -1 0 270 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3__1880_
timestamp 1727493435
transform -1 0 1410 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1883_
timestamp 1727493435
transform 1 0 1230 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1887_
timestamp 1727493435
transform -1 0 250 0 -1 4950
box -6 -8 26 272
use FILL  FILL_3__1891_
timestamp 1727493435
transform -1 0 230 0 1 4430
box -6 -8 26 272
use FILL  FILL_3__1894_
timestamp 1727493435
transform -1 0 870 0 1 4430
box -6 -8 26 272
use FILL  FILL_3__1898_
timestamp 1727493435
transform 1 0 3630 0 1 2870
box -6 -8 26 272
use FILL  FILL_3__1902_
timestamp 1727493435
transform -1 0 5150 0 1 3390
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert3
timestamp 1727493435
transform 1 0 3610 0 1 2350
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert6
timestamp 1727493435
transform 1 0 4390 0 -1 3390
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert10
timestamp 1727493435
transform 1 0 5070 0 -1 5990
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert18
timestamp 1727493435
transform 1 0 4250 0 1 3910
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert21
timestamp 1727493435
transform 1 0 3830 0 -1 2870
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert25
timestamp 1727493435
transform -1 0 4650 0 1 4950
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert29
timestamp 1727493435
transform -1 0 2310 0 -1 5470
box -6 -8 26 272
use FILL  FILL_3_BUFX2_insert32
timestamp 1727493435
transform -1 0 4150 0 1 5990
box -6 -8 26 272
use FILL  FILL_3_CLKBUF1_insert14
timestamp 1727493435
transform -1 0 3910 0 -1 4430
box -6 -8 26 272
<< labels >>
flabel metal1 s 6517 2 6577 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -57 2 3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s 2256 6556 2264 6564 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal3 s 2296 6556 2304 6564 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal3 s 3316 6556 3324 6564 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal3 s 3496 6556 3504 6564 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal3 s 3976 6556 3984 6564 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal2 s 6557 6077 6563 6083 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal2 s 6557 5597 6563 5603 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal2 s 6557 5377 6563 5383 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal3 s 2776 -24 2784 -16 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal3 s 3196 -24 3204 -16 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal3 s 3296 -24 3304 -16 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal3 s 3676 -24 3684 -16 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal3 s 3956 -24 3964 -16 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal2 s -23 5077 -17 5083 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal2 s -23 4597 -17 4603 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal2 s -23 4557 -17 4563 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal3 s 5176 -24 5184 -16 7 FreeSans 16 270 0 0 Done_o
port 18 nsew
flabel metal3 s 6236 6556 6244 6564 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal3 s 6196 6556 6204 6564 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal3 s 5936 6556 5944 6564 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s 4256 6556 4264 6564 3 FreeSans 16 90 0 0 clk
port 22 nsew
flabel metal3 s 5556 6556 5564 6564 3 FreeSans 16 90 0 0 reset
port 23 nsew
<< properties >>
string FIXED_BBOX -40 -40 6560 6560
<< end >>
