** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1_TB.sch
**.subckt INVX1_TB
Vdd VDD GND 5
VAin A GND pulse(0 5 0 1n 1n 5n 12n)
R1 VDD Y 1Mega m=1
x1 A Y VDD GND INVX1
**** begin user architecture code



.include ~/ETRI050_DesignKit/tech/05cmos_model_240201.lib
.tran 0.01 70n
.dc VAin 0 5 0.01
.save all



**** end user architecture code
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sym # of pins=4
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sym
** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/INVX1.sch
.subckt INVX1 A Y vdd gnd
*.ipin A
*.opin Y
*.iopin vdd
*.iopin gnd
M1 Y A gnd GND nfet w=3u l=0.6u m=1
M2 Y A vdd VDD pfet w=6u l=0.6u m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
