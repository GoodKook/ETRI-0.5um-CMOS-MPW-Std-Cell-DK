magic
tech scmos
magscale 1 3
timestamp 1569139307
<< checkpaint >>
rect -60 -60 1260 2566
<< metal3 >>
rect 0 2340 1200 2506
rect 0 2110 1200 2276
rect 0 1130 1200 1910
rect 0 0 1200 780
<< end >>
