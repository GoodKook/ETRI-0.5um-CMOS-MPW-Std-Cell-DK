* NGSPICE file created from AND2X2.ext - technology: scmos

.subckt AND2X2 A B Y vdd gnd
M1000 Y a_4_12# gnd gnd nfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=5.4p ps=7.8u
M1001 a_18_12# A a_4_12# gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=9p ps=15.000001u
M1002 vdd B a_4_12# vdd pfet w=6u l=0.6u
+  ad=9.720001p pd=13.8u as=5.4p ps=7.8u
M1003 Y a_4_12# vdd vdd pfet w=12u l=0.6u
+  ad=18p pd=27.000002u as=9.720001p ps=13.8u
M1004 gnd B a_18_12# gnd nfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=2.7p ps=6.9u
M1005 a_4_12# A vdd vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=9p ps=15.000001u
.ends

