magic
tech scmos
magscale 1 2
timestamp 1728304789
<< nwell >>
rect -12 134 72 252
<< ntransistor >>
rect 21 14 25 34
<< ptransistor >>
rect 21 186 25 226
<< ndiffusion >>
rect 19 14 21 34
rect 25 14 27 34
<< pdiffusion >>
rect 19 186 21 226
rect 25 186 27 226
<< ndcontact >>
rect 7 14 19 34
rect 27 14 39 34
<< pdcontact >>
rect 7 186 19 226
rect 27 186 39 226
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 234 66 246
<< polysilicon >>
rect 21 226 25 230
rect 21 103 25 186
rect 16 91 25 103
rect 21 34 25 91
rect 21 10 25 14
<< polycontact >>
rect 4 91 16 103
<< metal1 >>
rect -6 246 66 248
rect -6 232 66 234
rect 7 226 19 232
rect 26 103 34 186
rect 26 34 34 89
rect 7 8 19 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m2contact >>
rect 3 77 17 91
rect 23 89 37 103
<< metal2 >>
rect 23 103 37 117
rect 3 63 17 77
<< m1p >>
rect -6 232 66 248
rect -6 -8 66 8
<< m2p >>
rect 23 103 37 117
rect 3 63 17 77
<< labels >>
rlabel metal1 -6 -8 66 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 66 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 3 63 17 77 0 A
port 0 nsew signal input
rlabel metal2 23 103 37 117 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
