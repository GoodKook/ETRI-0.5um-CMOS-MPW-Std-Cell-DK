/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module ALU8_Mult(
    inout vdd,
    inout gnd,
    input [7:0] ABCmd_i,
    output [7:0] ACC_o,
    input Flag_i,
    input LoadA_i,
    input LoadB_i,
    input LoadCmd_i,
    input MulH_i,
    input MulL_i,
    input clk,
    input reset
);

wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _873_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire [7:0] ABCmd_i ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire LoadA_i ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _864_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _799_ ;
wire _379_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire BCD ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _793_ ;
wire _373_ ;
wire _849_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire HC ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire [3:0] alu_op ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _881_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire [7:0] BI ;
wire _784_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _878_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _840_ ;
wire _420_ ;
wire \u_ALU8.AI7  ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire MUL ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _775_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire [7:0] ACC_o ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire [7:0] _919_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _898_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _895_ ;
wire _475_ ;
wire _284_ ;
wire [7:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire _187_ ;
wire _913_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire MulH_i ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _904_ ;
wire _713_ ;
wire [7:0] ACC ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _883_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _786_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _842_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire Flag_i ;
wire [7:0] AI ;
wire AN ;
wire AV ;
wire AZ ;
wire _783_ ;
wire _363_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire LoadB_i ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire MUL_bF$buf0 ;
wire MUL_bF$buf1 ;
wire MUL_bF$buf2 ;
wire MUL_bF$buf3 ;
wire MUL_bF$buf4 ;
wire MUL_bF$buf5 ;
wire _874_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _774_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire LoadCmd_i ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _897_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire shr ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire MulL_i ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire _186_ ;
wire _912_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire CI ;
wire CO ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _879_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire reset ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire alu_op_2_bF$buf0 ;
wire alu_op_2_bF$buf1 ;
wire alu_op_2_bF$buf2 ;
wire alu_op_2_bF$buf3 ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert14 (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf0)
);

BUFX2 BUFX2_insert13 (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf1)
);

BUFX2 BUFX2_insert12 (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf2)
);

BUFX2 BUFX2_insert11 (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[2]),
    .Y(alu_op_2_bF$buf3)
);

BUFX2 BUFX2_insert10 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf3)
);

BUFX2 BUFX2_insert6 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf4)
);

BUFX2 BUFX2_insert5 (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL),
    .Y(MUL_bF$buf5)
);

CLKBUF1 CLKBUF1_insert4 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert3 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert2 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert0 (
    .vdd(vdd),
    .gnd(gnd),
    .A(clk),
    .Y(clk_bF$buf4)
);

NAND3X1 _1000_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[1]),
    .C(AI[5]),
    .Y(_92_)
);

NAND3X1 _1001_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(BI[0]),
    .C(AI[6]),
    .Y(_93_)
);

NOR2X1 _1002_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_92_),
    .B(_93_),
    .Y(_94_)
);

AND2X2 _1003_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_92_),
    .B(_93_),
    .Y(_95_)
);

NAND3X1 _1004_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[2]),
    .C(AI[4]),
    .Y(_96_)
);

INVX1 _1005_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_96_),
    .Y(_97_)
);

OAI21X1 _1006_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_94_),
    .B(_95_),
    .C(_97_),
    .Y(_98_)
);

OR2X2 _1007_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_92_),
    .B(_93_),
    .Y(_99_)
);

OAI21X1 _1008_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_36_),
    .B(_54_),
    .C(_93_),
    .Y(_100_)
);

NAND3X1 _1009_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_100_),
    .B(_96_),
    .C(_99_),
    .Y(_101_)
);

NAND3X1 _1010_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_91_),
    .B(_98_),
    .C(_101_),
    .Y(_102_)
);

OAI21X1 _1011_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_56_),
    .B(_60_),
    .C(_52_),
    .Y(_103_)
);

NAND3X1 _1012_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_100_),
    .B(_97_),
    .C(_99_),
    .Y(_104_)
);

OAI21X1 _1013_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_94_),
    .B(_95_),
    .C(_96_),
    .Y(_105_)
);

NAND3X1 _1014_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_106_)
);

NAND3X1 _1015_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(BI[5]),
    .C(AI[1]),
    .Y(_107_)
);

INVX1 _1016_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_107_),
    .Y(_108_)
);

NAND3X1 _1017_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(BI[4]),
    .C(AI[2]),
    .Y(_109_)
);

NAND3X1 _1018_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(BI[3]),
    .C(AI[3]),
    .Y(_110_)
);

NOR2X1 _1019_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_109_),
    .B(_110_),
    .Y(_111_)
);

OAI21X1 _1020_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_44_),
    .C(_110_),
    .Y(_112_)
);

INVX1 _1021_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_112_),
    .Y(_113_)
);

OAI21X1 _1022_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_111_),
    .B(_113_),
    .C(_108_),
    .Y(_114_)
);

INVX1 _1023_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_109_),
    .Y(_115_)
);

INVX1 _1024_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_110_),
    .Y(_116_)
);

NAND2X1 _1025_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_115_),
    .B(_116_),
    .Y(_117_)
);

NAND3X1 _1026_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_107_),
    .B(_112_),
    .C(_117_),
    .Y(_118_)
);

NAND2X1 _1027_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_118_),
    .B(_114_),
    .Y(_119_)
);

NAND3X1 _1028_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_102_),
    .B(_119_),
    .C(_106_),
    .Y(_120_)
);

AOI21X1 _1029_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_121_)
);

AOI21X1 _1030_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_101_),
    .B(_98_),
    .C(_91_),
    .Y(_122_)
);

AND2X2 _1031_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_114_),
    .B(_118_),
    .Y(_123_)
);

OAI21X1 _1032_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_122_),
    .B(_121_),
    .C(_123_),
    .Y(_124_)
);

AOI21X1 _1033_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_125_)
);

AOI21X1 _1034_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_79_),
    .B(_66_),
    .C(_81_),
    .Y(_126_)
);

OAI21X1 _1035_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_122_),
    .B(_121_),
    .C(_119_),
    .Y(_127_)
);

NAND3X1 _1036_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_102_),
    .B(_106_),
    .C(_123_),
    .Y(_128_)
);

AOI21X1 _1037_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_127_),
    .B(_128_),
    .C(_126_),
    .Y(_129_)
);

NAND2X1 _1038_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .B(_68_),
    .Y(_130_)
);

AOI21X1 _1039_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_70_),
    .B(_74_),
    .C(_73_),
    .Y(_131_)
);

OR2X2 _1040_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_131_),
    .B(_130_),
    .Y(_132_)
);

INVX1 _1041_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .Y(_133_)
);

NOR2X1 _1042_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_715_),
    .B(_133_),
    .Y(_134_)
);

INVX4 _1043_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_134_),
    .Y(_135_)
);

OAI21X1 _1044_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_43_),
    .B(_135_),
    .C(_131_),
    .Y(_136_)
);

NAND2X1 _1045_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_136_),
    .B(_132_),
    .Y(_137_)
);

INVX1 _1046_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_137_),
    .Y(_138_)
);

OAI21X1 _1047_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_129_),
    .B(_125_),
    .C(_138_),
    .Y(_139_)
);

NAND3X1 _1048_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_128_),
    .B(_127_),
    .C(_126_),
    .Y(_140_)
);

NAND3X1 _1049_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_120_),
    .B(_124_),
    .C(_90_),
    .Y(_141_)
);

NAND3X1 _1050_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_137_),
    .B(_141_),
    .C(_140_),
    .Y(_142_)
);

NAND2X1 _1051_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_142_),
    .B(_139_),
    .Y(_143_)
);

NAND2X1 _1052_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_89_),
    .B(_143_),
    .Y(_144_)
);

INVX1 _1053_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_144_),
    .Y(_145_)
);

INVX1 _1054_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .Y(_146_)
);

AOI21X1 _1055_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_138_),
    .B(_140_),
    .C(_129_),
    .Y(_147_)
);

OAI21X1 _1056_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_121_),
    .B(_123_),
    .C(_106_),
    .Y(_148_)
);

AOI21X1 _1057_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_100_),
    .B(_97_),
    .C(_94_),
    .Y(_149_)
);

NAND3X1 _1058_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[1]),
    .C(AI[6]),
    .Y(_150_)
);

NAND3X1 _1059_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(BI[0]),
    .C(\u_ALU8.AI7 ),
    .Y(_151_)
);

NOR2X1 _1060_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_150_),
    .B(_151_),
    .Y(_152_)
);

AND2X2 _1061_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_150_),
    .B(_151_),
    .Y(_153_)
);

NAND3X1 _1062_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[2]),
    .C(AI[5]),
    .Y(_154_)
);

INVX1 _1063_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_154_),
    .Y(_155_)
);

OAI21X1 _1064_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_152_),
    .B(_153_),
    .C(_155_),
    .Y(_156_)
);

OR2X2 _1065_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_150_),
    .B(_151_),
    .Y(_157_)
);

NAND2X1 _1066_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(AI[6]),
    .Y(_158_)
);

OAI21X1 _1067_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_36_),
    .B(_158_),
    .C(_151_),
    .Y(_159_)
);

NAND3X1 _1068_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_159_),
    .B(_154_),
    .C(_157_),
    .Y(_160_)
);

NAND3X1 _1069_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_149_),
    .B(_156_),
    .C(_160_),
    .Y(_161_)
);

OAI21X1 _1070_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_96_),
    .B(_95_),
    .C(_99_),
    .Y(_162_)
);

NAND3X1 _1071_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_159_),
    .B(_155_),
    .C(_157_),
    .Y(_163_)
);

OAI21X1 _1072_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_152_),
    .B(_153_),
    .C(_154_),
    .Y(_164_)
);

NAND3X1 _1073_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_164_),
    .B(_162_),
    .C(_163_),
    .Y(_165_)
);

NAND3X1 _1074_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(BI[5]),
    .C(AI[2]),
    .Y(_166_)
);

INVX1 _1075_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_166_),
    .Y(_167_)
);

NAND3X1 _1076_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(AI[4]),
    .C(BI[4]),
    .Y(_168_)
);

INVX1 _1077_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[4]),
    .Y(_169_)
);

NAND3X1 _1078_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[3]),
    .C(AI[4]),
    .Y(_170_)
);

OAI21X1 _1079_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_169_),
    .B(_37_),
    .C(_170_),
    .Y(_171_)
);

OAI21X1 _1080_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_110_),
    .B(_168_),
    .C(_171_),
    .Y(_172_)
);

NAND2X1 _1081_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_167_),
    .B(_172_),
    .Y(_173_)
);

INVX1 _1082_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_168_),
    .Y(_174_)
);

NAND2X1 _1083_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_116_),
    .B(_174_),
    .Y(_175_)
);

NAND3X1 _1084_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_166_),
    .B(_171_),
    .C(_175_),
    .Y(_176_)
);

NAND2X1 _1085_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_176_),
    .B(_173_),
    .Y(_177_)
);

NAND3X1 _1086_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_161_),
    .B(_177_),
    .C(_165_),
    .Y(_178_)
);

AOI21X1 _1087_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_163_),
    .B(_164_),
    .C(_162_),
    .Y(_179_)
);

AOI21X1 _1088_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_160_),
    .B(_156_),
    .C(_149_),
    .Y(_180_)
);

NAND3X1 _1089_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_167_),
    .B(_171_),
    .C(_175_),
    .Y(_181_)
);

NAND2X1 _1090_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(BI[5]),
    .Y(_182_)
);

OAI21X1 _1091_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_182_),
    .C(_172_),
    .Y(_183_)
);

NAND2X1 _1092_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_181_),
    .B(_183_),
    .Y(_184_)
);

OAI21X1 _1093_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_180_),
    .B(_179_),
    .C(_184_),
    .Y(_185_)
);

AOI21X1 _1094_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_186_)
);

AOI21X1 _1095_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_119_),
    .B(_102_),
    .C(_122_),
    .Y(_187_)
);

OAI21X1 _1096_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_180_),
    .B(_179_),
    .C(_177_),
    .Y(_188_)
);

NAND3X1 _1097_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_161_),
    .B(_165_),
    .C(_184_),
    .Y(_189_)
);

AOI21X1 _1098_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_188_),
    .B(_189_),
    .C(_187_),
    .Y(_190_)
);

NAND2X1 _1099_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(_68_),
    .Y(_191_)
);

INVX1 _1100_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_191_),
    .Y(_192_)
);

AOI21X1 _1101_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_108_),
    .B(_112_),
    .C(_111_),
    .Y(_193_)
);

INVX1 _1102_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_193_),
    .Y(_194_)
);

OAI21X1 _1103_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_716_),
    .B(_135_),
    .C(_194_),
    .Y(_195_)
);

NAND2X1 _1104_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(_134_),
    .Y(_196_)
);

INVX1 _1105_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_196_),
    .Y(_197_)
);

NAND2X1 _1106_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_193_),
    .B(_197_),
    .Y(_198_)
);

NAND3X1 _1107_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_192_),
    .B(_198_),
    .C(_195_),
    .Y(_199_)
);

NAND2X1 _1108_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_197_),
    .B(_194_),
    .Y(_200_)
);

OAI21X1 _1109_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_716_),
    .B(_135_),
    .C(_193_),
    .Y(_201_)
);

NAND3X1 _1110_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_191_),
    .B(_201_),
    .C(_200_),
    .Y(_202_)
);

NAND2X1 _1111_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_202_),
    .B(_199_),
    .Y(_203_)
);

OAI21X1 _1112_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_186_),
    .C(_203_),
    .Y(_204_)
);

NAND3X1 _1113_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_189_),
    .B(_187_),
    .C(_188_),
    .Y(_205_)
);

NAND3X1 _1114_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_178_),
    .B(_185_),
    .C(_148_),
    .Y(_206_)
);

AND2X2 _1115_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_199_),
    .B(_202_),
    .Y(_207_)
);

NAND3X1 _1116_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_205_),
    .B(_206_),
    .C(_207_),
    .Y(_208_)
);

NAND3X1 _1117_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_208_),
    .B(_204_),
    .C(_147_),
    .Y(_209_)
);

OAI21X1 _1118_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_137_),
    .B(_125_),
    .C(_141_),
    .Y(_210_)
);

NAND3X1 _1119_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_203_),
    .B(_205_),
    .C(_206_),
    .Y(_211_)
);

OAI21X1 _1120_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_190_),
    .B(_186_),
    .C(_207_),
    .Y(_212_)
);

NAND3X1 _1121_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_211_),
    .B(_210_),
    .C(_212_),
    .Y(_213_)
);

NAND3X1 _1122_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_146_),
    .B(_213_),
    .C(_209_),
    .Y(_214_)
);

AOI21X1 _1123_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_212_),
    .B(_211_),
    .C(_210_),
    .Y(_215_)
);

AOI21X1 _1124_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_204_),
    .B(_208_),
    .C(_147_),
    .Y(_216_)
);

OAI21X1 _1125_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_215_),
    .B(_216_),
    .C(_132_),
    .Y(_217_)
);

NAND3X1 _1126_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_145_),
    .B(_214_),
    .C(_217_),
    .Y(_218_)
);

AOI21X1 _1127_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_217_),
    .B(_214_),
    .C(_145_),
    .Y(_219_)
);

NOR2X1 _1128_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_714_),
    .B(_718_),
    .Y(_220_)
);

INVX1 _1129_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .Y(_221_)
);

AOI21X1 _1130_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_221_),
    .B(_27_),
    .C(_722_),
    .Y(_222_)
);

OAI21X1 _1131_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_34_),
    .B(_40_),
    .C(_31_),
    .Y(_223_)
);

NAND3X1 _1132_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_30_),
    .B(_38_),
    .C(_35_),
    .Y(_224_)
);

AOI21X1 _1133_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_224_),
    .B(_223_),
    .C(_222_),
    .Y(_225_)
);

AND2X2 _1134_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_718_),
    .B(_714_),
    .Y(_226_)
);

NOR2X1 _1135_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_220_),
    .B(_226_),
    .Y(_227_)
);

NAND3X1 _1136_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_222_),
    .B(_223_),
    .C(_224_),
    .Y(_228_)
);

AOI21X1 _1137_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_227_),
    .B(_228_),
    .C(_225_),
    .Y(_229_)
);

OAI21X1 _1138_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_81_),
    .B(_82_),
    .C(_79_),
    .Y(_230_)
);

NAND3X1 _1139_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_66_),
    .B(_62_),
    .C(_85_),
    .Y(_231_)
);

NAND3X1 _1140_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_231_),
    .B(_230_),
    .C(_229_),
    .Y(_232_)
);

NAND3X1 _1141_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_220_),
    .B(_87_),
    .C(_232_),
    .Y(_233_)
);

NAND3X1 _1142_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_42_),
    .B(_228_),
    .C(_227_),
    .Y(_234_)
);

NAND3X1 _1143_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_221_),
    .B(_27_),
    .C(_723_),
    .Y(_235_)
);

NAND3X1 _1144_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[0]),
    .C(AI[2]),
    .Y(_236_)
);

INVX1 _1145_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_236_),
    .Y(_237_)
);

NAND3X1 _1146_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(BI[1]),
    .C(AI[1]),
    .Y(_238_)
);

INVX1 _1147_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_238_),
    .Y(_239_)
);

NAND2X1 _1148_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_237_),
    .B(_239_),
    .Y(_240_)
);

NAND2X1 _1149_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[2]),
    .B(_68_),
    .Y(_241_)
);

OAI21X1 _1150_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_716_),
    .B(_26_),
    .C(_236_),
    .Y(_242_)
);

INVX1 _1151_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_242_),
    .Y(_243_)
);

OAI21X1 _1152_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_241_),
    .B(_243_),
    .C(_240_),
    .Y(_244_)
);

OAI21X1 _1153_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .B(_28_),
    .C(_724_),
    .Y(_245_)
);

NAND3X1 _1154_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_244_),
    .B(_245_),
    .C(_235_),
    .Y(_246_)
);

NAND2X1 _1155_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .B(_68_),
    .Y(_247_)
);

AOI21X1 _1156_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_235_),
    .B(_245_),
    .C(_244_),
    .Y(_248_)
);

OAI21X1 _1157_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_247_),
    .B(_248_),
    .C(_246_),
    .Y(_249_)
);

OAI21X1 _1158_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_225_),
    .B(_47_),
    .C(_46_),
    .Y(_250_)
);

NAND3X1 _1159_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_234_),
    .B(_249_),
    .C(_250_),
    .Y(_251_)
);

INVX1 _1160_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_251_),
    .Y(_252_)
);

AOI21X1 _1161_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_230_),
    .B(_231_),
    .C(_229_),
    .Y(_253_)
);

OAI21X1 _1162_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_88_),
    .B(_253_),
    .C(_719_),
    .Y(_254_)
);

NAND3X1 _1163_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_233_),
    .B(_252_),
    .C(_254_),
    .Y(_255_)
);

INVX1 _1164_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_255_),
    .Y(_256_)
);

INVX1 _1165_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_89_),
    .Y(_257_)
);

NAND3X1 _1166_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_139_),
    .B(_142_),
    .C(_257_),
    .Y(_258_)
);

AND2X2 _1167_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_258_),
    .B(_144_),
    .Y(_259_)
);

INVX1 _1168_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_247_),
    .Y(_260_)
);

INVX1 _1169_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_248_),
    .Y(_261_)
);

NAND3X1 _1170_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_246_),
    .B(_260_),
    .C(_261_),
    .Y(_262_)
);

NAND2X1 _1171_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_242_),
    .B(_240_),
    .Y(_263_)
);

OR2X2 _1172_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_263_),
    .B(_241_),
    .Y(_264_)
);

NAND2X1 _1173_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[1]),
    .B(_68_),
    .Y(_265_)
);

NAND2X1 _1174_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_717_),
    .Y(_266_)
);

NOR2X1 _1175_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_265_),
    .B(_266_),
    .Y(_267_)
);

INVX1 _1176_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[2]),
    .Y(_268_)
);

OAI21X1 _1177_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_268_),
    .B(_67_),
    .C(_263_),
    .Y(_269_)
);

NAND3X1 _1178_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_267_),
    .B(_269_),
    .C(_264_),
    .Y(_270_)
);

INVX1 _1179_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_270_),
    .Y(_271_)
);

INVX1 _1180_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_246_),
    .Y(_272_)
);

OAI21X1 _1181_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_248_),
    .B(_272_),
    .C(_247_),
    .Y(_273_)
);

NAND3X1 _1182_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_271_),
    .B(_262_),
    .C(_273_),
    .Y(_274_)
);

AOI21X1 _1183_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_250_),
    .B(_234_),
    .C(_249_),
    .Y(_275_)
);

NOR3X1 _1184_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_275_),
    .B(_274_),
    .C(_252_),
    .Y(_276_)
);

OAI21X1 _1185_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_88_),
    .B(_253_),
    .C(_220_),
    .Y(_277_)
);

NAND3X1 _1186_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_719_),
    .B(_87_),
    .C(_232_),
    .Y(_278_)
);

NAND3X1 _1187_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_251_),
    .B(_278_),
    .C(_277_),
    .Y(_279_)
);

NAND3X1 _1188_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_276_),
    .B(_255_),
    .C(_279_),
    .Y(_280_)
);

INVX1 _1189_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .Y(_281_)
);

OAI21X1 _1190_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_256_),
    .B(_281_),
    .C(_259_),
    .Y(_282_)
);

OAI21X1 _1191_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .B(_282_),
    .C(_218_),
    .Y(_283_)
);

AOI21X1 _1192_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_209_),
    .B(_146_),
    .C(_216_),
    .Y(_284_)
);

NOR2X1 _1193_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_197_),
    .B(_194_),
    .Y(_285_)
);

OAI21X1 _1194_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_191_),
    .B(_285_),
    .C(_200_),
    .Y(_286_)
);

OAI21X1 _1195_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_207_),
    .B(_186_),
    .C(_206_),
    .Y(_287_)
);

INVX1 _1196_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .Y(_288_)
);

NOR2X1 _1197_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_715_),
    .B(_288_),
    .Y(_289_)
);

NAND2X1 _1198_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(_289_),
    .Y(_290_)
);

INVX1 _1199_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_290_),
    .Y(_291_)
);

NAND2X1 _1200_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .B(_134_),
    .Y(_292_)
);

AOI22X1 _1201_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_116_),
    .B(_174_),
    .C(_171_),
    .D(_167_),
    .Y(_293_)
);

OR2X2 _1202_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_293_),
    .B(_292_),
    .Y(_294_)
);

OAI21X1 _1203_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_135_),
    .C(_293_),
    .Y(_295_)
);

NAND3X1 _1204_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_291_),
    .B(_295_),
    .C(_294_),
    .Y(_296_)
);

NOR2X1 _1205_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_292_),
    .B(_293_),
    .Y(_297_)
);

AND2X2 _1206_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_293_),
    .B(_292_),
    .Y(_298_)
);

OAI21X1 _1207_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_297_),
    .B(_298_),
    .C(_290_),
    .Y(_299_)
);

NAND2X1 _1208_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_299_),
    .B(_296_),
    .Y(_300_)
);

AOI21X1 _1209_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_161_),
    .B(_177_),
    .C(_180_),
    .Y(_301_)
);

NAND3X1 _1210_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(AI[3]),
    .C(BI[5]),
    .Y(_302_)
);

NAND3X1 _1211_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(AI[5]),
    .C(BI[3]),
    .Y(_303_)
);

NOR2X1 _1212_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_168_),
    .B(_303_),
    .Y(_304_)
);

AND2X2 _1213_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_168_),
    .B(_303_),
    .Y(_305_)
);

OAI21X1 _1214_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_304_),
    .B(_305_),
    .C(_302_),
    .Y(_306_)
);

INVX1 _1215_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_302_),
    .Y(_307_)
);

OR2X2 _1216_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_168_),
    .B(_303_),
    .Y(_308_)
);

INVX1 _1217_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .Y(_309_)
);

OAI21X1 _1218_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_309_),
    .B(_54_),
    .C(_168_),
    .Y(_310_)
);

NAND3X1 _1219_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_307_),
    .B(_310_),
    .C(_308_),
    .Y(_311_)
);

NAND2X1 _1220_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_306_),
    .B(_311_),
    .Y(_312_)
);

AOI21X1 _1221_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_159_),
    .B(_155_),
    .C(_152_),
    .Y(_313_)
);

NAND3X1 _1222_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(AI[6]),
    .C(BI[2]),
    .Y(_314_)
);

NAND3X1 _1223_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(\u_ALU8.AI7 ),
    .C(BI[1]),
    .Y(_315_)
);

NOR2X1 _1224_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_315_),
    .Y(_316_)
);

AND2X2 _1225_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_315_),
    .Y(_317_)
);

NOR2X1 _1226_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_317_),
    .Y(_318_)
);

NAND2X1 _1227_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_313_),
    .B(_318_),
    .Y(_319_)
);

OAI21X1 _1228_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_153_),
    .B(_154_),
    .C(_157_),
    .Y(_320_)
);

OAI21X1 _1229_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_317_),
    .C(_320_),
    .Y(_321_)
);

NAND3X1 _1230_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_319_),
    .B(_312_),
    .C(_321_),
    .Y(_322_)
);

AND2X2 _1231_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_311_),
    .B(_306_),
    .Y(_323_)
);

NAND2X1 _1232_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_320_),
    .B(_318_),
    .Y(_324_)
);

OAI21X1 _1233_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_317_),
    .C(_313_),
    .Y(_325_)
);

NAND3X1 _1234_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_324_),
    .B(_325_),
    .C(_323_),
    .Y(_326_)
);

NAND3X1 _1235_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_326_),
    .C(_301_),
    .Y(_327_)
);

OAI21X1 _1236_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_184_),
    .B(_179_),
    .C(_165_),
    .Y(_328_)
);

AOI22X1 _1237_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_306_),
    .B(_311_),
    .C(_324_),
    .D(_325_),
    .Y(_329_)
);

AOI21X1 _1238_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_321_),
    .B(_319_),
    .C(_312_),
    .Y(_330_)
);

OAI21X1 _1239_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_330_),
    .C(_328_),
    .Y(_331_)
);

NAND3X1 _1240_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_331_),
    .C(_327_),
    .Y(_332_)
);

AND2X2 _1241_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_296_),
    .B(_299_),
    .Y(_333_)
);

NAND3X1 _1242_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_334_)
);

OAI21X1 _1243_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_335_)
);

NAND3X1 _1244_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_335_),
    .C(_334_),
    .Y(_336_)
);

NAND3X1 _1245_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_337_)
);

AOI21X1 _1246_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_203_),
    .B(_205_),
    .C(_190_),
    .Y(_338_)
);

AOI21X1 _1247_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_334_),
    .B(_335_),
    .C(_333_),
    .Y(_339_)
);

AOI21X1 _1248_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_327_),
    .B(_331_),
    .C(_300_),
    .Y(_340_)
);

OAI21X1 _1249_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_339_),
    .B(_340_),
    .C(_338_),
    .Y(_341_)
);

AOI21X1 _1250_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_337_),
    .B(_341_),
    .C(_286_),
    .Y(_342_)
);

INVX1 _1251_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_286_),
    .Y(_343_)
);

NAND3X1 _1252_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_332_),
    .B(_336_),
    .C(_338_),
    .Y(_344_)
);

OAI21X1 _1253_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_339_),
    .B(_340_),
    .C(_287_),
    .Y(_345_)
);

AOI21X1 _1254_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_345_),
    .B(_344_),
    .C(_343_),
    .Y(_346_)
);

OAI21X1 _1255_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_346_),
    .B(_342_),
    .C(_284_),
    .Y(_347_)
);

OAI21X1 _1256_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_132_),
    .B(_215_),
    .C(_213_),
    .Y(_348_)
);

NAND3X1 _1257_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_344_),
    .C(_345_),
    .Y(_349_)
);

NAND3X1 _1258_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_286_),
    .B(_341_),
    .C(_337_),
    .Y(_350_)
);

NAND3X1 _1259_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_349_),
    .B(_350_),
    .C(_348_),
    .Y(_351_)
);

AND2X2 _1260_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_347_),
    .B(_351_),
    .Y(_352_)
);

NAND2X1 _1261_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_283_),
    .Y(_353_)
);

INVX1 _1262_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_218_),
    .Y(_354_)
);

INVX1 _1263_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .Y(_355_)
);

NAND2X1 _1264_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_144_),
    .B(_258_),
    .Y(_356_)
);

NAND3X1 _1265_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_144_),
    .B(_258_),
    .C(_256_),
    .Y(_357_)
);

OAI21X1 _1266_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_356_),
    .C(_357_),
    .Y(_358_)
);

AOI21X1 _1267_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_355_),
    .B(_358_),
    .C(_354_),
    .Y(_359_)
);

NAND2X1 _1268_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .B(_347_),
    .Y(_360_)
);

NAND2X1 _1269_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_360_),
    .B(_359_),
    .Y(_361_)
);

NAND2X1 _1270_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_353_),
    .B(_361_),
    .Y(_362_)
);

NOR2X1 _1271_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ACC[0]),
    .B(Flag_i),
    .Y(_363_)
);

INVX1 _1272_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .Y(_364_)
);

INVX2 _1273_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MulL_i),
    .Y(_365_)
);

OAI21X1 _1274_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_364_),
    .C(_365_),
    .Y(_366_)
);

NAND3X1 _1275_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(MulL_i),
    .C(_68_),
    .Y(_367_)
);

OAI21X1 _1276_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_363_),
    .B(_366_),
    .C(_367_),
    .Y(_368_)
);

NAND2X1 _1277_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_368_),
    .Y(_369_)
);

OAI21X1 _1278_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_362_),
    .C(_369_),
    .Y(_0_[0])
);

AND2X2 _1279_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_266_),
    .B(_265_),
    .Y(_370_)
);

OAI21X1 _1280_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_267_),
    .B(_370_),
    .C(MulL_i),
    .Y(_371_)
);

MUX2X1 _1281_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(ACC[1]),
    .S(Flag_i),
    .Y(_372_)
);

AOI21X1 _1282_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_372_),
    .B(_365_),
    .C(MulH_i),
    .Y(_373_)
);

NAND2X1 _1283_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_373_),
    .B(_371_),
    .Y(_374_)
);

NAND2X1 _1284_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_332_),
    .B(_336_),
    .Y(_375_)
);

NOR2X1 _1285_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_338_),
    .B(_375_),
    .Y(_376_)
);

AOI21X1 _1286_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_286_),
    .B(_341_),
    .C(_376_),
    .Y(_377_)
);

OAI21X1 _1287_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_290_),
    .B(_298_),
    .C(_294_),
    .Y(_378_)
);

INVX1 _1288_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_378_),
    .Y(_379_)
);

NOR3X1 _1289_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_329_),
    .B(_330_),
    .C(_301_),
    .Y(_380_)
);

AOI21X1 _1290_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_333_),
    .B(_335_),
    .C(_380_),
    .Y(_381_)
);

NAND2X1 _1291_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .B(_289_),
    .Y(_382_)
);

INVX1 _1292_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_382_),
    .Y(_383_)
);

INVX1 _1293_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_37_),
    .Y(_384_)
);

OAI21X1 _1294_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_302_),
    .B(_305_),
    .C(_308_),
    .Y(_385_)
);

NAND3X1 _1295_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_384_),
    .B(_134_),
    .C(_385_),
    .Y(_386_)
);

INVX1 _1296_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[3]),
    .Y(_387_)
);

AOI21X1 _1297_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_307_),
    .B(_310_),
    .C(_304_),
    .Y(_388_)
);

OAI21X1 _1298_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_387_),
    .B(_135_),
    .C(_388_),
    .Y(_389_)
);

NAND3X1 _1299_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_383_),
    .B(_389_),
    .C(_386_),
    .Y(_390_)
);

NAND2X1 _1300_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .B(_384_),
    .Y(_391_)
);

NOR2X1 _1301_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_391_),
    .B(_388_),
    .Y(_392_)
);

AND2X2 _1302_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_388_),
    .B(_391_),
    .Y(_393_)
);

OAI21X1 _1303_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_392_),
    .B(_393_),
    .C(_382_),
    .Y(_394_)
);

NAND2X1 _1304_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_390_),
    .B(_394_),
    .Y(_395_)
);

NAND3X1 _1305_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(AI[4]),
    .C(BI[5]),
    .Y(_396_)
);

INVX1 _1306_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_396_),
    .Y(_397_)
);

NAND3X1 _1307_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(AI[5]),
    .C(BI[4]),
    .Y(_398_)
);

NAND3X1 _1308_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(AI[6]),
    .C(BI[3]),
    .Y(_399_)
);

OR2X2 _1309_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

INVX1 _1310_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .Y(_401_)
);

OAI21X1 _1311_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_401_),
    .B(_44_),
    .C(_399_),
    .Y(_402_)
);

AOI21X1 _1312_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_400_),
    .B(_402_),
    .C(_397_),
    .Y(_403_)
);

NAND3X1 _1313_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_399_),
    .C(_713_),
    .Y(_404_)
);

AND2X2 _1314_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(AI[6]),
    .Y(_405_)
);

NAND3X1 _1315_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .B(_398_),
    .C(_405_),
    .Y(_406_)
);

AOI21X1 _1316_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_404_),
    .B(_406_),
    .C(_396_),
    .Y(_407_)
);

NAND3X1 _1317_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(\u_ALU8.AI7 ),
    .C(BI[2]),
    .Y(_408_)
);

OAI22X1 _1318_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_408_),
    .C(_407_),
    .D(_403_),
    .Y(_409_)
);

NAND3X1 _1319_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_396_),
    .B(_404_),
    .C(_406_),
    .Y(_410_)
);

NAND3X1 _1320_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_397_),
    .B(_402_),
    .C(_400_),
    .Y(_411_)
);

NOR2X1 _1321_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_408_),
    .B(_316_),
    .Y(_412_)
);

NAND3X1 _1322_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_410_),
    .B(_412_),
    .C(_411_),
    .Y(_413_)
);

NAND2X1 _1323_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_413_),
    .B(_409_),
    .Y(_414_)
);

AOI21X1 _1324_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_326_),
    .B(_324_),
    .C(_414_),
    .Y(_415_)
);

OR2X2 _1325_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_314_),
    .B(_315_),
    .Y(_416_)
);

INVX2 _1326_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .Y(_417_)
);

OAI21X1 _1327_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_26_),
    .C(_314_),
    .Y(_418_)
);

AOI21X1 _1328_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_416_),
    .B(_418_),
    .C(_320_),
    .Y(_419_)
);

OAI21X1 _1329_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_312_),
    .B(_419_),
    .C(_324_),
    .Y(_420_)
);

AOI21X1 _1330_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_409_),
    .B(_413_),
    .C(_420_),
    .Y(_421_)
);

OAI21X1 _1331_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_415_),
    .B(_421_),
    .C(_395_),
    .Y(_422_)
);

AND2X2 _1332_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_394_),
    .B(_390_),
    .Y(_423_)
);

AND2X2 _1333_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_318_),
    .B(_320_),
    .Y(_424_)
);

AND2X2 _1334_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_409_),
    .B(_413_),
    .Y(_425_)
);

OAI21X1 _1335_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_424_),
    .B(_330_),
    .C(_425_),
    .Y(_426_)
);

AOI21X1 _1336_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_323_),
    .B(_325_),
    .C(_424_),
    .Y(_427_)
);

NAND2X1 _1337_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_414_),
    .B(_427_),
    .Y(_428_)
);

NAND3X1 _1338_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_428_),
    .B(_423_),
    .C(_426_),
    .Y(_429_)
);

NAND3X1 _1339_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_422_),
    .B(_429_),
    .C(_381_),
    .Y(_430_)
);

AOI21X1 _1340_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_322_),
    .B(_326_),
    .C(_328_),
    .Y(_431_)
);

OAI21X1 _1341_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_300_),
    .B(_431_),
    .C(_334_),
    .Y(_432_)
);

AOI21X1 _1342_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_426_),
    .B(_428_),
    .C(_423_),
    .Y(_433_)
);

NAND2X1 _1343_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_427_),
    .B(_425_),
    .Y(_434_)
);

OAI21X1 _1344_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_424_),
    .B(_330_),
    .C(_414_),
    .Y(_435_)
);

AOI21X1 _1345_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_434_),
    .B(_435_),
    .C(_395_),
    .Y(_436_)
);

OAI21X1 _1346_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_436_),
    .B(_433_),
    .C(_432_),
    .Y(_437_)
);

AOI21X1 _1347_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_430_),
    .B(_437_),
    .C(_379_),
    .Y(_438_)
);

NAND3X1 _1348_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_429_),
    .B(_422_),
    .C(_432_),
    .Y(_439_)
);

OAI21X1 _1349_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_433_),
    .B(_436_),
    .C(_381_),
    .Y(_440_)
);

AOI21X1 _1350_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_440_),
    .B(_439_),
    .C(_378_),
    .Y(_441_)
);

OAI21X1 _1351_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_438_),
    .B(_441_),
    .C(_377_),
    .Y(_442_)
);

AOI21X1 _1352_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_332_),
    .B(_336_),
    .C(_287_),
    .Y(_443_)
);

OAI21X1 _1353_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_343_),
    .B(_443_),
    .C(_337_),
    .Y(_444_)
);

NAND3X1 _1354_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_378_),
    .B(_439_),
    .C(_440_),
    .Y(_445_)
);

NAND3X1 _1355_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_379_),
    .B(_437_),
    .C(_430_),
    .Y(_446_)
);

NAND3X1 _1356_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_445_),
    .B(_446_),
    .C(_444_),
    .Y(_447_)
);

NAND2X1 _1357_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_447_),
    .B(_442_),
    .Y(_448_)
);

AOI21X1 _1358_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_353_),
    .B(_351_),
    .C(_448_),
    .Y(_449_)
);

OAI21X1 _1359_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_360_),
    .B(_359_),
    .C(_351_),
    .Y(_450_)
);

AND2X2 _1360_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_442_),
    .B(_447_),
    .Y(_451_)
);

OAI21X1 _1361_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_451_),
    .B(_450_),
    .C(MulH_i),
    .Y(_452_)
);

OAI21X1 _1362_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_449_),
    .B(_452_),
    .C(_374_),
    .Y(_0_[1])
);

NAND2X1 _1363_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_352_),
    .B(_451_),
    .Y(_453_)
);

NAND2X1 _1364_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_447_),
    .B(_351_),
    .Y(_454_)
);

NAND2X1 _1365_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_442_),
    .B(_454_),
    .Y(_455_)
);

OAI21X1 _1366_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_453_),
    .B(_359_),
    .C(_455_),
    .Y(_456_)
);

OAI21X1 _1367_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_382_),
    .B(_393_),
    .C(_386_),
    .Y(_457_)
);

INVX1 _1368_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_457_),
    .Y(_458_)
);

AOI21X1 _1369_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_423_),
    .B(_428_),
    .C(_415_),
    .Y(_459_)
);

NAND2X1 _1370_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(_384_),
    .Y(_460_)
);

INVX1 _1371_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_460_),
    .Y(_461_)
);

NOR2X1 _1372_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_398_),
    .B(_399_),
    .Y(_462_)
);

INVX1 _1373_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .Y(_463_)
);

NOR2X1 _1374_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_715_),
    .B(_463_),
    .Y(_464_)
);

NAND2X1 _1375_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .B(_464_),
    .Y(_465_)
);

INVX1 _1376_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .Y(_466_)
);

OAI21X1 _1377_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_462_),
    .B(_407_),
    .C(_466_),
    .Y(_467_)
);

AOI21X1 _1378_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_397_),
    .B(_402_),
    .C(_462_),
    .Y(_468_)
);

OAI21X1 _1379_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_463_),
    .B(_135_),
    .C(_468_),
    .Y(_469_)
);

NAND3X1 _1380_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_461_),
    .B(_469_),
    .C(_467_),
    .Y(_470_)
);

NOR2X1 _1381_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_465_),
    .B(_468_),
    .Y(_471_)
);

AND2X2 _1382_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_468_),
    .B(_465_),
    .Y(_472_)
);

OAI21X1 _1383_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_471_),
    .B(_472_),
    .C(_460_),
    .Y(_473_)
);

NAND2X1 _1384_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_473_),
    .Y(_474_)
);

NAND3X1 _1385_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(AI[5]),
    .C(BI[5]),
    .Y(_475_)
);

INVX1 _1386_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_475_),
    .Y(_476_)
);

NAND3X1 _1387_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(AI[6]),
    .C(BI[4]),
    .Y(_477_)
);

NAND3X1 _1388_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(\u_ALU8.AI7 ),
    .C(BI[3]),
    .Y(_478_)
);

OR2X2 _1389_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_477_),
    .B(_478_),
    .Y(_479_)
);

INVX1 _1390_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[6]),
    .Y(_480_)
);

OAI21X1 _1391_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_480_),
    .B(_44_),
    .C(_478_),
    .Y(_481_)
);

NAND3X1 _1392_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_476_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

NOR2X1 _1393_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_477_),
    .B(_478_),
    .Y(_483_)
);

AND2X2 _1394_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_477_),
    .B(_478_),
    .Y(_484_)
);

OAI21X1 _1395_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_483_),
    .B(_484_),
    .C(_475_),
    .Y(_485_)
);

NAND2X1 _1396_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_485_),
    .B(_482_),
    .Y(_486_)
);

AOI21X1 _1397_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_413_),
    .B(_416_),
    .C(_486_),
    .Y(_487_)
);

NAND3X1 _1398_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_416_),
    .B(_486_),
    .C(_413_),
    .Y(_488_)
);

INVX1 _1399_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_488_),
    .Y(_489_)
);

OAI21X1 _1400_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_489_),
    .C(_474_),
    .Y(_490_)
);

AND2X2 _1401_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_473_),
    .B(_470_),
    .Y(_491_)
);

INVX1 _1402_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .Y(_492_)
);

NAND3X1 _1403_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_492_),
    .B(_488_),
    .C(_491_),
    .Y(_493_)
);

NAND3X1 _1404_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_490_),
    .B(_493_),
    .C(_459_),
    .Y(_494_)
);

OAI21X1 _1405_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_395_),
    .B(_421_),
    .C(_426_),
    .Y(_495_)
);

AOI22X1 _1406_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_470_),
    .B(_473_),
    .C(_492_),
    .D(_488_),
    .Y(_496_)
);

INVX1 _1407_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_486_),
    .Y(_497_)
);

NAND3X1 _1408_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_416_),
    .B(_413_),
    .C(_497_),
    .Y(_498_)
);

INVX1 _1409_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_413_),
    .Y(_499_)
);

OAI21X1 _1410_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_316_),
    .B(_499_),
    .C(_486_),
    .Y(_500_)
);

AOI21X1 _1411_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_498_),
    .B(_500_),
    .C(_474_),
    .Y(_501_)
);

OAI21X1 _1412_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_496_),
    .B(_501_),
    .C(_495_),
    .Y(_502_)
);

NAND3X1 _1413_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_458_),
    .B(_502_),
    .C(_494_),
    .Y(_503_)
);

NAND3X1 _1414_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_504_)
);

OAI21X1 _1415_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_505_)
);

NAND3X1 _1416_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_457_),
    .B(_504_),
    .C(_505_),
    .Y(_506_)
);

NAND2X1 _1417_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_503_),
    .B(_506_),
    .Y(_507_)
);

NAND3X1 _1418_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_439_),
    .B(_445_),
    .C(_507_),
    .Y(_508_)
);

AOI21X1 _1419_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_422_),
    .B(_429_),
    .C(_432_),
    .Y(_509_)
);

OAI21X1 _1420_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_379_),
    .B(_509_),
    .C(_439_),
    .Y(_510_)
);

NAND3X1 _1421_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_503_),
    .B(_506_),
    .C(_510_),
    .Y(_511_)
);

NAND2X1 _1422_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .B(_508_),
    .Y(_512_)
);

INVX1 _1423_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_512_),
    .Y(_513_)
);

NAND2X1 _1424_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_513_),
    .B(_456_),
    .Y(_514_)
);

OR2X2 _1425_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_456_),
    .B(_513_),
    .Y(_515_)
);

NAND2X1 _1426_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_514_),
    .B(_515_),
    .Y(_516_)
);

AND2X2 _1427_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_264_),
    .B(_269_),
    .Y(_517_)
);

NOR2X1 _1428_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_365_),
    .B(_271_),
    .Y(_518_)
);

OAI21X1 _1429_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_267_),
    .B(_517_),
    .C(_518_),
    .Y(_519_)
);

NOR2X1 _1430_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .B(ACC[2]),
    .Y(_520_)
);

OAI21X1 _1431_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AZ),
    .B(_364_),
    .C(_365_),
    .Y(_521_)
);

OAI21X1 _1432_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_520_),
    .B(_521_),
    .C(_519_),
    .Y(_522_)
);

NAND2X1 _1433_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_522_),
    .Y(_523_)
);

OAI21X1 _1434_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_516_),
    .C(_523_),
    .Y(_0_[2])
);

NOR3X1 _1435_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_496_),
    .B(_501_),
    .C(_459_),
    .Y(_524_)
);

AOI21X1 _1436_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_457_),
    .B(_505_),
    .C(_524_),
    .Y(_525_)
);

OAI21X1 _1437_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_460_),
    .B(_472_),
    .C(_467_),
    .Y(_526_)
);

INVX1 _1438_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_526_),
    .Y(_527_)
);

AOI21X1 _1439_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_491_),
    .B(_488_),
    .C(_487_),
    .Y(_528_)
);

NAND2X1 _1440_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[7]),
    .B(_464_),
    .Y(_529_)
);

INVX1 _1441_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .Y(_530_)
);

OAI21X1 _1442_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_475_),
    .B(_484_),
    .C(_479_),
    .Y(_531_)
);

NAND3X1 _1443_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_134_),
    .C(_531_),
    .Y(_532_)
);

AOI21X1 _1444_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_476_),
    .B(_481_),
    .C(_483_),
    .Y(_533_)
);

OAI21X1 _1445_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_401_),
    .B(_135_),
    .C(_533_),
    .Y(_534_)
);

NAND3X1 _1446_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_530_),
    .B(_534_),
    .C(_532_),
    .Y(_535_)
);

INVX1 _1447_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_535_),
    .Y(_536_)
);

AOI21X1 _1448_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_532_),
    .B(_534_),
    .C(_530_),
    .Y(_537_)
);

NAND2X1 _1449_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[5]),
    .B(_405_),
    .Y(_538_)
);

NAND2X1 _1450_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_713_),
    .Y(_539_)
);

OR2X2 _1451_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_538_),
    .B(_539_),
    .Y(_540_)
);

OAI21X1 _1452_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_44_),
    .C(_538_),
    .Y(_541_)
);

NAND2X1 _1453_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_541_),
    .B(_540_),
    .Y(_542_)
);

OAI21X1 _1454_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_537_),
    .B(_536_),
    .C(_542_),
    .Y(_543_)
);

INVX1 _1455_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_537_),
    .Y(_544_)
);

INVX1 _1456_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_542_),
    .Y(_545_)
);

NAND3X1 _1457_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_535_),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

NAND3X1 _1458_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_546_),
    .C(_528_),
    .Y(_547_)
);

NAND2X1 _1459_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_546_),
    .Y(_548_)
);

OAI21X1 _1460_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_487_),
    .B(_501_),
    .C(_548_),
    .Y(_549_)
);

NAND3X1 _1461_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_527_),
    .B(_549_),
    .C(_547_),
    .Y(_550_)
);

OAI21X1 _1462_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_489_),
    .B(_474_),
    .C(_492_),
    .Y(_551_)
);

NAND3X1 _1463_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_543_),
    .B(_546_),
    .C(_551_),
    .Y(_552_)
);

NAND2X1 _1464_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_548_),
    .B(_528_),
    .Y(_553_)
);

NAND3X1 _1465_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_526_),
    .B(_552_),
    .C(_553_),
    .Y(_554_)
);

NAND2X1 _1466_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_554_),
    .B(_550_),
    .Y(_555_)
);

NAND2X1 _1467_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_525_),
    .B(_555_),
    .Y(_556_)
);

AOI21X1 _1468_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_490_),
    .B(_493_),
    .C(_495_),
    .Y(_557_)
);

OAI21X1 _1469_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_458_),
    .B(_557_),
    .C(_504_),
    .Y(_558_)
);

NAND3X1 _1470_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_550_),
    .B(_554_),
    .C(_558_),
    .Y(_559_)
);

NAND2X1 _1471_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_559_),
    .B(_556_),
    .Y(_560_)
);

NAND3X1 _1472_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .B(_560_),
    .C(_514_),
    .Y(_561_)
);

INVX1 _1473_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_511_),
    .Y(_562_)
);

NOR2X1 _1474_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_360_),
    .B(_448_),
    .Y(_563_)
);

NAND2X1 _1475_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_283_),
    .B(_563_),
    .Y(_564_)
);

AOI21X1 _1476_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_564_),
    .B(_455_),
    .C(_512_),
    .Y(_565_)
);

INVX1 _1477_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_560_),
    .Y(_566_)
);

OAI21X1 _1478_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_562_),
    .B(_565_),
    .C(_566_),
    .Y(_567_)
);

NAND2X1 _1479_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_561_),
    .B(_567_),
    .Y(_568_)
);

NAND2X1 _1480_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_262_),
    .B(_273_),
    .Y(_569_)
);

OAI21X1 _1481_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_270_),
    .B(_569_),
    .C(MulL_i),
    .Y(_570_)
);

AOI21X1 _1482_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_270_),
    .B(_569_),
    .C(_570_),
    .Y(_571_)
);

INVX1 _1483_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AV),
    .Y(_572_)
);

OAI21X1 _1484_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .B(ACC[3]),
    .C(_365_),
    .Y(_573_)
);

AOI21X1 _1485_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

OAI21X1 _1486_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_574_),
    .B(_571_),
    .C(_712_),
    .Y(_575_)
);

OAI21X1 _1487_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_568_),
    .C(_575_),
    .Y(_0_[3])
);

OAI21X1 _1488_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_528_),
    .B(_548_),
    .C(_554_),
    .Y(_576_)
);

INVX1 _1489_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_576_),
    .Y(_577_)
);

NAND2X1 _1490_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_534_),
    .B(_532_),
    .Y(_578_)
);

OAI21X1 _1491_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_529_),
    .B(_578_),
    .C(_532_),
    .Y(_579_)
);

INVX1 _1492_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .Y(_580_)
);

NAND2X1 _1493_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_289_),
    .Y(_581_)
);

NAND2X1 _1494_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[6]),
    .B(_405_),
    .Y(_582_)
);

OAI21X1 _1495_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_538_),
    .B(_539_),
    .C(_582_),
    .Y(_583_)
);

OAI21X1 _1496_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_540_),
    .C(_583_),
    .Y(_584_)
);

OR2X2 _1497_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_584_),
    .B(_581_),
    .Y(_585_)
);

OAI21X1 _1498_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_288_),
    .B(_54_),
    .C(_584_),
    .Y(_586_)
);

NAND2X1 _1499_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_586_),
    .B(_585_),
    .Y(_587_)
);

OAI21X1 _1500_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_417_),
    .B(_182_),
    .C(_587_),
    .Y(_588_)
);

INVX1 _1501_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_182_),
    .Y(_589_)
);

NAND2X1 _1502_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_589_),
    .Y(_590_)
);

INVX1 _1503_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_590_),
    .Y(_591_)
);

NAND3X1 _1504_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_586_),
    .B(_591_),
    .C(_585_),
    .Y(_592_)
);

NAND2X1 _1505_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_592_),
    .B(_588_),
    .Y(_593_)
);

NOR2X1 _1506_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_546_),
    .B(_593_),
    .Y(_594_)
);

AND2X2 _1507_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_593_),
    .B(_546_),
    .Y(_595_)
);

OAI21X1 _1508_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_594_),
    .B(_595_),
    .C(_580_),
    .Y(_596_)
);

OR2X2 _1509_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_593_),
    .B(_546_),
    .Y(_597_)
);

NAND2X1 _1510_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_546_),
    .B(_593_),
    .Y(_598_)
);

NAND3X1 _1511_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .B(_598_),
    .C(_597_),
    .Y(_599_)
);

NAND2X1 _1512_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_596_),
    .B(_599_),
    .Y(_600_)
);

NAND2X1 _1513_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_577_),
    .B(_600_),
    .Y(_601_)
);

NAND3X1 _1514_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_576_),
    .B(_596_),
    .C(_599_),
    .Y(_602_)
);

NAND2X1 _1515_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .B(_601_),
    .Y(_603_)
);

INVX1 _1516_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_603_),
    .Y(_604_)
);

NAND2X1 _1517_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_508_),
    .Y(_605_)
);

OAI21X1 _1518_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_525_),
    .B(_555_),
    .C(_605_),
    .Y(_606_)
);

OAI21X1 _1519_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_525_),
    .B(_555_),
    .C(_511_),
    .Y(_607_)
);

AOI22X1 _1520_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_607_),
    .C(_454_),
    .D(_442_),
    .Y(_608_)
);

OAI21X1 _1521_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_453_),
    .B(_359_),
    .C(_608_),
    .Y(_609_)
);

NAND3X1 _1522_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_604_),
    .B(_606_),
    .C(_609_),
    .Y(_610_)
);

OAI21X1 _1523_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_351_),
    .B(_448_),
    .C(_447_),
    .Y(_611_)
);

NOR2X1 _1524_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_560_),
    .B(_512_),
    .Y(_612_)
);

AOI22X1 _1525_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_556_),
    .B(_607_),
    .C(_612_),
    .D(_611_),
    .Y(_613_)
);

NAND3X1 _1526_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_283_),
    .B(_612_),
    .C(_563_),
    .Y(_614_)
);

NAND3X1 _1527_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_603_),
    .B(_614_),
    .C(_613_),
    .Y(_615_)
);

NAND2X1 _1528_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_615_),
    .B(_610_),
    .Y(_616_)
);

INVX1 _1529_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_276_),
    .Y(_617_)
);

OAI21X1 _1530_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_275_),
    .B(_252_),
    .C(_274_),
    .Y(_618_)
);

NAND3X1 _1531_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MulL_i),
    .B(_618_),
    .C(_617_),
    .Y(_619_)
);

NOR2X1 _1532_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .B(ACC[4]),
    .Y(_620_)
);

OAI21X1 _1533_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_364_),
    .C(_365_),
    .Y(_621_)
);

OAI21X1 _1534_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_620_),
    .B(_621_),
    .C(_619_),
    .Y(_622_)
);

NAND2X1 _1535_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_622_),
    .Y(_623_)
);

OAI21X1 _1536_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_616_),
    .C(_623_),
    .Y(_0_[4])
);

NAND2X1 _1537_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_255_),
    .B(_279_),
    .Y(_624_)
);

OAI21X1 _1538_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_617_),
    .B(_624_),
    .C(MulL_i),
    .Y(_625_)
);

AOI21X1 _1539_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_617_),
    .B(_624_),
    .C(_625_),
    .Y(_626_)
);

NOR2X1 _1540_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(Flag_i),
    .B(MulL_i),
    .Y(_627_)
);

AND2X2 _1541_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_627_),
    .B(ACC[5]),
    .Y(_628_)
);

OAI21X1 _1542_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_628_),
    .B(_626_),
    .C(_712_),
    .Y(_629_)
);

AOI21X1 _1543_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_579_),
    .B(_598_),
    .C(_594_),
    .Y(_630_)
);

INVX1 _1544_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_581_),
    .Y(_631_)
);

NOR2X1 _1545_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_135_),
    .B(_540_),
    .Y(_632_)
);

AOI21X1 _1546_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_631_),
    .B(_583_),
    .C(_632_),
    .Y(_633_)
);

NAND2X1 _1547_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_289_),
    .Y(_634_)
);

OAI22X1 _1548_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_288_),
    .B(_158_),
    .C(_417_),
    .D(_135_),
    .Y(_635_)
);

OAI21X1 _1549_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_582_),
    .B(_634_),
    .C(_635_),
    .Y(_636_)
);

OR2X2 _1550_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_592_),
    .B(_636_),
    .Y(_637_)
);

OAI21X1 _1551_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_590_),
    .B(_587_),
    .C(_636_),
    .Y(_638_)
);

NAND2X1 _1552_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_638_),
    .B(_637_),
    .Y(_639_)
);

NAND2X1 _1553_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_633_),
    .B(_639_),
    .Y(_640_)
);

INVX1 _1554_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_633_),
    .Y(_641_)
);

NAND3X1 _1555_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_641_),
    .B(_638_),
    .C(_637_),
    .Y(_642_)
);

NAND2X1 _1556_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_642_),
    .B(_640_),
    .Y(_643_)
);

NAND2X1 _1557_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_630_),
    .B(_643_),
    .Y(_644_)
);

OR2X2 _1558_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_643_),
    .B(_630_),
    .Y(_645_)
);

NAND2X1 _1559_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_644_),
    .B(_645_),
    .Y(_646_)
);

NAND3X1 _1560_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .B(_646_),
    .C(_610_),
    .Y(_647_)
);

INVX1 _1561_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .Y(_648_)
);

AOI21X1 _1562_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_614_),
    .C(_603_),
    .Y(_649_)
);

AND2X2 _1563_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_645_),
    .B(_644_),
    .Y(_650_)
);

OAI21X1 _1564_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_648_),
    .B(_649_),
    .C(_650_),
    .Y(_651_)
);

NAND3X1 _1565_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MulH_i),
    .B(_647_),
    .C(_651_),
    .Y(_652_)
);

NAND2X1 _1566_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_629_),
    .B(_652_),
    .Y(_0_[5])
);

NAND2X1 _1567_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_255_),
    .B(_356_),
    .Y(_653_)
);

AOI21X1 _1568_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_653_),
    .B(_357_),
    .C(_281_),
    .Y(_654_)
);

OAI21X1 _1569_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_280_),
    .B(_356_),
    .C(MulL_i),
    .Y(_655_)
);

NAND2X1 _1570_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ACC[6]),
    .B(_627_),
    .Y(_656_)
);

OAI21X1 _1571_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_655_),
    .B(_654_),
    .C(_656_),
    .Y(_657_)
);

NAND2X1 _1572_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_657_),
    .Y(_658_)
);

NAND3X1 _1573_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_601_),
    .B(_602_),
    .C(_650_),
    .Y(_659_)
);

AOI21X1 _1574_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_613_),
    .B(_614_),
    .C(_659_),
    .Y(_660_)
);

OAI21X1 _1575_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_602_),
    .B(_646_),
    .C(_645_),
    .Y(_661_)
);

OAI21X1 _1576_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_592_),
    .B(_636_),
    .C(_642_),
    .Y(_662_)
);

AOI21X1 _1577_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_405_),
    .B(_134_),
    .C(_634_),
    .Y(_663_)
);

OR2X2 _1578_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_662_),
    .B(_663_),
    .Y(_664_)
);

NAND2X1 _1579_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_663_),
    .B(_662_),
    .Y(_665_)
);

NAND2X1 _1580_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_665_),
    .B(_664_),
    .Y(_666_)
);

INVX1 _1581_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_666_),
    .Y(_667_)
);

OAI21X1 _1582_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_661_),
    .B(_660_),
    .C(_667_),
    .Y(_668_)
);

NOR2X1 _1583_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_646_),
    .B(_603_),
    .Y(_669_)
);

NAND3X1 _1584_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_606_),
    .B(_669_),
    .C(_609_),
    .Y(_670_)
);

INVX1 _1585_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_661_),
    .Y(_671_)
);

NAND3X1 _1586_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_671_),
    .B(_666_),
    .C(_670_),
    .Y(_672_)
);

NAND3X1 _1587_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MulH_i),
    .B(_672_),
    .C(_668_),
    .Y(_673_)
);

NAND2X1 _1588_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_658_),
    .B(_673_),
    .Y(_0_[6])
);

OAI21X1 _1589_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_582_),
    .B(_634_),
    .C(_665_),
    .Y(_674_)
);

NOR2X1 _1590_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_712_),
    .B(_674_),
    .Y(_675_)
);

NOR2X1 _1591_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_219_),
    .B(_354_),
    .Y(_676_)
);

AOI21X1 _1592_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_676_),
    .B(_358_),
    .C(_365_),
    .Y(_677_)
);

OAI21X1 _1593_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_676_),
    .B(_358_),
    .C(_677_),
    .Y(_678_)
);

AOI21X1 _1594_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_627_),
    .B(AN),
    .C(MulH_i),
    .Y(_679_)
);

AOI22X1 _1595_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_678_),
    .B(_679_),
    .C(_668_),
    .D(_675_),
    .Y(_0_[7])
);

INVX4 _1596_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(reset),
    .Y(_1_)
);

INVX1 _1597_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .Y(_680_)
);

NAND2X1 _1598_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[0]),
    .B(LoadCmd_i),
    .Y(_681_)
);

OAI21X1 _1599_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_680_),
    .C(_681_),
    .Y(_2_)
);

INVX1 _1600_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .Y(_682_)
);

NAND2X1 _1601_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[1]),
    .Y(_683_)
);

OAI21X1 _1602_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_682_),
    .C(_683_),
    .Y(_3_)
);

INVX1 _1603_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .Y(_684_)
);

NAND2X1 _1604_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[2]),
    .Y(_685_)
);

OAI21X1 _1605_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_684_),
    .C(_685_),
    .Y(_4_)
);

INVX1 _1606_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .Y(_686_)
);

NAND2X1 _1607_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[3]),
    .Y(_687_)
);

OAI21X1 _1608_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_686_),
    .C(_687_),
    .Y(_5_)
);

INVX1 _1609_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CI),
    .Y(_688_)
);

NAND2X1 _1610_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[4]),
    .Y(_689_)
);

OAI21X1 _1611_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_688_),
    .C(_689_),
    .Y(_6_)
);

INVX1 _1612_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .Y(_690_)
);

NAND2X1 _1613_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[5]),
    .Y(_691_)
);

OAI21X1 _1614_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_690_),
    .C(_691_),
    .Y(_7_)
);

INVX1 _1615_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BCD),
    .Y(_692_)
);

NAND2X1 _1616_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[6]),
    .Y(_693_)
);

OAI21X1 _1617_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_692_),
    .C(_693_),
    .Y(_8_)
);

NAND2X1 _1618_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(ABCmd_i[7]),
    .Y(_694_)
);

OAI21X1 _1619_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadCmd_i),
    .B(_715_),
    .C(_694_),
    .Y(_9_)
);

NAND2X1 _1620_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[0]),
    .B(LoadA_i),
    .Y(_695_)
);

OAI21X1 _1621_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_43_),
    .C(_695_),
    .Y(_10_)
);

NAND2X1 _1622_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[1]),
    .B(LoadA_i),
    .Y(_696_)
);

OAI21X1 _1623_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_716_),
    .C(_696_),
    .Y(_11_)
);

NAND2X1 _1624_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[2]),
    .B(LoadA_i),
    .Y(_697_)
);

OAI21X1 _1625_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_725_),
    .C(_697_),
    .Y(_12_)
);

NAND2X1 _1626_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[3]),
    .B(LoadA_i),
    .Y(_698_)
);

OAI21X1 _1627_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_387_),
    .C(_698_),
    .Y(_13_)
);

NAND2X1 _1628_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[4]),
    .B(LoadA_i),
    .Y(_699_)
);

OAI21X1 _1629_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_463_),
    .C(_699_),
    .Y(_14_)
);

NAND2X1 _1630_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[5]),
    .B(LoadA_i),
    .Y(_700_)
);

OAI21X1 _1631_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_401_),
    .C(_700_),
    .Y(_15_)
);

NAND2X1 _1632_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[6]),
    .B(LoadA_i),
    .Y(_701_)
);

OAI21X1 _1633_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_480_),
    .C(_701_),
    .Y(_16_)
);

NAND2X1 _1634_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[7]),
    .B(LoadA_i),
    .Y(_702_)
);

OAI21X1 _1635_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadA_i),
    .B(_417_),
    .C(_702_),
    .Y(_17_)
);

NAND2X1 _1636_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[0]),
    .B(LoadB_i),
    .Y(_703_)
);

OAI21X1 _1637_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_53_),
    .C(_703_),
    .Y(_18_)
);

NAND2X1 _1638_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[1]),
    .B(LoadB_i),
    .Y(_704_)
);

OAI21X1 _1639_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_36_),
    .C(_704_),
    .Y(_19_)
);

NAND2X1 _1640_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[2]),
    .B(LoadB_i),
    .Y(_705_)
);

OAI21X1 _1641_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_268_),
    .C(_705_),
    .Y(_20_)
);

NAND2X1 _1642_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[3]),
    .B(LoadB_i),
    .Y(_706_)
);

OAI21X1 _1643_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_309_),
    .C(_706_),
    .Y(_21_)
);

NAND2X1 _1644_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[4]),
    .B(LoadB_i),
    .Y(_707_)
);

OAI21X1 _1645_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_169_),
    .C(_707_),
    .Y(_22_)
);

INVX1 _1646_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[5]),
    .Y(_708_)
);

NAND2X1 _1647_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[5]),
    .B(LoadB_i),
    .Y(_709_)
);

OAI21X1 _1648_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_708_),
    .C(_709_),
    .Y(_23_)
);

NAND2X1 _1649_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[6]),
    .B(LoadB_i),
    .Y(_710_)
);

OAI21X1 _1650_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_133_),
    .C(_710_),
    .Y(_24_)
);

NAND2X1 _1651_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ABCmd_i[7]),
    .B(LoadB_i),
    .Y(_711_)
);

OAI21X1 _1652_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(LoadB_i),
    .B(_288_),
    .C(_711_),
    .Y(_25_)
);

DFFPOSX1 _1653_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_2_),
    .Q(alu_op[0])
);

DFFPOSX1 _1654_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_3_),
    .Q(alu_op[1])
);

DFFPOSX1 _1655_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_4_),
    .Q(alu_op[2])
);

DFFPOSX1 _1656_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_5_),
    .Q(alu_op[3])
);

DFFPOSX1 _1657_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_6_),
    .Q(CI)
);

DFFPOSX1 _1658_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_7_),
    .Q(shr)
);

DFFPOSX1 _1659_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_8_),
    .Q(BCD)
);

DFFPOSX1 _1660_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_9_),
    .Q(MUL)
);

DFFSR _1661_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_0_[0]),
    .Q(_919_[0]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1662_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_0_[1]),
    .Q(_919_[1]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1663_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_0_[2]),
    .Q(_919_[2]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1664_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_0_[3]),
    .Q(_919_[3]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1665_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_0_[4]),
    .Q(_919_[4]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1666_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_0_[5]),
    .Q(_919_[5]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1667_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_0_[6]),
    .Q(_919_[6]),
    .R(_1_),
    .S(vdd)
);

DFFSR _1668_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_0_[7]),
    .Q(_919_[7]),
    .R(_1_),
    .S(vdd)
);

DFFPOSX1 _1669_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_10_),
    .Q(AI[0])
);

DFFPOSX1 _1670_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_11_),
    .Q(AI[1])
);

DFFPOSX1 _1671_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_12_),
    .Q(AI[2])
);

DFFPOSX1 _1672_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_13_),
    .Q(AI[3])
);

DFFPOSX1 _1673_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_14_),
    .Q(AI[4])
);

DFFPOSX1 _1674_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_15_),
    .Q(AI[5])
);

DFFPOSX1 _1675_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_16_),
    .Q(AI[6])
);

DFFPOSX1 _1676_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_17_),
    .Q(\u_ALU8.AI7 )
);

DFFPOSX1 _1677_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_18_),
    .Q(BI[0])
);

DFFPOSX1 _1678_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_19_),
    .Q(BI[1])
);

DFFPOSX1 _1679_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_20_),
    .Q(BI[2])
);

DFFPOSX1 _1680_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf2),
    .D(_21_),
    .Q(BI[3])
);

DFFPOSX1 _1681_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf1),
    .D(_22_),
    .Q(BI[4])
);

DFFPOSX1 _1682_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf0),
    .D(_23_),
    .Q(BI[5])
);

DFFPOSX1 _1683_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf4),
    .D(_24_),
    .Q(BI[6])
);

DFFPOSX1 _1684_ (
    .vdd(vdd),
    .gnd(gnd),
    .CLK(clk_bF$buf3),
    .D(_25_),
    .Q(BI[7])
);

INVX1 _1685_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .Y(_857_)
);

INVX4 _1686_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[3]),
    .Y(_858_)
);

OAI21X1 _1687_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_857_),
    .B(_858_),
    .C(CI),
    .Y(_859_)
);

NOR2X1 _1688_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(_859_),
    .Y(_860_)
);

INVX1 _1689_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_860_),
    .Y(_861_)
);

INVX2 _1690_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .Y(_862_)
);

NAND2X1 _1691_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_862_),
    .Y(_863_)
);

INVX2 _1692_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .Y(_864_)
);

NAND2X1 _1693_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_864_),
    .Y(_865_)
);

NAND2X1 _1694_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[0]),
    .B(alu_op[1]),
    .Y(_866_)
);

AOI22X1 _1695_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(_866_),
    .C(_863_),
    .D(_865_),
    .Y(_867_)
);

INVX2 _1696_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .Y(_868_)
);

INVX1 _1697_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .Y(_869_)
);

INVX1 _1698_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[0]),
    .Y(_870_)
);

OAI21X1 _1699_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_869_),
    .C(_870_),
    .Y(_871_)
);

NAND2X1 _1700_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_868_),
    .B(_871_),
    .Y(_872_)
);

NAND2X1 _1701_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(shr),
    .Y(_873_)
);

OAI21X1 _1702_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_867_),
    .B(_872_),
    .C(_873_),
    .Y(_874_)
);

OAI21X1 _1703_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(alu_op_2_bF$buf1),
    .C(_858_),
    .Y(_875_)
);

AOI21X1 _1704_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .B(alu_op_2_bF$buf0),
    .C(_875_),
    .Y(_876_)
);

NOR2X1 _1705_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .B(_858_),
    .Y(_877_)
);

OAI21X1 _1706_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_876_),
    .C(_874_),
    .Y(_878_)
);

OAI21X1 _1707_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_874_),
    .B(_876_),
    .C(_878_),
    .Y(_879_)
);

OR2X2 _1708_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_879_),
    .B(_861_),
    .Y(_880_)
);

OAI21X1 _1709_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(_859_),
    .C(_879_),
    .Y(_881_)
);

NAND2X1 _1710_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_881_),
    .B(_880_),
    .Y(_882_)
);

INVX1 _1711_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_882_),
    .Y(ACC[0])
);

NOR2X1 _1712_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_876_),
    .B(_874_),
    .Y(_883_)
);

OAI21X1 _1713_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_861_),
    .B(_883_),
    .C(_878_),
    .Y(_884_)
);

NAND2X1 _1714_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(AI[2]),
    .Y(_885_)
);

NAND3X1 _1715_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(BI[1]),
    .C(_864_),
    .Y(_886_)
);

AOI22X1 _1716_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[1]),
    .C(_886_),
    .D(_863_),
    .Y(_887_)
);

INVX1 _1717_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[1]),
    .Y(_888_)
);

NOR2X1 _1718_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_888_),
    .Y(_889_)
);

OAI21X1 _1719_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .B(_889_),
    .C(_868_),
    .Y(_890_)
);

OAI21X1 _1720_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_887_),
    .B(_890_),
    .C(_885_),
    .Y(_891_)
);

OAI21X1 _1721_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .B(BI[1]),
    .C(_858_),
    .Y(_892_)
);

AOI21X1 _1722_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf1),
    .B(BI[1]),
    .C(_892_),
    .Y(_893_)
);

INVX1 _1723_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .Y(_894_)
);

OAI21X1 _1724_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_894_),
    .Y(_895_)
);

MUX2X1 _1725_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_895_),
    .B(_894_),
    .S(_891_),
    .Y(_896_)
);

NAND2X1 _1726_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_896_),
    .B(_884_),
    .Y(_897_)
);

INVX1 _1727_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_876_),
    .Y(_898_)
);

OAI21X1 _1728_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .B(_858_),
    .C(_898_),
    .Y(_899_)
);

MUX2X1 _1729_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[1]),
    .B(_869_),
    .S(alu_op[0]),
    .Y(_900_)
);

OAI21X1 _1730_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_870_),
    .B(_862_),
    .C(BI[0]),
    .Y(_901_)
);

NAND2X1 _1731_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_901_),
    .B(_900_),
    .Y(_902_)
);

NAND3X1 _1732_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_868_),
    .B(_871_),
    .C(_902_),
    .Y(_903_)
);

NAND3X1 _1733_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_873_),
    .B(_898_),
    .C(_903_),
    .Y(_904_)
);

AOI22X1 _1734_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_874_),
    .B(_899_),
    .C(_904_),
    .D(_860_),
    .Y(_905_)
);

OAI21X1 _1735_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_893_),
    .C(_891_),
    .Y(_906_)
);

OAI21X1 _1736_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_891_),
    .B(_893_),
    .C(_906_),
    .Y(_907_)
);

NAND2X1 _1737_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_905_),
    .B(_907_),
    .Y(_908_)
);

NAND2X1 _1738_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_908_),
    .B(_897_),
    .Y(_909_)
);

INVX1 _1739_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_909_),
    .Y(ACC[1])
);

NOR2X1 _1740_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_893_),
    .B(_891_),
    .Y(_910_)
);

OAI21X1 _1741_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_910_),
    .B(_905_),
    .C(_906_),
    .Y(_911_)
);

NAND2X1 _1742_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(AI[3]),
    .Y(_912_)
);

INVX1 _1743_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[2]),
    .Y(_913_)
);

NOR2X1 _1744_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op[0]),
    .B(_913_),
    .Y(_914_)
);

NAND2X1 _1745_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .B(_914_),
    .Y(_915_)
);

AOI22X1 _1746_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[2]),
    .C(_915_),
    .D(_863_),
    .Y(_916_)
);

OAI21X1 _1747_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .B(_914_),
    .C(_868_),
    .Y(_917_)
);

OAI21X1 _1748_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_917_),
    .B(_916_),
    .C(_912_),
    .Y(_918_)
);

OAI21X1 _1749_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .B(BI[2]),
    .C(_858_),
    .Y(_726_)
);

AOI21X1 _1750_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf1),
    .B(BI[2]),
    .C(_726_),
    .Y(_727_)
);

INVX1 _1751_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_727_),
    .Y(_728_)
);

OAI21X1 _1752_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf0),
    .B(_858_),
    .C(_728_),
    .Y(_729_)
);

MUX2X1 _1753_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_729_),
    .B(_728_),
    .S(_918_),
    .Y(_730_)
);

NAND2X1 _1754_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_730_),
    .B(_911_),
    .Y(_731_)
);

OAI21X1 _1755_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_727_),
    .C(_918_),
    .Y(_732_)
);

OAI21X1 _1756_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_918_),
    .B(_727_),
    .C(_732_),
    .Y(_733_)
);

NAND3X1 _1757_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_906_),
    .B(_733_),
    .C(_897_),
    .Y(_734_)
);

NAND2X1 _1758_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_731_),
    .B(_734_),
    .Y(_735_)
);

INVX1 _1759_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_735_),
    .Y(ACC[2])
);

INVX1 _1760_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .Y(_736_)
);

AND2X2 _1761_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_911_),
    .B(_730_),
    .Y(_737_)
);

NAND2X1 _1762_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(AI[4]),
    .Y(_738_)
);

AND2X2 _1763_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(BI[3]),
    .Y(_739_)
);

NAND2X1 _1764_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[3]),
    .B(_739_),
    .Y(_740_)
);

AOI22X1 _1765_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[3]),
    .C(_740_),
    .D(_863_),
    .Y(_741_)
);

OAI21X1 _1766_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[3]),
    .B(_739_),
    .C(_868_),
    .Y(_742_)
);

OAI21X1 _1767_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_742_),
    .B(_741_),
    .C(_738_),
    .Y(_743_)
);

OAI21X1 _1768_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .B(BI[3]),
    .C(_858_),
    .Y(_744_)
);

AOI21X1 _1769_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .B(BI[3]),
    .C(_744_),
    .Y(_745_)
);

OAI21X1 _1770_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_745_),
    .C(_743_),
    .Y(_746_)
);

OAI21X1 _1771_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_743_),
    .B(_745_),
    .C(_746_),
    .Y(_747_)
);

INVX1 _1772_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_747_),
    .Y(_748_)
);

OAI21X1 _1773_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_736_),
    .B(_737_),
    .C(_748_),
    .Y(_749_)
);

NAND3X1 _1774_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_747_),
    .C(_731_),
    .Y(_750_)
);

NAND2X1 _1775_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_750_),
    .B(_749_),
    .Y(_751_)
);

INVX1 _1776_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .Y(ACC[3])
);

INVX1 _1777_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BCD),
    .Y(_752_)
);

AOI21X1 _1778_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_735_),
    .B(_909_),
    .C(_752_),
    .Y(_753_)
);

NAND3X1 _1779_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_749_),
    .B(_750_),
    .C(_753_),
    .Y(_754_)
);

NAND2X1 _1780_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_732_),
    .B(_731_),
    .Y(_755_)
);

INVX1 _1781_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_746_),
    .Y(_756_)
);

AOI21X1 _1782_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_755_),
    .B(_748_),
    .C(_756_),
    .Y(_757_)
);

NAND2X1 _1783_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(AI[5]),
    .Y(_758_)
);

AND2X2 _1784_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(BI[4]),
    .Y(_759_)
);

NAND2X1 _1785_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .B(_759_),
    .Y(_760_)
);

AOI22X1 _1786_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[4]),
    .C(_760_),
    .D(_863_),
    .Y(_761_)
);

OAI21X1 _1787_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[4]),
    .B(_759_),
    .C(_868_),
    .Y(_762_)
);

OAI21X1 _1788_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_762_),
    .B(_761_),
    .C(_758_),
    .Y(_763_)
);

OAI21X1 _1789_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf1),
    .B(BI[4]),
    .C(_858_),
    .Y(_764_)
);

AOI21X1 _1790_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf0),
    .B(BI[4]),
    .C(_764_),
    .Y(_765_)
);

OAI21X1 _1791_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_765_),
    .C(_763_),
    .Y(_766_)
);

OAI21X1 _1792_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_763_),
    .B(_765_),
    .C(_766_),
    .Y(_767_)
);

AOI21X1 _1793_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_754_),
    .B(_757_),
    .C(_767_),
    .Y(_768_)
);

NOR2X1 _1794_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_730_),
    .B(_911_),
    .Y(_769_)
);

OAI21X1 _1795_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_769_),
    .B(_737_),
    .C(_909_),
    .Y(_770_)
);

NAND2X1 _1796_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BCD),
    .B(_770_),
    .Y(_771_)
);

OAI21X1 _1797_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .B(_771_),
    .C(_757_),
    .Y(HC)
);

INVX1 _1798_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_767_),
    .Y(_772_)
);

NOR2X1 _1799_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_772_),
    .B(HC),
    .Y(_773_)
);

NOR2X1 _1800_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_768_),
    .B(_773_),
    .Y(ACC[4])
);

INVX1 _1801_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_766_),
    .Y(_774_)
);

NAND2X1 _1802_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(AI[6]),
    .Y(_775_)
);

AND2X2 _1803_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(BI[5]),
    .Y(_776_)
);

NAND2X1 _1804_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_776_),
    .Y(_777_)
);

AOI22X1 _1805_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[5]),
    .C(_777_),
    .D(_863_),
    .Y(_778_)
);

OAI21X1 _1806_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[5]),
    .B(_776_),
    .C(_868_),
    .Y(_779_)
);

OAI21X1 _1807_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_779_),
    .B(_778_),
    .C(_775_),
    .Y(_780_)
);

OAI21X1 _1808_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .B(BI[5]),
    .C(_858_),
    .Y(_781_)
);

AOI21X1 _1809_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .B(BI[5]),
    .C(_781_),
    .Y(_782_)
);

OAI21X1 _1810_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_782_),
    .C(_780_),
    .Y(_783_)
);

OAI21X1 _1811_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_780_),
    .B(_782_),
    .C(_783_),
    .Y(_784_)
);

INVX1 _1812_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_784_),
    .Y(_785_)
);

OAI21X1 _1813_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_774_),
    .B(_768_),
    .C(_785_),
    .Y(_786_)
);

AOI21X1 _1814_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(HC),
    .B(_772_),
    .C(_774_),
    .Y(_787_)
);

NAND2X1 _1815_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_784_),
    .B(_787_),
    .Y(_788_)
);

NAND2X1 _1816_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_786_),
    .B(_788_),
    .Y(_789_)
);

INVX1 _1817_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_789_),
    .Y(ACC[5])
);

OAI21X1 _1818_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_784_),
    .B(_787_),
    .C(_783_),
    .Y(_790_)
);

INVX1 _1819_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .Y(_791_)
);

AND2X2 _1820_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(BI[6]),
    .Y(_792_)
);

NAND2X1 _1821_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[6]),
    .B(_792_),
    .Y(_793_)
);

AOI22X1 _1822_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[6]),
    .C(_793_),
    .D(_863_),
    .Y(_794_)
);

OAI21X1 _1823_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[6]),
    .B(_792_),
    .C(_868_),
    .Y(_795_)
);

OAI22X1 _1824_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_868_),
    .B(_791_),
    .C(_795_),
    .D(_794_),
    .Y(_796_)
);

OAI21X1 _1825_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf1),
    .B(BI[6]),
    .C(_858_),
    .Y(_797_)
);

AOI21X1 _1826_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf0),
    .B(BI[6]),
    .C(_797_),
    .Y(_798_)
);

OAI21X1 _1827_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_798_),
    .C(_796_),
    .Y(_799_)
);

OAI21X1 _1828_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_796_),
    .B(_798_),
    .C(_799_),
    .Y(_800_)
);

INVX1 _1829_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_800_),
    .Y(_801_)
);

NAND2X1 _1830_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .B(_790_),
    .Y(_802_)
);

NAND3X1 _1831_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_783_),
    .B(_800_),
    .C(_786_),
    .Y(_803_)
);

NAND2X1 _1832_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_803_),
    .B(_802_),
    .Y(_804_)
);

INVX1 _1833_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_804_),
    .Y(ACC[6])
);

INVX1 _1834_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_799_),
    .Y(_805_)
);

AOI21X1 _1835_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_786_),
    .B(_783_),
    .C(_800_),
    .Y(_806_)
);

NAND2X1 _1836_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(shr),
    .B(CI),
    .Y(_807_)
);

AND2X2 _1837_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_864_),
    .B(BI[7]),
    .Y(_808_)
);

NAND2X1 _1838_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .Y(_809_)
);

AOI22X1 _1839_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_862_),
    .B(BI[7]),
    .C(_809_),
    .D(_863_),
    .Y(_810_)
);

OAI21X1 _1840_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_808_),
    .C(_868_),
    .Y(_811_)
);

OAI21X1 _1841_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_811_),
    .B(_810_),
    .C(_807_),
    .Y(_812_)
);

OAI21X1 _1842_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf3),
    .B(BI[7]),
    .C(_858_),
    .Y(_813_)
);

AOI21X1 _1843_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(alu_op_2_bF$buf2),
    .B(BI[7]),
    .C(_813_),
    .Y(_814_)
);

OAI21X1 _1844_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_814_),
    .C(_812_),
    .Y(_815_)
);

OAI21X1 _1845_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_812_),
    .B(_814_),
    .C(_815_),
    .Y(_816_)
);

INVX1 _1846_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_816_),
    .Y(_817_)
);

OAI21X1 _1847_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_805_),
    .B(_806_),
    .C(_817_),
    .Y(_818_)
);

NAND3X1 _1848_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_799_),
    .B(_816_),
    .C(_802_),
    .Y(_819_)
);

AND2X2 _1849_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_818_),
    .B(_819_),
    .Y(AN)
);

NOR2X1 _1850_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(ACC[0]),
    .B(_770_),
    .Y(_820_)
);

NAND2X1 _1851_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_751_),
    .B(_820_),
    .Y(_821_)
);

NOR2X1 _1852_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_821_),
    .B(ACC[4]),
    .Y(_822_)
);

NOR2X1 _1853_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_801_),
    .B(_790_),
    .Y(_823_)
);

OAI21X1 _1854_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_806_),
    .B(_823_),
    .C(_789_),
    .Y(_824_)
);

NOR2X1 _1855_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_824_),
    .B(AN),
    .Y(_825_)
);

AND2X2 _1856_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_825_),
    .B(_822_),
    .Y(AZ)
);

NAND2X1 _1857_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_819_),
    .B(_818_),
    .Y(_826_)
);

NAND2X1 _1858_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BCD),
    .B(_824_),
    .Y(_827_)
);

OAI21X1 _1859_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_799_),
    .B(_816_),
    .C(_815_),
    .Y(_828_)
);

INVX1 _1860_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_828_),
    .Y(_829_)
);

NOR2X1 _1861_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_816_),
    .B(_800_),
    .Y(_830_)
);

NAND2X1 _1862_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_830_),
    .B(_790_),
    .Y(_831_)
);

NOR2X1 _1863_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_870_),
    .B(_868_),
    .Y(_832_)
);

NAND3X1 _1864_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_829_),
    .B(_832_),
    .C(_831_),
    .Y(_833_)
);

INVX1 _1865_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_830_),
    .Y(_834_)
);

AOI21X1 _1866_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_786_),
    .B(_783_),
    .C(_834_),
    .Y(_835_)
);

INVX1 _1867_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_832_),
    .Y(_836_)
);

OAI21X1 _1868_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_828_),
    .B(_835_),
    .C(_836_),
    .Y(_837_)
);

AND2X2 _1869_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_837_),
    .B(_833_),
    .Y(_838_)
);

OAI21X1 _1870_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_826_),
    .B(_827_),
    .C(_838_),
    .Y(CO)
);

AOI21X1 _1871_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_804_),
    .B(_789_),
    .C(_752_),
    .Y(_839_)
);

NAND2X1 _1872_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_833_),
    .B(_837_),
    .Y(_840_)
);

AOI21X1 _1873_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AN),
    .B(_839_),
    .C(_840_),
    .Y(_841_)
);

AOI21X1 _1874_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_790_),
    .B(_801_),
    .C(_805_),
    .Y(_842_)
);

NOR2X1 _1875_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_816_),
    .B(_842_),
    .Y(_843_)
);

AND2X2 _1876_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_842_),
    .B(_816_),
    .Y(_844_)
);

INVX1 _1877_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_814_),
    .Y(_845_)
);

NAND2X1 _1878_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_877_),
    .B(_812_),
    .Y(_846_)
);

NAND2X1 _1879_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_845_),
    .B(_846_),
    .Y(_847_)
);

NAND2X1 _1880_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(\u_ALU8.AI7 ),
    .B(_847_),
    .Y(_848_)
);

OR2X2 _1881_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_847_),
    .B(\u_ALU8.AI7 ),
    .Y(_849_)
);

NAND2X1 _1882_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_848_),
    .B(_849_),
    .Y(_850_)
);

INVX1 _1883_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .Y(_851_)
);

OAI21X1 _1884_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_843_),
    .B(_844_),
    .C(_851_),
    .Y(_852_)
);

NAND3X1 _1885_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_850_),
    .B(_819_),
    .C(_818_),
    .Y(_853_)
);

NAND3X1 _1886_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_852_),
    .B(_853_),
    .C(_841_),
    .Y(_854_)
);

NAND2X1 _1887_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_853_),
    .B(_852_),
    .Y(_855_)
);

NAND2X1 _1888_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(CO),
    .B(_855_),
    .Y(_856_)
);

AND2X2 _1889_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_854_),
    .B(_856_),
    .Y(AV)
);

BUFX2 _1890_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[0]),
    .Y(ACC_o[0])
);

BUFX2 _1891_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[1]),
    .Y(ACC_o[1])
);

BUFX2 _1892_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[2]),
    .Y(ACC_o[2])
);

BUFX2 _1893_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[3]),
    .Y(ACC_o[3])
);

BUFX2 _1894_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[4]),
    .Y(ACC_o[4])
);

BUFX2 _1895_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[5]),
    .Y(ACC_o[5])
);

BUFX2 _1896_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[6]),
    .Y(ACC_o[6])
);

BUFX2 _1897_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_919_[7]),
    .Y(ACC_o[7])
);

INVX2 _920_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MulH_i),
    .Y(_712_)
);

AND2X2 _921_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(BI[4]),
    .Y(_713_)
);

NAND2X1 _922_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[0]),
    .B(_713_),
    .Y(_714_)
);

INVX1 _923_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .Y(_715_)
);

INVX2 _924_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[1]),
    .Y(_716_)
);

NOR2X1 _925_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_715_),
    .B(_716_),
    .Y(_717_)
);

NAND2X1 _926_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[3]),
    .B(_717_),
    .Y(_718_)
);

OR2X2 _927_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_718_),
    .B(_714_),
    .Y(_719_)
);

NAND3X1 _928_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[0]),
    .C(AI[3]),
    .Y(_720_)
);

NAND3X1 _929_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(BI[1]),
    .C(AI[2]),
    .Y(_721_)
);

NOR2X1 _930_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_720_),
    .B(_721_),
    .Y(_722_)
);

INVX1 _931_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_722_),
    .Y(_723_)
);

NAND3X1 _932_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[2]),
    .C(AI[1]),
    .Y(_724_)
);

INVX2 _933_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[2]),
    .Y(_725_)
);

NAND2X1 _934_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(BI[1]),
    .Y(_26_)
);

OAI21X1 _935_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_725_),
    .B(_26_),
    .C(_720_),
    .Y(_27_)
);

INVX1 _936_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_27_),
    .Y(_28_)
);

OAI21X1 _937_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_724_),
    .B(_28_),
    .C(_723_),
    .Y(_29_)
);

NAND3X1 _938_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(BI[2]),
    .C(AI[2]),
    .Y(_30_)
);

INVX1 _939_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_30_),
    .Y(_31_)
);

NAND3X1 _940_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(BI[0]),
    .C(AI[4]),
    .Y(_32_)
);

NAND3X1 _941_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[1]),
    .C(AI[3]),
    .Y(_33_)
);

NOR2X1 _942_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_32_),
    .B(_33_),
    .Y(_34_)
);

INVX1 _943_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_34_),
    .Y(_35_)
);

INVX1 _944_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[1]),
    .Y(_36_)
);

NAND2X1 _945_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(AI[3]),
    .Y(_37_)
);

OAI21X1 _946_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_36_),
    .B(_37_),
    .C(_32_),
    .Y(_38_)
);

NAND3X1 _947_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_31_),
    .B(_38_),
    .C(_35_),
    .Y(_39_)
);

INVX1 _948_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_38_),
    .Y(_40_)
);

OAI21X1 _949_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_34_),
    .B(_40_),
    .C(_30_),
    .Y(_41_)
);

NAND3X1 _950_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_41_),
    .B(_29_),
    .C(_39_),
    .Y(_42_)
);

INVX1 _951_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(AI[0]),
    .Y(_43_)
);

NAND2X1 _952_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[4]),
    .Y(_44_)
);

OAI21X1 _953_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_43_),
    .B(_44_),
    .C(_718_),
    .Y(_45_)
);

NAND2X1 _954_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_45_),
    .B(_719_),
    .Y(_46_)
);

AOI21X1 _955_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_39_),
    .B(_41_),
    .C(_29_),
    .Y(_47_)
);

OAI21X1 _956_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_46_),
    .B(_47_),
    .C(_42_),
    .Y(_48_)
);

OAI21X1 _957_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_30_),
    .B(_40_),
    .C(_35_),
    .Y(_49_)
);

NAND3X1 _958_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(BI[1]),
    .C(AI[4]),
    .Y(_50_)
);

NAND3X1 _959_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf1),
    .B(BI[0]),
    .C(AI[5]),
    .Y(_51_)
);

OR2X2 _960_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_50_),
    .B(_51_),
    .Y(_52_)
);

INVX1 _961_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[0]),
    .Y(_53_)
);

NAND2X1 _962_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf0),
    .B(AI[5]),
    .Y(_54_)
);

OAI21X1 _963_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_53_),
    .B(_54_),
    .C(_50_),
    .Y(_55_)
);

NAND3X1 _964_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf5),
    .B(BI[2]),
    .C(AI[3]),
    .Y(_56_)
);

INVX1 _965_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_56_),
    .Y(_57_)
);

NAND3X1 _966_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_55_),
    .B(_57_),
    .C(_52_),
    .Y(_58_)
);

NOR2X1 _967_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_50_),
    .B(_51_),
    .Y(_59_)
);

INVX1 _968_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_55_),
    .Y(_60_)
);

OAI21X1 _969_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_59_),
    .B(_60_),
    .C(_56_),
    .Y(_61_)
);

NAND3X1 _970_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_62_)
);

AOI21X1 _971_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_31_),
    .B(_38_),
    .C(_34_),
    .Y(_63_)
);

OAI21X1 _972_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_59_),
    .B(_60_),
    .C(_57_),
    .Y(_64_)
);

NAND3X1 _973_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_55_),
    .B(_56_),
    .C(_52_),
    .Y(_65_)
);

NAND3X1 _974_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_63_),
    .B(_65_),
    .C(_64_),
    .Y(_66_)
);

NAND2X1 _975_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf4),
    .B(AI[0]),
    .Y(_67_)
);

INVX2 _976_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_67_),
    .Y(_68_)
);

NAND2X1 _977_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(BI[5]),
    .B(_68_),
    .Y(_69_)
);

INVX1 _978_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_69_),
    .Y(_70_)
);

NAND3X1 _979_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf3),
    .B(BI[4]),
    .C(AI[1]),
    .Y(_71_)
);

NAND3X1 _980_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(MUL_bF$buf2),
    .B(BI[3]),
    .C(AI[2]),
    .Y(_72_)
);

NOR2X1 _981_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_71_),
    .B(_72_),
    .Y(_73_)
);

OAI21X1 _982_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_716_),
    .B(_44_),
    .C(_72_),
    .Y(_74_)
);

INVX1 _983_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .Y(_75_)
);

OAI21X1 _984_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_73_),
    .B(_75_),
    .C(_70_),
    .Y(_76_)
);

INVX1 _985_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_73_),
    .Y(_77_)
);

NAND3X1 _986_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_69_),
    .B(_74_),
    .C(_77_),
    .Y(_78_)
);

NAND2X1 _987_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_78_),
    .B(_76_),
    .Y(_79_)
);

NAND3X1 _988_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_66_),
    .B(_62_),
    .C(_79_),
    .Y(_80_)
);

AOI21X1 _989_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_64_),
    .B(_65_),
    .C(_63_),
    .Y(_81_)
);

AOI21X1 _990_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_58_),
    .B(_61_),
    .C(_49_),
    .Y(_82_)
);

NAND3X1 _991_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_74_),
    .B(_77_),
    .C(_70_),
    .Y(_83_)
);

OAI21X1 _992_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_73_),
    .B(_75_),
    .C(_69_),
    .Y(_84_)
);

NAND2X1 _993_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_84_),
    .B(_83_),
    .Y(_85_)
);

OAI21X1 _994_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_81_),
    .B(_82_),
    .C(_85_),
    .Y(_86_)
);

NAND3X1 _995_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_80_),
    .B(_86_),
    .C(_48_),
    .Y(_87_)
);

AOI21X1 _996_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_86_),
    .B(_80_),
    .C(_48_),
    .Y(_88_)
);

OAI21X1 _997_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_719_),
    .B(_88_),
    .C(_87_),
    .Y(_89_)
);

OAI21X1 _998_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_85_),
    .B(_82_),
    .C(_62_),
    .Y(_90_)
);

AOI21X1 _999_ (
    .vdd(vdd),
    .gnd(gnd),
    .A(_55_),
    .B(_57_),
    .C(_59_),
    .Y(_91_)
);

endmodule
