magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -140 -140 2539 912
<< nwell >>
rect -20 -20 2419 352
<< psubstratepdiff >>
rect 0 756 2400 792
rect 0 496 40 756
rect 2360 496 2400 756
rect 0 460 2400 496
<< nsubstratendiff >>
rect 0 296 2400 332
rect 0 36 40 296
rect 2360 36 2400 296
rect 0 0 2400 36
<< metal1 >>
rect 0 756 2400 792
rect 0 496 40 756
rect 2360 496 2400 756
rect 0 460 2400 496
rect 0 296 2400 332
rect 0 36 40 296
rect 2360 36 2400 296
rect 0 0 2400 36
<< metal2 >>
rect 0 460 40 792
rect 2360 460 2400 792
rect 0 0 40 332
rect 2360 0 2400 332
<< metal3 >>
rect 0 460 40 792
rect 2360 460 2400 792
rect 0 0 40 332
rect 2360 0 2400 332
use CONT  CONT_0
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 508
box -6 -6 6 6
use CONT  CONT_1
array 0 95 24 0 0 0
timestamp 1537935238
transform 1 0 56 0 1 314
box -6 -6 6 6
use CONT  CONT_2
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 48
box -6 -6 6 6
use CONT  CONT_3
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 48
box -6 -6 6 6
use CONT  CONT_4
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 508
box -6 -6 6 6
use CONT  CONT_5
array 0 95 24 0 0 0
timestamp 1537935238
transform 1 0 56 0 1 18
box -6 -6 6 6
use CONT  CONT_6
array 0 95 24 0 0 0
timestamp 1537935238
transform 1 0 56 0 1 478
box -6 -6 6 6
use CONT  CONT_7
array 0 95 24 0 0 0
timestamp 1537935238
transform 1 0 56 0 1 774
box -6 -6 6 6
use VIA1  VIA1_0
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 20
box -8 -8 8 8
use VIA1  VIA1_1
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 20
box -8 -8 8 8
use VIA1  VIA1_2
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 480
box -8 -8 8 8
use VIA1  VIA1_3
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 480
box -8 -8 8 8
use VIA2  VIA2_0
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 48
box -8 -8 8 8
use VIA2  VIA2_1
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 48
box -8 -8 8 8
use VIA2  VIA2_2
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 2380 0 1 508
box -8 -8 8 8
use VIA2  VIA2_3
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 20 0 1 508
box -8 -8 8 8
<< end >>
