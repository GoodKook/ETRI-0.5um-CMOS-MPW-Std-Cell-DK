magic
tech scmos
magscale 1 2
timestamp 1739349528
<< metal1 >>
rect 100 451 148 475
rect 192 474 193 475
rect 160 473 176 474
rect 178 473 181 474
rect 160 470 177 473
rect 171 469 175 470
rect 168 467 171 469
rect 172 467 175 469
rect 162 466 165 467
rect 161 465 166 466
rect 161 464 167 465
rect 160 463 167 464
rect 168 464 175 467
rect 168 463 172 464
rect 160 462 163 463
rect 164 462 172 463
rect 159 458 162 462
rect 165 460 172 462
rect 165 459 175 460
rect 178 459 182 473
rect 189 472 193 474
rect 189 471 191 472
rect 192 471 193 472
rect 194 473 195 474
rect 194 471 196 473
rect 189 469 195 471
rect 191 468 194 469
rect 189 467 191 468
rect 194 467 196 468
rect 187 465 195 467
rect 188 464 194 465
rect 189 462 195 463
rect 189 461 196 462
rect 194 460 195 461
rect 194 459 196 460
rect 165 458 182 459
rect 159 457 163 458
rect 164 457 182 458
rect 189 458 196 459
rect 189 457 195 458
rect 160 456 172 457
rect 160 455 167 456
rect 161 454 167 455
rect 162 453 166 454
rect 168 452 172 456
rect 176 455 182 457
rect 194 456 195 457
rect 189 455 191 456
rect 194 455 196 456
rect 187 454 196 455
rect 187 453 195 454
rect 189 452 191 453
rect 169 451 172 452
rect 186 449 188 451
rect 189 450 196 451
rect 189 449 195 450
rect 194 448 195 449
rect 189 447 191 448
rect 194 447 196 448
rect 187 446 196 447
rect 188 445 195 446
rect 189 444 191 445
rect 189 442 191 443
rect 192 442 195 444
rect 150 440 152 442
rect 189 441 196 442
rect 149 439 152 440
rect 148 438 152 439
rect 147 436 152 438
rect 146 435 152 436
rect 145 434 152 435
rect 106 433 126 434
rect 144 433 152 434
rect 105 432 126 433
rect 143 432 152 433
rect 104 431 126 432
rect 103 430 126 431
rect 142 430 152 432
rect 102 429 126 430
rect 141 429 152 430
rect 101 426 126 429
rect 140 428 152 429
rect 139 427 152 428
rect 100 412 126 426
rect 138 425 152 427
rect 137 424 152 425
rect 136 423 152 424
rect 135 422 152 423
rect 134 420 152 422
rect 133 419 152 420
rect 161 437 166 438
rect 161 436 169 437
rect 170 436 173 441
rect 189 440 193 441
rect 194 440 196 441
rect 190 439 192 440
rect 194 439 195 440
rect 190 438 191 439
rect 161 433 173 436
rect 161 419 164 433
rect 170 430 173 433
rect 189 437 196 438
rect 189 436 195 437
rect 189 434 191 436
rect 189 433 196 434
rect 189 432 195 433
rect 187 430 195 431
rect 170 426 182 430
rect 187 429 196 430
rect 187 428 195 429
rect 132 418 152 419
rect 162 418 163 419
rect 131 417 152 418
rect 130 416 152 417
rect 170 416 173 426
rect 189 423 196 424
rect 189 421 191 423
rect 192 422 195 423
rect 186 420 195 421
rect 186 419 196 420
rect 189 417 190 418
rect 194 417 195 418
rect 129 414 152 416
rect 189 415 191 417
rect 194 416 196 417
rect 193 415 195 416
rect 189 414 195 415
rect 128 413 151 414
rect 190 413 195 414
rect 127 412 150 413
rect 100 411 149 412
rect 189 411 191 413
rect 100 410 148 411
rect 60 400 73 401
rect 57 399 77 400
rect 55 398 79 399
rect 53 397 81 398
rect 51 396 83 397
rect 50 395 62 396
rect 72 395 84 396
rect 13 394 14 395
rect 49 394 57 395
rect 77 394 85 395
rect 12 393 16 394
rect 49 393 54 394
rect 80 393 85 394
rect 12 392 18 393
rect 49 392 52 393
rect 82 392 85 393
rect 13 391 20 392
rect 15 390 22 391
rect 18 389 24 390
rect 20 388 26 389
rect 66 388 72 389
rect 22 387 28 388
rect 54 387 59 388
rect 64 387 74 388
rect 13 386 28 387
rect 52 386 60 387
rect 63 386 75 387
rect 12 384 28 386
rect 51 385 61 386
rect 63 385 76 386
rect 50 384 76 385
rect 13 383 18 384
rect 50 383 77 384
rect 14 382 21 383
rect 49 382 55 383
rect 58 382 66 383
rect 72 382 77 383
rect 16 381 23 382
rect 18 380 25 381
rect 20 379 27 380
rect 22 378 28 379
rect 13 377 28 378
rect 49 377 54 382
rect 59 381 65 382
rect 60 378 64 381
rect 73 378 77 382
rect 59 377 65 378
rect 72 377 77 378
rect 12 375 28 377
rect 50 376 66 377
rect 71 376 77 377
rect 50 375 77 376
rect 100 376 111 410
rect 125 409 148 410
rect 189 410 196 411
rect 189 409 195 410
rect 125 408 147 409
rect 125 407 146 408
rect 189 407 195 408
rect 125 406 145 407
rect 189 406 196 407
rect 125 405 144 406
rect 125 403 143 405
rect 161 404 175 405
rect 178 404 181 405
rect 189 404 193 406
rect 194 405 195 406
rect 194 404 196 405
rect 125 402 142 403
rect 125 401 141 402
rect 125 400 140 401
rect 160 400 176 404
rect 125 398 139 400
rect 125 397 138 398
rect 162 397 166 400
rect 167 397 170 400
rect 125 396 137 397
rect 125 395 136 396
rect 162 395 170 397
rect 125 393 135 395
rect 162 394 171 395
rect 161 393 171 394
rect 125 392 134 393
rect 161 392 165 393
rect 167 392 172 393
rect 125 391 133 392
rect 161 391 164 392
rect 168 391 172 392
rect 125 390 132 391
rect 160 390 164 391
rect 125 389 131 390
rect 160 389 163 390
rect 125 387 130 389
rect 160 388 164 389
rect 169 388 172 391
rect 178 390 182 404
rect 189 403 191 404
rect 192 403 196 404
rect 192 402 195 403
rect 191 401 193 402
rect 189 399 193 401
rect 189 398 191 399
rect 192 398 193 399
rect 194 400 195 401
rect 194 398 196 400
rect 189 397 196 398
rect 189 396 195 397
rect 191 395 194 396
rect 189 394 190 395
rect 192 394 195 395
rect 189 393 191 394
rect 192 393 196 394
rect 189 391 193 393
rect 194 391 196 393
rect 191 390 192 391
rect 161 387 164 388
rect 168 387 172 388
rect 125 386 129 387
rect 161 386 165 387
rect 167 386 172 387
rect 174 386 182 390
rect 190 389 193 390
rect 189 388 193 389
rect 189 386 191 388
rect 192 386 193 388
rect 194 389 195 391
rect 194 386 196 389
rect 125 385 128 386
rect 161 385 171 386
rect 189 385 195 386
rect 126 384 127 385
rect 162 384 170 385
rect 190 384 195 385
rect 163 383 169 384
rect 192 383 193 384
rect 194 383 195 384
rect 187 382 191 383
rect 192 382 195 383
rect 187 381 195 382
rect 187 380 189 381
rect 190 380 193 381
rect 187 379 188 380
rect 190 379 192 380
rect 187 378 195 379
rect 187 377 196 378
rect 50 374 76 375
rect 51 373 61 374
rect 63 373 75 374
rect 14 372 19 373
rect 52 372 60 373
rect 64 372 74 373
rect 13 370 21 372
rect 54 371 58 372
rect 65 371 73 372
rect 13 369 16 370
rect 18 369 22 370
rect 12 365 15 369
rect 12 364 18 365
rect 19 364 22 369
rect 76 368 77 369
rect 74 367 77 368
rect 54 366 60 367
rect 73 366 77 367
rect 52 365 62 366
rect 71 365 77 366
rect 12 363 23 364
rect 51 363 63 365
rect 69 364 77 365
rect 68 363 77 364
rect 13 362 27 363
rect 16 361 28 362
rect 50 361 64 363
rect 67 362 77 363
rect 66 361 76 362
rect 21 360 28 361
rect 25 359 28 360
rect 49 360 56 361
rect 59 360 74 361
rect 13 358 14 359
rect 49 358 55 360
rect 60 359 73 360
rect 60 358 72 359
rect 12 357 20 358
rect 12 356 25 357
rect 12 355 28 356
rect 13 354 19 355
rect 20 354 28 355
rect 14 353 20 354
rect 25 353 28 354
rect 16 352 23 353
rect 18 351 25 352
rect 20 350 27 351
rect 49 350 54 358
rect 60 357 70 358
rect 60 356 69 357
rect 60 355 67 356
rect 60 352 66 355
rect 100 352 148 376
rect 189 372 190 373
rect 189 371 191 372
rect 192 371 195 373
rect 179 370 181 371
rect 189 370 196 371
rect 160 366 176 370
rect 170 363 171 364
rect 169 361 173 363
rect 168 360 172 361
rect 167 359 172 360
rect 166 358 171 359
rect 160 356 170 358
rect 160 355 169 356
rect 178 355 182 370
rect 189 369 193 370
rect 194 369 196 370
rect 190 368 192 369
rect 194 368 195 369
rect 189 366 196 367
rect 189 365 195 366
rect 189 364 191 365
rect 189 363 192 364
rect 194 363 195 364
rect 189 362 196 363
rect 189 361 192 362
rect 193 361 195 362
rect 192 360 193 361
rect 189 358 195 360
rect 189 356 191 358
rect 194 357 196 358
rect 194 356 195 357
rect 189 355 195 356
rect 160 354 170 355
rect 164 353 171 354
rect 174 353 182 355
rect 190 354 195 355
rect 167 352 172 353
rect 174 352 181 353
rect 60 351 65 352
rect 168 351 172 352
rect 186 351 188 353
rect 189 351 195 353
rect 60 350 66 351
rect 169 350 173 351
rect 22 349 28 350
rect 13 348 28 349
rect 12 347 28 348
rect 12 346 19 347
rect 12 345 22 346
rect 13 344 27 345
rect 49 344 77 350
rect 170 348 173 350
rect 189 350 190 351
rect 194 350 195 351
rect 189 349 191 350
rect 194 349 196 350
rect 171 347 172 348
rect 187 347 195 349
rect 189 346 191 347
rect 194 345 195 346
rect 189 344 196 345
rect 17 343 28 344
rect 22 342 28 343
rect 26 341 28 342
rect 189 343 195 344
rect 189 342 193 343
rect 194 342 196 343
rect 189 341 196 342
rect 19 334 23 335
rect 17 333 25 334
rect 49 333 77 339
rect 17 332 26 333
rect 16 331 27 332
rect 16 330 19 331
rect 24 330 28 331
rect 16 329 18 330
rect 25 329 28 330
rect 17 328 19 329
rect 26 328 28 329
rect 17 327 20 328
rect 25 327 28 328
rect 16 326 27 327
rect 16 325 28 326
rect 17 324 32 325
rect 22 323 32 324
rect 13 322 15 323
rect 26 322 32 323
rect 12 320 15 322
rect 17 321 20 322
rect 16 320 24 321
rect 13 319 15 320
rect 17 319 28 320
rect 18 318 28 319
rect 23 317 28 318
rect 49 316 54 329
rect 60 316 65 327
rect 19 315 20 316
rect 17 314 25 315
rect 16 312 28 314
rect 16 311 19 312
rect 23 311 28 312
rect 13 309 15 310
rect 17 309 19 311
rect 49 310 77 316
rect 100 314 111 341
rect 189 340 191 341
rect 192 340 195 341
rect 193 339 194 340
rect 172 337 173 338
rect 167 334 169 335
rect 160 320 163 334
rect 164 320 166 334
rect 167 327 170 334
rect 171 328 174 337
rect 189 336 191 339
rect 194 338 195 339
rect 194 337 196 338
rect 193 336 195 337
rect 189 335 195 336
rect 177 334 180 335
rect 190 334 194 335
rect 176 333 181 334
rect 187 333 188 334
rect 192 333 193 334
rect 194 333 195 334
rect 176 332 182 333
rect 175 331 182 332
rect 186 331 188 333
rect 189 332 196 333
rect 189 331 195 332
rect 175 328 178 331
rect 179 329 182 331
rect 189 329 196 330
rect 171 327 177 328
rect 167 323 177 327
rect 167 320 170 323
rect 160 316 170 320
rect 171 322 177 323
rect 12 308 20 309
rect 12 307 24 308
rect 13 306 28 307
rect 18 305 28 306
rect 23 304 28 305
rect 49 305 51 306
rect 83 305 85 306
rect 49 304 54 305
rect 80 304 85 305
rect 49 303 56 304
rect 78 303 85 304
rect 15 302 17 303
rect 49 302 60 303
rect 73 302 84 303
rect 14 301 18 302
rect 13 300 18 301
rect 23 301 25 302
rect 51 301 83 302
rect 23 300 26 301
rect 52 300 81 301
rect 12 299 16 300
rect 23 299 27 300
rect 54 299 80 300
rect 12 296 15 299
rect 24 298 28 299
rect 56 298 77 299
rect 12 295 16 296
rect 13 294 16 295
rect 25 294 28 298
rect 59 297 74 298
rect 65 296 68 297
rect 13 293 18 294
rect 24 293 28 294
rect 14 292 28 293
rect 15 291 27 292
rect 16 290 26 291
rect 100 290 148 314
rect 171 313 174 322
rect 175 321 177 322
rect 180 322 183 329
rect 189 328 195 329
rect 189 327 191 328
rect 189 326 192 327
rect 194 326 195 327
rect 189 325 196 326
rect 189 324 195 325
rect 189 322 195 323
rect 180 321 182 322
rect 189 321 196 322
rect 175 320 178 321
rect 179 320 182 321
rect 175 318 182 320
rect 194 319 195 321
rect 189 318 196 319
rect 175 317 181 318
rect 189 317 195 318
rect 176 316 181 317
rect 177 315 180 316
rect 190 315 195 316
rect 189 314 195 315
rect 172 312 173 313
rect 189 312 191 314
rect 189 311 196 312
rect 189 310 195 311
rect 189 309 191 310
rect 189 308 195 309
rect 189 307 196 308
rect 190 306 191 307
rect 194 306 195 307
rect 190 305 195 306
rect 189 304 196 305
rect 169 303 171 304
rect 189 303 195 304
rect 168 300 172 303
rect 189 302 191 303
rect 189 301 195 302
rect 189 300 196 301
rect 160 297 182 300
rect 189 298 191 300
rect 189 297 196 298
rect 161 296 181 297
rect 189 296 195 297
rect 192 295 193 296
rect 175 294 176 295
rect 190 294 195 295
rect 19 289 24 290
rect 65 282 68 283
rect 16 281 19 282
rect 61 281 69 282
rect 16 280 21 281
rect 60 280 69 281
rect 17 279 23 280
rect 59 279 69 280
rect 18 278 25 279
rect 58 278 69 279
rect 71 281 73 282
rect 71 280 75 281
rect 71 278 76 280
rect 20 277 27 278
rect 57 277 69 278
rect 70 277 77 278
rect 22 276 28 277
rect 57 276 63 277
rect 23 275 30 276
rect 57 275 61 276
rect 17 274 31 275
rect 16 273 32 274
rect 16 272 24 273
rect 29 272 32 273
rect 17 271 18 272
rect 30 270 32 272
rect 56 271 61 275
rect 57 270 62 271
rect 65 270 69 277
rect 71 276 77 277
rect 73 272 77 276
rect 72 270 77 272
rect 12 269 17 270
rect 57 269 77 270
rect 12 268 22 269
rect 12 267 27 268
rect 58 267 76 269
rect 12 266 28 267
rect 59 266 75 267
rect 13 265 19 266
rect 22 265 28 266
rect 60 265 74 266
rect 15 264 21 265
rect 27 264 28 265
rect 62 264 72 265
rect 17 263 24 264
rect 100 263 111 290
rect 162 289 165 294
rect 174 293 177 294
rect 189 293 195 294
rect 173 292 178 293
rect 173 291 177 292
rect 189 291 191 293
rect 194 291 196 293
rect 171 290 176 291
rect 189 290 195 291
rect 169 289 176 290
rect 190 289 195 290
rect 162 288 175 289
rect 191 288 192 289
rect 193 288 195 289
rect 162 286 173 288
rect 189 286 191 288
rect 194 286 196 288
rect 162 285 175 286
rect 162 280 165 285
rect 167 284 176 285
rect 189 284 195 286
rect 171 283 177 284
rect 191 283 194 284
rect 172 282 178 283
rect 190 282 193 283
rect 173 281 178 282
rect 174 280 178 281
rect 164 279 165 280
rect 175 279 178 280
rect 189 281 193 282
rect 189 280 191 281
rect 192 280 193 281
rect 189 279 193 280
rect 194 281 195 283
rect 194 279 196 281
rect 176 278 177 279
rect 189 278 195 279
rect 190 277 195 278
rect 186 274 195 276
rect 190 272 193 273
rect 189 271 193 272
rect 189 270 191 271
rect 192 270 193 271
rect 194 272 195 273
rect 194 270 196 272
rect 189 269 196 270
rect 189 268 195 269
rect 179 267 181 268
rect 160 263 176 267
rect 19 262 26 263
rect 21 261 28 262
rect 65 261 68 262
rect 13 260 28 261
rect 61 260 72 261
rect 164 260 168 263
rect 12 258 28 260
rect 60 259 74 260
rect 161 259 168 260
rect 170 260 171 261
rect 170 259 172 260
rect 59 258 75 259
rect 12 257 19 258
rect 58 257 76 258
rect 12 256 25 257
rect 57 256 77 257
rect 14 255 28 256
rect 57 255 64 256
rect 70 255 77 256
rect 19 254 28 255
rect 24 253 28 254
rect 56 254 62 255
rect 72 254 77 255
rect 56 252 61 254
rect 57 249 61 252
rect 73 250 77 254
rect 161 255 164 259
rect 169 258 173 259
rect 168 256 172 258
rect 166 255 171 256
rect 161 254 171 255
rect 161 252 170 254
rect 178 253 182 267
rect 187 266 188 268
rect 190 267 194 268
rect 187 265 195 266
rect 187 264 196 265
rect 187 263 189 264
rect 187 261 188 263
rect 186 257 195 258
rect 186 255 196 257
rect 161 251 171 252
rect 72 249 76 250
rect 58 248 62 249
rect 71 248 76 249
rect 59 247 65 248
rect 68 247 75 248
rect 15 245 19 246
rect 22 245 24 246
rect 14 244 20 245
rect 21 244 26 245
rect 13 243 27 244
rect 13 240 16 243
rect 18 242 27 243
rect 57 242 85 247
rect 18 241 22 242
rect 19 240 21 241
rect 13 239 18 240
rect 25 239 28 242
rect 14 238 18 239
rect 24 238 28 239
rect 81 239 84 240
rect 15 237 18 238
rect 23 236 27 238
rect 23 235 25 236
rect 21 228 24 234
rect 13 226 17 227
rect 22 226 24 227
rect 13 225 21 226
rect 22 225 25 226
rect 13 224 26 225
rect 14 223 28 224
rect 15 222 19 223
rect 21 222 28 223
rect 16 221 20 222
rect 18 220 21 221
rect 22 220 25 222
rect 26 221 28 222
rect 19 219 25 220
rect 20 218 25 219
rect 21 217 25 218
rect 22 216 25 217
rect 57 218 59 219
rect 81 218 85 239
rect 57 216 62 218
rect 81 217 84 218
rect 16 215 18 216
rect 14 214 20 215
rect 56 214 62 216
rect 13 213 21 214
rect 13 212 22 213
rect 13 210 16 212
rect 19 211 23 212
rect 20 210 24 211
rect 25 210 28 214
rect 57 213 62 214
rect 57 212 63 213
rect 58 211 65 212
rect 13 209 17 210
rect 21 209 28 210
rect 13 208 18 209
rect 22 208 28 209
rect 14 207 18 208
rect 23 207 28 208
rect 16 206 18 207
rect 24 206 28 207
rect 57 206 77 211
rect 25 205 28 206
rect 16 203 21 204
rect 14 202 24 203
rect 13 201 26 202
rect 13 198 16 201
rect 19 200 27 201
rect 23 199 27 200
rect 13 197 17 198
rect 14 196 20 197
rect 25 196 28 199
rect 15 195 28 196
rect 49 195 54 201
rect 57 195 77 201
rect 100 197 111 250
rect 119 199 129 250
rect 119 198 130 199
rect 138 198 148 250
rect 161 246 164 251
rect 166 250 172 251
rect 167 249 172 250
rect 174 250 182 253
rect 189 254 191 255
rect 194 254 196 255
rect 189 252 195 254
rect 191 251 194 252
rect 190 250 195 251
rect 174 249 181 250
rect 189 249 196 250
rect 168 248 173 249
rect 169 247 173 248
rect 170 246 173 247
rect 189 248 195 249
rect 189 247 191 248
rect 189 246 195 247
rect 170 245 172 246
rect 189 245 196 246
rect 190 243 195 244
rect 189 242 196 243
rect 189 241 195 242
rect 189 240 193 241
rect 194 240 196 241
rect 189 239 195 240
rect 189 238 191 239
rect 192 238 195 239
rect 169 234 171 235
rect 161 231 163 232
rect 168 231 172 234
rect 189 232 191 234
rect 192 233 195 234
rect 192 232 196 233
rect 160 227 172 231
rect 160 213 164 227
rect 168 223 172 227
rect 174 227 182 231
rect 189 230 193 232
rect 194 230 196 232
rect 190 229 192 230
rect 189 228 190 229
rect 194 228 195 230
rect 174 223 178 227
rect 189 226 191 228
rect 194 227 196 228
rect 193 226 195 227
rect 189 225 195 226
rect 190 224 194 225
rect 168 220 178 223
rect 186 221 188 223
rect 189 221 195 223
rect 161 212 163 213
rect 168 210 172 220
rect 174 213 178 220
rect 189 219 196 220
rect 189 218 195 219
rect 189 216 191 218
rect 189 215 196 216
rect 189 214 195 215
rect 175 212 177 213
rect 190 212 195 213
rect 189 211 195 212
rect 169 209 170 210
rect 189 209 191 211
rect 194 209 196 211
rect 189 208 195 209
rect 190 207 195 208
rect 189 206 194 207
rect 189 205 191 206
rect 189 204 195 205
rect 189 203 196 204
rect 189 202 195 203
rect 189 201 190 202
rect 194 201 195 202
rect 112 197 117 198
rect 118 197 136 198
rect 137 197 148 198
rect 166 197 169 200
rect 187 199 195 201
rect 188 198 194 199
rect 179 197 181 198
rect 189 197 190 198
rect 16 194 27 195
rect 19 193 26 194
rect 49 193 52 194
rect 15 191 19 192
rect 14 190 20 191
rect 25 190 27 191
rect 13 189 21 190
rect 13 186 16 189
rect 18 188 22 189
rect 19 187 23 188
rect 20 186 24 187
rect 25 186 28 190
rect 49 189 53 193
rect 57 189 61 193
rect 49 186 77 189
rect 13 185 18 186
rect 21 185 28 186
rect 14 184 18 185
rect 22 184 28 185
rect 50 184 77 186
rect 15 183 18 184
rect 23 183 28 184
rect 52 183 77 184
rect 16 182 17 183
rect 24 182 28 183
rect 26 181 28 182
rect 57 180 61 183
rect 100 180 148 197
rect 160 194 176 197
rect 163 191 165 192
rect 100 178 147 180
rect 160 179 162 188
rect 163 187 166 191
rect 169 190 172 191
rect 168 189 173 190
rect 167 187 174 189
rect 163 185 170 187
rect 171 185 174 187
rect 163 182 169 185
rect 172 182 174 185
rect 178 184 182 197
rect 189 194 191 197
rect 194 195 196 197
rect 193 194 195 195
rect 189 193 195 194
rect 191 192 194 193
rect 191 191 193 192
rect 189 189 193 191
rect 189 188 191 189
rect 192 188 193 189
rect 194 190 195 192
rect 194 188 196 190
rect 189 187 195 188
rect 190 186 195 187
rect 176 183 182 184
rect 186 183 195 185
rect 163 181 170 182
rect 171 181 174 182
rect 100 177 146 178
rect 100 176 145 177
rect 163 176 166 181
rect 167 179 174 181
rect 175 180 182 183
rect 176 179 181 180
rect 187 179 188 182
rect 190 179 192 182
rect 194 181 196 182
rect 194 179 195 181
rect 167 178 173 179
rect 168 177 173 178
rect 187 178 195 179
rect 187 177 196 178
rect 170 176 171 177
rect 187 176 195 177
rect 100 175 144 176
rect 100 174 142 175
rect 174 167 178 168
rect 161 165 165 167
rect 175 166 179 167
rect 167 165 172 166
rect 176 165 179 166
rect 161 163 163 165
rect 167 164 173 165
rect 177 164 179 165
rect 168 163 171 164
rect 161 160 162 163
rect 169 160 171 163
rect 178 161 179 164
rect 177 160 179 161
rect 161 155 179 160
rect 161 153 162 155
rect 178 153 179 155
rect 174 150 177 151
rect 40 149 46 150
rect 162 149 165 150
rect 174 149 179 150
rect 35 148 50 149
rect 32 147 50 148
rect 161 148 166 149
rect 176 148 179 149
rect 30 146 49 147
rect 161 146 163 148
rect 167 147 173 148
rect 177 147 179 148
rect 168 146 172 147
rect 29 145 47 146
rect 28 144 46 145
rect 27 143 44 144
rect 161 143 162 146
rect 169 143 171 146
rect 178 143 179 147
rect 26 142 43 143
rect 54 142 64 143
rect 161 142 163 143
rect 168 142 171 143
rect 177 142 179 143
rect 21 141 22 142
rect 26 141 42 142
rect 51 141 69 142
rect 18 140 22 141
rect 25 140 41 141
rect 49 140 71 141
rect 17 139 21 140
rect 16 138 21 139
rect 25 138 40 140
rect 48 139 73 140
rect 47 138 74 139
rect 161 138 179 142
rect 15 137 20 138
rect 14 136 20 137
rect 24 137 39 138
rect 46 137 75 138
rect 24 136 38 137
rect 45 136 71 137
rect 161 136 162 138
rect 178 136 179 138
rect 13 135 19 136
rect 12 134 19 135
rect 11 133 19 134
rect 23 134 37 136
rect 45 135 68 136
rect 187 135 188 136
rect 44 134 65 135
rect 187 134 190 135
rect 23 133 36 134
rect 43 133 63 134
rect 189 133 195 134
rect 11 132 18 133
rect 10 131 18 132
rect 9 130 18 131
rect 22 131 35 133
rect 42 132 61 133
rect 81 132 82 133
rect 83 132 92 133
rect 41 131 60 132
rect 79 131 97 132
rect 161 131 162 133
rect 178 132 179 133
rect 190 132 195 133
rect 177 131 179 132
rect 22 130 34 131
rect 41 130 58 131
rect 80 130 100 131
rect 8 128 17 130
rect 7 126 17 128
rect 21 129 34 130
rect 40 129 57 130
rect 81 129 102 130
rect 21 127 33 129
rect 39 128 56 129
rect 82 128 104 129
rect 39 127 55 128
rect 83 127 106 128
rect 161 127 179 131
rect 187 131 196 132
rect 187 130 190 131
rect 187 129 188 130
rect 20 126 33 127
rect 38 126 54 127
rect 66 126 71 127
rect 84 126 108 127
rect 161 126 163 127
rect 168 126 171 127
rect 177 126 179 127
rect 6 124 16 126
rect 20 124 32 126
rect 38 125 53 126
rect 64 125 74 126
rect 85 125 109 126
rect 5 121 16 124
rect 4 118 16 121
rect 19 123 32 124
rect 37 124 53 125
rect 62 124 75 125
rect 86 124 110 125
rect 161 124 162 126
rect 19 120 31 123
rect 37 121 52 124
rect 60 123 77 124
rect 86 123 112 124
rect 59 122 78 123
rect 87 122 113 123
rect 58 121 79 122
rect 88 121 114 122
rect 18 119 31 120
rect 36 119 51 121
rect 57 120 80 121
rect 88 120 115 121
rect 161 120 162 122
rect 168 120 170 126
rect 178 124 179 126
rect 186 124 189 125
rect 187 122 188 124
rect 189 122 193 123
rect 194 122 195 123
rect 178 120 179 122
rect 187 121 195 122
rect 187 120 196 121
rect 57 119 81 120
rect 89 119 116 120
rect 161 119 164 120
rect 168 119 171 120
rect 177 119 179 120
rect 4 113 15 118
rect 18 116 30 119
rect 36 117 50 119
rect 56 118 81 119
rect 90 118 117 119
rect 56 117 82 118
rect 90 117 118 118
rect 35 116 50 117
rect 18 113 29 116
rect 35 113 49 116
rect 55 115 83 117
rect 91 116 119 117
rect 91 115 120 116
rect 4 108 14 113
rect 18 111 28 113
rect 34 112 49 113
rect 54 113 84 115
rect 92 114 120 115
rect 161 115 179 119
rect 187 118 188 119
rect 187 117 189 118
rect 161 114 163 115
rect 92 113 121 114
rect 161 113 162 114
rect 178 113 179 115
rect 187 113 188 114
rect 194 113 195 114
rect 54 112 85 113
rect 34 111 48 112
rect 18 110 27 111
rect 33 110 48 111
rect 17 109 27 110
rect 4 105 13 108
rect 17 106 26 109
rect 32 108 48 110
rect 53 111 85 112
rect 93 112 122 113
rect 53 109 86 111
rect 93 110 123 112
rect 187 111 196 113
rect 187 110 188 111
rect 31 107 48 108
rect 30 106 48 107
rect 52 108 81 109
rect 84 108 86 109
rect 94 109 124 110
rect 94 108 125 109
rect 52 107 76 108
rect 94 107 126 108
rect 52 106 72 107
rect 95 106 127 107
rect 187 106 189 107
rect 191 106 194 107
rect 16 105 26 106
rect 27 105 47 106
rect 4 102 12 105
rect 16 103 47 105
rect 52 105 70 106
rect 95 105 128 106
rect 52 104 68 105
rect 95 104 129 105
rect 51 103 67 104
rect 95 103 131 104
rect 170 103 172 105
rect 186 103 188 106
rect 190 105 195 106
rect 190 104 193 105
rect 189 103 192 104
rect 195 103 196 105
rect 5 101 12 102
rect 4 100 12 101
rect 15 101 46 103
rect 51 102 66 103
rect 96 102 132 103
rect 161 102 166 103
rect 51 101 65 102
rect 79 101 92 102
rect 96 101 110 102
rect 111 101 134 102
rect 15 100 45 101
rect 51 100 64 101
rect 76 100 111 101
rect 113 100 134 101
rect 161 101 165 102
rect 161 100 164 101
rect 170 100 179 103
rect 187 102 191 103
rect 194 102 196 103
rect 188 101 190 102
rect 193 101 195 102
rect 5 98 12 100
rect 14 99 44 100
rect 14 98 43 99
rect 50 98 63 100
rect 74 99 111 100
rect 117 99 130 100
rect 160 99 163 100
rect 170 99 180 100
rect 72 98 112 99
rect 5 97 13 98
rect 14 97 42 98
rect 50 97 62 98
rect 70 97 113 98
rect 5 96 40 97
rect 49 96 62 97
rect 69 96 114 97
rect 5 95 38 96
rect 5 94 36 95
rect 48 94 62 96
rect 68 95 115 96
rect 160 95 162 99
rect 170 97 172 99
rect 170 96 171 97
rect 178 95 180 99
rect 194 97 196 98
rect 69 94 116 95
rect 6 93 35 94
rect 47 93 62 94
rect 71 93 118 94
rect 147 93 148 94
rect 6 92 33 93
rect 45 92 62 93
rect 73 92 120 93
rect 145 92 148 93
rect 161 93 163 95
rect 177 94 180 95
rect 187 96 191 97
rect 193 96 196 97
rect 187 95 195 96
rect 177 93 179 94
rect 161 92 164 93
rect 175 92 179 93
rect 6 91 32 92
rect 44 91 62 92
rect 75 91 122 92
rect 142 91 148 92
rect 162 91 166 92
rect 173 91 179 92
rect 187 93 188 95
rect 190 94 194 95
rect 191 93 192 94
rect 195 93 196 94
rect 187 91 196 93
rect 6 90 31 91
rect 42 90 63 91
rect 78 90 125 91
rect 138 90 147 91
rect 162 90 178 91
rect 187 90 188 91
rect 6 89 30 90
rect 39 89 64 90
rect 80 89 147 90
rect 163 89 177 90
rect 7 88 29 89
rect 37 88 67 89
rect 81 88 146 89
rect 164 88 176 89
rect 7 86 28 88
rect 36 87 70 88
rect 83 87 146 88
rect 165 87 175 88
rect 34 86 72 87
rect 84 86 145 87
rect 168 86 172 87
rect 188 86 189 87
rect 193 86 195 87
rect 7 85 27 86
rect 33 85 74 86
rect 85 85 103 86
rect 105 85 145 86
rect 187 85 189 86
rect 8 83 26 85
rect 32 84 76 85
rect 86 84 103 85
rect 106 84 144 85
rect 161 84 162 85
rect 187 84 188 85
rect 32 83 77 84
rect 87 83 104 84
rect 108 83 143 84
rect 161 83 163 84
rect 190 83 192 86
rect 194 85 196 86
rect 195 83 196 84
rect 8 82 25 83
rect 31 82 78 83
rect 8 81 16 82
rect 21 81 24 82
rect 31 81 79 82
rect 88 81 105 83
rect 109 82 142 83
rect 161 82 179 83
rect 187 82 196 83
rect 111 81 141 82
rect 161 81 180 82
rect 187 81 195 82
rect 8 79 15 81
rect 31 80 80 81
rect 89 80 106 81
rect 112 80 140 81
rect 161 80 163 81
rect 172 80 179 81
rect 187 80 188 81
rect 194 80 196 81
rect 31 79 81 80
rect 90 79 106 80
rect 113 79 139 80
rect 8 77 14 79
rect 31 78 82 79
rect 90 78 107 79
rect 115 78 137 79
rect 161 78 162 80
rect 171 79 178 80
rect 170 78 176 79
rect 31 77 37 78
rect 38 77 83 78
rect 91 77 108 78
rect 117 77 136 78
rect 169 77 175 78
rect 8 73 13 77
rect 20 76 23 77
rect 31 76 34 77
rect 46 76 84 77
rect 92 76 108 77
rect 120 76 134 77
rect 168 76 174 77
rect 18 75 25 76
rect 49 75 85 76
rect 92 75 109 76
rect 124 75 130 76
rect 166 75 173 76
rect 187 75 189 76
rect 18 74 26 75
rect 52 74 86 75
rect 7 70 13 73
rect 17 72 27 74
rect 54 73 86 74
rect 93 74 110 75
rect 165 74 171 75
rect 187 74 192 75
rect 93 73 111 74
rect 164 73 170 74
rect 191 73 194 74
rect 55 72 87 73
rect 94 72 112 73
rect 163 72 169 73
rect 6 69 13 70
rect 16 71 28 72
rect 57 71 88 72
rect 94 71 113 72
rect 162 71 168 72
rect 178 71 179 73
rect 192 72 196 73
rect 16 70 29 71
rect 36 70 44 71
rect 58 70 88 71
rect 95 70 114 71
rect 161 70 167 71
rect 177 70 179 71
rect 16 69 31 70
rect 32 69 47 70
rect 59 69 89 70
rect 95 69 116 70
rect 6 67 14 69
rect 17 68 48 69
rect 61 68 89 69
rect 96 68 118 69
rect 161 68 179 70
rect 187 71 188 72
rect 189 71 195 72
rect 187 70 192 71
rect 187 69 190 70
rect 187 68 188 69
rect 17 67 50 68
rect 6 65 15 67
rect 17 66 51 67
rect 62 66 90 68
rect 96 67 121 68
rect 131 67 135 68
rect 161 67 163 68
rect 177 67 179 68
rect 97 66 134 67
rect 7 64 15 65
rect 18 65 53 66
rect 63 65 91 66
rect 18 64 54 65
rect 64 64 91 65
rect 98 65 133 66
rect 161 65 162 67
rect 178 66 179 67
rect 98 64 132 65
rect 8 63 16 64
rect 19 63 56 64
rect 65 63 91 64
rect 99 63 131 64
rect 8 62 15 63
rect 10 61 15 62
rect 19 62 57 63
rect 19 61 58 62
rect 66 61 92 63
rect 100 62 131 63
rect 161 63 162 64
rect 161 62 163 63
rect 187 62 195 64
rect 100 61 130 62
rect 161 61 166 62
rect 173 61 174 62
rect 187 61 188 62
rect 194 61 196 62
rect 12 60 13 61
rect 19 60 59 61
rect 18 59 60 60
rect 67 59 93 61
rect 101 60 129 61
rect 102 59 129 60
rect 161 60 177 61
rect 161 59 178 60
rect 17 58 61 59
rect 16 57 62 58
rect 68 57 94 59
rect 103 58 128 59
rect 161 58 163 59
rect 175 58 179 59
rect 105 57 127 58
rect 16 56 27 57
rect 28 56 62 57
rect 69 56 95 57
rect 106 56 126 57
rect 161 56 162 58
rect 176 57 179 58
rect 15 55 27 56
rect 15 51 28 55
rect 29 54 63 56
rect 69 55 96 56
rect 108 55 124 56
rect 70 54 96 55
rect 110 54 123 55
rect 30 52 64 54
rect 70 53 97 54
rect 113 53 121 54
rect 177 53 180 57
rect 187 56 196 57
rect 187 55 190 56
rect 191 55 196 56
rect 191 54 194 55
rect 190 53 193 54
rect 70 52 99 53
rect 161 52 162 53
rect 176 52 180 53
rect 189 52 192 53
rect 31 51 65 52
rect 16 49 29 51
rect 32 50 65 51
rect 71 51 101 52
rect 161 51 163 52
rect 175 51 179 52
rect 71 50 103 51
rect 33 49 65 50
rect 72 49 109 50
rect 161 49 179 51
rect 187 51 191 52
rect 187 50 190 51
rect 194 50 196 51
rect 187 49 196 50
rect 17 48 29 49
rect 35 48 66 49
rect 72 48 114 49
rect 161 48 178 49
rect 19 47 30 48
rect 36 47 51 48
rect 53 47 66 48
rect 20 46 30 47
rect 34 46 50 47
rect 22 45 31 46
rect 23 44 31 45
rect 33 45 50 46
rect 54 46 66 47
rect 73 47 113 48
rect 161 47 176 48
rect 73 46 112 47
rect 161 46 172 47
rect 33 44 51 45
rect 24 43 32 44
rect 33 43 52 44
rect 54 43 67 46
rect 74 45 111 46
rect 74 44 110 45
rect 161 44 162 46
rect 187 44 189 45
rect 75 43 109 44
rect 187 43 195 44
rect 25 42 52 43
rect 26 40 53 42
rect 27 39 53 40
rect 28 37 53 39
rect 55 40 68 43
rect 76 42 108 43
rect 194 42 196 43
rect 77 41 106 42
rect 161 41 162 42
rect 195 41 196 42
rect 78 40 104 41
rect 161 40 163 41
rect 194 40 196 41
rect 55 37 69 40
rect 80 39 102 40
rect 161 39 164 40
rect 187 39 188 40
rect 193 39 196 40
rect 82 38 100 39
rect 161 38 165 39
rect 187 38 195 39
rect 85 37 96 38
rect 161 37 167 38
rect 29 36 54 37
rect 30 34 54 36
rect 31 32 54 34
rect 56 36 68 37
rect 161 36 162 37
rect 165 36 169 37
rect 178 36 179 38
rect 187 37 194 38
rect 56 35 66 36
rect 167 35 179 36
rect 56 34 64 35
rect 169 34 179 35
rect 56 33 62 34
rect 167 33 179 34
rect 56 32 60 33
rect 161 32 162 33
rect 165 32 179 33
rect 32 31 53 32
rect 32 30 40 31
rect 41 30 53 31
rect 161 31 179 32
rect 161 30 170 31
rect 33 28 41 30
rect 42 29 52 30
rect 161 29 168 30
rect 178 29 179 31
rect 43 28 51 29
rect 161 28 166 29
rect 34 26 42 28
rect 44 27 49 28
rect 161 27 164 28
rect 45 26 47 27
rect 161 26 163 27
rect 35 25 42 26
rect 161 25 162 26
rect 36 24 42 25
rect 38 23 40 24
rect 161 21 162 23
rect 178 22 179 23
rect 177 21 179 22
rect 161 19 163 21
rect 176 20 179 21
rect 175 19 179 20
rect 161 18 164 19
rect 174 18 179 19
rect 161 17 165 18
rect 172 17 179 18
rect 161 15 162 17
rect 163 16 166 17
rect 171 16 178 17
rect 165 15 167 16
rect 169 15 177 16
rect 166 14 175 15
rect 167 13 174 14
rect 161 12 162 13
rect 168 12 172 13
rect 178 12 179 13
rect 161 11 163 12
rect 169 11 171 12
rect 177 11 179 12
rect 161 7 179 11
rect 161 6 163 7
rect 177 6 179 7
rect 161 5 162 6
rect 178 5 179 6
<< metal2 >>
rect 102 453 150 477
rect 194 476 195 477
rect 162 475 178 476
rect 180 475 183 476
rect 162 472 179 475
rect 173 471 177 472
rect 170 469 173 471
rect 174 469 177 471
rect 164 468 167 469
rect 163 467 168 468
rect 163 466 169 467
rect 162 465 169 466
rect 170 466 177 469
rect 170 465 174 466
rect 162 464 165 465
rect 166 464 174 465
rect 161 460 164 464
rect 167 462 174 464
rect 167 461 177 462
rect 180 461 184 475
rect 191 474 195 476
rect 191 473 193 474
rect 194 473 195 474
rect 196 475 197 476
rect 196 473 198 475
rect 191 471 197 473
rect 193 470 196 471
rect 191 469 193 470
rect 196 469 198 470
rect 189 467 197 469
rect 190 466 196 467
rect 191 464 197 465
rect 191 463 198 464
rect 196 462 197 463
rect 196 461 198 462
rect 167 460 184 461
rect 161 459 165 460
rect 166 459 184 460
rect 191 460 198 461
rect 191 459 197 460
rect 162 458 174 459
rect 162 457 169 458
rect 163 456 169 457
rect 164 455 168 456
rect 170 454 174 458
rect 178 457 184 459
rect 196 458 197 459
rect 191 457 193 458
rect 196 457 198 458
rect 189 456 198 457
rect 189 455 197 456
rect 191 454 193 455
rect 171 453 174 454
rect 188 451 190 453
rect 191 452 198 453
rect 191 451 197 452
rect 196 450 197 451
rect 191 449 193 450
rect 196 449 198 450
rect 189 448 198 449
rect 190 447 197 448
rect 191 446 193 447
rect 191 444 193 445
rect 194 444 197 446
rect 152 442 154 444
rect 191 443 198 444
rect 151 441 154 442
rect 150 440 154 441
rect 149 438 154 440
rect 148 437 154 438
rect 147 436 154 437
rect 108 435 128 436
rect 146 435 154 436
rect 107 434 128 435
rect 145 434 154 435
rect 106 433 128 434
rect 105 432 128 433
rect 144 432 154 434
rect 104 431 128 432
rect 143 431 154 432
rect 103 428 128 431
rect 142 430 154 431
rect 141 429 154 430
rect 102 414 128 428
rect 140 427 154 429
rect 139 426 154 427
rect 138 425 154 426
rect 137 424 154 425
rect 136 422 154 424
rect 135 421 154 422
rect 163 439 168 440
rect 163 438 171 439
rect 172 438 175 443
rect 191 442 195 443
rect 196 442 198 443
rect 192 441 194 442
rect 196 441 197 442
rect 192 440 193 441
rect 163 435 175 438
rect 163 421 166 435
rect 172 432 175 435
rect 191 439 198 440
rect 191 438 197 439
rect 191 436 193 438
rect 191 435 198 436
rect 191 434 197 435
rect 189 432 197 433
rect 172 428 184 432
rect 189 431 198 432
rect 189 430 197 431
rect 134 420 154 421
rect 164 420 165 421
rect 133 419 154 420
rect 132 418 154 419
rect 172 418 175 428
rect 191 425 198 426
rect 191 423 193 425
rect 194 424 197 425
rect 188 422 197 423
rect 188 421 198 422
rect 191 419 192 420
rect 196 419 197 420
rect 131 416 154 418
rect 191 417 193 419
rect 196 418 198 419
rect 195 417 197 418
rect 191 416 197 417
rect 130 415 153 416
rect 192 415 197 416
rect 129 414 152 415
rect 102 413 151 414
rect 191 413 193 415
rect 102 412 150 413
rect 62 402 75 403
rect 59 401 79 402
rect 57 400 81 401
rect 55 399 83 400
rect 53 398 85 399
rect 52 397 64 398
rect 74 397 86 398
rect 15 396 16 397
rect 51 396 59 397
rect 79 396 87 397
rect 14 395 18 396
rect 51 395 56 396
rect 82 395 87 396
rect 14 394 20 395
rect 51 394 54 395
rect 84 394 87 395
rect 15 393 22 394
rect 17 392 24 393
rect 20 391 26 392
rect 22 390 28 391
rect 68 390 74 391
rect 24 389 30 390
rect 56 389 61 390
rect 66 389 76 390
rect 15 388 30 389
rect 54 388 62 389
rect 65 388 77 389
rect 14 386 30 388
rect 53 387 63 388
rect 65 387 78 388
rect 52 386 78 387
rect 15 385 20 386
rect 52 385 79 386
rect 16 384 23 385
rect 51 384 57 385
rect 60 384 68 385
rect 74 384 79 385
rect 18 383 25 384
rect 20 382 27 383
rect 22 381 29 382
rect 24 380 30 381
rect 15 379 30 380
rect 51 379 56 384
rect 61 383 67 384
rect 62 380 66 383
rect 75 380 79 384
rect 61 379 67 380
rect 74 379 79 380
rect 14 377 30 379
rect 52 378 68 379
rect 73 378 79 379
rect 52 377 79 378
rect 102 378 113 412
rect 127 411 150 412
rect 191 412 198 413
rect 191 411 197 412
rect 127 410 149 411
rect 127 409 148 410
rect 191 409 197 410
rect 127 408 147 409
rect 191 408 198 409
rect 127 407 146 408
rect 127 405 145 407
rect 163 406 177 407
rect 180 406 183 407
rect 191 406 195 408
rect 196 407 197 408
rect 196 406 198 407
rect 127 404 144 405
rect 127 403 143 404
rect 127 402 142 403
rect 162 402 178 406
rect 127 400 141 402
rect 127 399 140 400
rect 164 399 168 402
rect 169 399 172 402
rect 127 398 139 399
rect 127 397 138 398
rect 164 397 172 399
rect 127 395 137 397
rect 164 396 173 397
rect 163 395 173 396
rect 127 394 136 395
rect 163 394 167 395
rect 169 394 174 395
rect 127 393 135 394
rect 163 393 166 394
rect 170 393 174 394
rect 127 392 134 393
rect 162 392 166 393
rect 127 391 133 392
rect 162 391 165 392
rect 127 389 132 391
rect 162 390 166 391
rect 171 390 174 393
rect 180 392 184 406
rect 191 405 193 406
rect 194 405 198 406
rect 194 404 197 405
rect 193 403 195 404
rect 191 401 195 403
rect 191 400 193 401
rect 194 400 195 401
rect 196 402 197 403
rect 196 400 198 402
rect 191 399 198 400
rect 191 398 197 399
rect 193 397 196 398
rect 191 396 192 397
rect 194 396 197 397
rect 191 395 193 396
rect 194 395 198 396
rect 191 393 195 395
rect 196 393 198 395
rect 193 392 194 393
rect 163 389 166 390
rect 170 389 174 390
rect 127 388 131 389
rect 163 388 167 389
rect 169 388 174 389
rect 176 388 184 392
rect 192 391 195 392
rect 191 390 195 391
rect 191 388 193 390
rect 194 388 195 390
rect 196 391 197 393
rect 196 388 198 391
rect 127 387 130 388
rect 163 387 173 388
rect 191 387 197 388
rect 128 386 129 387
rect 164 386 172 387
rect 192 386 197 387
rect 165 385 171 386
rect 194 385 195 386
rect 196 385 197 386
rect 189 384 193 385
rect 194 384 197 385
rect 189 383 197 384
rect 189 382 191 383
rect 192 382 195 383
rect 189 381 190 382
rect 192 381 194 382
rect 189 380 197 381
rect 189 379 198 380
rect 52 376 78 377
rect 53 375 63 376
rect 65 375 77 376
rect 16 374 21 375
rect 54 374 62 375
rect 66 374 76 375
rect 15 372 23 374
rect 56 373 60 374
rect 67 373 75 374
rect 15 371 18 372
rect 20 371 24 372
rect 14 367 17 371
rect 14 366 20 367
rect 21 366 24 371
rect 78 370 79 371
rect 76 369 79 370
rect 56 368 62 369
rect 75 368 79 369
rect 54 367 64 368
rect 73 367 79 368
rect 14 365 25 366
rect 53 365 65 367
rect 71 366 79 367
rect 70 365 79 366
rect 15 364 29 365
rect 18 363 30 364
rect 52 363 66 365
rect 69 364 79 365
rect 68 363 78 364
rect 23 362 30 363
rect 27 361 30 362
rect 51 362 58 363
rect 61 362 76 363
rect 15 360 16 361
rect 51 360 57 362
rect 62 361 75 362
rect 62 360 74 361
rect 14 359 22 360
rect 14 358 27 359
rect 14 357 30 358
rect 15 356 21 357
rect 22 356 30 357
rect 16 355 22 356
rect 27 355 30 356
rect 18 354 25 355
rect 20 353 27 354
rect 22 352 29 353
rect 51 352 56 360
rect 62 359 72 360
rect 62 358 71 359
rect 62 357 69 358
rect 62 354 68 357
rect 102 354 150 378
rect 191 374 192 375
rect 191 373 193 374
rect 194 373 197 375
rect 181 372 183 373
rect 191 372 198 373
rect 162 368 178 372
rect 172 365 173 366
rect 171 363 175 365
rect 170 362 174 363
rect 169 361 174 362
rect 168 360 173 361
rect 162 358 172 360
rect 162 357 171 358
rect 180 357 184 372
rect 191 371 195 372
rect 196 371 198 372
rect 192 370 194 371
rect 196 370 197 371
rect 191 368 198 369
rect 191 367 197 368
rect 191 366 193 367
rect 191 365 194 366
rect 196 365 197 366
rect 191 364 198 365
rect 191 363 194 364
rect 195 363 197 364
rect 194 362 195 363
rect 191 360 197 362
rect 191 358 193 360
rect 196 359 198 360
rect 196 358 197 359
rect 191 357 197 358
rect 162 356 172 357
rect 166 355 173 356
rect 176 355 184 357
rect 192 356 197 357
rect 169 354 174 355
rect 176 354 183 355
rect 62 353 67 354
rect 170 353 174 354
rect 188 353 190 355
rect 191 353 197 355
rect 62 352 68 353
rect 171 352 175 353
rect 24 351 30 352
rect 15 350 30 351
rect 14 349 30 350
rect 14 348 21 349
rect 14 347 24 348
rect 15 346 29 347
rect 51 346 79 352
rect 172 350 175 352
rect 191 352 192 353
rect 196 352 197 353
rect 191 351 193 352
rect 196 351 198 352
rect 173 349 174 350
rect 189 349 197 351
rect 191 348 193 349
rect 196 347 197 348
rect 191 346 198 347
rect 19 345 30 346
rect 24 344 30 345
rect 28 343 30 344
rect 191 345 197 346
rect 191 344 195 345
rect 196 344 198 345
rect 191 343 198 344
rect 21 336 25 337
rect 19 335 27 336
rect 51 335 79 341
rect 19 334 28 335
rect 18 333 29 334
rect 18 332 21 333
rect 26 332 30 333
rect 18 331 20 332
rect 27 331 30 332
rect 19 330 21 331
rect 28 330 30 331
rect 19 329 22 330
rect 27 329 30 330
rect 18 328 29 329
rect 18 327 30 328
rect 19 326 34 327
rect 24 325 34 326
rect 15 324 17 325
rect 28 324 34 325
rect 14 322 17 324
rect 19 323 22 324
rect 18 322 26 323
rect 15 321 17 322
rect 19 321 30 322
rect 20 320 30 321
rect 25 319 30 320
rect 51 318 56 331
rect 62 318 67 329
rect 21 317 22 318
rect 19 316 27 317
rect 18 314 30 316
rect 18 313 21 314
rect 25 313 30 314
rect 15 311 17 312
rect 19 311 21 313
rect 51 312 79 318
rect 102 316 113 343
rect 191 342 193 343
rect 194 342 197 343
rect 195 341 196 342
rect 174 339 175 340
rect 169 336 171 337
rect 162 322 165 336
rect 166 322 168 336
rect 169 329 172 336
rect 173 330 176 339
rect 191 338 193 341
rect 196 340 197 341
rect 196 339 198 340
rect 195 338 197 339
rect 191 337 197 338
rect 179 336 182 337
rect 192 336 196 337
rect 178 335 183 336
rect 189 335 190 336
rect 194 335 195 336
rect 196 335 197 336
rect 178 334 184 335
rect 177 333 184 334
rect 188 333 190 335
rect 191 334 198 335
rect 191 333 197 334
rect 177 330 180 333
rect 181 331 184 333
rect 191 331 198 332
rect 173 329 179 330
rect 169 325 179 329
rect 169 322 172 325
rect 162 318 172 322
rect 173 324 179 325
rect 14 310 22 311
rect 14 309 26 310
rect 15 308 30 309
rect 20 307 30 308
rect 25 306 30 307
rect 51 307 53 308
rect 85 307 87 308
rect 51 306 56 307
rect 82 306 87 307
rect 51 305 58 306
rect 80 305 87 306
rect 17 304 19 305
rect 51 304 62 305
rect 75 304 86 305
rect 16 303 20 304
rect 15 302 20 303
rect 25 303 27 304
rect 53 303 85 304
rect 25 302 28 303
rect 54 302 83 303
rect 14 301 18 302
rect 25 301 29 302
rect 56 301 82 302
rect 14 298 17 301
rect 26 300 30 301
rect 58 300 79 301
rect 14 297 18 298
rect 15 296 18 297
rect 27 296 30 300
rect 61 299 76 300
rect 67 298 70 299
rect 15 295 20 296
rect 26 295 30 296
rect 16 294 30 295
rect 17 293 29 294
rect 18 292 28 293
rect 102 292 150 316
rect 173 315 176 324
rect 177 323 179 324
rect 182 324 185 331
rect 191 330 197 331
rect 191 329 193 330
rect 191 328 194 329
rect 196 328 197 329
rect 191 327 198 328
rect 191 326 197 327
rect 191 324 197 325
rect 182 323 184 324
rect 191 323 198 324
rect 177 322 180 323
rect 181 322 184 323
rect 177 320 184 322
rect 196 321 197 323
rect 191 320 198 321
rect 177 319 183 320
rect 191 319 197 320
rect 178 318 183 319
rect 179 317 182 318
rect 192 317 197 318
rect 191 316 197 317
rect 174 314 175 315
rect 191 314 193 316
rect 191 313 198 314
rect 191 312 197 313
rect 191 311 193 312
rect 191 310 197 311
rect 191 309 198 310
rect 192 308 193 309
rect 196 308 197 309
rect 192 307 197 308
rect 191 306 198 307
rect 171 305 173 306
rect 191 305 197 306
rect 170 302 174 305
rect 191 304 193 305
rect 191 303 197 304
rect 191 302 198 303
rect 162 299 184 302
rect 191 300 193 302
rect 191 299 198 300
rect 163 298 183 299
rect 191 298 197 299
rect 194 297 195 298
rect 177 296 178 297
rect 192 296 197 297
rect 21 291 26 292
rect 67 284 70 285
rect 18 283 21 284
rect 63 283 71 284
rect 18 282 23 283
rect 62 282 71 283
rect 19 281 25 282
rect 61 281 71 282
rect 20 280 27 281
rect 60 280 71 281
rect 73 283 75 284
rect 73 282 77 283
rect 73 280 78 282
rect 22 279 29 280
rect 59 279 71 280
rect 72 279 79 280
rect 24 278 30 279
rect 59 278 65 279
rect 25 277 32 278
rect 59 277 63 278
rect 19 276 33 277
rect 18 275 34 276
rect 18 274 26 275
rect 31 274 34 275
rect 19 273 20 274
rect 32 272 34 274
rect 58 273 63 277
rect 59 272 64 273
rect 67 272 71 279
rect 73 278 79 279
rect 75 274 79 278
rect 74 272 79 274
rect 14 271 19 272
rect 59 271 79 272
rect 14 270 24 271
rect 14 269 29 270
rect 60 269 78 271
rect 14 268 30 269
rect 61 268 77 269
rect 15 267 21 268
rect 24 267 30 268
rect 62 267 76 268
rect 17 266 23 267
rect 29 266 30 267
rect 64 266 74 267
rect 19 265 26 266
rect 102 265 113 292
rect 164 291 167 296
rect 176 295 179 296
rect 191 295 197 296
rect 175 294 180 295
rect 175 293 179 294
rect 191 293 193 295
rect 196 293 198 295
rect 173 292 178 293
rect 191 292 197 293
rect 171 291 178 292
rect 192 291 197 292
rect 164 290 177 291
rect 193 290 194 291
rect 195 290 197 291
rect 164 288 175 290
rect 191 288 193 290
rect 196 288 198 290
rect 164 287 177 288
rect 164 282 167 287
rect 169 286 178 287
rect 191 286 197 288
rect 173 285 179 286
rect 193 285 196 286
rect 174 284 180 285
rect 192 284 195 285
rect 175 283 180 284
rect 176 282 180 283
rect 166 281 167 282
rect 177 281 180 282
rect 191 283 195 284
rect 191 282 193 283
rect 194 282 195 283
rect 191 281 195 282
rect 196 283 197 285
rect 196 281 198 283
rect 178 280 179 281
rect 191 280 197 281
rect 192 279 197 280
rect 188 276 197 278
rect 192 274 195 275
rect 191 273 195 274
rect 191 272 193 273
rect 194 272 195 273
rect 196 274 197 275
rect 196 272 198 274
rect 191 271 198 272
rect 191 270 197 271
rect 181 269 183 270
rect 162 265 178 269
rect 21 264 28 265
rect 23 263 30 264
rect 67 263 70 264
rect 15 262 30 263
rect 63 262 74 263
rect 166 262 170 265
rect 14 260 30 262
rect 62 261 76 262
rect 163 261 170 262
rect 172 262 173 263
rect 172 261 174 262
rect 61 260 77 261
rect 14 259 21 260
rect 60 259 78 260
rect 14 258 27 259
rect 59 258 79 259
rect 16 257 30 258
rect 59 257 66 258
rect 72 257 79 258
rect 21 256 30 257
rect 26 255 30 256
rect 58 256 64 257
rect 74 256 79 257
rect 58 254 63 256
rect 59 251 63 254
rect 75 252 79 256
rect 163 257 166 261
rect 171 260 175 261
rect 170 258 174 260
rect 168 257 173 258
rect 163 256 173 257
rect 163 254 172 256
rect 180 255 184 269
rect 189 268 190 270
rect 192 269 196 270
rect 189 267 197 268
rect 189 266 198 267
rect 189 265 191 266
rect 189 263 190 265
rect 188 259 197 260
rect 188 257 198 259
rect 163 253 173 254
rect 74 251 78 252
rect 60 250 64 251
rect 73 250 78 251
rect 61 249 67 250
rect 70 249 77 250
rect 17 247 21 248
rect 24 247 26 248
rect 16 246 22 247
rect 23 246 28 247
rect 15 245 29 246
rect 15 242 18 245
rect 20 244 29 245
rect 59 244 87 249
rect 20 243 24 244
rect 21 242 23 243
rect 15 241 20 242
rect 27 241 30 244
rect 16 240 20 241
rect 26 240 30 241
rect 83 241 86 242
rect 17 239 20 240
rect 25 238 29 240
rect 25 237 27 238
rect 23 230 26 236
rect 15 228 19 229
rect 24 228 26 229
rect 15 227 23 228
rect 24 227 27 228
rect 15 226 28 227
rect 16 225 30 226
rect 17 224 21 225
rect 23 224 30 225
rect 18 223 22 224
rect 20 222 23 223
rect 24 222 27 224
rect 28 223 30 224
rect 21 221 27 222
rect 22 220 27 221
rect 23 219 27 220
rect 24 218 27 219
rect 59 220 61 221
rect 83 220 87 241
rect 59 218 64 220
rect 83 219 86 220
rect 18 217 20 218
rect 16 216 22 217
rect 58 216 64 218
rect 15 215 23 216
rect 15 214 24 215
rect 15 212 18 214
rect 21 213 25 214
rect 22 212 26 213
rect 27 212 30 216
rect 59 215 64 216
rect 59 214 65 215
rect 60 213 67 214
rect 15 211 19 212
rect 23 211 30 212
rect 15 210 20 211
rect 24 210 30 211
rect 16 209 20 210
rect 25 209 30 210
rect 18 208 20 209
rect 26 208 30 209
rect 59 208 79 213
rect 27 207 30 208
rect 18 205 23 206
rect 16 204 26 205
rect 15 203 28 204
rect 15 200 18 203
rect 21 202 29 203
rect 25 201 29 202
rect 15 199 19 200
rect 16 198 22 199
rect 27 198 30 201
rect 17 197 30 198
rect 51 197 56 203
rect 59 197 79 203
rect 102 199 113 252
rect 121 201 131 252
rect 121 200 132 201
rect 140 200 150 252
rect 163 248 166 253
rect 168 252 174 253
rect 169 251 174 252
rect 176 252 184 255
rect 191 256 193 257
rect 196 256 198 257
rect 191 254 197 256
rect 193 253 196 254
rect 192 252 197 253
rect 176 251 183 252
rect 191 251 198 252
rect 170 250 175 251
rect 171 249 175 250
rect 172 248 175 249
rect 191 250 197 251
rect 191 249 193 250
rect 191 248 197 249
rect 172 247 174 248
rect 191 247 198 248
rect 192 245 197 246
rect 191 244 198 245
rect 191 243 197 244
rect 191 242 195 243
rect 196 242 198 243
rect 191 241 197 242
rect 191 240 193 241
rect 194 240 197 241
rect 171 236 173 237
rect 163 233 165 234
rect 170 233 174 236
rect 191 234 193 236
rect 194 235 197 236
rect 194 234 198 235
rect 162 229 174 233
rect 162 215 166 229
rect 170 225 174 229
rect 176 229 184 233
rect 191 232 195 234
rect 196 232 198 234
rect 192 231 194 232
rect 191 230 192 231
rect 196 230 197 232
rect 176 225 180 229
rect 191 228 193 230
rect 196 229 198 230
rect 195 228 197 229
rect 191 227 197 228
rect 192 226 196 227
rect 170 222 180 225
rect 188 223 190 225
rect 191 223 197 225
rect 163 214 165 215
rect 170 212 174 222
rect 176 215 180 222
rect 191 221 198 222
rect 191 220 197 221
rect 191 218 193 220
rect 191 217 198 218
rect 191 216 197 217
rect 177 214 179 215
rect 192 214 197 215
rect 191 213 197 214
rect 171 211 172 212
rect 191 211 193 213
rect 196 211 198 213
rect 191 210 197 211
rect 192 209 197 210
rect 191 208 196 209
rect 191 207 193 208
rect 191 206 197 207
rect 191 205 198 206
rect 191 204 197 205
rect 191 203 192 204
rect 196 203 197 204
rect 114 199 119 200
rect 120 199 138 200
rect 139 199 150 200
rect 168 199 171 202
rect 189 201 197 203
rect 190 200 196 201
rect 181 199 183 200
rect 191 199 192 200
rect 18 196 29 197
rect 21 195 28 196
rect 51 195 54 196
rect 17 193 21 194
rect 16 192 22 193
rect 27 192 29 193
rect 15 191 23 192
rect 15 188 18 191
rect 20 190 24 191
rect 21 189 25 190
rect 22 188 26 189
rect 27 188 30 192
rect 51 191 55 195
rect 59 191 63 195
rect 51 188 79 191
rect 15 187 20 188
rect 23 187 30 188
rect 16 186 20 187
rect 24 186 30 187
rect 52 186 79 188
rect 17 185 20 186
rect 25 185 30 186
rect 54 185 79 186
rect 18 184 19 185
rect 26 184 30 185
rect 28 183 30 184
rect 59 182 63 185
rect 102 182 150 199
rect 162 196 178 199
rect 165 193 167 194
rect 102 180 149 182
rect 162 181 164 190
rect 165 189 168 193
rect 171 192 174 193
rect 170 191 175 192
rect 169 189 176 191
rect 165 187 172 189
rect 173 187 176 189
rect 165 184 171 187
rect 174 184 176 187
rect 180 186 184 199
rect 191 196 193 199
rect 196 197 198 199
rect 195 196 197 197
rect 191 195 197 196
rect 193 194 196 195
rect 193 193 195 194
rect 191 191 195 193
rect 191 190 193 191
rect 194 190 195 191
rect 196 192 197 194
rect 196 190 198 192
rect 191 189 197 190
rect 192 188 197 189
rect 178 185 184 186
rect 188 185 197 187
rect 165 183 172 184
rect 173 183 176 184
rect 102 179 148 180
rect 102 178 147 179
rect 165 178 168 183
rect 169 181 176 183
rect 177 182 184 185
rect 178 181 183 182
rect 189 181 190 184
rect 192 181 194 184
rect 196 183 198 184
rect 196 181 197 183
rect 169 180 175 181
rect 170 179 175 180
rect 189 180 197 181
rect 189 179 198 180
rect 172 178 173 179
rect 189 178 197 179
rect 102 177 146 178
rect 102 176 144 177
rect 176 169 180 170
rect 163 167 167 169
rect 177 168 181 169
rect 169 167 174 168
rect 178 167 181 168
rect 163 165 165 167
rect 169 166 175 167
rect 179 166 181 167
rect 170 165 173 166
rect 163 162 164 165
rect 171 162 173 165
rect 180 163 181 166
rect 179 162 181 163
rect 163 157 181 162
rect 163 155 164 157
rect 180 155 181 157
rect 176 152 179 153
rect 42 151 48 152
rect 164 151 167 152
rect 176 151 181 152
rect 37 150 52 151
rect 34 149 52 150
rect 163 150 168 151
rect 178 150 181 151
rect 32 148 51 149
rect 163 148 165 150
rect 169 149 175 150
rect 179 149 181 150
rect 170 148 174 149
rect 31 147 49 148
rect 30 146 48 147
rect 29 145 46 146
rect 163 145 164 148
rect 171 145 173 148
rect 180 145 181 149
rect 28 144 45 145
rect 56 144 66 145
rect 163 144 165 145
rect 170 144 173 145
rect 179 144 181 145
rect 23 143 24 144
rect 28 143 44 144
rect 53 143 71 144
rect 20 142 24 143
rect 27 142 43 143
rect 51 142 73 143
rect 19 141 23 142
rect 18 140 23 141
rect 27 140 42 142
rect 50 141 75 142
rect 49 140 76 141
rect 163 140 181 144
rect 17 139 22 140
rect 16 138 22 139
rect 26 139 41 140
rect 48 139 77 140
rect 26 138 40 139
rect 47 138 73 139
rect 163 138 164 140
rect 180 138 181 140
rect 15 137 21 138
rect 14 136 21 137
rect 13 135 21 136
rect 25 136 39 138
rect 47 137 70 138
rect 189 137 190 138
rect 46 136 67 137
rect 189 136 192 137
rect 25 135 38 136
rect 45 135 65 136
rect 191 135 197 136
rect 13 134 20 135
rect 12 133 20 134
rect 11 132 20 133
rect 24 133 37 135
rect 44 134 63 135
rect 83 134 84 135
rect 85 134 94 135
rect 43 133 62 134
rect 81 133 99 134
rect 163 133 164 135
rect 180 134 181 135
rect 192 134 197 135
rect 179 133 181 134
rect 24 132 36 133
rect 43 132 60 133
rect 82 132 102 133
rect 10 130 19 132
rect 9 128 19 130
rect 23 131 36 132
rect 42 131 59 132
rect 83 131 104 132
rect 23 129 35 131
rect 41 130 58 131
rect 84 130 106 131
rect 41 129 57 130
rect 85 129 108 130
rect 163 129 181 133
rect 189 133 198 134
rect 189 132 192 133
rect 189 131 190 132
rect 22 128 35 129
rect 40 128 56 129
rect 68 128 73 129
rect 86 128 110 129
rect 163 128 165 129
rect 170 128 173 129
rect 179 128 181 129
rect 8 126 18 128
rect 22 126 34 128
rect 40 127 55 128
rect 66 127 76 128
rect 87 127 111 128
rect 7 123 18 126
rect 6 120 18 123
rect 21 125 34 126
rect 39 126 55 127
rect 64 126 77 127
rect 88 126 112 127
rect 163 126 164 128
rect 21 122 33 125
rect 39 123 54 126
rect 62 125 79 126
rect 88 125 114 126
rect 61 124 80 125
rect 89 124 115 125
rect 60 123 81 124
rect 90 123 116 124
rect 20 121 33 122
rect 38 121 53 123
rect 59 122 82 123
rect 90 122 117 123
rect 163 122 164 124
rect 170 122 172 128
rect 180 126 181 128
rect 188 126 191 127
rect 189 124 190 126
rect 191 124 195 125
rect 196 124 197 125
rect 180 122 181 124
rect 189 123 197 124
rect 189 122 198 123
rect 59 121 83 122
rect 91 121 118 122
rect 163 121 166 122
rect 170 121 173 122
rect 179 121 181 122
rect 6 115 17 120
rect 20 118 32 121
rect 38 119 52 121
rect 58 120 83 121
rect 92 120 119 121
rect 58 119 84 120
rect 92 119 120 120
rect 37 118 52 119
rect 20 115 31 118
rect 37 115 51 118
rect 57 117 85 119
rect 93 118 121 119
rect 93 117 122 118
rect 6 110 16 115
rect 20 113 30 115
rect 36 114 51 115
rect 56 115 86 117
rect 94 116 122 117
rect 163 117 181 121
rect 189 120 190 121
rect 189 119 191 120
rect 163 116 165 117
rect 94 115 123 116
rect 163 115 164 116
rect 180 115 181 117
rect 189 115 190 116
rect 196 115 197 116
rect 56 114 87 115
rect 36 113 50 114
rect 20 112 29 113
rect 35 112 50 113
rect 19 111 29 112
rect 6 107 15 110
rect 19 108 28 111
rect 34 110 50 112
rect 55 113 87 114
rect 95 114 124 115
rect 55 111 88 113
rect 95 112 125 114
rect 189 113 198 115
rect 189 112 190 113
rect 33 109 50 110
rect 32 108 50 109
rect 54 110 83 111
rect 86 110 88 111
rect 96 111 126 112
rect 96 110 127 111
rect 54 109 78 110
rect 96 109 128 110
rect 54 108 74 109
rect 97 108 129 109
rect 189 108 191 109
rect 193 108 196 109
rect 18 107 28 108
rect 29 107 49 108
rect 6 104 14 107
rect 18 105 49 107
rect 54 107 72 108
rect 97 107 130 108
rect 54 106 70 107
rect 97 106 131 107
rect 53 105 69 106
rect 97 105 133 106
rect 172 105 174 107
rect 188 105 190 108
rect 192 107 197 108
rect 192 106 195 107
rect 191 105 194 106
rect 197 105 198 107
rect 7 103 14 104
rect 6 102 14 103
rect 17 103 48 105
rect 53 104 68 105
rect 98 104 134 105
rect 163 104 168 105
rect 53 103 67 104
rect 81 103 94 104
rect 98 103 112 104
rect 113 103 136 104
rect 17 102 47 103
rect 53 102 66 103
rect 78 102 113 103
rect 115 102 136 103
rect 163 103 167 104
rect 163 102 166 103
rect 172 102 181 105
rect 189 104 193 105
rect 196 104 198 105
rect 190 103 192 104
rect 195 103 197 104
rect 7 100 14 102
rect 16 101 46 102
rect 16 100 45 101
rect 52 100 65 102
rect 76 101 113 102
rect 119 101 132 102
rect 162 101 165 102
rect 172 101 182 102
rect 74 100 114 101
rect 7 99 15 100
rect 16 99 44 100
rect 52 99 64 100
rect 72 99 115 100
rect 7 98 42 99
rect 51 98 64 99
rect 71 98 116 99
rect 7 97 40 98
rect 7 96 38 97
rect 50 96 64 98
rect 70 97 117 98
rect 162 97 164 101
rect 172 99 174 101
rect 172 98 173 99
rect 180 97 182 101
rect 196 99 198 100
rect 71 96 118 97
rect 8 95 37 96
rect 49 95 64 96
rect 73 95 120 96
rect 149 95 150 96
rect 8 94 35 95
rect 47 94 64 95
rect 75 94 122 95
rect 147 94 150 95
rect 163 95 165 97
rect 179 96 182 97
rect 189 98 193 99
rect 195 98 198 99
rect 189 97 197 98
rect 179 95 181 96
rect 163 94 166 95
rect 177 94 181 95
rect 8 93 34 94
rect 46 93 64 94
rect 77 93 124 94
rect 144 93 150 94
rect 164 93 168 94
rect 175 93 181 94
rect 189 95 190 97
rect 192 96 196 97
rect 193 95 194 96
rect 197 95 198 96
rect 189 93 198 95
rect 8 92 33 93
rect 44 92 65 93
rect 80 92 127 93
rect 140 92 149 93
rect 164 92 180 93
rect 189 92 190 93
rect 8 91 32 92
rect 41 91 66 92
rect 82 91 149 92
rect 165 91 179 92
rect 9 90 31 91
rect 39 90 69 91
rect 83 90 148 91
rect 166 90 178 91
rect 9 88 30 90
rect 38 89 72 90
rect 85 89 148 90
rect 167 89 177 90
rect 36 88 74 89
rect 86 88 147 89
rect 170 88 174 89
rect 190 88 191 89
rect 195 88 197 89
rect 9 87 29 88
rect 35 87 76 88
rect 87 87 105 88
rect 107 87 147 88
rect 189 87 191 88
rect 10 85 28 87
rect 34 86 78 87
rect 88 86 105 87
rect 108 86 146 87
rect 163 86 164 87
rect 189 86 190 87
rect 34 85 79 86
rect 89 85 106 86
rect 110 85 145 86
rect 163 85 165 86
rect 192 85 194 88
rect 196 87 198 88
rect 197 85 198 86
rect 10 84 27 85
rect 33 84 80 85
rect 10 83 18 84
rect 23 83 26 84
rect 33 83 81 84
rect 90 83 107 85
rect 111 84 144 85
rect 163 84 181 85
rect 189 84 198 85
rect 113 83 143 84
rect 163 83 182 84
rect 189 83 197 84
rect 10 81 17 83
rect 33 82 82 83
rect 91 82 108 83
rect 114 82 142 83
rect 163 82 165 83
rect 174 82 181 83
rect 189 82 190 83
rect 196 82 198 83
rect 33 81 83 82
rect 92 81 108 82
rect 115 81 141 82
rect 10 79 16 81
rect 33 80 84 81
rect 92 80 109 81
rect 117 80 139 81
rect 163 80 164 82
rect 173 81 180 82
rect 172 80 178 81
rect 33 79 39 80
rect 40 79 85 80
rect 93 79 110 80
rect 119 79 138 80
rect 171 79 177 80
rect 10 75 15 79
rect 22 78 25 79
rect 33 78 36 79
rect 48 78 86 79
rect 94 78 110 79
rect 122 78 136 79
rect 170 78 176 79
rect 20 77 27 78
rect 51 77 87 78
rect 94 77 111 78
rect 126 77 132 78
rect 168 77 175 78
rect 189 77 191 78
rect 20 76 28 77
rect 54 76 88 77
rect 9 72 15 75
rect 19 74 29 76
rect 56 75 88 76
rect 95 76 112 77
rect 167 76 173 77
rect 189 76 194 77
rect 95 75 113 76
rect 166 75 172 76
rect 193 75 196 76
rect 57 74 89 75
rect 96 74 114 75
rect 165 74 171 75
rect 8 71 15 72
rect 18 73 30 74
rect 59 73 90 74
rect 96 73 115 74
rect 164 73 170 74
rect 180 73 181 75
rect 194 74 198 75
rect 18 72 31 73
rect 38 72 46 73
rect 60 72 90 73
rect 97 72 116 73
rect 163 72 169 73
rect 179 72 181 73
rect 18 71 33 72
rect 34 71 49 72
rect 61 71 91 72
rect 97 71 118 72
rect 8 69 16 71
rect 19 70 50 71
rect 63 70 91 71
rect 98 70 120 71
rect 163 70 181 72
rect 189 73 190 74
rect 191 73 197 74
rect 189 72 194 73
rect 189 71 192 72
rect 189 70 190 71
rect 19 69 52 70
rect 8 67 17 69
rect 19 68 53 69
rect 64 68 92 70
rect 98 69 123 70
rect 133 69 137 70
rect 163 69 165 70
rect 179 69 181 70
rect 99 68 136 69
rect 9 66 17 67
rect 20 67 55 68
rect 65 67 93 68
rect 20 66 56 67
rect 66 66 93 67
rect 100 67 135 68
rect 163 67 164 69
rect 180 68 181 69
rect 100 66 134 67
rect 10 65 18 66
rect 21 65 58 66
rect 67 65 93 66
rect 101 65 133 66
rect 10 64 17 65
rect 12 63 17 64
rect 21 64 59 65
rect 21 63 60 64
rect 68 63 94 65
rect 102 64 133 65
rect 163 65 164 66
rect 163 64 165 65
rect 189 64 197 66
rect 102 63 132 64
rect 163 63 168 64
rect 175 63 176 64
rect 189 63 190 64
rect 196 63 198 64
rect 14 62 15 63
rect 21 62 61 63
rect 20 61 62 62
rect 69 61 95 63
rect 103 62 131 63
rect 104 61 131 62
rect 163 62 179 63
rect 163 61 180 62
rect 19 60 63 61
rect 18 59 64 60
rect 70 59 96 61
rect 105 60 130 61
rect 163 60 165 61
rect 177 60 181 61
rect 107 59 129 60
rect 18 58 29 59
rect 30 58 64 59
rect 71 58 97 59
rect 108 58 128 59
rect 163 58 164 60
rect 178 59 181 60
rect 17 57 29 58
rect 17 53 30 57
rect 31 56 65 58
rect 71 57 98 58
rect 110 57 126 58
rect 72 56 98 57
rect 112 56 125 57
rect 32 54 66 56
rect 72 55 99 56
rect 115 55 123 56
rect 179 55 182 59
rect 189 58 198 59
rect 189 57 192 58
rect 193 57 198 58
rect 193 56 196 57
rect 192 55 195 56
rect 72 54 101 55
rect 163 54 164 55
rect 178 54 182 55
rect 191 54 194 55
rect 33 53 67 54
rect 18 51 31 53
rect 34 52 67 53
rect 73 53 103 54
rect 163 53 165 54
rect 177 53 181 54
rect 73 52 105 53
rect 35 51 67 52
rect 74 51 111 52
rect 163 51 181 53
rect 189 53 193 54
rect 189 52 192 53
rect 196 52 198 53
rect 189 51 198 52
rect 19 50 31 51
rect 37 50 68 51
rect 74 50 116 51
rect 163 50 180 51
rect 21 49 32 50
rect 38 49 53 50
rect 55 49 68 50
rect 22 48 32 49
rect 36 48 52 49
rect 24 47 33 48
rect 25 46 33 47
rect 35 47 52 48
rect 56 48 68 49
rect 75 49 115 50
rect 163 49 178 50
rect 75 48 114 49
rect 163 48 174 49
rect 35 46 53 47
rect 26 45 34 46
rect 35 45 54 46
rect 56 45 69 48
rect 76 47 113 48
rect 76 46 112 47
rect 163 46 164 48
rect 189 46 191 47
rect 77 45 111 46
rect 189 45 197 46
rect 27 44 54 45
rect 28 42 55 44
rect 29 41 55 42
rect 30 39 55 41
rect 57 42 70 45
rect 78 44 110 45
rect 196 44 198 45
rect 79 43 108 44
rect 163 43 164 44
rect 197 43 198 44
rect 80 42 106 43
rect 163 42 165 43
rect 196 42 198 43
rect 57 39 71 42
rect 82 41 104 42
rect 163 41 166 42
rect 189 41 190 42
rect 195 41 198 42
rect 84 40 102 41
rect 163 40 167 41
rect 189 40 197 41
rect 87 39 98 40
rect 163 39 169 40
rect 31 38 56 39
rect 32 36 56 38
rect 33 34 56 36
rect 58 38 70 39
rect 163 38 164 39
rect 167 38 171 39
rect 180 38 181 40
rect 189 39 196 40
rect 58 37 68 38
rect 169 37 181 38
rect 58 36 66 37
rect 171 36 181 37
rect 58 35 64 36
rect 169 35 181 36
rect 58 34 62 35
rect 163 34 164 35
rect 167 34 181 35
rect 34 33 55 34
rect 34 32 42 33
rect 43 32 55 33
rect 163 33 181 34
rect 163 32 172 33
rect 35 30 43 32
rect 44 31 54 32
rect 163 31 170 32
rect 180 31 181 33
rect 45 30 53 31
rect 163 30 168 31
rect 36 28 44 30
rect 46 29 51 30
rect 163 29 166 30
rect 47 28 49 29
rect 163 28 165 29
rect 37 27 44 28
rect 163 27 164 28
rect 38 26 44 27
rect 40 25 42 26
rect 163 23 164 25
rect 180 24 181 25
rect 179 23 181 24
rect 163 21 165 23
rect 178 22 181 23
rect 177 21 181 22
rect 163 20 166 21
rect 176 20 181 21
rect 163 19 167 20
rect 174 19 181 20
rect 163 17 164 19
rect 165 18 168 19
rect 173 18 180 19
rect 167 17 169 18
rect 171 17 179 18
rect 168 16 177 17
rect 169 15 176 16
rect 163 14 164 15
rect 170 14 174 15
rect 180 14 181 15
rect 163 13 165 14
rect 171 13 173 14
rect 179 13 181 14
rect 163 9 181 13
rect 163 8 165 9
rect 179 8 181 9
rect 163 7 164 8
rect 180 7 181 8
<< metal3 >>
rect 104 455 152 479
rect 196 478 197 479
rect 164 477 180 478
rect 182 477 185 478
rect 164 474 181 477
rect 175 473 179 474
rect 172 471 175 473
rect 176 471 179 473
rect 166 470 169 471
rect 165 469 170 470
rect 165 468 171 469
rect 164 467 171 468
rect 172 468 179 471
rect 172 467 176 468
rect 164 466 167 467
rect 168 466 176 467
rect 163 462 166 466
rect 169 464 176 466
rect 169 463 179 464
rect 182 463 186 477
rect 193 476 197 478
rect 193 475 195 476
rect 196 475 197 476
rect 198 477 199 478
rect 198 475 200 477
rect 193 473 199 475
rect 195 472 198 473
rect 193 471 195 472
rect 198 471 200 472
rect 191 469 199 471
rect 192 468 198 469
rect 193 466 199 467
rect 193 465 200 466
rect 198 464 199 465
rect 198 463 200 464
rect 169 462 186 463
rect 163 461 167 462
rect 168 461 186 462
rect 193 462 200 463
rect 193 461 199 462
rect 164 460 176 461
rect 164 459 171 460
rect 165 458 171 459
rect 166 457 170 458
rect 172 456 176 460
rect 180 459 186 461
rect 198 460 199 461
rect 193 459 195 460
rect 198 459 200 460
rect 191 458 200 459
rect 191 457 199 458
rect 193 456 195 457
rect 173 455 176 456
rect 190 453 192 455
rect 193 454 200 455
rect 193 453 199 454
rect 198 452 199 453
rect 193 451 195 452
rect 198 451 200 452
rect 191 450 200 451
rect 192 449 199 450
rect 193 448 195 449
rect 193 446 195 447
rect 196 446 199 448
rect 154 444 156 446
rect 193 445 200 446
rect 153 443 156 444
rect 152 442 156 443
rect 151 440 156 442
rect 150 439 156 440
rect 149 438 156 439
rect 110 437 130 438
rect 148 437 156 438
rect 109 436 130 437
rect 147 436 156 437
rect 108 435 130 436
rect 107 434 130 435
rect 146 434 156 436
rect 106 433 130 434
rect 145 433 156 434
rect 105 430 130 433
rect 144 432 156 433
rect 143 431 156 432
rect 104 416 130 430
rect 142 429 156 431
rect 141 428 156 429
rect 140 427 156 428
rect 139 426 156 427
rect 138 424 156 426
rect 137 423 156 424
rect 165 441 170 442
rect 165 440 173 441
rect 174 440 177 445
rect 193 444 197 445
rect 198 444 200 445
rect 194 443 196 444
rect 198 443 199 444
rect 194 442 195 443
rect 165 437 177 440
rect 165 423 168 437
rect 174 434 177 437
rect 193 441 200 442
rect 193 440 199 441
rect 193 438 195 440
rect 193 437 200 438
rect 193 436 199 437
rect 191 434 199 435
rect 174 430 186 434
rect 191 433 200 434
rect 191 432 199 433
rect 136 422 156 423
rect 166 422 167 423
rect 135 421 156 422
rect 134 420 156 421
rect 174 420 177 430
rect 193 427 200 428
rect 193 425 195 427
rect 196 426 199 427
rect 190 424 199 425
rect 190 423 200 424
rect 193 421 194 422
rect 198 421 199 422
rect 133 418 156 420
rect 193 419 195 421
rect 198 420 200 421
rect 197 419 199 420
rect 193 418 199 419
rect 132 417 155 418
rect 194 417 199 418
rect 131 416 154 417
rect 104 415 153 416
rect 193 415 195 417
rect 104 414 152 415
rect 64 404 77 405
rect 61 403 81 404
rect 59 402 83 403
rect 57 401 85 402
rect 55 400 87 401
rect 54 399 66 400
rect 76 399 88 400
rect 17 398 18 399
rect 53 398 61 399
rect 81 398 89 399
rect 16 397 20 398
rect 53 397 58 398
rect 84 397 89 398
rect 16 396 22 397
rect 53 396 56 397
rect 86 396 89 397
rect 17 395 24 396
rect 19 394 26 395
rect 22 393 28 394
rect 24 392 30 393
rect 70 392 76 393
rect 26 391 32 392
rect 58 391 63 392
rect 68 391 78 392
rect 17 390 32 391
rect 56 390 64 391
rect 67 390 79 391
rect 16 388 32 390
rect 55 389 65 390
rect 67 389 80 390
rect 54 388 80 389
rect 17 387 22 388
rect 54 387 81 388
rect 18 386 25 387
rect 53 386 59 387
rect 62 386 70 387
rect 76 386 81 387
rect 20 385 27 386
rect 22 384 29 385
rect 24 383 31 384
rect 26 382 32 383
rect 17 381 32 382
rect 53 381 58 386
rect 63 385 69 386
rect 64 382 68 385
rect 77 382 81 386
rect 63 381 69 382
rect 76 381 81 382
rect 16 379 32 381
rect 54 380 70 381
rect 75 380 81 381
rect 54 379 81 380
rect 104 380 115 414
rect 129 413 152 414
rect 193 414 200 415
rect 193 413 199 414
rect 129 412 151 413
rect 129 411 150 412
rect 193 411 199 412
rect 129 410 149 411
rect 193 410 200 411
rect 129 409 148 410
rect 129 407 147 409
rect 165 408 179 409
rect 182 408 185 409
rect 193 408 197 410
rect 198 409 199 410
rect 198 408 200 409
rect 129 406 146 407
rect 129 405 145 406
rect 129 404 144 405
rect 164 404 180 408
rect 129 402 143 404
rect 129 401 142 402
rect 166 401 170 404
rect 171 401 174 404
rect 129 400 141 401
rect 129 399 140 400
rect 166 399 174 401
rect 129 397 139 399
rect 166 398 175 399
rect 165 397 175 398
rect 129 396 138 397
rect 165 396 169 397
rect 171 396 176 397
rect 129 395 137 396
rect 165 395 168 396
rect 172 395 176 396
rect 129 394 136 395
rect 164 394 168 395
rect 129 393 135 394
rect 164 393 167 394
rect 129 391 134 393
rect 164 392 168 393
rect 173 392 176 395
rect 182 394 186 408
rect 193 407 195 408
rect 196 407 200 408
rect 196 406 199 407
rect 195 405 197 406
rect 193 403 197 405
rect 193 402 195 403
rect 196 402 197 403
rect 198 404 199 405
rect 198 402 200 404
rect 193 401 200 402
rect 193 400 199 401
rect 195 399 198 400
rect 193 398 194 399
rect 196 398 199 399
rect 193 397 195 398
rect 196 397 200 398
rect 193 395 197 397
rect 198 395 200 397
rect 195 394 196 395
rect 165 391 168 392
rect 172 391 176 392
rect 129 390 133 391
rect 165 390 169 391
rect 171 390 176 391
rect 178 390 186 394
rect 194 393 197 394
rect 193 392 197 393
rect 193 390 195 392
rect 196 390 197 392
rect 198 393 199 395
rect 198 390 200 393
rect 129 389 132 390
rect 165 389 175 390
rect 193 389 199 390
rect 130 388 131 389
rect 166 388 174 389
rect 194 388 199 389
rect 167 387 173 388
rect 196 387 197 388
rect 198 387 199 388
rect 191 386 195 387
rect 196 386 199 387
rect 191 385 199 386
rect 191 384 193 385
rect 194 384 197 385
rect 191 383 192 384
rect 194 383 196 384
rect 191 382 199 383
rect 191 381 200 382
rect 54 378 80 379
rect 55 377 65 378
rect 67 377 79 378
rect 18 376 23 377
rect 56 376 64 377
rect 68 376 78 377
rect 17 374 25 376
rect 58 375 62 376
rect 69 375 77 376
rect 17 373 20 374
rect 22 373 26 374
rect 16 369 19 373
rect 16 368 22 369
rect 23 368 26 373
rect 80 372 81 373
rect 78 371 81 372
rect 58 370 64 371
rect 77 370 81 371
rect 56 369 66 370
rect 75 369 81 370
rect 16 367 27 368
rect 55 367 67 369
rect 73 368 81 369
rect 72 367 81 368
rect 17 366 31 367
rect 20 365 32 366
rect 54 365 68 367
rect 71 366 81 367
rect 70 365 80 366
rect 25 364 32 365
rect 29 363 32 364
rect 53 364 60 365
rect 63 364 78 365
rect 17 362 18 363
rect 53 362 59 364
rect 64 363 77 364
rect 64 362 76 363
rect 16 361 24 362
rect 16 360 29 361
rect 16 359 32 360
rect 17 358 23 359
rect 24 358 32 359
rect 18 357 24 358
rect 29 357 32 358
rect 20 356 27 357
rect 22 355 29 356
rect 24 354 31 355
rect 53 354 58 362
rect 64 361 74 362
rect 64 360 73 361
rect 64 359 71 360
rect 64 356 70 359
rect 104 356 152 380
rect 193 376 194 377
rect 193 375 195 376
rect 196 375 199 377
rect 183 374 185 375
rect 193 374 200 375
rect 164 370 180 374
rect 174 367 175 368
rect 173 365 177 367
rect 172 364 176 365
rect 171 363 176 364
rect 170 362 175 363
rect 164 360 174 362
rect 164 359 173 360
rect 182 359 186 374
rect 193 373 197 374
rect 198 373 200 374
rect 194 372 196 373
rect 198 372 199 373
rect 193 370 200 371
rect 193 369 199 370
rect 193 368 195 369
rect 193 367 196 368
rect 198 367 199 368
rect 193 366 200 367
rect 193 365 196 366
rect 197 365 199 366
rect 196 364 197 365
rect 193 362 199 364
rect 193 360 195 362
rect 198 361 200 362
rect 198 360 199 361
rect 193 359 199 360
rect 164 358 174 359
rect 168 357 175 358
rect 178 357 186 359
rect 194 358 199 359
rect 171 356 176 357
rect 178 356 185 357
rect 64 355 69 356
rect 172 355 176 356
rect 190 355 192 357
rect 193 355 199 357
rect 64 354 70 355
rect 173 354 177 355
rect 26 353 32 354
rect 17 352 32 353
rect 16 351 32 352
rect 16 350 23 351
rect 16 349 26 350
rect 17 348 31 349
rect 53 348 81 354
rect 174 352 177 354
rect 193 354 194 355
rect 198 354 199 355
rect 193 353 195 354
rect 198 353 200 354
rect 175 351 176 352
rect 191 351 199 353
rect 193 350 195 351
rect 198 349 199 350
rect 193 348 200 349
rect 21 347 32 348
rect 26 346 32 347
rect 30 345 32 346
rect 193 347 199 348
rect 193 346 197 347
rect 198 346 200 347
rect 193 345 200 346
rect 23 338 27 339
rect 21 337 29 338
rect 53 337 81 343
rect 21 336 30 337
rect 20 335 31 336
rect 20 334 23 335
rect 28 334 32 335
rect 20 333 22 334
rect 29 333 32 334
rect 21 332 23 333
rect 30 332 32 333
rect 21 331 24 332
rect 29 331 32 332
rect 20 330 31 331
rect 20 329 32 330
rect 21 328 36 329
rect 26 327 36 328
rect 17 326 19 327
rect 30 326 36 327
rect 16 324 19 326
rect 21 325 24 326
rect 20 324 28 325
rect 17 323 19 324
rect 21 323 32 324
rect 22 322 32 323
rect 27 321 32 322
rect 53 320 58 333
rect 64 320 69 331
rect 23 319 24 320
rect 21 318 29 319
rect 20 316 32 318
rect 20 315 23 316
rect 27 315 32 316
rect 17 313 19 314
rect 21 313 23 315
rect 53 314 81 320
rect 104 318 115 345
rect 193 344 195 345
rect 196 344 199 345
rect 197 343 198 344
rect 176 341 177 342
rect 171 338 173 339
rect 164 324 167 338
rect 168 324 170 338
rect 171 331 174 338
rect 175 332 178 341
rect 193 340 195 343
rect 198 342 199 343
rect 198 341 200 342
rect 197 340 199 341
rect 193 339 199 340
rect 181 338 184 339
rect 194 338 198 339
rect 180 337 185 338
rect 191 337 192 338
rect 196 337 197 338
rect 198 337 199 338
rect 180 336 186 337
rect 179 335 186 336
rect 190 335 192 337
rect 193 336 200 337
rect 193 335 199 336
rect 179 332 182 335
rect 183 333 186 335
rect 193 333 200 334
rect 175 331 181 332
rect 171 327 181 331
rect 171 324 174 327
rect 164 320 174 324
rect 175 326 181 327
rect 16 312 24 313
rect 16 311 28 312
rect 17 310 32 311
rect 22 309 32 310
rect 27 308 32 309
rect 53 309 55 310
rect 87 309 89 310
rect 53 308 58 309
rect 84 308 89 309
rect 53 307 60 308
rect 82 307 89 308
rect 19 306 21 307
rect 53 306 64 307
rect 77 306 88 307
rect 18 305 22 306
rect 17 304 22 305
rect 27 305 29 306
rect 55 305 87 306
rect 27 304 30 305
rect 56 304 85 305
rect 16 303 20 304
rect 27 303 31 304
rect 58 303 84 304
rect 16 300 19 303
rect 28 302 32 303
rect 60 302 81 303
rect 16 299 20 300
rect 17 298 20 299
rect 29 298 32 302
rect 63 301 78 302
rect 69 300 72 301
rect 17 297 22 298
rect 28 297 32 298
rect 18 296 32 297
rect 19 295 31 296
rect 20 294 30 295
rect 104 294 152 318
rect 175 317 178 326
rect 179 325 181 326
rect 184 326 187 333
rect 193 332 199 333
rect 193 331 195 332
rect 193 330 196 331
rect 198 330 199 331
rect 193 329 200 330
rect 193 328 199 329
rect 193 326 199 327
rect 184 325 186 326
rect 193 325 200 326
rect 179 324 182 325
rect 183 324 186 325
rect 179 322 186 324
rect 198 323 199 325
rect 193 322 200 323
rect 179 321 185 322
rect 193 321 199 322
rect 180 320 185 321
rect 181 319 184 320
rect 194 319 199 320
rect 193 318 199 319
rect 176 316 177 317
rect 193 316 195 318
rect 193 315 200 316
rect 193 314 199 315
rect 193 313 195 314
rect 193 312 199 313
rect 193 311 200 312
rect 194 310 195 311
rect 198 310 199 311
rect 194 309 199 310
rect 193 308 200 309
rect 173 307 175 308
rect 193 307 199 308
rect 172 304 176 307
rect 193 306 195 307
rect 193 305 199 306
rect 193 304 200 305
rect 164 301 186 304
rect 193 302 195 304
rect 193 301 200 302
rect 165 300 185 301
rect 193 300 199 301
rect 196 299 197 300
rect 179 298 180 299
rect 194 298 199 299
rect 23 293 28 294
rect 69 286 72 287
rect 20 285 23 286
rect 65 285 73 286
rect 20 284 25 285
rect 64 284 73 285
rect 21 283 27 284
rect 63 283 73 284
rect 22 282 29 283
rect 62 282 73 283
rect 75 285 77 286
rect 75 284 79 285
rect 75 282 80 284
rect 24 281 31 282
rect 61 281 73 282
rect 74 281 81 282
rect 26 280 32 281
rect 61 280 67 281
rect 27 279 34 280
rect 61 279 65 280
rect 21 278 35 279
rect 20 277 36 278
rect 20 276 28 277
rect 33 276 36 277
rect 21 275 22 276
rect 34 274 36 276
rect 60 275 65 279
rect 61 274 66 275
rect 69 274 73 281
rect 75 280 81 281
rect 77 276 81 280
rect 76 274 81 276
rect 16 273 21 274
rect 61 273 81 274
rect 16 272 26 273
rect 16 271 31 272
rect 62 271 80 273
rect 16 270 32 271
rect 63 270 79 271
rect 17 269 23 270
rect 26 269 32 270
rect 64 269 78 270
rect 19 268 25 269
rect 31 268 32 269
rect 66 268 76 269
rect 21 267 28 268
rect 104 267 115 294
rect 166 293 169 298
rect 178 297 181 298
rect 193 297 199 298
rect 177 296 182 297
rect 177 295 181 296
rect 193 295 195 297
rect 198 295 200 297
rect 175 294 180 295
rect 193 294 199 295
rect 173 293 180 294
rect 194 293 199 294
rect 166 292 179 293
rect 195 292 196 293
rect 197 292 199 293
rect 166 290 177 292
rect 193 290 195 292
rect 198 290 200 292
rect 166 289 179 290
rect 166 284 169 289
rect 171 288 180 289
rect 193 288 199 290
rect 175 287 181 288
rect 195 287 198 288
rect 176 286 182 287
rect 194 286 197 287
rect 177 285 182 286
rect 178 284 182 285
rect 168 283 169 284
rect 179 283 182 284
rect 193 285 197 286
rect 193 284 195 285
rect 196 284 197 285
rect 193 283 197 284
rect 198 285 199 287
rect 198 283 200 285
rect 180 282 181 283
rect 193 282 199 283
rect 194 281 199 282
rect 190 278 199 280
rect 194 276 197 277
rect 193 275 197 276
rect 193 274 195 275
rect 196 274 197 275
rect 198 276 199 277
rect 198 274 200 276
rect 193 273 200 274
rect 193 272 199 273
rect 183 271 185 272
rect 164 267 180 271
rect 23 266 30 267
rect 25 265 32 266
rect 69 265 72 266
rect 17 264 32 265
rect 65 264 76 265
rect 168 264 172 267
rect 16 262 32 264
rect 64 263 78 264
rect 165 263 172 264
rect 174 264 175 265
rect 174 263 176 264
rect 63 262 79 263
rect 16 261 23 262
rect 62 261 80 262
rect 16 260 29 261
rect 61 260 81 261
rect 18 259 32 260
rect 61 259 68 260
rect 74 259 81 260
rect 23 258 32 259
rect 28 257 32 258
rect 60 258 66 259
rect 76 258 81 259
rect 60 256 65 258
rect 61 253 65 256
rect 77 254 81 258
rect 165 259 168 263
rect 173 262 177 263
rect 172 260 176 262
rect 170 259 175 260
rect 165 258 175 259
rect 165 256 174 258
rect 182 257 186 271
rect 191 270 192 272
rect 194 271 198 272
rect 191 269 199 270
rect 191 268 200 269
rect 191 267 193 268
rect 191 265 192 267
rect 190 261 199 262
rect 190 259 200 261
rect 165 255 175 256
rect 76 253 80 254
rect 62 252 66 253
rect 75 252 80 253
rect 63 251 69 252
rect 72 251 79 252
rect 19 249 23 250
rect 26 249 28 250
rect 18 248 24 249
rect 25 248 30 249
rect 17 247 31 248
rect 17 244 20 247
rect 22 246 31 247
rect 61 246 89 251
rect 22 245 26 246
rect 23 244 25 245
rect 17 243 22 244
rect 29 243 32 246
rect 18 242 22 243
rect 28 242 32 243
rect 85 243 88 244
rect 19 241 22 242
rect 27 240 31 242
rect 27 239 29 240
rect 25 232 28 238
rect 17 230 21 231
rect 26 230 28 231
rect 17 229 25 230
rect 26 229 29 230
rect 17 228 30 229
rect 18 227 32 228
rect 19 226 23 227
rect 25 226 32 227
rect 20 225 24 226
rect 22 224 25 225
rect 26 224 29 226
rect 30 225 32 226
rect 23 223 29 224
rect 24 222 29 223
rect 25 221 29 222
rect 26 220 29 221
rect 61 222 63 223
rect 85 222 89 243
rect 61 220 66 222
rect 85 221 88 222
rect 20 219 22 220
rect 18 218 24 219
rect 60 218 66 220
rect 17 217 25 218
rect 17 216 26 217
rect 17 214 20 216
rect 23 215 27 216
rect 24 214 28 215
rect 29 214 32 218
rect 61 217 66 218
rect 61 216 67 217
rect 62 215 69 216
rect 17 213 21 214
rect 25 213 32 214
rect 17 212 22 213
rect 26 212 32 213
rect 18 211 22 212
rect 27 211 32 212
rect 20 210 22 211
rect 28 210 32 211
rect 61 210 81 215
rect 29 209 32 210
rect 20 207 25 208
rect 18 206 28 207
rect 17 205 30 206
rect 17 202 20 205
rect 23 204 31 205
rect 27 203 31 204
rect 17 201 21 202
rect 18 200 24 201
rect 29 200 32 203
rect 19 199 32 200
rect 53 199 58 205
rect 61 199 81 205
rect 104 201 115 254
rect 123 203 133 254
rect 123 202 134 203
rect 142 202 152 254
rect 165 250 168 255
rect 170 254 176 255
rect 171 253 176 254
rect 178 254 186 257
rect 193 258 195 259
rect 198 258 200 259
rect 193 256 199 258
rect 195 255 198 256
rect 194 254 199 255
rect 178 253 185 254
rect 193 253 200 254
rect 172 252 177 253
rect 173 251 177 252
rect 174 250 177 251
rect 193 252 199 253
rect 193 251 195 252
rect 193 250 199 251
rect 174 249 176 250
rect 193 249 200 250
rect 194 247 199 248
rect 193 246 200 247
rect 193 245 199 246
rect 193 244 197 245
rect 198 244 200 245
rect 193 243 199 244
rect 193 242 195 243
rect 196 242 199 243
rect 173 238 175 239
rect 165 235 167 236
rect 172 235 176 238
rect 193 236 195 238
rect 196 237 199 238
rect 196 236 200 237
rect 164 231 176 235
rect 164 217 168 231
rect 172 227 176 231
rect 178 231 186 235
rect 193 234 197 236
rect 198 234 200 236
rect 194 233 196 234
rect 193 232 194 233
rect 198 232 199 234
rect 178 227 182 231
rect 193 230 195 232
rect 198 231 200 232
rect 197 230 199 231
rect 193 229 199 230
rect 194 228 198 229
rect 172 224 182 227
rect 190 225 192 227
rect 193 225 199 227
rect 165 216 167 217
rect 172 214 176 224
rect 178 217 182 224
rect 193 223 200 224
rect 193 222 199 223
rect 193 220 195 222
rect 193 219 200 220
rect 193 218 199 219
rect 179 216 181 217
rect 194 216 199 217
rect 193 215 199 216
rect 173 213 174 214
rect 193 213 195 215
rect 198 213 200 215
rect 193 212 199 213
rect 194 211 199 212
rect 193 210 198 211
rect 193 209 195 210
rect 193 208 199 209
rect 193 207 200 208
rect 193 206 199 207
rect 193 205 194 206
rect 198 205 199 206
rect 116 201 121 202
rect 122 201 140 202
rect 141 201 152 202
rect 170 201 173 204
rect 191 203 199 205
rect 192 202 198 203
rect 183 201 185 202
rect 193 201 194 202
rect 20 198 31 199
rect 23 197 30 198
rect 53 197 56 198
rect 19 195 23 196
rect 18 194 24 195
rect 29 194 31 195
rect 17 193 25 194
rect 17 190 20 193
rect 22 192 26 193
rect 23 191 27 192
rect 24 190 28 191
rect 29 190 32 194
rect 53 193 57 197
rect 61 193 65 197
rect 53 190 81 193
rect 17 189 22 190
rect 25 189 32 190
rect 18 188 22 189
rect 26 188 32 189
rect 54 188 81 190
rect 19 187 22 188
rect 27 187 32 188
rect 56 187 81 188
rect 20 186 21 187
rect 28 186 32 187
rect 30 185 32 186
rect 61 184 65 187
rect 104 184 152 201
rect 164 198 180 201
rect 167 195 169 196
rect 104 182 151 184
rect 164 183 166 192
rect 167 191 170 195
rect 173 194 176 195
rect 172 193 177 194
rect 171 191 178 193
rect 167 189 174 191
rect 175 189 178 191
rect 167 186 173 189
rect 176 186 178 189
rect 182 188 186 201
rect 193 198 195 201
rect 198 199 200 201
rect 197 198 199 199
rect 193 197 199 198
rect 195 196 198 197
rect 195 195 197 196
rect 193 193 197 195
rect 193 192 195 193
rect 196 192 197 193
rect 198 194 199 196
rect 198 192 200 194
rect 193 191 199 192
rect 194 190 199 191
rect 180 187 186 188
rect 190 187 199 189
rect 167 185 174 186
rect 175 185 178 186
rect 104 181 150 182
rect 104 180 149 181
rect 167 180 170 185
rect 171 183 178 185
rect 179 184 186 187
rect 180 183 185 184
rect 191 183 192 186
rect 194 183 196 186
rect 198 185 200 186
rect 198 183 199 185
rect 171 182 177 183
rect 172 181 177 182
rect 191 182 199 183
rect 191 181 200 182
rect 174 180 175 181
rect 191 180 199 181
rect 104 179 148 180
rect 104 178 146 179
rect 178 171 182 172
rect 165 169 169 171
rect 179 170 183 171
rect 171 169 176 170
rect 180 169 183 170
rect 165 167 167 169
rect 171 168 177 169
rect 181 168 183 169
rect 172 167 175 168
rect 165 164 166 167
rect 173 164 175 167
rect 182 165 183 168
rect 181 164 183 165
rect 165 159 183 164
rect 165 157 166 159
rect 182 157 183 159
rect 178 154 181 155
rect 44 153 50 154
rect 166 153 169 154
rect 178 153 183 154
rect 39 152 54 153
rect 36 151 54 152
rect 165 152 170 153
rect 180 152 183 153
rect 34 150 53 151
rect 165 150 167 152
rect 171 151 177 152
rect 181 151 183 152
rect 172 150 176 151
rect 33 149 51 150
rect 32 148 50 149
rect 31 147 48 148
rect 165 147 166 150
rect 173 147 175 150
rect 182 147 183 151
rect 30 146 47 147
rect 58 146 68 147
rect 165 146 167 147
rect 172 146 175 147
rect 181 146 183 147
rect 25 145 26 146
rect 30 145 46 146
rect 55 145 73 146
rect 22 144 26 145
rect 29 144 45 145
rect 53 144 75 145
rect 21 143 25 144
rect 20 142 25 143
rect 29 142 44 144
rect 52 143 77 144
rect 51 142 78 143
rect 165 142 183 146
rect 19 141 24 142
rect 18 140 24 141
rect 28 141 43 142
rect 50 141 79 142
rect 28 140 42 141
rect 49 140 75 141
rect 165 140 166 142
rect 182 140 183 142
rect 17 139 23 140
rect 16 138 23 139
rect 15 137 23 138
rect 27 138 41 140
rect 49 139 72 140
rect 191 139 192 140
rect 48 138 69 139
rect 191 138 194 139
rect 27 137 40 138
rect 47 137 67 138
rect 193 137 199 138
rect 15 136 22 137
rect 14 135 22 136
rect 13 134 22 135
rect 26 135 39 137
rect 46 136 65 137
rect 85 136 86 137
rect 87 136 96 137
rect 45 135 64 136
rect 83 135 101 136
rect 165 135 166 137
rect 182 136 183 137
rect 194 136 199 137
rect 181 135 183 136
rect 26 134 38 135
rect 45 134 62 135
rect 84 134 104 135
rect 12 132 21 134
rect 11 130 21 132
rect 25 133 38 134
rect 44 133 61 134
rect 85 133 106 134
rect 25 131 37 133
rect 43 132 60 133
rect 86 132 108 133
rect 43 131 59 132
rect 87 131 110 132
rect 165 131 183 135
rect 191 135 200 136
rect 191 134 194 135
rect 191 133 192 134
rect 24 130 37 131
rect 42 130 58 131
rect 70 130 75 131
rect 88 130 112 131
rect 165 130 167 131
rect 172 130 175 131
rect 181 130 183 131
rect 10 128 20 130
rect 24 128 36 130
rect 42 129 57 130
rect 68 129 78 130
rect 89 129 113 130
rect 9 125 20 128
rect 8 122 20 125
rect 23 127 36 128
rect 41 128 57 129
rect 66 128 79 129
rect 90 128 114 129
rect 165 128 166 130
rect 23 124 35 127
rect 41 125 56 128
rect 64 127 81 128
rect 90 127 116 128
rect 63 126 82 127
rect 91 126 117 127
rect 62 125 83 126
rect 92 125 118 126
rect 22 123 35 124
rect 40 123 55 125
rect 61 124 84 125
rect 92 124 119 125
rect 165 124 166 126
rect 172 124 174 130
rect 182 128 183 130
rect 190 128 193 129
rect 191 126 192 128
rect 193 126 197 127
rect 198 126 199 127
rect 182 124 183 126
rect 191 125 199 126
rect 191 124 200 125
rect 61 123 85 124
rect 93 123 120 124
rect 165 123 168 124
rect 172 123 175 124
rect 181 123 183 124
rect 8 117 19 122
rect 22 120 34 123
rect 40 121 54 123
rect 60 122 85 123
rect 94 122 121 123
rect 60 121 86 122
rect 94 121 122 122
rect 39 120 54 121
rect 22 117 33 120
rect 39 117 53 120
rect 59 119 87 121
rect 95 120 123 121
rect 95 119 124 120
rect 8 112 18 117
rect 22 115 32 117
rect 38 116 53 117
rect 58 117 88 119
rect 96 118 124 119
rect 165 119 183 123
rect 191 122 192 123
rect 191 121 193 122
rect 165 118 167 119
rect 96 117 125 118
rect 165 117 166 118
rect 182 117 183 119
rect 191 117 192 118
rect 198 117 199 118
rect 58 116 89 117
rect 38 115 52 116
rect 22 114 31 115
rect 37 114 52 115
rect 21 113 31 114
rect 8 109 17 112
rect 21 110 30 113
rect 36 112 52 114
rect 57 115 89 116
rect 97 116 126 117
rect 57 113 90 115
rect 97 114 127 116
rect 191 115 200 117
rect 191 114 192 115
rect 35 111 52 112
rect 34 110 52 111
rect 56 112 85 113
rect 88 112 90 113
rect 98 113 128 114
rect 98 112 129 113
rect 56 111 80 112
rect 98 111 130 112
rect 56 110 76 111
rect 99 110 131 111
rect 191 110 193 111
rect 195 110 198 111
rect 20 109 30 110
rect 31 109 51 110
rect 8 106 16 109
rect 20 107 51 109
rect 56 109 74 110
rect 99 109 132 110
rect 56 108 72 109
rect 99 108 133 109
rect 55 107 71 108
rect 99 107 135 108
rect 174 107 176 109
rect 190 107 192 110
rect 194 109 199 110
rect 194 108 197 109
rect 193 107 196 108
rect 199 107 200 109
rect 9 105 16 106
rect 8 104 16 105
rect 19 105 50 107
rect 55 106 70 107
rect 100 106 136 107
rect 165 106 170 107
rect 55 105 69 106
rect 83 105 96 106
rect 100 105 114 106
rect 115 105 138 106
rect 19 104 49 105
rect 55 104 68 105
rect 80 104 115 105
rect 117 104 138 105
rect 165 105 169 106
rect 165 104 168 105
rect 174 104 183 107
rect 191 106 195 107
rect 198 106 200 107
rect 192 105 194 106
rect 197 105 199 106
rect 9 102 16 104
rect 18 103 48 104
rect 18 102 47 103
rect 54 102 67 104
rect 78 103 115 104
rect 121 103 134 104
rect 164 103 167 104
rect 174 103 184 104
rect 76 102 116 103
rect 9 101 17 102
rect 18 101 46 102
rect 54 101 66 102
rect 74 101 117 102
rect 9 100 44 101
rect 53 100 66 101
rect 73 100 118 101
rect 9 99 42 100
rect 9 98 40 99
rect 52 98 66 100
rect 72 99 119 100
rect 164 99 166 103
rect 174 101 176 103
rect 174 100 175 101
rect 182 99 184 103
rect 198 101 200 102
rect 73 98 120 99
rect 10 97 39 98
rect 51 97 66 98
rect 75 97 122 98
rect 151 97 152 98
rect 10 96 37 97
rect 49 96 66 97
rect 77 96 124 97
rect 149 96 152 97
rect 165 97 167 99
rect 181 98 184 99
rect 191 100 195 101
rect 197 100 200 101
rect 191 99 199 100
rect 181 97 183 98
rect 165 96 168 97
rect 179 96 183 97
rect 10 95 36 96
rect 48 95 66 96
rect 79 95 126 96
rect 146 95 152 96
rect 166 95 170 96
rect 177 95 183 96
rect 191 97 192 99
rect 194 98 198 99
rect 195 97 196 98
rect 199 97 200 98
rect 191 95 200 97
rect 10 94 35 95
rect 46 94 67 95
rect 82 94 129 95
rect 142 94 151 95
rect 166 94 182 95
rect 191 94 192 95
rect 10 93 34 94
rect 43 93 68 94
rect 84 93 151 94
rect 167 93 181 94
rect 11 92 33 93
rect 41 92 71 93
rect 85 92 150 93
rect 168 92 180 93
rect 11 90 32 92
rect 40 91 74 92
rect 87 91 150 92
rect 169 91 179 92
rect 38 90 76 91
rect 88 90 149 91
rect 172 90 176 91
rect 192 90 193 91
rect 197 90 199 91
rect 11 89 31 90
rect 37 89 78 90
rect 89 89 107 90
rect 109 89 149 90
rect 191 89 193 90
rect 12 87 30 89
rect 36 88 80 89
rect 90 88 107 89
rect 110 88 148 89
rect 165 88 166 89
rect 191 88 192 89
rect 36 87 81 88
rect 91 87 108 88
rect 112 87 147 88
rect 165 87 167 88
rect 194 87 196 90
rect 198 89 200 90
rect 199 87 200 88
rect 12 86 29 87
rect 35 86 82 87
rect 12 85 20 86
rect 25 85 28 86
rect 35 85 83 86
rect 92 85 109 87
rect 113 86 146 87
rect 165 86 183 87
rect 191 86 200 87
rect 115 85 145 86
rect 165 85 184 86
rect 191 85 199 86
rect 12 83 19 85
rect 35 84 84 85
rect 93 84 110 85
rect 116 84 144 85
rect 165 84 167 85
rect 176 84 183 85
rect 191 84 192 85
rect 198 84 200 85
rect 35 83 85 84
rect 94 83 110 84
rect 117 83 143 84
rect 12 81 18 83
rect 35 82 86 83
rect 94 82 111 83
rect 119 82 141 83
rect 165 82 166 84
rect 175 83 182 84
rect 174 82 180 83
rect 35 81 41 82
rect 42 81 87 82
rect 95 81 112 82
rect 121 81 140 82
rect 173 81 179 82
rect 12 77 17 81
rect 24 80 27 81
rect 35 80 38 81
rect 50 80 88 81
rect 96 80 112 81
rect 124 80 138 81
rect 172 80 178 81
rect 22 79 29 80
rect 53 79 89 80
rect 96 79 113 80
rect 128 79 134 80
rect 170 79 177 80
rect 191 79 193 80
rect 22 78 30 79
rect 56 78 90 79
rect 11 74 17 77
rect 21 76 31 78
rect 58 77 90 78
rect 97 78 114 79
rect 169 78 175 79
rect 191 78 196 79
rect 97 77 115 78
rect 168 77 174 78
rect 195 77 198 78
rect 59 76 91 77
rect 98 76 116 77
rect 167 76 173 77
rect 10 73 17 74
rect 20 75 32 76
rect 61 75 92 76
rect 98 75 117 76
rect 166 75 172 76
rect 182 75 183 77
rect 196 76 200 77
rect 20 74 33 75
rect 40 74 48 75
rect 62 74 92 75
rect 99 74 118 75
rect 165 74 171 75
rect 181 74 183 75
rect 20 73 35 74
rect 36 73 51 74
rect 63 73 93 74
rect 99 73 120 74
rect 10 71 18 73
rect 21 72 52 73
rect 65 72 93 73
rect 100 72 122 73
rect 165 72 183 74
rect 191 75 192 76
rect 193 75 199 76
rect 191 74 196 75
rect 191 73 194 74
rect 191 72 192 73
rect 21 71 54 72
rect 10 69 19 71
rect 21 70 55 71
rect 66 70 94 72
rect 100 71 125 72
rect 135 71 139 72
rect 165 71 167 72
rect 181 71 183 72
rect 101 70 138 71
rect 11 68 19 69
rect 22 69 57 70
rect 67 69 95 70
rect 22 68 58 69
rect 68 68 95 69
rect 102 69 137 70
rect 165 69 166 71
rect 182 70 183 71
rect 102 68 136 69
rect 12 67 20 68
rect 23 67 60 68
rect 69 67 95 68
rect 103 67 135 68
rect 12 66 19 67
rect 14 65 19 66
rect 23 66 61 67
rect 23 65 62 66
rect 70 65 96 67
rect 104 66 135 67
rect 165 67 166 68
rect 165 66 167 67
rect 191 66 199 68
rect 104 65 134 66
rect 165 65 170 66
rect 177 65 178 66
rect 191 65 192 66
rect 198 65 200 66
rect 16 64 17 65
rect 23 64 63 65
rect 22 63 64 64
rect 71 63 97 65
rect 105 64 133 65
rect 106 63 133 64
rect 165 64 181 65
rect 165 63 182 64
rect 21 62 65 63
rect 20 61 66 62
rect 72 61 98 63
rect 107 62 132 63
rect 165 62 167 63
rect 179 62 183 63
rect 109 61 131 62
rect 20 60 31 61
rect 32 60 66 61
rect 73 60 99 61
rect 110 60 130 61
rect 165 60 166 62
rect 180 61 183 62
rect 19 59 31 60
rect 19 55 32 59
rect 33 58 67 60
rect 73 59 100 60
rect 112 59 128 60
rect 74 58 100 59
rect 114 58 127 59
rect 34 56 68 58
rect 74 57 101 58
rect 117 57 125 58
rect 181 57 184 61
rect 191 60 200 61
rect 191 59 194 60
rect 195 59 200 60
rect 195 58 198 59
rect 194 57 197 58
rect 74 56 103 57
rect 165 56 166 57
rect 180 56 184 57
rect 193 56 196 57
rect 35 55 69 56
rect 20 53 33 55
rect 36 54 69 55
rect 75 55 105 56
rect 165 55 167 56
rect 179 55 183 56
rect 75 54 107 55
rect 37 53 69 54
rect 76 53 113 54
rect 165 53 183 55
rect 191 55 195 56
rect 191 54 194 55
rect 198 54 200 55
rect 191 53 200 54
rect 21 52 33 53
rect 39 52 70 53
rect 76 52 118 53
rect 165 52 182 53
rect 23 51 34 52
rect 40 51 55 52
rect 57 51 70 52
rect 24 50 34 51
rect 38 50 54 51
rect 26 49 35 50
rect 27 48 35 49
rect 37 49 54 50
rect 58 50 70 51
rect 77 51 117 52
rect 165 51 180 52
rect 77 50 116 51
rect 165 50 176 51
rect 37 48 55 49
rect 28 47 36 48
rect 37 47 56 48
rect 58 47 71 50
rect 78 49 115 50
rect 78 48 114 49
rect 165 48 166 50
rect 191 48 193 49
rect 79 47 113 48
rect 191 47 199 48
rect 29 46 56 47
rect 30 44 57 46
rect 31 43 57 44
rect 32 41 57 43
rect 59 44 72 47
rect 80 46 112 47
rect 198 46 200 47
rect 81 45 110 46
rect 165 45 166 46
rect 199 45 200 46
rect 82 44 108 45
rect 165 44 167 45
rect 198 44 200 45
rect 59 41 73 44
rect 84 43 106 44
rect 165 43 168 44
rect 191 43 192 44
rect 197 43 200 44
rect 86 42 104 43
rect 165 42 169 43
rect 191 42 199 43
rect 89 41 100 42
rect 165 41 171 42
rect 33 40 58 41
rect 34 38 58 40
rect 35 36 58 38
rect 60 40 72 41
rect 165 40 166 41
rect 169 40 173 41
rect 182 40 183 42
rect 191 41 198 42
rect 60 39 70 40
rect 171 39 183 40
rect 60 38 68 39
rect 173 38 183 39
rect 60 37 66 38
rect 171 37 183 38
rect 60 36 64 37
rect 165 36 166 37
rect 169 36 183 37
rect 36 35 57 36
rect 36 34 44 35
rect 45 34 57 35
rect 165 35 183 36
rect 165 34 174 35
rect 37 32 45 34
rect 46 33 56 34
rect 165 33 172 34
rect 182 33 183 35
rect 47 32 55 33
rect 165 32 170 33
rect 38 30 46 32
rect 48 31 53 32
rect 165 31 168 32
rect 49 30 51 31
rect 165 30 167 31
rect 39 29 46 30
rect 165 29 166 30
rect 40 28 46 29
rect 42 27 44 28
rect 165 25 166 27
rect 182 26 183 27
rect 181 25 183 26
rect 165 23 167 25
rect 180 24 183 25
rect 179 23 183 24
rect 165 22 168 23
rect 178 22 183 23
rect 165 21 169 22
rect 176 21 183 22
rect 165 19 166 21
rect 167 20 170 21
rect 175 20 182 21
rect 169 19 171 20
rect 173 19 181 20
rect 170 18 179 19
rect 171 17 178 18
rect 165 16 166 17
rect 172 16 176 17
rect 182 16 183 17
rect 165 15 167 16
rect 173 15 175 16
rect 181 15 183 16
rect 165 11 183 15
rect 165 10 167 11
rect 181 10 183 11
rect 165 9 166 10
rect 182 9 183 10
<< end >>
