magic
tech scmos
magscale 1 2
timestamp 1727918344
<< nwell >>
rect -13 134 252 252
rect -13 132 51 134
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 34
rect 52 14 56 34
rect 72 14 76 34
rect 82 14 86 34
rect 104 14 108 34
rect 148 14 152 34
rect 158 14 162 34
rect 178 14 182 34
rect 188 14 192 34
rect 208 14 212 54
<< ptransistor >>
rect 20 146 24 226
rect 40 186 44 226
rect 52 186 56 226
rect 72 186 76 226
rect 84 186 88 226
rect 104 186 108 226
rect 148 186 152 226
rect 158 186 162 226
rect 178 206 182 226
rect 188 206 192 226
rect 208 146 212 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 34 35 54
rect 197 34 208 54
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 52 34
rect 56 14 58 34
rect 70 14 72 34
rect 76 14 82 34
rect 86 14 88 34
rect 100 14 104 34
rect 108 14 110 34
rect 146 14 148 34
rect 152 14 158 34
rect 162 14 164 34
rect 176 14 178 34
rect 182 14 188 34
rect 192 14 194 34
rect 206 14 208 34
rect 212 14 214 54
<< pdiffusion >>
rect 18 146 20 226
rect 24 186 26 226
rect 38 186 40 226
rect 44 186 52 226
rect 56 186 58 226
rect 70 186 72 226
rect 76 186 84 226
rect 88 186 90 226
rect 102 186 104 226
rect 108 186 110 226
rect 146 186 148 226
rect 152 186 158 226
rect 162 206 164 226
rect 176 206 178 226
rect 182 206 188 226
rect 192 206 194 226
rect 206 206 208 226
rect 162 186 172 206
rect 24 146 35 186
rect 197 146 208 206
rect 212 146 214 226
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 34
rect 58 14 70 34
rect 88 14 100 34
rect 110 14 122 34
rect 134 14 146 34
rect 164 14 176 34
rect 194 14 206 34
rect 214 14 226 54
<< pdcontact >>
rect 6 146 18 226
rect 26 186 38 226
rect 58 186 70 226
rect 90 186 102 226
rect 110 186 122 226
rect 134 186 146 226
rect 164 206 176 226
rect 194 206 206 226
rect 214 146 226 226
<< psubstratepcontact >>
rect -6 -6 246 6
<< nsubstratencontact >>
rect -6 234 246 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 52 226 56 230
rect 72 226 76 230
rect 84 226 88 230
rect 104 226 108 230
rect 148 226 152 230
rect 158 226 162 230
rect 178 226 182 230
rect 188 226 192 230
rect 208 226 212 230
rect 20 137 24 146
rect 12 131 24 137
rect 12 76 16 131
rect 40 123 44 186
rect 52 142 56 186
rect 72 180 76 186
rect 84 180 88 186
rect 64 130 76 134
rect 36 111 44 123
rect 12 64 19 76
rect 20 54 24 64
rect 40 34 44 111
rect 52 34 56 60
rect 72 34 76 130
rect 84 54 88 168
rect 104 128 108 186
rect 148 182 152 186
rect 82 52 88 54
rect 82 40 84 52
rect 82 34 86 40
rect 104 34 108 116
rect 116 180 152 182
rect 128 178 152 180
rect 158 177 162 186
rect 156 172 162 177
rect 116 42 120 168
rect 134 50 138 148
rect 156 70 160 172
rect 178 164 182 206
rect 180 152 182 164
rect 188 143 192 206
rect 158 60 160 70
rect 180 139 192 143
rect 180 81 184 139
rect 158 58 182 60
rect 146 54 182 58
rect 134 46 162 50
rect 116 38 152 42
rect 148 34 152 38
rect 158 34 162 46
rect 178 34 182 54
rect 188 34 192 69
rect 208 54 212 146
rect 20 10 24 14
rect 40 10 44 14
rect 52 10 56 14
rect 72 10 76 14
rect 82 10 86 14
rect 104 10 108 14
rect 148 10 152 14
rect 158 10 162 14
rect 178 10 182 14
rect 188 10 192 14
rect 208 10 212 14
<< polycontact >>
rect 64 168 76 180
rect 84 168 96 180
rect 52 130 64 142
rect 24 111 36 123
rect 19 64 31 76
rect 52 60 64 72
rect 96 116 108 128
rect 84 40 96 52
rect 116 168 128 180
rect 134 148 146 160
rect 168 152 180 164
rect 146 58 158 70
rect 196 112 208 124
rect 180 69 192 81
<< metal1 >>
rect -6 246 246 248
rect -6 232 246 234
rect 26 226 38 232
rect 90 226 102 232
rect 134 226 146 232
rect 194 226 206 232
rect 46 186 58 194
rect 164 186 176 206
rect 46 182 57 186
rect 110 180 122 186
rect 96 172 116 180
rect 64 162 76 168
rect 146 152 168 160
rect 6 142 18 146
rect 134 142 140 148
rect 6 134 52 142
rect 6 54 12 134
rect 64 134 140 142
rect 57 116 96 124
rect 176 112 196 120
rect 31 74 63 76
rect 214 83 222 146
rect 77 74 103 76
rect 31 72 103 74
rect 31 68 52 72
rect 64 69 103 72
rect 117 70 158 76
rect 117 69 146 70
rect 64 68 146 69
rect 192 69 203 81
rect 217 69 222 83
rect 214 54 222 69
rect 96 40 118 48
rect 46 34 57 40
rect 110 34 118 40
rect 46 27 58 34
rect 162 28 164 34
rect 26 8 38 14
rect 88 8 100 14
rect 134 8 146 14
rect 194 8 206 14
rect -6 6 246 8
rect -6 -8 246 -6
<< m2contact >>
rect 43 168 57 182
rect 162 172 176 186
rect 63 148 77 162
rect 23 97 37 111
rect 43 110 57 124
rect 162 110 176 124
rect 63 74 77 88
rect 103 69 117 83
rect 203 69 217 83
rect 43 40 57 54
rect 162 34 176 48
<< metal2 >>
rect 47 124 54 168
rect 23 83 37 97
rect 47 54 54 110
rect 67 88 76 148
rect 162 124 170 172
rect 103 83 117 97
rect 162 48 170 110
rect 203 83 217 97
<< m2p >>
rect 23 83 37 97
rect 103 83 117 97
rect 203 83 217 97
<< labels >>
rlabel metal1 -6 -8 246 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 246 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 23 83 37 97 0 D
port 0 nsew signal input
rlabel metal2 203 83 217 97 0 Q
port 2 nsew signal output
rlabel metal2 103 83 117 97 0 CLK
port 1 nsew clock input
<< properties >>
string FIXED_BBOX 0 0 240 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
