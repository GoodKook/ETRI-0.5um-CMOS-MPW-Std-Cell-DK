magic
tech scmos
magscale 1 6
timestamp 1555589239
<< checkpaint >>
rect -140 -1950 2540 5180
<< metal2 >>
rect 2260 5032 2324 5060
use CMD_TR  CMD_TR_0
timestamp 1555589239
transform 1 0 1524 0 1 4798
box 10 -35 254 178
use DOUBLE_GUARD  DOUBLE_GUARD_0
timestamp 1555589239
transform 1 0 0 0 1 1660
box -20 -20 2419 500
use GUARD  GUARD_0
timestamp 1555589239
transform 1 0 0 0 1 4220
box -20 -20 2419 792
use INV2  INV2_0
timestamp 1555589239
transform 1 0 1914 0 1 4314
box -2 -42 426 646
use INV  INV_0
timestamp 1555589239
transform 1 0 1738 0 1 4314
box -2 -42 186 614
use METAL_RING  METAL_RING_0
timestamp 1555589239
transform 1 0 0 0 1 0
box 0 0 2400 5012
use NDRV  NDRV_0
timestamp 1555589239
transform 1 0 0 0 1 0
box 0 0 2400 1560
use PAD_80  PAD_80_0
timestamp 1555589239
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_PIC  PAD_METAL_PIC_0
timestamp 1555589239
transform 1 0 0 0 1 0
box 0 0 2400 5060
use PDRV  PDRV_0
timestamp 1555589239
transform 1 0 0 0 1 2260
box -20 -20 2420 1580
use SINGLE_GUARD  SINGLE_GUARD_0
timestamp 1555589239
transform 1 0 0 0 1 3920
box 0 0 2400 200
<< labels >>
flabel m2p s 2292 5060 2292 5060 0 FreeSans 400 0 0 0 Y
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 PAD
flabel m3p s 0 3018 0 3018 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4339 0 4339 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4788 0 4788 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 752 0 752 0 FreeSans 1000 0 0 0 VSS
<< end >>
