magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -58 -120 2457 5180
<< metal1 >>
rect 433 4706 985 4874
rect 433 4369 977 4486
rect 62 1960 102 2160
rect 2297 1660 2337 1860
<< metal2 >>
rect 433 4766 985 5060
rect 1076 4616 2020 5060
rect 380 4340 2020 4616
rect 250 2354 290 3774
rect 62 1924 102 2160
rect 62 1891 290 1924
rect 250 71 290 1891
rect 380 0 580 4340
rect 670 2354 710 3774
rect 730 2354 770 3774
rect 670 71 710 1491
rect 730 71 770 1491
rect 860 0 1060 4340
rect 1150 2354 1190 3774
rect 1210 2354 1250 3774
rect 1150 71 1190 1491
rect 1210 71 1250 1491
rect 1340 0 1540 4340
rect 1630 2354 1670 3774
rect 1690 2354 1730 3774
rect 1630 71 1670 1491
rect 1690 71 1730 1491
rect 1820 0 2020 4340
rect 2110 1937 2150 3774
rect 2110 1900 2337 1937
rect 2297 1660 2337 1900
rect 2110 71 2150 1491
use M2_M1_CDNS_704676826050  M2_M1_CDNS_704676826050_0
timestamp 1537935238
transform 1 0 2317 0 1 1760
box -20 -96 20 96
use M2_M1_CDNS_704676826050  M2_M1_CDNS_704676826050_1
timestamp 1537935238
transform 1 0 82 0 1 2060
box -20 -96 20 96
use p2res_CDNS_704676826058  p2res_CDNS_704676826058_0
array 0 0 0 0 9 56
timestamp 1537935238
transform 0 -1 993 1 0 4446
box 16 16 264 56
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_0
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_1
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_2
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_3
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_4
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 202
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_5
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_6
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 202
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_7
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_8
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_9
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 682
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_10
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_11
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 682
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_12
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 1162
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_13
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_14
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_15
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_16
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 1162
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_17
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_18
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_19
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 1162
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_20
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_21
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 202
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_22
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 202
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_23
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_24
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_25
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 682
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_26
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_27
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_28
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 682
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_29
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 621
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_30
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_31
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 1162
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_32
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_33
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 141
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_34
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_35
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 1101
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_36
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_37
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_38
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_39
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 2965
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_40
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_41
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_42
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_43
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_44
array 0 16 32 0 2 32
timestamp 1537935238
transform 1 0 433 0 1 4766
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_45
array 0 16 32 0 2 32
timestamp 1537935238
transform 1 0 433 0 1 4369
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_46
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 3445
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_47
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_48
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 3445
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_49
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 2965
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_50
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 2965
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_51
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_52
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 3445
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_53
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_54
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_55
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 2965
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_56
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_57
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 2904
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_58
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_59
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_60
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 3445
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_61
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 3384
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_62
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1822 0 1 2485
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_63
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_64
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_65
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 862 0 1 2485
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_66
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_67
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_68
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 382 0 1 2485
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_69
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_70
array 0 3 52 0 3 53
timestamp 1537935238
transform 1 0 1342 0 1 2485
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_71
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_72
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 2424
box 0 0 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_73
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 2424
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_0
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_1
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_2
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_3
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_4
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_5
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_6
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_7
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_8
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_9
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_10
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_11
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_12
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_13
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_14
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_15
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_16
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_17
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_18
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_19
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 593
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_20
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_21
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_22
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 1073
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_23
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 113
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_24
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_25
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_26
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_27
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_28
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_29
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_30
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_31
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_32
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_33
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_34
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_35
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_36
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_37
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 3356
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_38
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_39
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 2876
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_40
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1210 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_41
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1690 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_42
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1150 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_43
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 730 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_44
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 670 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_45
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 1630 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_46
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 2110 0 1 2396
box 0 0 40 40
use via2_array_CDNS_704676826052  via2_array_CDNS_704676826052_47
array 0 0 0 0 6 56
timestamp 1537935238
transform 1 0 250 0 1 2396
box 0 0 40 40
<< end >>
